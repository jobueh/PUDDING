VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DAC2U128OUT4IN
CLASS BLOCK ;
  FOREIGN DAC2U128OUT4IN ;
  ORIGIN 2.210 5.110 ;
  SIZE 134.420 BY 26.590 ;
PIN ON[64]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 128.130 18.805 128.420 21.280 ;
    END
  END ON[64]
PIN ONB[64]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 127.580 18.805 127.870 21.280 ;
    END
  END ONB[64]
PIN ON[65]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 126.130 18.805 126.420 21.280 ;
    END
  END ON[65]
PIN ONB[65]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 125.580 18.805 125.870 21.280 ;
    END
  END ONB[65]
PIN ON[66]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 124.130 18.805 124.420 21.280 ;
    END
  END ON[66]
PIN ONB[66]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 123.580 18.805 123.870 21.280 ;
    END
  END ONB[66]
PIN ON[67]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 122.130 18.805 122.420 21.280 ;
    END
  END ON[67]
PIN ONB[67]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 121.580 18.805 121.870 21.280 ;
    END
  END ONB[67]
PIN ON[68]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 120.130 18.805 120.420 21.280 ;
    END
  END ON[68]
PIN ONB[68]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 119.580 18.805 119.870 21.280 ;
    END
  END ONB[68]
PIN ON[69]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.130 18.805 118.420 21.280 ;
    END
  END ON[69]
PIN ONB[69]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.580 18.805 117.870 21.280 ;
    END
  END ONB[69]
PIN ON[70]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 116.130 18.805 116.420 21.280 ;
    END
  END ON[70]
PIN ONB[70]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 115.580 18.805 115.870 21.280 ;
    END
  END ONB[70]
PIN ON[71]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 114.130 18.805 114.420 21.280 ;
    END
  END ON[71]
PIN ONB[71]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 113.580 18.805 113.870 21.280 ;
    END
  END ONB[71]
PIN ON[72]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 112.130 18.805 112.420 21.280 ;
    END
  END ON[72]
PIN ONB[72]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 111.580 18.805 111.870 21.280 ;
    END
  END ONB[72]
PIN ON[73]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.130 18.805 110.420 21.280 ;
    END
  END ON[73]
PIN ONB[73]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 109.580 18.805 109.870 21.280 ;
    END
  END ONB[73]
PIN ON[74]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 108.130 18.805 108.420 21.280 ;
    END
  END ON[74]
PIN ONB[74]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 107.580 18.805 107.870 21.280 ;
    END
  END ONB[74]
PIN ON[75]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 106.130 18.805 106.420 21.280 ;
    END
  END ON[75]
PIN ONB[75]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 105.580 18.805 105.870 21.280 ;
    END
  END ONB[75]
PIN ON[76]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 104.130 18.805 104.420 21.280 ;
    END
  END ON[76]
PIN ONB[76]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 103.580 18.805 103.870 21.280 ;
    END
  END ONB[76]
PIN ON[77]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 102.130 18.805 102.420 21.280 ;
    END
  END ON[77]
PIN ONB[77]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 101.580 18.805 101.870 21.280 ;
    END
  END ONB[77]
PIN ON[78]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 100.130 18.805 100.420 21.280 ;
    END
  END ON[78]
PIN ONB[78]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 99.580 18.805 99.870 21.280 ;
    END
  END ONB[78]
PIN ON[79]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 98.130 18.805 98.420 21.280 ;
    END
  END ON[79]
PIN ONB[79]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 97.580 18.805 97.870 21.280 ;
    END
  END ONB[79]
PIN ON[80]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 96.130 18.805 96.420 21.280 ;
    END
  END ON[80]
PIN ONB[80]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 95.580 18.805 95.870 21.280 ;
    END
  END ONB[80]
PIN ON[81]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 94.130 18.805 94.420 21.280 ;
    END
  END ON[81]
PIN ONB[81]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 93.580 18.805 93.870 21.280 ;
    END
  END ONB[81]
PIN ON[82]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 92.130 18.805 92.420 21.280 ;
    END
  END ON[82]
PIN ONB[82]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 91.580 18.805 91.870 21.280 ;
    END
  END ONB[82]
PIN ON[83]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 90.130 18.805 90.420 21.280 ;
    END
  END ON[83]
PIN ONB[83]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 89.580 18.805 89.870 21.280 ;
    END
  END ONB[83]
PIN ON[84]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 88.130 18.805 88.420 21.280 ;
    END
  END ON[84]
PIN ONB[84]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 87.580 18.805 87.870 21.280 ;
    END
  END ONB[84]
PIN ON[85]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 86.130 18.805 86.420 21.280 ;
    END
  END ON[85]
PIN ONB[85]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 85.580 18.805 85.870 21.280 ;
    END
  END ONB[85]
PIN ON[86]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 84.130 18.805 84.420 21.280 ;
    END
  END ON[86]
PIN ONB[86]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 83.580 18.805 83.870 21.280 ;
    END
  END ONB[86]
PIN ON[87]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 82.130 18.805 82.420 21.280 ;
    END
  END ON[87]
PIN ONB[87]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 81.580 18.805 81.870 21.280 ;
    END
  END ONB[87]
PIN ON[88]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 80.130 18.805 80.420 21.280 ;
    END
  END ON[88]
PIN ONB[88]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 79.580 18.805 79.870 21.280 ;
    END
  END ONB[88]
PIN ON[89]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 78.130 18.805 78.420 21.280 ;
    END
  END ON[89]
PIN ONB[89]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.580 18.805 77.870 21.280 ;
    END
  END ONB[89]
PIN ON[90]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 76.130 18.805 76.420 21.280 ;
    END
  END ON[90]
PIN ONB[90]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 75.580 18.805 75.870 21.280 ;
    END
  END ONB[90]
PIN ON[91]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 74.130 18.805 74.420 21.280 ;
    END
  END ON[91]
PIN ONB[91]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 73.580 18.805 73.870 21.280 ;
    END
  END ONB[91]
PIN ON[92]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 72.130 18.805 72.420 21.280 ;
    END
  END ON[92]
PIN ONB[92]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 71.580 18.805 71.870 21.280 ;
    END
  END ONB[92]
PIN ON[93]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.130 18.805 70.420 21.280 ;
    END
  END ON[93]
PIN ONB[93]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.580 18.805 69.870 21.280 ;
    END
  END ONB[93]
PIN ON[94]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.130 18.805 68.420 21.280 ;
    END
  END ON[94]
PIN ONB[94]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 67.580 18.805 67.870 21.280 ;
    END
  END ONB[94]
PIN ON[95]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 66.130 18.805 66.420 21.280 ;
    END
  END ON[95]
PIN ONB[95]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 65.580 18.805 65.870 21.280 ;
    END
  END ONB[95]
PIN EN[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 130.130 18.805 130.420 21.280 ;
    END
  END EN[2]
PIN ENB[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 129.580 18.805 129.870 21.280 ;
    END
  END ENB[2]
PIN ON[97]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 62.130 18.805 62.420 21.280 ;
    END
  END ON[97]
PIN ONB[97]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 61.580 18.805 61.870 21.280 ;
    END
  END ONB[97]
PIN ON[98]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 60.130 18.805 60.420 21.280 ;
    END
  END ON[98]
PIN ONB[98]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 59.580 18.805 59.870 21.280 ;
    END
  END ONB[98]
PIN ON[99]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 58.130 18.805 58.420 21.280 ;
    END
  END ON[99]
PIN ONB[99]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.580 18.805 57.870 21.280 ;
    END
  END ONB[99]
PIN ON[100]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 56.130 18.805 56.420 21.280 ;
    END
  END ON[100]
PIN ONB[100]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 55.580 18.805 55.870 21.280 ;
    END
  END ONB[100]
PIN ON[101]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 54.130 18.805 54.420 21.280 ;
    END
  END ON[101]
PIN ONB[101]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 53.580 18.805 53.870 21.280 ;
    END
  END ONB[101]
PIN ON[102]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 52.130 18.805 52.420 21.280 ;
    END
  END ON[102]
PIN ONB[102]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 51.580 18.805 51.870 21.280 ;
    END
  END ONB[102]
PIN ON[103]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 50.130 18.805 50.420 21.280 ;
    END
  END ON[103]
PIN ONB[103]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 49.580 18.805 49.870 21.280 ;
    END
  END ONB[103]
PIN ON[104]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 48.130 18.805 48.420 21.280 ;
    END
  END ON[104]
PIN ONB[104]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 47.580 18.805 47.870 21.280 ;
    END
  END ONB[104]
PIN ON[105]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 46.130 18.805 46.420 21.280 ;
    END
  END ON[105]
PIN ONB[105]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 45.580 18.805 45.870 21.280 ;
    END
  END ONB[105]
PIN ON[106]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 44.130 18.805 44.420 21.280 ;
    END
  END ON[106]
PIN ONB[106]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 43.580 18.805 43.870 21.280 ;
    END
  END ONB[106]
PIN ON[107]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 42.130 18.805 42.420 21.280 ;
    END
  END ON[107]
PIN ONB[107]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 41.580 18.805 41.870 21.280 ;
    END
  END ONB[107]
PIN ON[108]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 40.130 18.805 40.420 21.280 ;
    END
  END ON[108]
PIN ONB[108]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 39.580 18.805 39.870 21.280 ;
    END
  END ONB[108]
PIN ON[109]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 38.130 18.805 38.420 21.280 ;
    END
  END ON[109]
PIN ONB[109]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 37.580 18.805 37.870 21.280 ;
    END
  END ONB[109]
PIN ON[110]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.130 18.805 36.420 21.280 ;
    END
  END ON[110]
PIN ONB[110]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 35.580 18.805 35.870 21.280 ;
    END
  END ONB[110]
PIN ON[111]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 34.130 18.805 34.420 21.280 ;
    END
  END ON[111]
PIN ONB[111]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 33.580 18.805 33.870 21.280 ;
    END
  END ONB[111]
PIN ON[112]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 32.130 18.805 32.420 21.280 ;
    END
  END ON[112]
PIN ONB[112]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 31.580 18.805 31.870 21.280 ;
    END
  END ONB[112]
PIN ON[113]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.130 18.805 30.420 21.280 ;
    END
  END ON[113]
PIN ONB[113]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 29.580 18.805 29.870 21.280 ;
    END
  END ONB[113]
PIN ON[114]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.130 18.805 28.420 21.280 ;
    END
  END ON[114]
PIN ONB[114]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 27.580 18.805 27.870 21.280 ;
    END
  END ONB[114]
PIN ON[115]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 26.130 18.805 26.420 21.280 ;
    END
  END ON[115]
PIN ONB[115]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.580 18.805 25.870 21.280 ;
    END
  END ONB[115]
PIN ON[116]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 24.130 18.805 24.420 21.280 ;
    END
  END ON[116]
PIN ONB[116]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 23.580 18.805 23.870 21.280 ;
    END
  END ONB[116]
PIN ON[117]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 22.130 18.805 22.420 21.280 ;
    END
  END ON[117]
PIN ONB[117]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.580 18.805 21.870 21.280 ;
    END
  END ONB[117]
PIN ON[118]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 20.130 18.805 20.420 21.280 ;
    END
  END ON[118]
PIN ONB[118]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 19.580 18.805 19.870 21.280 ;
    END
  END ONB[118]
PIN ON[119]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 18.130 18.805 18.420 21.280 ;
    END
  END ON[119]
PIN ONB[119]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.580 18.805 17.870 21.280 ;
    END
  END ONB[119]
PIN ON[120]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.130 18.805 16.420 21.280 ;
    END
  END ON[120]
PIN ONB[120]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 15.580 18.805 15.870 21.280 ;
    END
  END ONB[120]
PIN ON[121]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.130 18.805 14.420 21.280 ;
    END
  END ON[121]
PIN ONB[121]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.580 18.805 13.870 21.280 ;
    END
  END ONB[121]
PIN ON[122]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.130 18.805 12.420 21.280 ;
    END
  END ON[122]
PIN ONB[122]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.580 18.805 11.870 21.280 ;
    END
  END ONB[122]
PIN ON[123]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.130 18.805 10.420 21.280 ;
    END
  END ON[123]
PIN ONB[123]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.580 18.805 9.870 21.280 ;
    END
  END ONB[123]
PIN ON[124]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 8.130 18.805 8.420 21.280 ;
    END
  END ON[124]
PIN ONB[124]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.580 18.805 7.870 21.280 ;
    END
  END ONB[124]
PIN ON[125]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 6.130 18.805 6.420 21.280 ;
    END
  END ON[125]
PIN ONB[125]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.580 18.805 5.870 21.280 ;
    END
  END ONB[125]
PIN ON[126]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 4.130 18.805 4.420 21.280 ;
    END
  END ON[126]
PIN ONB[126]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.580 18.805 3.870 21.280 ;
    END
  END ONB[126]
PIN ON[127]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.130 18.805 2.420 21.280 ;
    END
  END ON[127]
PIN ONB[127]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.580 18.805 1.870 21.280 ;
    END
  END ONB[127]
PIN ON[96]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.130 18.805 64.420 21.280 ;
    END
  END ON[96]
PIN ONB[96]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.580 18.805 63.870 21.280 ;
    END
  END ONB[96]
PIN EN[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.130 18.805 0.420 21.280 ;
    END
  END EN[3]
PIN ENB[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT -0.420 18.805 -0.130 21.280 ;
    END
  END ENB[3]
PIN ON[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.580 -4.910 1.870 -2.435 ;
    END
  END ON[0]
PIN ONB[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.130 -4.910 2.420 -2.435 ;
    END
  END ONB[0]
PIN ON[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.580 -4.910 3.870 -2.435 ;
    END
  END ON[1]
PIN ONB[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 4.130 -4.910 4.420 -2.435 ;
    END
  END ONB[1]
PIN ON[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.580 -4.910 5.870 -2.435 ;
    END
  END ON[2]
PIN ONB[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 6.130 -4.910 6.420 -2.435 ;
    END
  END ONB[2]
PIN ON[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.580 -4.910 7.870 -2.435 ;
    END
  END ON[3]
PIN ONB[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 8.130 -4.910 8.420 -2.435 ;
    END
  END ONB[3]
PIN ON[4]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.580 -4.910 9.870 -2.435 ;
    END
  END ON[4]
PIN ONB[4]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.130 -4.910 10.420 -2.435 ;
    END
  END ONB[4]
PIN ON[5]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.580 -4.910 11.870 -2.435 ;
    END
  END ON[5]
PIN ONB[5]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.130 -4.910 12.420 -2.435 ;
    END
  END ONB[5]
PIN ON[6]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.580 -4.910 13.870 -2.435 ;
    END
  END ON[6]
PIN ONB[6]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.130 -4.910 14.420 -2.435 ;
    END
  END ONB[6]
PIN ON[7]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 15.580 -4.910 15.870 -2.435 ;
    END
  END ON[7]
PIN ONB[7]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.130 -4.910 16.420 -2.435 ;
    END
  END ONB[7]
PIN ON[8]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.580 -4.910 17.870 -2.435 ;
    END
  END ON[8]
PIN ONB[8]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 18.130 -4.910 18.420 -2.435 ;
    END
  END ONB[8]
PIN ON[9]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 19.580 -4.910 19.870 -2.435 ;
    END
  END ON[9]
PIN ONB[9]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 20.130 -4.910 20.420 -2.435 ;
    END
  END ONB[9]
PIN ON[10]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.580 -4.910 21.870 -2.435 ;
    END
  END ON[10]
PIN ONB[10]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 22.130 -4.910 22.420 -2.435 ;
    END
  END ONB[10]
PIN ON[11]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 23.580 -4.910 23.870 -2.435 ;
    END
  END ON[11]
PIN ONB[11]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 24.130 -4.910 24.420 -2.435 ;
    END
  END ONB[11]
PIN ON[12]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.580 -4.910 25.870 -2.435 ;
    END
  END ON[12]
PIN ONB[12]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 26.130 -4.910 26.420 -2.435 ;
    END
  END ONB[12]
PIN ON[13]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 27.580 -4.910 27.870 -2.435 ;
    END
  END ON[13]
PIN ONB[13]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.130 -4.910 28.420 -2.435 ;
    END
  END ONB[13]
PIN ON[14]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 29.580 -4.910 29.870 -2.435 ;
    END
  END ON[14]
PIN ONB[14]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.130 -4.910 30.420 -2.435 ;
    END
  END ONB[14]
PIN ON[15]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 31.580 -4.910 31.870 -2.435 ;
    END
  END ON[15]
PIN ONB[15]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 32.130 -4.910 32.420 -2.435 ;
    END
  END ONB[15]
PIN ON[16]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 33.580 -4.910 33.870 -2.435 ;
    END
  END ON[16]
PIN ONB[16]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 34.130 -4.910 34.420 -2.435 ;
    END
  END ONB[16]
PIN ON[17]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 35.580 -4.910 35.870 -2.435 ;
    END
  END ON[17]
PIN ONB[17]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.130 -4.910 36.420 -2.435 ;
    END
  END ONB[17]
PIN ON[18]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 37.580 -4.910 37.870 -2.435 ;
    END
  END ON[18]
PIN ONB[18]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 38.130 -4.910 38.420 -2.435 ;
    END
  END ONB[18]
PIN ON[19]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 39.580 -4.910 39.870 -2.435 ;
    END
  END ON[19]
PIN ONB[19]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 40.130 -4.910 40.420 -2.435 ;
    END
  END ONB[19]
PIN ON[20]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 41.580 -4.910 41.870 -2.435 ;
    END
  END ON[20]
PIN ONB[20]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 42.130 -4.910 42.420 -2.435 ;
    END
  END ONB[20]
PIN ON[21]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 43.580 -4.910 43.870 -2.435 ;
    END
  END ON[21]
PIN ONB[21]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 44.130 -4.910 44.420 -2.435 ;
    END
  END ONB[21]
PIN ON[22]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 45.580 -4.910 45.870 -2.435 ;
    END
  END ON[22]
PIN ONB[22]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 46.130 -4.910 46.420 -2.435 ;
    END
  END ONB[22]
PIN ON[23]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 47.580 -4.910 47.870 -2.435 ;
    END
  END ON[23]
PIN ONB[23]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 48.130 -4.910 48.420 -2.435 ;
    END
  END ONB[23]
PIN ON[24]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 49.580 -4.910 49.870 -2.435 ;
    END
  END ON[24]
PIN ONB[24]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 50.130 -4.910 50.420 -2.435 ;
    END
  END ONB[24]
PIN ON[25]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 51.580 -4.910 51.870 -2.435 ;
    END
  END ON[25]
PIN ONB[25]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 52.130 -4.910 52.420 -2.435 ;
    END
  END ONB[25]
PIN ON[26]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 53.580 -4.910 53.870 -2.435 ;
    END
  END ON[26]
PIN ONB[26]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 54.130 -4.910 54.420 -2.435 ;
    END
  END ONB[26]
PIN ON[27]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 55.580 -4.910 55.870 -2.435 ;
    END
  END ON[27]
PIN ONB[27]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 56.130 -4.910 56.420 -2.435 ;
    END
  END ONB[27]
PIN ON[28]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.580 -4.910 57.870 -2.435 ;
    END
  END ON[28]
PIN ONB[28]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 58.130 -4.910 58.420 -2.435 ;
    END
  END ONB[28]
PIN ON[29]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 59.580 -4.910 59.870 -2.435 ;
    END
  END ON[29]
PIN ONB[29]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 60.130 -4.910 60.420 -2.435 ;
    END
  END ONB[29]
PIN ON[30]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 61.580 -4.910 61.870 -2.435 ;
    END
  END ON[30]
PIN ONB[30]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 62.130 -4.910 62.420 -2.435 ;
    END
  END ONB[30]
PIN ON[31]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.580 -4.910 63.870 -2.435 ;
    END
  END ON[31]
PIN ONB[31]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.130 -4.910 64.420 -2.435 ;
    END
  END ONB[31]
PIN EN[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT -0.420 -4.910 -0.130 -2.435 ;
    END
  END EN[0]
PIN ENB[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.130 -4.910 0.420 -2.435 ;
    END
  END ENB[0]
PIN ON[33]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 67.580 -4.910 67.870 -2.435 ;
    END
  END ON[33]
PIN ONB[33]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.130 -4.910 68.420 -2.435 ;
    END
  END ONB[33]
PIN ON[34]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.580 -4.910 69.870 -2.435 ;
    END
  END ON[34]
PIN ONB[34]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.130 -4.910 70.420 -2.435 ;
    END
  END ONB[34]
PIN ON[35]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 71.580 -4.910 71.870 -2.435 ;
    END
  END ON[35]
PIN ONB[35]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 72.130 -4.910 72.420 -2.435 ;
    END
  END ONB[35]
PIN ON[36]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 73.580 -4.910 73.870 -2.435 ;
    END
  END ON[36]
PIN ONB[36]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 74.130 -4.910 74.420 -2.435 ;
    END
  END ONB[36]
PIN ON[37]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 75.580 -4.910 75.870 -2.435 ;
    END
  END ON[37]
PIN ONB[37]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 76.130 -4.910 76.420 -2.435 ;
    END
  END ONB[37]
PIN ON[38]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.580 -4.910 77.870 -2.435 ;
    END
  END ON[38]
PIN ONB[38]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 78.130 -4.910 78.420 -2.435 ;
    END
  END ONB[38]
PIN ON[39]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 79.580 -4.910 79.870 -2.435 ;
    END
  END ON[39]
PIN ONB[39]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 80.130 -4.910 80.420 -2.435 ;
    END
  END ONB[39]
PIN ON[40]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 81.580 -4.910 81.870 -2.435 ;
    END
  END ON[40]
PIN ONB[40]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 82.130 -4.910 82.420 -2.435 ;
    END
  END ONB[40]
PIN ON[41]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 83.580 -4.910 83.870 -2.435 ;
    END
  END ON[41]
PIN ONB[41]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 84.130 -4.910 84.420 -2.435 ;
    END
  END ONB[41]
PIN ON[42]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 85.580 -4.910 85.870 -2.435 ;
    END
  END ON[42]
PIN ONB[42]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 86.130 -4.910 86.420 -2.435 ;
    END
  END ONB[42]
PIN ON[43]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 87.580 -4.910 87.870 -2.435 ;
    END
  END ON[43]
PIN ONB[43]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 88.130 -4.910 88.420 -2.435 ;
    END
  END ONB[43]
PIN ON[44]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 89.580 -4.910 89.870 -2.435 ;
    END
  END ON[44]
PIN ONB[44]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 90.130 -4.910 90.420 -2.435 ;
    END
  END ONB[44]
PIN ON[45]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 91.580 -4.910 91.870 -2.435 ;
    END
  END ON[45]
PIN ONB[45]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 92.130 -4.910 92.420 -2.435 ;
    END
  END ONB[45]
PIN ON[46]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 93.580 -4.910 93.870 -2.435 ;
    END
  END ON[46]
PIN ONB[46]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 94.130 -4.910 94.420 -2.435 ;
    END
  END ONB[46]
PIN ON[47]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 95.580 -4.910 95.870 -2.435 ;
    END
  END ON[47]
PIN ONB[47]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 96.130 -4.910 96.420 -2.435 ;
    END
  END ONB[47]
PIN ON[48]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 97.580 -4.910 97.870 -2.435 ;
    END
  END ON[48]
PIN ONB[48]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 98.130 -4.910 98.420 -2.435 ;
    END
  END ONB[48]
PIN ON[49]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 99.580 -4.910 99.870 -2.435 ;
    END
  END ON[49]
PIN ONB[49]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 100.130 -4.910 100.420 -2.435 ;
    END
  END ONB[49]
PIN ON[50]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 101.580 -4.910 101.870 -2.435 ;
    END
  END ON[50]
PIN ONB[50]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 102.130 -4.910 102.420 -2.435 ;
    END
  END ONB[50]
PIN ON[51]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 103.580 -4.910 103.870 -2.435 ;
    END
  END ON[51]
PIN ONB[51]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 104.130 -4.910 104.420 -2.435 ;
    END
  END ONB[51]
PIN ON[52]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 105.580 -4.910 105.870 -2.435 ;
    END
  END ON[52]
PIN ONB[52]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 106.130 -4.910 106.420 -2.435 ;
    END
  END ONB[52]
PIN ON[53]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 107.580 -4.910 107.870 -2.435 ;
    END
  END ON[53]
PIN ONB[53]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 108.130 -4.910 108.420 -2.435 ;
    END
  END ONB[53]
PIN ON[54]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 109.580 -4.910 109.870 -2.435 ;
    END
  END ON[54]
PIN ONB[54]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.130 -4.910 110.420 -2.435 ;
    END
  END ONB[54]
PIN ON[55]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 111.580 -4.910 111.870 -2.435 ;
    END
  END ON[55]
PIN ONB[55]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 112.130 -4.910 112.420 -2.435 ;
    END
  END ONB[55]
PIN ON[56]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 113.580 -4.910 113.870 -2.435 ;
    END
  END ON[56]
PIN ONB[56]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 114.130 -4.910 114.420 -2.435 ;
    END
  END ONB[56]
PIN ON[57]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 115.580 -4.910 115.870 -2.435 ;
    END
  END ON[57]
PIN ONB[57]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 116.130 -4.910 116.420 -2.435 ;
    END
  END ONB[57]
PIN ON[58]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.580 -4.910 117.870 -2.435 ;
    END
  END ON[58]
PIN ONB[58]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.130 -4.910 118.420 -2.435 ;
    END
  END ONB[58]
PIN ON[59]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 119.580 -4.910 119.870 -2.435 ;
    END
  END ON[59]
PIN ONB[59]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 120.130 -4.910 120.420 -2.435 ;
    END
  END ONB[59]
PIN ON[60]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 121.580 -4.910 121.870 -2.435 ;
    END
  END ON[60]
PIN ONB[60]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 122.130 -4.910 122.420 -2.435 ;
    END
  END ONB[60]
PIN ON[61]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 123.580 -4.910 123.870 -2.435 ;
    END
  END ON[61]
PIN ONB[61]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 124.130 -4.910 124.420 -2.435 ;
    END
  END ONB[61]
PIN ON[62]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 125.580 -4.910 125.870 -2.435 ;
    END
  END ON[62]
PIN ONB[62]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 126.130 -4.910 126.420 -2.435 ;
    END
  END ONB[62]
PIN ON[63]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 127.580 -4.910 127.870 -2.435 ;
    END
  END ON[63]
PIN ONB[63]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 128.130 -4.910 128.420 -2.435 ;
    END
  END ONB[63]
PIN ON[32]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 65.580 -4.910 65.870 -2.435 ;
    END
  END ON[32]
PIN ONB[32]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 66.130 -4.910 66.420 -2.435 ;
    END
  END ONB[32]
PIN EN[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 129.580 -4.910 129.870 -2.435 ;
    END
  END EN[1]
PIN ENB[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 130.130 -4.910 130.420 -2.435 ;
    END
  END ENB[1]
PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal2 ;
        RECT 2.210 30.700 4.210 31.700 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal2 ;
        RECT 134.630 5.110 136.630 6.110 ;
    END
  END VSS
  PIN Iout
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 68.420 30.700 70.420 31.700 ;
    END
  END Iout
  PIN VcascP[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2.210 17.905 4.210 18.905 ;
    END
  END VcascP[0]
  PIN VcascP[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.630 17.905 136.630 18.905 ;
    END
  END VcascP[1]
OBS
    LAYER Metal1 ;
      RECT 2.210 5.110 136.630 31.700 ;
    LAYER Metal2 ;
      RECT 2.210 5.110 136.630 31.700 ;
    LAYER Metal3 ;
      RECT 2.210 5.110 136.630 31.700 ;
  END
END DAC2U128OUT4IN
