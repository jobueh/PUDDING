* Extracted by KLayout with SG13G2 LVS runset on : 24/08/2025 22:56

.SUBCKT non_overlap
X$1 4 7 1 5 sg13g2_dlygate4sd1_1
X$2 8 4 3 1 2 sg13g2_nor2_1
X$3 4 7 1 sg13g2_buf_1
X$4 4 8 9 2 sg13g2_dlygate4sd1_1
X$5 7 4 6 3 sg13g2_inv_1
X$6 7 4 10 6 5 sg13g2_nor2_1
X$7 4 8 9 sg13g2_buf_1
.ENDS non_overlap

.SUBCKT sg13g2_inv_1 1 2 3 4
M$1 2 3 4 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.2516p PS=2.16u PD=2.16u
M$2 1 3 4 1 sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.3808p PS=2.92u PD=2.92u
.ENDS sg13g2_inv_1

.SUBCKT sg13g2_nor2_1 1 2 3 4 5
M$1 2 4 5 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.1406p PS=2.16u PD=1.12u
M$2 5 3 2 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.1406p AD=0.2516p PS=1.12u PD=2.16u
M$3 1 4 6 1 sg13_lv_pmos L=0.13u W=1.12u AS=0.4032p AD=0.1176p PS=2.96u PD=1.33u
M$4 6 3 5 1 sg13_lv_pmos L=0.13u W=1.12u AS=0.1176p AD=0.3808p PS=1.33u PD=2.92u
.ENDS sg13g2_nor2_1

.SUBCKT sg13g2_buf_1 2 4 5
M$1 2 5 1 2 sg13_lv_nmos L=0.13u W=0.55u AS=0.14875p AD=0.187p PS=1.16u PD=1.78u
M$2 2 1 3 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.14875p AD=0.2886p PS=1.16u
+ PD=2.26u
M$3 4 5 1 4 sg13_lv_pmos L=0.13u W=0.84u AS=0.2114p AD=0.2856p PS=1.54u PD=2.36u
M$4 4 1 3 4 sg13_lv_pmos L=0.13u W=1.12u AS=0.2114p AD=0.42p PS=1.54u PD=2.99u
.ENDS sg13g2_buf_1

.SUBCKT sg13g2_dlygate4sd1_1 2 3 5 7
M$1 1 7 2 2 sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.1428p PS=1.52u PD=1.1u
M$2 2 1 4 2 sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.1428p PS=1.1u PD=1.52u
M$3 2 4 6 2 sg13_lv_nmos L=0.13u W=0.42u AS=0.1405p AD=0.2373p PS=1.15u PD=1.97u
M$4 2 6 5 2 sg13_lv_nmos L=0.13u W=0.74u AS=0.1405p AD=0.2516p PS=1.15u PD=2.16u
M$5 6 4 3 3 sg13_lv_pmos L=0.13u W=1u AS=0.565p AD=0.2245p PS=3.13u PD=1.53u
M$6 3 6 5 3 sg13_lv_pmos L=0.13u W=1.12u AS=0.2245p AD=0.3808p PS=1.53u PD=2.92u
M$7 3 7 1 3 sg13_lv_pmos L=0.13u W=0.42u AS=0.2931p AD=0.1428p PS=1.65u PD=1.52u
M$8 3 1 4 3 sg13_lv_pmos L=0.13u W=1u AS=0.2931p AD=0.37p PS=1.65u PD=2.74u
.ENDS sg13g2_dlygate4sd1_1
