* Extracted by KLayout with SG13G2 LVS runset on : 28/10/2025 12:49

.SUBCKT dac128module VSS EN[0]|INP|ON ENB[0]|INN|ONB INP|ON|ON[0]
+ INN|ONB|ONB[0] INP|ON|ON[1] INN|ONB|ONB[1] INP|ON|ON[2] INN|ONB|ONB[2]
+ INP|ON|ON[3] INN|ONB|ONB[3] VDD INP|ON|ON[4] INN|ONB|ONB[4] INP|ON|ON[5]
+ INN|ONB|ONB[5] INP|ON|ON[6] INN|ONB|ONB[6] INP|ON|ON[7] INN|ONB|ONB[7]
+ INP|ON|ON[8] INN|ONB|ONB[8] INP|ON|ON[9] INN|ONB|ONB[9] INP|ON|ON[10]
+ INN|ONB|ONB[10] INP|ON|ON[11] INN|ONB|ONB[11] INP|ON|ON[12] INN|ONB|ONB[12]
+ INP|ON|ON[13] INN|ONB|ONB[13] INP|ON|ON[14] INN|ONB|ONB[14] INP|ON|ON[15]
+ INN|ONB|ONB[15] INP|ON|ON[16] INN|ONB|ONB[16] INP|ON|ON[17] INN|ONB|ONB[17]
+ INP|ON|ON[18] INN|ONB|ONB[18] INP|ON|ON[19] INN|ONB|ONB[19] INP|ON|ON[20]
+ INN|ONB|ONB[20] INP|ON|ON[21] INN|ONB|ONB[21] INP|ON|ON[22] INN|ONB|ONB[22]
+ INP|ON|ON[23] INN|ONB|ONB[23] INP|ON|ON[24] INN|ONB|ONB[24] INP|ON|ON[25]
+ INN|ONB|ONB[25] INP|ON|ON[26] INN|ONB|ONB[26] INP|ON|ON[27] INN|ONB|ONB[27]
+ INP|ON|ON[28] INN|ONB|ONB[28] INP|ON|ON[29] INN|ONB|ONB[29] INP|ON|ON[30]
+ INN|ONB|ONB[30] INP|ON|ON[31] INN|ONB|ONB[31] INP|ON|ON[32] INN|ONB|ONB[32]
+ INP|ON|ON[33] INN|ONB|ONB[33] INP|ON|ON[34] INN|ONB|ONB[34] INP|ON|ON[35]
+ INN|ONB|ONB[35] INP|ON|ON[36] INN|ONB|ONB[36] INP|ON|ON[37] INN|ONB|ONB[37]
+ INP|ON|ON[38] INN|ONB|ONB[38] INP|ON|ON[39] INN|ONB|ONB[39] INP|ON|ON[40]
+ INN|ONB|ONB[40] INP|ON|ON[41] INN|ONB|ONB[41] INP|ON|ON[42] INN|ONB|ONB[42]
+ INP|ON|ON[43] INN|ONB|ONB[43] INP|ON|ON[44] INN|ONB|ONB[44] INP|ON|ON[45]
+ INN|ONB|ONB[45] INP|ON|ON[46] INN|ONB|ONB[46] INP|ON|ON[47] INN|ONB|ONB[47]
+ INP|ON|ON[48] INN|ONB|ONB[48] INP|ON|ON[49] INN|ONB|ONB[49] INP|ON|ON[50]
+ INN|ONB|ONB[50] INP|ON|ON[51] INN|ONB|ONB[51] INP|ON|ON[52] INN|ONB|ONB[52]
+ INP|ON|ON[53] INN|ONB|ONB[53] INP|ON|ON[54] INN|ONB|ONB[54] INP|ON|ON[55]
+ INN|ONB|ONB[55] INP|ON|ON[56] INN|ONB|ONB[56] INP|ON|ON[57] INN|ONB|ONB[57]
+ INP|ON|ON[58] INN|ONB|ONB[58] INP|ON|ON[59] INN|ONB|ONB[59] INP|ON|ON[60]
+ INN|ONB|ONB[60] INP|ON|ON[61] INN|ONB|ONB[61] INP|ON|ON[62] INN|ONB|ONB[62]
+ INP|ON|ON[63] INN|ONB|ONB[63] EN[1]|INP|ON ENB[1]|INN|ONB OUTN OUTP OUTN$1
+ OUTP$1 OUTN$2 OUTP$2 OUTN$3 OUTP$3 OUTN$4 OUTP$4 OUTN$5 OUTP$5 OUTN$6 OUTP$6
+ OUTN$7 OUTP$7 OUTN$8 OUTP$8 OUTN$9 OUTP$9 OUTN$10 OUTP$10 OUTN$11 OUTP$11
+ OUTN$12 OUTP$12 OUTN$13 OUTP$13 OUTN$14 OUTP$14 OUTN$15 OUTP$15 OUTN$16
+ OUTP$16 OUTN$17 OUTP$17 OUTN$18 OUTP$18 OUTN$19 OUTP$19 OUTN$20 OUTP$20
+ OUTN$21 OUTP$21 OUTN$22 OUTP$22 OUTN$23 OUTP$23 OUTN$24 OUTP$24 OUTN$25
+ OUTP$25 OUTN$26 OUTP$26 OUTN$27 OUTP$27 OUTN$28 OUTP$28 OUTN$29 OUTP$29
+ OUTN$30 OUTP$30 OUTN$31 OUTP$31 OUTN$32 OUTP$32 OUTN$33 OUTP$33 OUTN$34
+ OUTP$34 OUTN$35 OUTP$35 OUTN$36 OUTP$36 OUTN$37 OUTP$37 OUTN$38 OUTP$38
+ OUTN$39 OUTP$39 OUTN$40 OUTP$40 OUTN$41 OUTP$41 OUTN$42 OUTP$42 OUTN$43
+ OUTP$43 OUTN$44 OUTP$44 OUTN$45 OUTP$45 OUTN$46 OUTP$46 OUTN$47 OUTP$47
+ OUTN$48 OUTP$48 OUTN$49 OUTP$49 OUTN$50 OUTP$50 OUTN$51 OUTP$51 OUTN$52
+ OUTP$52 OUTN$53 OUTP$53 OUTN$54 OUTP$54 OUTN$55 OUTP$55 OUTN$56 OUTP$56
+ OUTN$57 OUTP$57 OUTN$58 OUTP$58 OUTN$59 OUTP$59 OUTN$60 OUTP$60 OUTN$61
+ OUTP$61 OUTN$62 OUTP$62 OUTN$63 OUTP$63 OUTN$64 OUTP$64 OUTN$65 OUTP$65
+ VcascP|VcascP[0] VcascodeP VcascodeP$1 VcascodeP$2 VcascodeP$3 VcascodeP$4
+ VcascodeP$5 VcascodeP$6 VcascodeP$7 VcascodeP$8 VcascodeP$9 VcascodeP$10
+ VcascodeP$11 VcascodeP$12 VcascodeP$13 VcascodeP$14 VcascodeP$15 VcascodeP$16
+ VcascodeP$17 VcascodeP$18 VcascodeP$19 VcascodeP$20 VcascodeP$21 VcascodeP$22
+ VcascodeP$23 VcascodeP$24 VcascodeP$25 VcascodeP$26 VcascodeP$27 VcascodeP$28
+ VcascodeP$29 VcascodeP$30 VcascodeP$31 VcascodeP$32 VcascodeP$33 VcascodeP$34
+ VcascodeP$35 VcascodeP$36 VcascodeP$37 VcascodeP$38 VcascodeP$39 VcascodeP$40
+ VcascodeP$41 VcascodeP$42 VcascodeP$43 VcascodeP$44 VcascodeP$45 VcascodeP$46
+ VcascodeP$47 VcascodeP$48 VcascodeP$49 VcascodeP$50 VcascodeP$51 VcascodeP$52
+ VcascodeP$53 VcascodeP$54 VcascodeP$55 VcascodeP$56 VcascodeP$57 VcascodeP$58
+ VcascodeP$59 VcascodeP$60 VcascodeP$61 VcascodeP$62 VcascodeP$63 VcascodeP$64
+ VcascodeP$65 Iout|VbiasP|VbiasP[0] Iout Iout|VbiasP|VbiasP[1]
+ VcascP|VcascP[1] VcascodeP$66 VcascodeP$67 VcascodeP$68 VcascodeP$69
+ VcascodeP$70 VcascodeP$71 VcascodeP$72 VcascodeP$73 VcascodeP$74 VcascodeP$75
+ VcascodeP$76 VcascodeP$77 VcascodeP$78 VcascodeP$79 VcascodeP$80 VcascodeP$81
+ VcascodeP$82 VcascodeP$83 VcascodeP$84 VcascodeP$85 VcascodeP$86 VcascodeP$87
+ VcascodeP$88 VcascodeP$89 VcascodeP$90 VcascodeP$91 VcascodeP$92 VcascodeP$93
+ VcascodeP$94 VcascodeP$95 VcascodeP$96 VcascodeP$97 VcascodeP$98 VcascodeP$99
+ VcascodeP$100 VcascodeP$101 VcascodeP$102 VcascodeP$103 VcascodeP$104
+ VcascodeP$105 VcascodeP$106 VcascodeP$107 VcascodeP$108 VcascodeP$109
+ VcascodeP$110 VcascodeP$111 VcascodeP$112 VcascodeP$113 VcascodeP$114
+ VcascodeP$115 VcascodeP$116 VcascodeP$117 VcascodeP$118 VcascodeP$119
+ VcascodeP$120 VcascodeP$121 VcascodeP$122 VcascodeP$123 VcascodeP$124
+ VcascodeP$125 VcascodeP$126 VcascodeP$127 VcascodeP$128 VcascodeP$129
+ VcascodeP$130 VcascodeP$131 OUTP$66 OUTN$66 OUTP$67 OUTN$67 OUTP$68 OUTN$68
+ OUTP$69 OUTN$69 OUTP$70 OUTN$70 OUTP$71 OUTN$71 OUTP$72 OUTN$72 OUTP$73
+ OUTN$73 OUTP$74 OUTN$74 OUTP$75 OUTN$75 OUTP$76 OUTN$76 OUTP$77 OUTN$77
+ OUTP$78 OUTN$78 OUTP$79 OUTN$79 OUTP$80 OUTN$80 OUTP$81 OUTN$81 OUTP$82
+ OUTN$82 OUTP$83 OUTN$83 OUTP$84 OUTN$84 OUTP$85 OUTN$85 OUTP$86 OUTN$86
+ OUTP$87 OUTN$87 OUTP$88 OUTN$88 OUTP$89 OUTN$89 OUTP$90 OUTN$90 OUTP$91
+ OUTN$91 OUTP$92 OUTN$92 OUTP$93 OUTN$93 OUTP$94 OUTN$94 OUTP$95 OUTN$95
+ OUTP$96 OUTN$96 OUTP$97 OUTN$97 OUTP$98 OUTN$98 OUTP$99 OUTN$99 OUTP$100
+ OUTN$100 OUTP$101 OUTN$101 OUTP$102 OUTN$102 OUTP$103 OUTN$103 OUTP$104
+ OUTN$104 OUTP$105 OUTN$105 OUTP$106 OUTN$106 OUTP$107 OUTN$107 OUTP$108
+ OUTN$108 OUTP$109 OUTN$109 OUTP$110 OUTN$110 OUTP$111 OUTN$111 OUTP$112
+ OUTN$112 OUTP$113 OUTN$113 OUTP$114 OUTN$114 OUTP$115 OUTN$115 OUTP$116
+ OUTN$116 OUTP$117 OUTN$117 OUTP$118 OUTN$118 OUTP$119 OUTN$119 OUTP$120
+ OUTN$120 OUTP$121 OUTN$121 OUTP$122 OUTN$122 OUTP$123 OUTN$123 OUTP$124
+ OUTN$124 OUTP$125 OUTN$125 OUTP$126 OUTN$126 OUTP$127 OUTN$127 OUTP$128
+ OUTN$128 OUTP$129 OUTN$129 OUTP$130 OUTN$130 OUTP$131 OUTN$131
+ ENB[1]|ENB[3]|INN|ONB EN[1]|EN[3]|INP|ON INN|ONB|ONB[127]|ONB[63]
+ INP|ON|ON[127]|ON[63] INN|ONB|ONB[126]|ONB[62] INP|ON|ON[126]|ON[62]
+ INN|ONB|ONB[125]|ONB[61] INP|ON|ON[125]|ON[61] INN|ONB|ONB[124]|ONB[60]
+ INP|ON|ON[124]|ON[60] INN|ONB|ONB[123]|ONB[59] INP|ON|ON[123]|ON[59]
+ INN|ONB|ONB[122]|ONB[58] INP|ON|ON[122]|ON[58] INN|ONB|ONB[121]|ONB[57]
+ INP|ON|ON[121]|ON[57] INN|ONB|ONB[120]|ONB[56] INP|ON|ON[120]|ON[56]
+ INN|ONB|ONB[119]|ONB[55] INP|ON|ON[119]|ON[55] INN|ONB|ONB[118]|ONB[54]
+ INP|ON|ON[118]|ON[54] INN|ONB|ONB[117]|ONB[53] INP|ON|ON[117]|ON[53]
+ INN|ONB|ONB[116]|ONB[52] INP|ON|ON[116]|ON[52] INN|ONB|ONB[115]|ONB[51]
+ INP|ON|ON[115]|ON[51] INN|ONB|ONB[114]|ONB[50] INP|ON|ON[114]|ON[50]
+ INN|ONB|ONB[113]|ONB[49] INP|ON|ON[113]|ON[49] INN|ONB|ONB[112]|ONB[48]
+ INP|ON|ON[112]|ON[48] INN|ONB|ONB[111]|ONB[47] INP|ON|ON[111]|ON[47]
+ INN|ONB|ONB[110]|ONB[46] INP|ON|ON[110]|ON[46] INN|ONB|ONB[109]|ONB[45]
+ INP|ON|ON[109]|ON[45] INN|ONB|ONB[108]|ONB[44] INP|ON|ON[108]|ON[44]
+ INN|ONB|ONB[107]|ONB[43] INP|ON|ON[107]|ON[43] INN|ONB|ONB[106]|ONB[42]
+ INP|ON|ON[106]|ON[42] INN|ONB|ONB[105]|ONB[41] INP|ON|ON[105]|ON[41]
+ INN|ONB|ONB[104]|ONB[40] INP|ON|ON[104]|ON[40] INN|ONB|ONB[103]|ONB[39]
+ INP|ON|ON[103]|ON[39] INN|ONB|ONB[102]|ONB[38] INP|ON|ON[102]|ON[38]
+ INN|ONB|ONB[101]|ONB[37] INP|ON|ON[101]|ON[37] INN|ONB|ONB[100]|ONB[36]
+ INP|ON|ON[100]|ON[36] INN|ONB|ONB[35]|ONB[99] INP|ON|ON[35]|ON[99]
+ INN|ONB|ONB[34]|ONB[98] INP|ON|ON[34]|ON[98] INN|ONB|ONB[33]|ONB[97]
+ INP|ON|ON[33]|ON[97] INN|ONB|ONB[32]|ONB[96] INP|ON|ON[32]|ON[96]
+ INN|ONB|ONB[31]|ONB[95] INP|ON|ON[31]|ON[95] INN|ONB|ONB[30]|ONB[94]
+ INP|ON|ON[30]|ON[94] INN|ONB|ONB[29]|ONB[93] INP|ON|ON[29]|ON[93]
+ INN|ONB|ONB[28]|ONB[92] INP|ON|ON[28]|ON[92] INN|ONB|ONB[27]|ONB[91]
+ INP|ON|ON[27]|ON[91] INN|ONB|ONB[26]|ONB[90] INP|ON|ON[26]|ON[90]
+ INN|ONB|ONB[25]|ONB[89] INP|ON|ON[25]|ON[89] INN|ONB|ONB[24]|ONB[88]
+ INP|ON|ON[24]|ON[88] INN|ONB|ONB[23]|ONB[87] INP|ON|ON[23]|ON[87]
+ INN|ONB|ONB[22]|ONB[86] INP|ON|ON[22]|ON[86] INN|ONB|ONB[21]|ONB[85]
+ INP|ON|ON[21]|ON[85] INN|ONB|ONB[20]|ONB[84] INP|ON|ON[20]|ON[84]
+ INN|ONB|ONB[19]|ONB[83] INP|ON|ON[19]|ON[83] INN|ONB|ONB[18]|ONB[82]
+ INP|ON|ON[18]|ON[82] INN|ONB|ONB[17]|ONB[81] INP|ON|ON[17]|ON[81]
+ INN|ONB|ONB[16]|ONB[80] INP|ON|ON[16]|ON[80] INN|ONB|ONB[15]|ONB[79]
+ INP|ON|ON[15]|ON[79] INN|ONB|ONB[14]|ONB[78] INP|ON|ON[14]|ON[78]
+ INN|ONB|ONB[13]|ONB[77] INP|ON|ON[13]|ON[77] INN|ONB|ONB[12]|ONB[76]
+ INP|ON|ON[12]|ON[76] INN|ONB|ONB[11]|ONB[75] INP|ON|ON[11]|ON[75]
+ INN|ONB|ONB[10]|ONB[74] INP|ON|ON[10]|ON[74] INN|ONB|ONB[73]|ONB[9]
+ INP|ON|ON[73]|ON[9] INN|ONB|ONB[72]|ONB[8] INP|ON|ON[72]|ON[8]
+ INN|ONB|ONB[71]|ONB[7] INP|ON|ON[71]|ON[7] INN|ONB|ONB[6]|ONB[70]
+ INP|ON|ON[6]|ON[70] INN|ONB|ONB[5]|ONB[69] INP|ON|ON[5]|ON[69]
+ INN|ONB|ONB[4]|ONB[68] INP|ON|ON[4]|ON[68] INN|ONB|ONB[3]|ONB[67]
+ INP|ON|ON[3]|ON[67] INN|ONB|ONB[2]|ONB[66] INP|ON|ON[2]|ON[66]
+ INN|ONB|ONB[1]|ONB[65] INP|ON|ON[1]|ON[65] INN|ONB|ONB[0]|ONB[64]
+ INP|ON|ON[0]|ON[64] ENB[0]|ENB[2]|INN|ONB EN[0]|EN[2]|INP|ON
M$1 OUTP$66 OUTN$66 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$2 VSS OUTP$66 OUTN$66 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$3 OUTN OUTP VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$4 VSS OUTN OUTP VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$5 OUTP$67 OUTN$67 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$6 VSS OUTP$67 OUTN$67 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$7 OUTN$1 OUTP$1 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$8 VSS OUTN$1 OUTP$1 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$9 OUTP$68 OUTN$68 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$10 VSS OUTP$68 OUTN$68 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$11 OUTN$2 OUTP$2 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$12 VSS OUTN$2 OUTP$2 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$13 OUTP$69 OUTN$69 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$14 VSS OUTP$69 OUTN$69 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$15 OUTN$3 OUTP$3 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$16 VSS OUTN$3 OUTP$3 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$17 OUTN$4 OUTP$4 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$18 VSS OUTN$4 OUTP$4 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$19 OUTP$70 OUTN$70 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$20 VSS OUTP$70 OUTN$70 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$21 OUTN$5 OUTP$5 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$22 VSS OUTN$5 OUTP$5 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$23 OUTP$71 OUTN$71 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$24 VSS OUTP$71 OUTN$71 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$25 OUTN$6 OUTP$6 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$26 VSS OUTN$6 OUTP$6 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$27 OUTP$72 OUTN$72 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$28 VSS OUTP$72 OUTN$72 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$29 OUTN$7 OUTP$7 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$30 VSS OUTN$7 OUTP$7 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$31 OUTP$73 OUTN$73 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$32 VSS OUTP$73 OUTN$73 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$33 OUTN$8 OUTP$8 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$34 VSS OUTN$8 OUTP$8 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$35 OUTP$74 OUTN$74 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$36 VSS OUTP$74 OUTN$74 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$37 OUTN$9 OUTP$9 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$38 VSS OUTN$9 OUTP$9 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$39 OUTP$75 OUTN$75 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$40 VSS OUTP$75 OUTN$75 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$41 OUTP$76 OUTN$76 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$42 VSS OUTP$76 OUTN$76 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$43 OUTN$10 OUTP$10 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$44 VSS OUTN$10 OUTP$10 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$45 OUTP$77 OUTN$77 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$46 VSS OUTP$77 OUTN$77 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$47 OUTN$11 OUTP$11 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$48 VSS OUTN$11 OUTP$11 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$49 OUTN$12 OUTP$12 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$50 VSS OUTN$12 OUTP$12 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$51 OUTP$78 OUTN$78 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$52 VSS OUTP$78 OUTN$78 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$53 OUTP$79 OUTN$79 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$54 VSS OUTP$79 OUTN$79 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$55 OUTN$13 OUTP$13 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$56 VSS OUTN$13 OUTP$13 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$57 OUTP$80 OUTN$80 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$58 VSS OUTP$80 OUTN$80 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$59 OUTN$14 OUTP$14 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$60 VSS OUTN$14 OUTP$14 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$61 OUTN$15 OUTP$15 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$62 VSS OUTN$15 OUTP$15 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$63 OUTP$81 OUTN$81 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$64 VSS OUTP$81 OUTN$81 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$65 OUTN$16 OUTP$16 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$66 VSS OUTN$16 OUTP$16 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$67 OUTP$82 OUTN$82 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$68 VSS OUTP$82 OUTN$82 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$69 OUTP$83 OUTN$83 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$70 VSS OUTP$83 OUTN$83 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$71 OUTN$17 OUTP$17 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$72 VSS OUTN$17 OUTP$17 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$73 OUTP$84 OUTN$84 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$74 VSS OUTP$84 OUTN$84 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$75 OUTN$18 OUTP$18 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$76 VSS OUTN$18 OUTP$18 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$77 OUTP$85 OUTN$85 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$78 VSS OUTP$85 OUTN$85 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$79 OUTN$19 OUTP$19 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$80 VSS OUTN$19 OUTP$19 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$81 OUTP$86 OUTN$86 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$82 VSS OUTP$86 OUTN$86 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$83 OUTN$20 OUTP$20 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$84 VSS OUTN$20 OUTP$20 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$85 OUTN$21 OUTP$21 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$86 VSS OUTN$21 OUTP$21 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$87 OUTP$87 OUTN$87 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$88 VSS OUTP$87 OUTN$87 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$89 OUTN$22 OUTP$22 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$90 VSS OUTN$22 OUTP$22 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$91 OUTP$88 OUTN$88 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$92 VSS OUTP$88 OUTN$88 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$93 OUTN$23 OUTP$23 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$94 VSS OUTN$23 OUTP$23 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$95 OUTP$89 OUTN$89 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$96 VSS OUTP$89 OUTN$89 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$97 OUTP$90 OUTN$90 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$98 VSS OUTP$90 OUTN$90 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$99 OUTN$24 OUTP$24 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$100 VSS OUTN$24 OUTP$24 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$101 OUTP$91 OUTN$91 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$102 VSS OUTP$91 OUTN$91 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$103 OUTN$25 OUTP$25 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$104 VSS OUTN$25 OUTP$25 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$105 OUTN$26 OUTP$26 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$106 VSS OUTN$26 OUTP$26 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$107 OUTP$92 OUTN$92 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$108 VSS OUTP$92 OUTN$92 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$109 OUTP$93 OUTN$93 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$110 VSS OUTP$93 OUTN$93 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$111 OUTN$27 OUTP$27 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$112 VSS OUTN$27 OUTP$27 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$113 OUTN$28 OUTP$28 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$114 VSS OUTN$28 OUTP$28 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$115 OUTP$94 OUTN$94 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$116 VSS OUTP$94 OUTN$94 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$117 OUTP$95 OUTN$95 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$118 VSS OUTP$95 OUTN$95 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$119 OUTN$29 OUTP$29 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$120 VSS OUTN$29 OUTP$29 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$121 OUTN$30 OUTP$30 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$122 VSS OUTN$30 OUTP$30 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$123 OUTP$96 OUTN$96 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$124 VSS OUTP$96 OUTN$96 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$125 OUTP$97 OUTN$97 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$126 VSS OUTP$97 OUTN$97 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$127 OUTN$31 OUTP$31 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$128 VSS OUTN$31 OUTP$31 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$129 OUTP$98 OUTN$98 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$130 VSS OUTP$98 OUTN$98 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$131 OUTN$32 OUTP$32 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$132 VSS OUTN$32 OUTP$32 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$133 OUTN$33 OUTP$33 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$134 VSS OUTN$33 OUTP$33 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$135 OUTP$99 OUTN$99 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$136 VSS OUTP$99 OUTN$99 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$137 OUTP$100 OUTN$100 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$138 VSS OUTP$100 OUTN$100 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$139 OUTN$34 OUTP$34 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$140 VSS OUTN$34 OUTP$34 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$141 OUTN$35 OUTP$35 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$142 VSS OUTN$35 OUTP$35 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$143 OUTP$101 OUTN$101 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$144 VSS OUTP$101 OUTN$101 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$145 OUTP$102 OUTN$102 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$146 VSS OUTP$102 OUTN$102 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$147 OUTN$36 OUTP$36 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$148 VSS OUTN$36 OUTP$36 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$149 OUTP$103 OUTN$103 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$150 VSS OUTP$103 OUTN$103 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$151 OUTN$37 OUTP$37 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$152 VSS OUTN$37 OUTP$37 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$153 OUTN$38 OUTP$38 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$154 VSS OUTN$38 OUTP$38 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$155 OUTP$104 OUTN$104 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$156 VSS OUTP$104 OUTN$104 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$157 OUTN$39 OUTP$39 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$158 VSS OUTN$39 OUTP$39 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$159 OUTP$105 OUTN$105 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$160 VSS OUTP$105 OUTN$105 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$161 OUTP$106 OUTN$106 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$162 VSS OUTP$106 OUTN$106 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$163 OUTN$40 OUTP$40 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$164 VSS OUTN$40 OUTP$40 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$165 OUTP$107 OUTN$107 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$166 VSS OUTP$107 OUTN$107 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$167 OUTN$41 OUTP$41 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$168 VSS OUTN$41 OUTP$41 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$169 OUTN$42 OUTP$42 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$170 VSS OUTN$42 OUTP$42 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$171 OUTP$108 OUTN$108 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$172 VSS OUTP$108 OUTN$108 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$173 OUTP$109 OUTN$109 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$174 VSS OUTP$109 OUTN$109 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$175 OUTN$43 OUTP$43 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$176 VSS OUTN$43 OUTP$43 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$177 OUTN$44 OUTP$44 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$178 VSS OUTN$44 OUTP$44 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$179 OUTP$110 OUTN$110 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$180 VSS OUTP$110 OUTN$110 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$181 OUTN$45 OUTP$45 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$182 VSS OUTN$45 OUTP$45 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$183 OUTP$111 OUTN$111 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$184 VSS OUTP$111 OUTN$111 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$185 OUTP$112 OUTN$112 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$186 VSS OUTP$112 OUTN$112 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$187 OUTN$46 OUTP$46 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$188 VSS OUTN$46 OUTP$46 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$189 OUTP$113 OUTN$113 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$190 VSS OUTP$113 OUTN$113 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$191 OUTN$47 OUTP$47 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$192 VSS OUTN$47 OUTP$47 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$193 OUTN$48 OUTP$48 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$194 VSS OUTN$48 OUTP$48 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$195 OUTP$114 OUTN$114 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$196 VSS OUTP$114 OUTN$114 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$197 OUTP$115 OUTN$115 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$198 VSS OUTP$115 OUTN$115 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$199 OUTN$49 OUTP$49 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$200 VSS OUTN$49 OUTP$49 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$201 OUTP$116 OUTN$116 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$202 VSS OUTP$116 OUTN$116 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$203 OUTN$50 OUTP$50 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$204 VSS OUTN$50 OUTP$50 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$205 OUTN$51 OUTP$51 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$206 VSS OUTN$51 OUTP$51 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$207 OUTP$117 OUTN$117 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$208 VSS OUTP$117 OUTN$117 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$209 OUTN$52 OUTP$52 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$210 VSS OUTN$52 OUTP$52 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$211 OUTP$118 OUTN$118 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$212 VSS OUTP$118 OUTN$118 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$213 OUTN$53 OUTP$53 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$214 VSS OUTN$53 OUTP$53 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$215 OUTP$119 OUTN$119 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$216 VSS OUTP$119 OUTN$119 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$217 OUTP$120 OUTN$120 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$218 VSS OUTP$120 OUTN$120 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$219 OUTN$54 OUTP$54 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$220 VSS OUTN$54 OUTP$54 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$221 OUTN$55 OUTP$55 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$222 VSS OUTN$55 OUTP$55 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$223 OUTP$121 OUTN$121 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$224 VSS OUTP$121 OUTN$121 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$225 OUTP$122 OUTN$122 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$226 VSS OUTP$122 OUTN$122 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$227 OUTN$56 OUTP$56 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$228 VSS OUTN$56 OUTP$56 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$229 OUTN$57 OUTP$57 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$230 VSS OUTN$57 OUTP$57 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$231 OUTP$123 OUTN$123 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$232 VSS OUTP$123 OUTN$123 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$233 OUTP$124 OUTN$124 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$234 VSS OUTP$124 OUTN$124 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$235 OUTN$58 OUTP$58 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$236 VSS OUTN$58 OUTP$58 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$237 OUTN$59 OUTP$59 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$238 VSS OUTN$59 OUTP$59 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$239 OUTP$125 OUTN$125 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$240 VSS OUTP$125 OUTN$125 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$241 OUTP$126 OUTN$126 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$242 VSS OUTP$126 OUTN$126 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$243 OUTN$60 OUTP$60 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$244 VSS OUTN$60 OUTP$60 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$245 OUTP$127 OUTN$127 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$246 VSS OUTP$127 OUTN$127 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$247 OUTN$61 OUTP$61 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$248 VSS OUTN$61 OUTP$61 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$249 OUTN$62 OUTP$62 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$250 VSS OUTN$62 OUTP$62 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$251 OUTP$128 OUTN$128 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$252 VSS OUTP$128 OUTN$128 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$253 OUTN$63 OUTP$63 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$254 VSS OUTN$63 OUTP$63 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$255 OUTP$129 OUTN$129 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$256 VSS OUTP$129 OUTN$129 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$257 OUTN$64 OUTP$64 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$258 VSS OUTN$64 OUTP$64 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$259 OUTP$130 OUTN$130 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$260 VSS OUTP$130 OUTN$130 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$261 OUTN$65 OUTP$65 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$262 VSS OUTN$65 OUTP$65 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$263 OUTP$131 OUTN$131 VSS VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.162p
+ AD=0.0855p PS=2.16u PD=1.14u
M$264 VSS OUTP$131 OUTN$131 VSS sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p
+ AD=0.162p PS=1.14u PD=2.16u
M$265 OUTN EN[0]|INP|ON VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$266 VDD ENB[0]|INN|ONB OUTP VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$267 OUTN$1 INP|ON|ON[0] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$268 VDD INN|ONB|ONB[0] OUTP$1 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$269 OUTN$2 INP|ON|ON[1] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$270 VDD INN|ONB|ONB[1] OUTP$2 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$271 OUTN$3 INP|ON|ON[2] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$272 VDD INN|ONB|ONB[2] OUTP$3 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$273 OUTN$4 INP|ON|ON[3] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$274 VDD INN|ONB|ONB[3] OUTP$4 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$275 OUTN$5 INP|ON|ON[4] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$276 VDD INN|ONB|ONB[4] OUTP$5 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$277 OUTN$6 INP|ON|ON[5] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$278 VDD INN|ONB|ONB[5] OUTP$6 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$279 OUTN$7 INP|ON|ON[6] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$280 VDD INN|ONB|ONB[6] OUTP$7 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$281 OUTN$8 INP|ON|ON[7] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$282 VDD INN|ONB|ONB[7] OUTP$8 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$283 OUTN$9 INP|ON|ON[8] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$284 VDD INN|ONB|ONB[8] OUTP$9 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$285 OUTN$10 INP|ON|ON[9] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$286 VDD INN|ONB|ONB[9] OUTP$10 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$287 OUTN$11 INP|ON|ON[10] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$288 VDD INN|ONB|ONB[10] OUTP$11 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$289 OUTN$12 INP|ON|ON[11] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$290 VDD INN|ONB|ONB[11] OUTP$12 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$291 OUTN$13 INP|ON|ON[12] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$292 VDD INN|ONB|ONB[12] OUTP$13 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$293 OUTN$14 INP|ON|ON[13] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$294 VDD INN|ONB|ONB[13] OUTP$14 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$295 OUTN$15 INP|ON|ON[14] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$296 VDD INN|ONB|ONB[14] OUTP$15 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$297 OUTN$16 INP|ON|ON[15] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$298 VDD INN|ONB|ONB[15] OUTP$16 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$299 OUTN$17 INP|ON|ON[16] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$300 VDD INN|ONB|ONB[16] OUTP$17 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$301 OUTN$18 INP|ON|ON[17] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$302 VDD INN|ONB|ONB[17] OUTP$18 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$303 OUTN$19 INP|ON|ON[18] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$304 VDD INN|ONB|ONB[18] OUTP$19 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$305 OUTN$20 INP|ON|ON[19] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$306 VDD INN|ONB|ONB[19] OUTP$20 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$307 OUTN$21 INP|ON|ON[20] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$308 VDD INN|ONB|ONB[20] OUTP$21 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$309 OUTN$22 INP|ON|ON[21] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$310 VDD INN|ONB|ONB[21] OUTP$22 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$311 OUTN$23 INP|ON|ON[22] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$312 VDD INN|ONB|ONB[22] OUTP$23 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$313 OUTN$24 INP|ON|ON[23] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$314 VDD INN|ONB|ONB[23] OUTP$24 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$315 OUTN$25 INP|ON|ON[24] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$316 VDD INN|ONB|ONB[24] OUTP$25 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$317 OUTN$26 INP|ON|ON[25] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$318 VDD INN|ONB|ONB[25] OUTP$26 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$319 OUTN$27 INP|ON|ON[26] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$320 VDD INN|ONB|ONB[26] OUTP$27 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$321 OUTN$28 INP|ON|ON[27] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$322 VDD INN|ONB|ONB[27] OUTP$28 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$323 OUTN$29 INP|ON|ON[28] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$324 VDD INN|ONB|ONB[28] OUTP$29 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$325 OUTN$30 INP|ON|ON[29] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$326 VDD INN|ONB|ONB[29] OUTP$30 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$327 OUTN$31 INP|ON|ON[30] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$328 VDD INN|ONB|ONB[30] OUTP$31 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$329 OUTN$32 INP|ON|ON[31] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$330 VDD INN|ONB|ONB[31] OUTP$32 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$331 OUTN$33 INP|ON|ON[32] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$332 VDD INN|ONB|ONB[32] OUTP$33 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$333 OUTN$34 INP|ON|ON[33] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$334 VDD INN|ONB|ONB[33] OUTP$34 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$335 OUTN$35 INP|ON|ON[34] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$336 VDD INN|ONB|ONB[34] OUTP$35 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$337 OUTN$36 INP|ON|ON[35] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$338 VDD INN|ONB|ONB[35] OUTP$36 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$339 OUTN$37 INP|ON|ON[36] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$340 VDD INN|ONB|ONB[36] OUTP$37 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$341 OUTN$38 INP|ON|ON[37] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$342 VDD INN|ONB|ONB[37] OUTP$38 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$343 OUTN$39 INP|ON|ON[38] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$344 VDD INN|ONB|ONB[38] OUTP$39 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$345 OUTN$40 INP|ON|ON[39] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$346 VDD INN|ONB|ONB[39] OUTP$40 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$347 OUTN$41 INP|ON|ON[40] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$348 VDD INN|ONB|ONB[40] OUTP$41 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$349 OUTN$42 INP|ON|ON[41] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$350 VDD INN|ONB|ONB[41] OUTP$42 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$351 OUTN$43 INP|ON|ON[42] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$352 VDD INN|ONB|ONB[42] OUTP$43 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$353 OUTN$44 INP|ON|ON[43] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$354 VDD INN|ONB|ONB[43] OUTP$44 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$355 OUTN$45 INP|ON|ON[44] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$356 VDD INN|ONB|ONB[44] OUTP$45 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$357 OUTN$46 INP|ON|ON[45] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$358 VDD INN|ONB|ONB[45] OUTP$46 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$359 OUTN$47 INP|ON|ON[46] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$360 VDD INN|ONB|ONB[46] OUTP$47 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$361 OUTN$48 INP|ON|ON[47] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$362 VDD INN|ONB|ONB[47] OUTP$48 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$363 OUTN$49 INP|ON|ON[48] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$364 VDD INN|ONB|ONB[48] OUTP$49 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$365 OUTN$50 INP|ON|ON[49] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$366 VDD INN|ONB|ONB[49] OUTP$50 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$367 OUTN$51 INP|ON|ON[50] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$368 VDD INN|ONB|ONB[50] OUTP$51 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$369 OUTN$52 INP|ON|ON[51] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$370 VDD INN|ONB|ONB[51] OUTP$52 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$371 OUTN$53 INP|ON|ON[52] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$372 VDD INN|ONB|ONB[52] OUTP$53 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$373 OUTN$54 INP|ON|ON[53] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$374 VDD INN|ONB|ONB[53] OUTP$54 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$375 OUTN$55 INP|ON|ON[54] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$376 VDD INN|ONB|ONB[54] OUTP$55 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$377 OUTN$56 INP|ON|ON[55] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$378 VDD INN|ONB|ONB[55] OUTP$56 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$379 OUTN$57 INP|ON|ON[56] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$380 VDD INN|ONB|ONB[56] OUTP$57 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$381 OUTN$58 INP|ON|ON[57] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$382 VDD INN|ONB|ONB[57] OUTP$58 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$383 OUTN$59 INP|ON|ON[58] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$384 VDD INN|ONB|ONB[58] OUTP$59 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$385 OUTN$60 INP|ON|ON[59] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$386 VDD INN|ONB|ONB[59] OUTP$60 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$387 OUTN$61 INP|ON|ON[60] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$388 VDD INN|ONB|ONB[60] OUTP$61 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$389 OUTN$62 INP|ON|ON[61] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$390 VDD INN|ONB|ONB[61] OUTP$62 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$391 OUTN$63 INP|ON|ON[62] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$392 VDD INN|ONB|ONB[62] OUTP$63 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$393 OUTN$64 INP|ON|ON[63] VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$394 VDD INN|ONB|ONB[63] OUTP$64 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$395 OUTN$65 EN[1]|INP|ON VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p
+ AD=0.057p PS=1.75u PD=0.68u
M$396 VDD ENB[1]|INN|ONB OUTP$65 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$397 VcascP|VcascP[0] OUTN VcascodeP VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$398 VcascodeP OUTP VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$399 VcascP|VcascP[0] OUTN$1 VcascodeP$1 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$400 VcascodeP$1 OUTP$1 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$401 VcascP|VcascP[0] OUTN$2 VcascodeP$2 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$402 VcascodeP$2 OUTP$2 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$403 VcascP|VcascP[0] OUTN$3 VcascodeP$3 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$404 VcascodeP$3 OUTP$3 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$405 VcascP|VcascP[0] OUTN$4 VcascodeP$4 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$406 VcascodeP$4 OUTP$4 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$407 VcascP|VcascP[0] OUTN$5 VcascodeP$5 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$408 VcascodeP$5 OUTP$5 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$409 VcascP|VcascP[0] OUTN$6 VcascodeP$6 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$410 VcascodeP$6 OUTP$6 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$411 VcascP|VcascP[0] OUTN$7 VcascodeP$7 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$412 VcascodeP$7 OUTP$7 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$413 VcascP|VcascP[0] OUTN$8 VcascodeP$8 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$414 VcascodeP$8 OUTP$8 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$415 VcascP|VcascP[0] OUTN$9 VcascodeP$9 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$416 VcascodeP$9 OUTP$9 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$417 VcascP|VcascP[0] OUTN$10 VcascodeP$10 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$418 VcascodeP$10 OUTP$10 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$419 VcascP|VcascP[0] OUTN$11 VcascodeP$11 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$420 VcascodeP$11 OUTP$11 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$421 VcascP|VcascP[0] OUTN$12 VcascodeP$12 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$422 VcascodeP$12 OUTP$12 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$423 VcascP|VcascP[0] OUTN$13 VcascodeP$13 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$424 VcascodeP$13 OUTP$13 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$425 VcascP|VcascP[0] OUTN$14 VcascodeP$14 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$426 VcascodeP$14 OUTP$14 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$427 VcascP|VcascP[0] OUTN$15 VcascodeP$15 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$428 VcascodeP$15 OUTP$15 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$429 VcascP|VcascP[0] OUTN$16 VcascodeP$16 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$430 VcascodeP$16 OUTP$16 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$431 VcascP|VcascP[0] OUTN$17 VcascodeP$17 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$432 VcascodeP$17 OUTP$17 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$433 VcascP|VcascP[0] OUTN$18 VcascodeP$18 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$434 VcascodeP$18 OUTP$18 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$435 VcascP|VcascP[0] OUTN$19 VcascodeP$19 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$436 VcascodeP$19 OUTP$19 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$437 VcascP|VcascP[0] OUTN$20 VcascodeP$20 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$438 VcascodeP$20 OUTP$20 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$439 VcascP|VcascP[0] OUTN$21 VcascodeP$21 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$440 VcascodeP$21 OUTP$21 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$441 VcascP|VcascP[0] OUTN$22 VcascodeP$22 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$442 VcascodeP$22 OUTP$22 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$443 VcascP|VcascP[0] OUTN$23 VcascodeP$23 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$444 VcascodeP$23 OUTP$23 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$445 VcascP|VcascP[0] OUTN$24 VcascodeP$24 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$446 VcascodeP$24 OUTP$24 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$447 VcascP|VcascP[0] OUTN$25 VcascodeP$25 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$448 VcascodeP$25 OUTP$25 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$449 VcascP|VcascP[0] OUTN$26 VcascodeP$26 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$450 VcascodeP$26 OUTP$26 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$451 VcascP|VcascP[0] OUTN$27 VcascodeP$27 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$452 VcascodeP$27 OUTP$27 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$453 VcascP|VcascP[0] OUTN$28 VcascodeP$28 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$454 VcascodeP$28 OUTP$28 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$455 VcascP|VcascP[0] OUTN$29 VcascodeP$29 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$456 VcascodeP$29 OUTP$29 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$457 VcascP|VcascP[0] OUTN$30 VcascodeP$30 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$458 VcascodeP$30 OUTP$30 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$459 VcascP|VcascP[0] OUTN$31 VcascodeP$31 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$460 VcascodeP$31 OUTP$31 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$461 VcascP|VcascP[0] OUTN$32 VcascodeP$32 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$462 VcascodeP$32 OUTP$32 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$463 VcascP|VcascP[0] OUTN$33 VcascodeP$33 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$464 VcascodeP$33 OUTP$33 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$465 VcascP|VcascP[0] OUTN$34 VcascodeP$34 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$466 VcascodeP$34 OUTP$34 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$467 VcascP|VcascP[0] OUTN$35 VcascodeP$35 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$468 VcascodeP$35 OUTP$35 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$469 VcascP|VcascP[0] OUTN$36 VcascodeP$36 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$470 VcascodeP$36 OUTP$36 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$471 VcascP|VcascP[0] OUTN$37 VcascodeP$37 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$472 VcascodeP$37 OUTP$37 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$473 VcascP|VcascP[0] OUTN$38 VcascodeP$38 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$474 VcascodeP$38 OUTP$38 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$475 VcascP|VcascP[0] OUTN$39 VcascodeP$39 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$476 VcascodeP$39 OUTP$39 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$477 VcascP|VcascP[0] OUTN$40 VcascodeP$40 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$478 VcascodeP$40 OUTP$40 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$479 VcascP|VcascP[0] OUTN$41 VcascodeP$41 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$480 VcascodeP$41 OUTP$41 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$481 VcascP|VcascP[0] OUTN$42 VcascodeP$42 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$482 VcascodeP$42 OUTP$42 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$483 VcascP|VcascP[0] OUTN$43 VcascodeP$43 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$484 VcascodeP$43 OUTP$43 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$485 VcascP|VcascP[0] OUTN$44 VcascodeP$44 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$486 VcascodeP$44 OUTP$44 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$487 VcascP|VcascP[0] OUTN$45 VcascodeP$45 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$488 VcascodeP$45 OUTP$45 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$489 VcascP|VcascP[0] OUTN$46 VcascodeP$46 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$490 VcascodeP$46 OUTP$46 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$491 VcascP|VcascP[0] OUTN$47 VcascodeP$47 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$492 VcascodeP$47 OUTP$47 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$493 VcascP|VcascP[0] OUTN$48 VcascodeP$48 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$494 VcascodeP$48 OUTP$48 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$495 VcascP|VcascP[0] OUTN$49 VcascodeP$49 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$496 VcascodeP$49 OUTP$49 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$497 VcascP|VcascP[0] OUTN$50 VcascodeP$50 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$498 VcascodeP$50 OUTP$50 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$499 VcascP|VcascP[0] OUTN$51 VcascodeP$51 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$500 VcascodeP$51 OUTP$51 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$501 VcascP|VcascP[0] OUTN$52 VcascodeP$52 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$502 VcascodeP$52 OUTP$52 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$503 VcascP|VcascP[0] OUTN$53 VcascodeP$53 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$504 VcascodeP$53 OUTP$53 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$505 VcascP|VcascP[0] OUTN$54 VcascodeP$54 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$506 VcascodeP$54 OUTP$54 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$507 VcascP|VcascP[0] OUTN$55 VcascodeP$55 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$508 VcascodeP$55 OUTP$55 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$509 VcascP|VcascP[0] OUTN$56 VcascodeP$56 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$510 VcascodeP$56 OUTP$56 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$511 VcascP|VcascP[0] OUTN$57 VcascodeP$57 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$512 VcascodeP$57 OUTP$57 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$513 VcascP|VcascP[0] OUTN$58 VcascodeP$58 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$514 VcascodeP$58 OUTP$58 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$515 VcascP|VcascP[0] OUTN$59 VcascodeP$59 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$516 VcascodeP$59 OUTP$59 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$517 VcascP|VcascP[0] OUTN$60 VcascodeP$60 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$518 VcascodeP$60 OUTP$60 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$519 VcascP|VcascP[0] OUTN$61 VcascodeP$61 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$520 VcascodeP$61 OUTP$61 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$521 VcascP|VcascP[0] OUTN$62 VcascodeP$62 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$522 VcascodeP$62 OUTP$62 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$523 VcascP|VcascP[0] OUTN$63 VcascodeP$63 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$524 VcascodeP$63 OUTP$63 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$525 VcascP|VcascP[0] OUTN$64 VcascodeP$64 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$526 VcascodeP$64 OUTP$64 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$527 VcascP|VcascP[0] OUTN$65 VcascodeP$65 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.102p AD=0.057p PS=1.28u PD=0.68u
M$528 VcascodeP$65 OUTP$65 VDD VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.102p PS=0.68u PD=1.28u
M$529 VcascP|VcascP[0] VcascP|VcascP[0] Iout|VbiasP|VbiasP[0] VDD sg13_lv_pmos
+ L=0.15u W=11.7u AS=3.978p AD=3.978p PS=24.76u PD=24.76u
M$530 VDD Iout|VbiasP|VbiasP[0] \$340 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$531 \$340 VcascodeP Iout|VbiasP|VbiasP[0] VDD sg13_lv_pmos L=0.6u W=1.2u
+ AS=0.20875p AD=0.516p PS=1.75u PD=3.26u
M$532 VDD Iout|VbiasP|VbiasP[0] \$336 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$533 \$336 VcascodeP$1 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$534 VDD Iout|VbiasP|VbiasP[0] \$342 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$535 \$342 VcascodeP$2 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$536 VDD Iout|VbiasP|VbiasP[0] \$350 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$537 \$350 VcascodeP$3 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$538 VDD Iout|VbiasP|VbiasP[0] \$355 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$539 \$355 VcascodeP$4 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$540 VDD Iout|VbiasP|VbiasP[0] \$359 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$541 \$359 VcascodeP$5 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$542 VDD Iout|VbiasP|VbiasP[0] \$361 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$543 \$361 VcascodeP$6 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$544 VDD Iout|VbiasP|VbiasP[0] \$374 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$545 \$374 VcascodeP$7 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$546 VDD Iout|VbiasP|VbiasP[0] \$368 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$547 \$368 VcascodeP$8 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$548 VDD Iout|VbiasP|VbiasP[0] \$375 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$549 \$375 VcascodeP$9 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$550 VDD Iout|VbiasP|VbiasP[0] \$384 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$551 \$384 VcascodeP$10 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$552 VDD Iout|VbiasP|VbiasP[0] \$377 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$553 \$377 VcascodeP$11 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$554 VDD Iout|VbiasP|VbiasP[0] \$385 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$555 \$385 VcascodeP$12 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$556 VDD Iout|VbiasP|VbiasP[0] \$392 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$557 \$392 VcascodeP$13 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$558 VDD Iout|VbiasP|VbiasP[0] \$397 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$559 \$397 VcascodeP$14 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$560 VDD Iout|VbiasP|VbiasP[0] \$395 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$561 \$395 VcascodeP$15 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$562 VDD Iout|VbiasP|VbiasP[0] \$400 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$563 \$400 VcascodeP$16 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$564 VDD Iout|VbiasP|VbiasP[0] \$398 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$565 \$398 VcascodeP$17 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$566 VDD Iout|VbiasP|VbiasP[0] \$399 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$567 \$399 VcascodeP$18 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$568 VDD Iout|VbiasP|VbiasP[0] \$396 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$569 \$396 VcascodeP$19 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$570 VDD Iout|VbiasP|VbiasP[0] \$394 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$571 \$394 VcascodeP$20 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$572 VDD Iout|VbiasP|VbiasP[0] \$393 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$573 \$393 VcascodeP$21 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$574 VDD Iout|VbiasP|VbiasP[0] \$390 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$575 \$390 VcascodeP$22 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$576 VDD Iout|VbiasP|VbiasP[0] \$391 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$577 \$391 VcascodeP$23 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$578 VDD Iout|VbiasP|VbiasP[0] \$389 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$579 \$389 VcascodeP$24 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$580 VDD Iout|VbiasP|VbiasP[0] \$387 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$581 \$387 VcascodeP$25 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$582 VDD Iout|VbiasP|VbiasP[0] \$388 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$583 \$388 VcascodeP$26 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$584 VDD Iout|VbiasP|VbiasP[0] \$386 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$585 \$386 VcascodeP$27 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$586 VDD Iout|VbiasP|VbiasP[0] \$383 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$587 \$383 VcascodeP$28 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$588 VDD Iout|VbiasP|VbiasP[0] \$381 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$589 \$381 VcascodeP$29 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$590 VDD Iout|VbiasP|VbiasP[0] \$382 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$591 \$382 VcascodeP$30 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$592 VDD Iout|VbiasP|VbiasP[0] \$379 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$593 \$379 VcascodeP$31 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$594 VDD Iout|VbiasP|VbiasP[0] \$380 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$595 \$380 VcascodeP$32 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$596 VDD Iout|VbiasP|VbiasP[0] \$378 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$597 \$378 VcascodeP$33 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$598 VDD Iout|VbiasP|VbiasP[0] \$376 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$599 \$376 VcascodeP$34 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$600 VDD Iout|VbiasP|VbiasP[0] \$373 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$601 \$373 VcascodeP$35 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$602 VDD Iout|VbiasP|VbiasP[0] \$372 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$603 \$372 VcascodeP$36 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$604 VDD Iout|VbiasP|VbiasP[0] \$370 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$605 \$370 VcascodeP$37 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$606 VDD Iout|VbiasP|VbiasP[0] \$371 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$607 \$371 VcascodeP$38 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$608 VDD Iout|VbiasP|VbiasP[0] \$369 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$609 \$369 VcascodeP$39 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$610 VDD Iout|VbiasP|VbiasP[0] \$366 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$611 \$366 VcascodeP$40 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$612 VDD Iout|VbiasP|VbiasP[0] \$367 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$613 \$367 VcascodeP$41 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$614 VDD Iout|VbiasP|VbiasP[0] \$365 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$615 \$365 VcascodeP$42 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$616 VDD Iout|VbiasP|VbiasP[0] \$364 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$617 \$364 VcascodeP$43 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$618 VDD Iout|VbiasP|VbiasP[0] \$362 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$619 \$362 VcascodeP$44 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$620 VDD Iout|VbiasP|VbiasP[0] \$363 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$621 \$363 VcascodeP$45 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$622 VDD Iout|VbiasP|VbiasP[0] \$358 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$623 \$358 VcascodeP$46 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$624 VDD Iout|VbiasP|VbiasP[0] \$360 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$625 \$360 VcascodeP$47 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$626 VDD Iout|VbiasP|VbiasP[0] \$357 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$627 \$357 VcascodeP$48 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$628 VDD Iout|VbiasP|VbiasP[0] \$356 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$629 \$356 VcascodeP$49 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$630 VDD Iout|VbiasP|VbiasP[0] \$354 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$631 \$354 VcascodeP$50 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$632 VDD Iout|VbiasP|VbiasP[0] \$353 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$633 \$353 VcascodeP$51 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$634 VDD Iout|VbiasP|VbiasP[0] \$351 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$635 \$351 VcascodeP$52 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$636 VDD Iout|VbiasP|VbiasP[0] \$352 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$637 \$352 VcascodeP$53 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$638 VDD Iout|VbiasP|VbiasP[0] \$349 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$639 \$349 VcascodeP$54 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$640 VDD Iout|VbiasP|VbiasP[0] \$347 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$641 \$347 VcascodeP$55 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$642 VDD Iout|VbiasP|VbiasP[0] \$348 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$643 \$348 VcascodeP$56 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$644 VDD Iout|VbiasP|VbiasP[0] \$346 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$645 \$346 VcascodeP$57 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$646 VDD Iout|VbiasP|VbiasP[0] \$345 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$647 \$345 VcascodeP$58 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$648 VDD Iout|VbiasP|VbiasP[0] \$343 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$649 \$343 VcascodeP$59 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$650 VDD Iout|VbiasP|VbiasP[0] \$344 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$651 \$344 VcascodeP$60 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$652 VDD Iout|VbiasP|VbiasP[0] \$339 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$653 \$339 VcascodeP$61 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$654 VDD Iout|VbiasP|VbiasP[0] \$341 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$655 \$341 VcascodeP$62 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$656 VDD Iout|VbiasP|VbiasP[0] \$338 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$657 \$338 VcascodeP$63 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$658 VDD Iout|VbiasP|VbiasP[0] \$337 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$659 \$337 VcascodeP$64 Iout VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p
+ AD=0.516p PS=1.75u PD=3.26u
M$660 VDD Iout|VbiasP|VbiasP[0] \$335 VDD sg13_lv_pmos L=5u W=1.45u AS=0.493p
+ AD=0.20875p PS=3.58u PD=1.75u
M$661 \$335 VcascodeP$65 Iout|VbiasP|VbiasP[0] VDD sg13_lv_pmos L=0.6u W=1.2u
+ AS=0.20875p AD=0.516p PS=1.75u PD=3.26u
M$663 VcascP|VcascP[1] VcascP|VcascP[1] Iout|VbiasP|VbiasP[1] VDD sg13_lv_pmos
+ L=0.15u W=11.7u AS=3.978p AD=3.978p PS=24.76u PD=24.76u
M$664 Iout|VbiasP|VbiasP[1] VcascodeP$66 \$470 VDD sg13_lv_pmos L=0.6u W=1.2u
+ AS=0.516p AD=0.20875p PS=3.26u PD=1.75u
M$665 \$470 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$666 Iout VcascodeP$69 \$475 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$667 \$475 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$668 Iout VcascodeP$72 \$479 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$669 \$479 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$670 Iout VcascodeP$73 \$480 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$671 \$480 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$672 Iout VcascodeP$74 \$482 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$673 \$482 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$674 Iout VcascodeP$75 \$483 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$675 \$483 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$676 Iout VcascodeP$76 \$484 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$677 \$484 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$678 Iout VcascodeP$80 \$489 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$679 \$489 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$680 Iout VcascodeP$81 \$490 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$681 \$490 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$682 Iout VcascodeP$83 \$492 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$683 \$492 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$684 Iout VcascodeP$85 \$495 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$685 \$495 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$686 Iout VcascodeP$86 \$497 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$687 \$497 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$688 Iout VcascodeP$87 \$496 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$689 \$496 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$690 Iout VcascodeP$91 \$501 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$691 \$501 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$692 Iout VcascodeP$92 \$503 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$693 \$503 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$694 Iout VcascodeP$93 \$504 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$695 \$504 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$696 Iout VcascodeP$95 \$507 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$697 \$507 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$698 Iout VcascodeP$96 \$508 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$699 \$508 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$700 Iout VcascodeP$97 \$510 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$701 \$510 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$702 Iout VcascodeP$99 \$513 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$703 \$513 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$704 Iout VcascodeP$101 \$516 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$705 \$516 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$706 Iout VcascodeP$102 \$515 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$707 \$515 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$708 Iout VcascodeP$103 \$518 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$709 \$518 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$710 Iout VcascodeP$104 \$520 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$711 \$520 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$712 Iout VcascodeP$105 \$521 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$713 \$521 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$714 Iout VcascodeP$107 \$523 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$715 \$523 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$716 Iout VcascodeP$108 \$524 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$717 \$524 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$718 Iout VcascodeP$109 \$526 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$719 \$526 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$720 Iout VcascodeP$112 \$530 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$721 \$530 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$722 Iout VcascodeP$113 \$532 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$723 \$532 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$724 Iout VcascodeP$114 \$533 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$725 \$533 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$726 Iout VcascodeP$115 \$535 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$727 \$535 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$728 Iout VcascodeP$117 \$534 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$729 \$534 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$730 Iout VcascodeP$119 \$525 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$731 \$525 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$732 Iout VcascodeP$121 \$517 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$733 \$517 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$734 Iout VcascodeP$122 \$511 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$735 \$511 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$736 Iout VcascodeP$123 \$509 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$737 \$509 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$738 Iout VcascodeP$124 \$506 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$739 \$506 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$740 Iout VcascodeP$127 \$487 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$741 \$487 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$742 Iout VcascodeP$128 \$481 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$743 \$481 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$744 Iout VcascodeP$130 \$473 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$745 \$473 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$746 Iout|VbiasP|VbiasP[1] VcascodeP$131 \$471 VDD sg13_lv_pmos L=0.6u W=1.2u
+ AS=0.516p AD=0.20875p PS=3.26u PD=1.75u
M$747 \$471 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$749 Iout VcascodeP$67 \$472 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$750 \$472 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$751 Iout VcascodeP$68 \$474 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$752 \$474 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$753 Iout VcascodeP$70 \$476 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$754 \$476 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$755 Iout VcascodeP$71 \$478 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$756 \$478 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$757 Iout VcascodeP$77 \$485 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$758 \$485 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$759 Iout VcascodeP$78 \$486 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$760 \$486 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$761 Iout VcascodeP$79 \$488 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$762 \$488 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$763 Iout VcascodeP$82 \$491 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$764 \$491 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$765 Iout VcascodeP$84 \$494 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$766 \$494 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$767 Iout VcascodeP$88 \$498 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$768 \$498 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$769 Iout VcascodeP$89 \$499 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$770 \$499 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$771 Iout VcascodeP$90 \$500 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$772 \$500 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$773 Iout VcascodeP$94 \$505 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$774 \$505 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$775 Iout VcascodeP$98 \$512 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$776 \$512 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$777 Iout VcascodeP$100 \$514 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$778 \$514 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$779 Iout VcascodeP$106 \$522 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$780 \$522 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$781 Iout VcascodeP$110 \$527 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$782 \$527 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$783 Iout VcascodeP$111 \$529 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$784 \$529 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$785 Iout VcascodeP$116 \$531 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$786 \$531 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$787 Iout VcascodeP$118 \$528 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$788 \$528 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$789 Iout VcascodeP$120 \$519 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$790 \$519 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$791 Iout VcascodeP$125 \$502 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$792 \$502 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$793 Iout VcascodeP$126 \$493 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$794 \$493 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$795 Iout VcascodeP$129 \$477 VDD sg13_lv_pmos L=0.6u W=1.2u AS=0.516p
+ AD=0.20875p PS=3.26u PD=1.75u
M$796 \$477 Iout|VbiasP|VbiasP[1] VDD VDD sg13_lv_pmos L=5u W=1.45u AS=0.20875p
+ AD=0.493p PS=1.75u PD=3.58u
M$797 VDD OUTP$66 VcascodeP$66 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$798 VcascodeP$66 OUTN$66 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$799 VDD OUTP$67 VcascodeP$67 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$800 VcascodeP$67 OUTN$67 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$801 VDD OUTP$68 VcascodeP$68 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$802 VcascodeP$68 OUTN$68 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$803 VDD OUTP$69 VcascodeP$69 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$804 VcascodeP$69 OUTN$69 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$805 VDD OUTP$70 VcascodeP$70 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$806 VcascodeP$70 OUTN$70 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$807 VDD OUTP$71 VcascodeP$71 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$808 VcascodeP$71 OUTN$71 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$809 VDD OUTP$72 VcascodeP$72 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$810 VcascodeP$72 OUTN$72 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$811 VDD OUTP$73 VcascodeP$73 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$812 VcascodeP$73 OUTN$73 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$813 VDD OUTP$74 VcascodeP$74 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$814 VcascodeP$74 OUTN$74 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$815 VDD OUTP$75 VcascodeP$75 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$816 VcascodeP$75 OUTN$75 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$817 VDD OUTP$76 VcascodeP$76 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$818 VcascodeP$76 OUTN$76 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$819 VDD OUTP$77 VcascodeP$77 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$820 VcascodeP$77 OUTN$77 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$821 VDD OUTP$78 VcascodeP$78 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$822 VcascodeP$78 OUTN$78 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$823 VDD OUTP$79 VcascodeP$79 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$824 VcascodeP$79 OUTN$79 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$825 VDD OUTP$80 VcascodeP$80 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$826 VcascodeP$80 OUTN$80 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$827 VDD OUTP$81 VcascodeP$81 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$828 VcascodeP$81 OUTN$81 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$829 VDD OUTP$82 VcascodeP$82 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$830 VcascodeP$82 OUTN$82 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$831 VDD OUTP$83 VcascodeP$83 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$832 VcascodeP$83 OUTN$83 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$833 VDD OUTP$84 VcascodeP$84 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$834 VcascodeP$84 OUTN$84 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$835 VDD OUTP$85 VcascodeP$85 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$836 VcascodeP$85 OUTN$85 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$837 VDD OUTP$86 VcascodeP$86 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$838 VcascodeP$86 OUTN$86 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$839 VDD OUTP$87 VcascodeP$87 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$840 VcascodeP$87 OUTN$87 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$841 VDD OUTP$88 VcascodeP$88 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$842 VcascodeP$88 OUTN$88 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$843 VDD OUTP$89 VcascodeP$89 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$844 VcascodeP$89 OUTN$89 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$845 VDD OUTP$90 VcascodeP$90 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$846 VcascodeP$90 OUTN$90 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$847 VDD OUTP$91 VcascodeP$91 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$848 VcascodeP$91 OUTN$91 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$849 VDD OUTP$92 VcascodeP$92 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$850 VcascodeP$92 OUTN$92 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$851 VDD OUTP$93 VcascodeP$93 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$852 VcascodeP$93 OUTN$93 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$853 VDD OUTP$94 VcascodeP$94 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$854 VcascodeP$94 OUTN$94 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$855 VDD OUTP$95 VcascodeP$95 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$856 VcascodeP$95 OUTN$95 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$857 VDD OUTP$96 VcascodeP$96 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$858 VcascodeP$96 OUTN$96 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$859 VDD OUTP$97 VcascodeP$97 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$860 VcascodeP$97 OUTN$97 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$861 VDD OUTP$98 VcascodeP$98 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$862 VcascodeP$98 OUTN$98 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$863 VDD OUTP$99 VcascodeP$99 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$864 VcascodeP$99 OUTN$99 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$865 VDD OUTP$100 VcascodeP$100 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$866 VcascodeP$100 OUTN$100 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$867 VDD OUTP$101 VcascodeP$101 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$868 VcascodeP$101 OUTN$101 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$869 VDD OUTP$102 VcascodeP$102 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$870 VcascodeP$102 OUTN$102 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$871 VDD OUTP$103 VcascodeP$103 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$872 VcascodeP$103 OUTN$103 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$873 VDD OUTP$104 VcascodeP$104 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$874 VcascodeP$104 OUTN$104 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$875 VDD OUTP$105 VcascodeP$105 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$876 VcascodeP$105 OUTN$105 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$877 VDD OUTP$106 VcascodeP$106 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$878 VcascodeP$106 OUTN$106 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$879 VDD OUTP$107 VcascodeP$107 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$880 VcascodeP$107 OUTN$107 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$881 VDD OUTP$108 VcascodeP$108 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$882 VcascodeP$108 OUTN$108 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$883 VDD OUTP$109 VcascodeP$109 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$884 VcascodeP$109 OUTN$109 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$885 VDD OUTP$110 VcascodeP$110 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$886 VcascodeP$110 OUTN$110 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$887 VDD OUTP$111 VcascodeP$111 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$888 VcascodeP$111 OUTN$111 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$889 VDD OUTP$112 VcascodeP$112 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$890 VcascodeP$112 OUTN$112 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$891 VDD OUTP$113 VcascodeP$113 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$892 VcascodeP$113 OUTN$113 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$893 VDD OUTP$114 VcascodeP$114 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$894 VcascodeP$114 OUTN$114 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$895 VDD OUTP$115 VcascodeP$115 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$896 VcascodeP$115 OUTN$115 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$897 VDD OUTP$116 VcascodeP$116 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$898 VcascodeP$116 OUTN$116 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$899 VDD OUTP$117 VcascodeP$117 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$900 VcascodeP$117 OUTN$117 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$901 VDD OUTP$118 VcascodeP$118 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$902 VcascodeP$118 OUTN$118 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$903 VDD OUTP$119 VcascodeP$119 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$904 VcascodeP$119 OUTN$119 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$905 VDD OUTP$120 VcascodeP$120 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$906 VcascodeP$120 OUTN$120 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$907 VDD OUTP$121 VcascodeP$121 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$908 VcascodeP$121 OUTN$121 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$909 VDD OUTP$122 VcascodeP$122 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$910 VcascodeP$122 OUTN$122 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$911 VDD OUTP$123 VcascodeP$123 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$912 VcascodeP$123 OUTN$123 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$913 VDD OUTP$124 VcascodeP$124 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$914 VcascodeP$124 OUTN$124 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$915 VDD OUTP$125 VcascodeP$125 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$916 VcascodeP$125 OUTN$125 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$917 VDD OUTP$126 VcascodeP$126 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$918 VcascodeP$126 OUTN$126 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$919 VDD OUTP$127 VcascodeP$127 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$920 VcascodeP$127 OUTN$127 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$921 VDD OUTP$128 VcascodeP$128 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$922 VcascodeP$128 OUTN$128 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$923 VDD OUTP$129 VcascodeP$129 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$924 VcascodeP$129 OUTN$129 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$925 VDD OUTP$130 VcascodeP$130 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$926 VcascodeP$130 OUTN$130 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$927 VDD OUTP$131 VcascodeP$131 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.102p
+ AD=0.057p PS=1.28u PD=0.68u
M$928 VcascodeP$131 OUTN$131 VcascP|VcascP[1] VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.102p PS=0.68u PD=1.28u
M$929 OUTP$66 ENB[1]|ENB[3]|INN|ONB VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$930 VDD EN[1]|EN[3]|INP|ON OUTN$66 VDD sg13_lv_pmos L=0.13u W=0.3u AS=0.057p
+ AD=0.1725p PS=0.68u PD=1.75u
M$931 OUTP$67 INN|ONB|ONB[127]|ONB[63] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$932 VDD INP|ON|ON[127]|ON[63] OUTN$67 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$933 OUTP$68 INN|ONB|ONB[126]|ONB[62] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$934 VDD INP|ON|ON[126]|ON[62] OUTN$68 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$935 OUTP$69 INN|ONB|ONB[125]|ONB[61] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$936 VDD INP|ON|ON[125]|ON[61] OUTN$69 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$937 OUTP$70 INN|ONB|ONB[124]|ONB[60] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$938 VDD INP|ON|ON[124]|ON[60] OUTN$70 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$939 OUTP$71 INN|ONB|ONB[123]|ONB[59] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$940 VDD INP|ON|ON[123]|ON[59] OUTN$71 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$941 OUTP$72 INN|ONB|ONB[122]|ONB[58] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$942 VDD INP|ON|ON[122]|ON[58] OUTN$72 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$943 OUTP$73 INN|ONB|ONB[121]|ONB[57] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$944 VDD INP|ON|ON[121]|ON[57] OUTN$73 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$945 OUTP$74 INN|ONB|ONB[120]|ONB[56] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$946 VDD INP|ON|ON[120]|ON[56] OUTN$74 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$947 OUTP$75 INN|ONB|ONB[119]|ONB[55] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$948 VDD INP|ON|ON[119]|ON[55] OUTN$75 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$949 OUTP$76 INN|ONB|ONB[118]|ONB[54] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$950 VDD INP|ON|ON[118]|ON[54] OUTN$76 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$951 OUTP$77 INN|ONB|ONB[117]|ONB[53] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$952 VDD INP|ON|ON[117]|ON[53] OUTN$77 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$953 OUTP$78 INN|ONB|ONB[116]|ONB[52] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$954 VDD INP|ON|ON[116]|ON[52] OUTN$78 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$955 OUTP$79 INN|ONB|ONB[115]|ONB[51] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$956 VDD INP|ON|ON[115]|ON[51] OUTN$79 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$957 OUTP$80 INN|ONB|ONB[114]|ONB[50] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$958 VDD INP|ON|ON[114]|ON[50] OUTN$80 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$959 OUTP$81 INN|ONB|ONB[113]|ONB[49] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$960 VDD INP|ON|ON[113]|ON[49] OUTN$81 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$961 OUTP$82 INN|ONB|ONB[112]|ONB[48] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$962 VDD INP|ON|ON[112]|ON[48] OUTN$82 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$963 OUTP$83 INN|ONB|ONB[111]|ONB[47] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$964 VDD INP|ON|ON[111]|ON[47] OUTN$83 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$965 OUTP$84 INN|ONB|ONB[110]|ONB[46] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$966 VDD INP|ON|ON[110]|ON[46] OUTN$84 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$967 OUTP$85 INN|ONB|ONB[109]|ONB[45] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$968 VDD INP|ON|ON[109]|ON[45] OUTN$85 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$969 OUTP$86 INN|ONB|ONB[108]|ONB[44] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$970 VDD INP|ON|ON[108]|ON[44] OUTN$86 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$971 OUTP$87 INN|ONB|ONB[107]|ONB[43] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$972 VDD INP|ON|ON[107]|ON[43] OUTN$87 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$973 OUTP$88 INN|ONB|ONB[106]|ONB[42] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$974 VDD INP|ON|ON[106]|ON[42] OUTN$88 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$975 OUTP$89 INN|ONB|ONB[105]|ONB[41] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$976 VDD INP|ON|ON[105]|ON[41] OUTN$89 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$977 OUTP$90 INN|ONB|ONB[104]|ONB[40] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$978 VDD INP|ON|ON[104]|ON[40] OUTN$90 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$979 OUTP$91 INN|ONB|ONB[103]|ONB[39] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$980 VDD INP|ON|ON[103]|ON[39] OUTN$91 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$981 OUTP$92 INN|ONB|ONB[102]|ONB[38] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$982 VDD INP|ON|ON[102]|ON[38] OUTN$92 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$983 OUTP$93 INN|ONB|ONB[101]|ONB[37] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$984 VDD INP|ON|ON[101]|ON[37] OUTN$93 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$985 OUTP$94 INN|ONB|ONB[100]|ONB[36] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$986 VDD INP|ON|ON[100]|ON[36] OUTN$94 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$987 OUTP$95 INN|ONB|ONB[35]|ONB[99] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$988 VDD INP|ON|ON[35]|ON[99] OUTN$95 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$989 OUTP$96 INN|ONB|ONB[34]|ONB[98] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$990 VDD INP|ON|ON[34]|ON[98] OUTN$96 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$991 OUTP$97 INN|ONB|ONB[33]|ONB[97] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$992 VDD INP|ON|ON[33]|ON[97] OUTN$97 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$993 OUTP$98 INN|ONB|ONB[32]|ONB[96] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$994 VDD INP|ON|ON[32]|ON[96] OUTN$98 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$995 OUTP$99 INN|ONB|ONB[31]|ONB[95] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$996 VDD INP|ON|ON[31]|ON[95] OUTN$99 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$997 OUTP$100 INN|ONB|ONB[30]|ONB[94] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$998 VDD INP|ON|ON[30]|ON[94] OUTN$100 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$999 OUTP$101 INN|ONB|ONB[29]|ONB[93] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1000 VDD INP|ON|ON[29]|ON[93] OUTN$101 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1001 OUTP$102 INN|ONB|ONB[28]|ONB[92] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1002 VDD INP|ON|ON[28]|ON[92] OUTN$102 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1003 OUTP$103 INN|ONB|ONB[27]|ONB[91] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1004 VDD INP|ON|ON[27]|ON[91] OUTN$103 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1005 OUTP$104 INN|ONB|ONB[26]|ONB[90] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1006 VDD INP|ON|ON[26]|ON[90] OUTN$104 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1007 OUTP$105 INN|ONB|ONB[25]|ONB[89] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1008 VDD INP|ON|ON[25]|ON[89] OUTN$105 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1009 OUTP$106 INN|ONB|ONB[24]|ONB[88] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1010 VDD INP|ON|ON[24]|ON[88] OUTN$106 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1011 OUTP$107 INN|ONB|ONB[23]|ONB[87] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1012 VDD INP|ON|ON[23]|ON[87] OUTN$107 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1013 OUTP$108 INN|ONB|ONB[22]|ONB[86] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1014 VDD INP|ON|ON[22]|ON[86] OUTN$108 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1015 OUTP$109 INN|ONB|ONB[21]|ONB[85] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1016 VDD INP|ON|ON[21]|ON[85] OUTN$109 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1017 OUTP$110 INN|ONB|ONB[20]|ONB[84] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1018 VDD INP|ON|ON[20]|ON[84] OUTN$110 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1019 OUTP$111 INN|ONB|ONB[19]|ONB[83] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1020 VDD INP|ON|ON[19]|ON[83] OUTN$111 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1021 OUTP$112 INN|ONB|ONB[18]|ONB[82] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1022 VDD INP|ON|ON[18]|ON[82] OUTN$112 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1023 OUTP$113 INN|ONB|ONB[17]|ONB[81] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1024 VDD INP|ON|ON[17]|ON[81] OUTN$113 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1025 OUTP$114 INN|ONB|ONB[16]|ONB[80] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1026 VDD INP|ON|ON[16]|ON[80] OUTN$114 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1027 OUTP$115 INN|ONB|ONB[15]|ONB[79] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1028 VDD INP|ON|ON[15]|ON[79] OUTN$115 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1029 OUTP$116 INN|ONB|ONB[14]|ONB[78] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1030 VDD INP|ON|ON[14]|ON[78] OUTN$116 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1031 OUTP$117 INN|ONB|ONB[13]|ONB[77] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1032 VDD INP|ON|ON[13]|ON[77] OUTN$117 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1033 OUTP$118 INN|ONB|ONB[12]|ONB[76] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1034 VDD INP|ON|ON[12]|ON[76] OUTN$118 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1035 OUTP$119 INN|ONB|ONB[11]|ONB[75] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1036 VDD INP|ON|ON[11]|ON[75] OUTN$119 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1037 OUTP$120 INN|ONB|ONB[10]|ONB[74] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1038 VDD INP|ON|ON[10]|ON[74] OUTN$120 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1039 OUTP$121 INN|ONB|ONB[73]|ONB[9] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1040 VDD INP|ON|ON[73]|ON[9] OUTN$121 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1041 OUTP$122 INN|ONB|ONB[72]|ONB[8] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1042 VDD INP|ON|ON[72]|ON[8] OUTN$122 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1043 OUTP$123 INN|ONB|ONB[71]|ONB[7] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1044 VDD INP|ON|ON[71]|ON[7] OUTN$123 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1045 OUTP$124 INN|ONB|ONB[6]|ONB[70] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1046 VDD INP|ON|ON[6]|ON[70] OUTN$124 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1047 OUTP$125 INN|ONB|ONB[5]|ONB[69] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1048 VDD INP|ON|ON[5]|ON[69] OUTN$125 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1049 OUTP$126 INN|ONB|ONB[4]|ONB[68] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1050 VDD INP|ON|ON[4]|ON[68] OUTN$126 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1051 OUTP$127 INN|ONB|ONB[3]|ONB[67] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1052 VDD INP|ON|ON[3]|ON[67] OUTN$127 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1053 OUTP$128 INN|ONB|ONB[2]|ONB[66] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1054 VDD INP|ON|ON[2]|ON[66] OUTN$128 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1055 OUTP$129 INN|ONB|ONB[1]|ONB[65] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1056 VDD INP|ON|ON[1]|ON[65] OUTN$129 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1057 OUTP$130 INN|ONB|ONB[0]|ONB[64] VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1058 VDD INP|ON|ON[0]|ON[64] OUTN$130 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
M$1059 OUTP$131 ENB[0]|ENB[2]|INN|ONB VDD VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.1725p AD=0.057p PS=1.75u PD=0.68u
M$1060 VDD EN[0]|EN[2]|INP|ON OUTN$131 VDD sg13_lv_pmos L=0.13u W=0.3u
+ AS=0.057p AD=0.1725p PS=0.68u PD=1.75u
.ENDS dac128module
