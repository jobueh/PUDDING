magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757158256
<< metal1 >>
rect 576 38576 99360 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 8352 38576
rect 8392 38536 8434 38576
rect 8474 38536 8516 38576
rect 8556 38536 8598 38576
rect 8638 38536 8680 38576
rect 8720 38536 12352 38576
rect 12392 38536 12434 38576
rect 12474 38536 12516 38576
rect 12556 38536 12598 38576
rect 12638 38536 12680 38576
rect 12720 38536 16352 38576
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16720 38536 20352 38576
rect 20392 38536 20434 38576
rect 20474 38536 20516 38576
rect 20556 38536 20598 38576
rect 20638 38536 20680 38576
rect 20720 38536 24352 38576
rect 24392 38536 24434 38576
rect 24474 38536 24516 38576
rect 24556 38536 24598 38576
rect 24638 38536 24680 38576
rect 24720 38536 28352 38576
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28720 38536 32352 38576
rect 32392 38536 32434 38576
rect 32474 38536 32516 38576
rect 32556 38536 32598 38576
rect 32638 38536 32680 38576
rect 32720 38536 36352 38576
rect 36392 38536 36434 38576
rect 36474 38536 36516 38576
rect 36556 38536 36598 38576
rect 36638 38536 36680 38576
rect 36720 38536 40352 38576
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40720 38536 44352 38576
rect 44392 38536 44434 38576
rect 44474 38536 44516 38576
rect 44556 38536 44598 38576
rect 44638 38536 44680 38576
rect 44720 38536 48352 38576
rect 48392 38536 48434 38576
rect 48474 38536 48516 38576
rect 48556 38536 48598 38576
rect 48638 38536 48680 38576
rect 48720 38536 52352 38576
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52720 38536 56352 38576
rect 56392 38536 56434 38576
rect 56474 38536 56516 38576
rect 56556 38536 56598 38576
rect 56638 38536 56680 38576
rect 56720 38536 60352 38576
rect 60392 38536 60434 38576
rect 60474 38536 60516 38576
rect 60556 38536 60598 38576
rect 60638 38536 60680 38576
rect 60720 38536 64352 38576
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64720 38536 68352 38576
rect 68392 38536 68434 38576
rect 68474 38536 68516 38576
rect 68556 38536 68598 38576
rect 68638 38536 68680 38576
rect 68720 38536 72352 38576
rect 72392 38536 72434 38576
rect 72474 38536 72516 38576
rect 72556 38536 72598 38576
rect 72638 38536 72680 38576
rect 72720 38536 76352 38576
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76720 38536 80352 38576
rect 80392 38536 80434 38576
rect 80474 38536 80516 38576
rect 80556 38536 80598 38576
rect 80638 38536 80680 38576
rect 80720 38536 84352 38576
rect 84392 38536 84434 38576
rect 84474 38536 84516 38576
rect 84556 38536 84598 38576
rect 84638 38536 84680 38576
rect 84720 38536 88352 38576
rect 88392 38536 88434 38576
rect 88474 38536 88516 38576
rect 88556 38536 88598 38576
rect 88638 38536 88680 38576
rect 88720 38536 92352 38576
rect 92392 38536 92434 38576
rect 92474 38536 92516 38576
rect 92556 38536 92598 38576
rect 92638 38536 92680 38576
rect 92720 38536 96352 38576
rect 96392 38536 96434 38576
rect 96474 38536 96516 38576
rect 96556 38536 96598 38576
rect 96638 38536 96680 38576
rect 96720 38536 99360 38576
rect 576 38512 99360 38536
rect 576 37820 99516 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 7112 37820
rect 7152 37780 7194 37820
rect 7234 37780 7276 37820
rect 7316 37780 7358 37820
rect 7398 37780 7440 37820
rect 7480 37780 11112 37820
rect 11152 37780 11194 37820
rect 11234 37780 11276 37820
rect 11316 37780 11358 37820
rect 11398 37780 11440 37820
rect 11480 37780 15112 37820
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15480 37780 19112 37820
rect 19152 37780 19194 37820
rect 19234 37780 19276 37820
rect 19316 37780 19358 37820
rect 19398 37780 19440 37820
rect 19480 37780 23112 37820
rect 23152 37780 23194 37820
rect 23234 37780 23276 37820
rect 23316 37780 23358 37820
rect 23398 37780 23440 37820
rect 23480 37780 27112 37820
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27480 37780 31112 37820
rect 31152 37780 31194 37820
rect 31234 37780 31276 37820
rect 31316 37780 31358 37820
rect 31398 37780 31440 37820
rect 31480 37780 35112 37820
rect 35152 37780 35194 37820
rect 35234 37780 35276 37820
rect 35316 37780 35358 37820
rect 35398 37780 35440 37820
rect 35480 37780 39112 37820
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39480 37780 43112 37820
rect 43152 37780 43194 37820
rect 43234 37780 43276 37820
rect 43316 37780 43358 37820
rect 43398 37780 43440 37820
rect 43480 37780 47112 37820
rect 47152 37780 47194 37820
rect 47234 37780 47276 37820
rect 47316 37780 47358 37820
rect 47398 37780 47440 37820
rect 47480 37780 51112 37820
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51480 37780 55112 37820
rect 55152 37780 55194 37820
rect 55234 37780 55276 37820
rect 55316 37780 55358 37820
rect 55398 37780 55440 37820
rect 55480 37780 59112 37820
rect 59152 37780 59194 37820
rect 59234 37780 59276 37820
rect 59316 37780 59358 37820
rect 59398 37780 59440 37820
rect 59480 37780 63112 37820
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63480 37780 67112 37820
rect 67152 37780 67194 37820
rect 67234 37780 67276 37820
rect 67316 37780 67358 37820
rect 67398 37780 67440 37820
rect 67480 37780 71112 37820
rect 71152 37780 71194 37820
rect 71234 37780 71276 37820
rect 71316 37780 71358 37820
rect 71398 37780 71440 37820
rect 71480 37780 75112 37820
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75480 37780 79112 37820
rect 79152 37780 79194 37820
rect 79234 37780 79276 37820
rect 79316 37780 79358 37820
rect 79398 37780 79440 37820
rect 79480 37780 83112 37820
rect 83152 37780 83194 37820
rect 83234 37780 83276 37820
rect 83316 37780 83358 37820
rect 83398 37780 83440 37820
rect 83480 37780 87112 37820
rect 87152 37780 87194 37820
rect 87234 37780 87276 37820
rect 87316 37780 87358 37820
rect 87398 37780 87440 37820
rect 87480 37780 91112 37820
rect 91152 37780 91194 37820
rect 91234 37780 91276 37820
rect 91316 37780 91358 37820
rect 91398 37780 91440 37820
rect 91480 37780 95112 37820
rect 95152 37780 95194 37820
rect 95234 37780 95276 37820
rect 95316 37780 95358 37820
rect 95398 37780 95440 37820
rect 95480 37780 99112 37820
rect 99152 37780 99194 37820
rect 99234 37780 99276 37820
rect 99316 37780 99358 37820
rect 99398 37780 99440 37820
rect 99480 37780 99516 37820
rect 576 37756 99516 37780
rect 576 37064 99360 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 8352 37064
rect 8392 37024 8434 37064
rect 8474 37024 8516 37064
rect 8556 37024 8598 37064
rect 8638 37024 8680 37064
rect 8720 37024 12352 37064
rect 12392 37024 12434 37064
rect 12474 37024 12516 37064
rect 12556 37024 12598 37064
rect 12638 37024 12680 37064
rect 12720 37024 16352 37064
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16720 37024 20352 37064
rect 20392 37024 20434 37064
rect 20474 37024 20516 37064
rect 20556 37024 20598 37064
rect 20638 37024 20680 37064
rect 20720 37024 24352 37064
rect 24392 37024 24434 37064
rect 24474 37024 24516 37064
rect 24556 37024 24598 37064
rect 24638 37024 24680 37064
rect 24720 37024 28352 37064
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28720 37024 32352 37064
rect 32392 37024 32434 37064
rect 32474 37024 32516 37064
rect 32556 37024 32598 37064
rect 32638 37024 32680 37064
rect 32720 37024 36352 37064
rect 36392 37024 36434 37064
rect 36474 37024 36516 37064
rect 36556 37024 36598 37064
rect 36638 37024 36680 37064
rect 36720 37024 40352 37064
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40720 37024 44352 37064
rect 44392 37024 44434 37064
rect 44474 37024 44516 37064
rect 44556 37024 44598 37064
rect 44638 37024 44680 37064
rect 44720 37024 48352 37064
rect 48392 37024 48434 37064
rect 48474 37024 48516 37064
rect 48556 37024 48598 37064
rect 48638 37024 48680 37064
rect 48720 37024 52352 37064
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52720 37024 56352 37064
rect 56392 37024 56434 37064
rect 56474 37024 56516 37064
rect 56556 37024 56598 37064
rect 56638 37024 56680 37064
rect 56720 37024 60352 37064
rect 60392 37024 60434 37064
rect 60474 37024 60516 37064
rect 60556 37024 60598 37064
rect 60638 37024 60680 37064
rect 60720 37024 64352 37064
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64720 37024 68352 37064
rect 68392 37024 68434 37064
rect 68474 37024 68516 37064
rect 68556 37024 68598 37064
rect 68638 37024 68680 37064
rect 68720 37024 72352 37064
rect 72392 37024 72434 37064
rect 72474 37024 72516 37064
rect 72556 37024 72598 37064
rect 72638 37024 72680 37064
rect 72720 37024 76352 37064
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76720 37024 80352 37064
rect 80392 37024 80434 37064
rect 80474 37024 80516 37064
rect 80556 37024 80598 37064
rect 80638 37024 80680 37064
rect 80720 37024 84352 37064
rect 84392 37024 84434 37064
rect 84474 37024 84516 37064
rect 84556 37024 84598 37064
rect 84638 37024 84680 37064
rect 84720 37024 88352 37064
rect 88392 37024 88434 37064
rect 88474 37024 88516 37064
rect 88556 37024 88598 37064
rect 88638 37024 88680 37064
rect 88720 37024 92352 37064
rect 92392 37024 92434 37064
rect 92474 37024 92516 37064
rect 92556 37024 92598 37064
rect 92638 37024 92680 37064
rect 92720 37024 96352 37064
rect 96392 37024 96434 37064
rect 96474 37024 96516 37064
rect 96556 37024 96598 37064
rect 96638 37024 96680 37064
rect 96720 37024 99360 37064
rect 576 37000 99360 37024
rect 576 36308 99516 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 7112 36308
rect 7152 36268 7194 36308
rect 7234 36268 7276 36308
rect 7316 36268 7358 36308
rect 7398 36268 7440 36308
rect 7480 36268 11112 36308
rect 11152 36268 11194 36308
rect 11234 36268 11276 36308
rect 11316 36268 11358 36308
rect 11398 36268 11440 36308
rect 11480 36268 15112 36308
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15480 36268 19112 36308
rect 19152 36268 19194 36308
rect 19234 36268 19276 36308
rect 19316 36268 19358 36308
rect 19398 36268 19440 36308
rect 19480 36268 23112 36308
rect 23152 36268 23194 36308
rect 23234 36268 23276 36308
rect 23316 36268 23358 36308
rect 23398 36268 23440 36308
rect 23480 36268 27112 36308
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27480 36268 31112 36308
rect 31152 36268 31194 36308
rect 31234 36268 31276 36308
rect 31316 36268 31358 36308
rect 31398 36268 31440 36308
rect 31480 36268 35112 36308
rect 35152 36268 35194 36308
rect 35234 36268 35276 36308
rect 35316 36268 35358 36308
rect 35398 36268 35440 36308
rect 35480 36268 39112 36308
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39480 36268 43112 36308
rect 43152 36268 43194 36308
rect 43234 36268 43276 36308
rect 43316 36268 43358 36308
rect 43398 36268 43440 36308
rect 43480 36268 47112 36308
rect 47152 36268 47194 36308
rect 47234 36268 47276 36308
rect 47316 36268 47358 36308
rect 47398 36268 47440 36308
rect 47480 36268 51112 36308
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51480 36268 55112 36308
rect 55152 36268 55194 36308
rect 55234 36268 55276 36308
rect 55316 36268 55358 36308
rect 55398 36268 55440 36308
rect 55480 36268 59112 36308
rect 59152 36268 59194 36308
rect 59234 36268 59276 36308
rect 59316 36268 59358 36308
rect 59398 36268 59440 36308
rect 59480 36268 63112 36308
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63480 36268 67112 36308
rect 67152 36268 67194 36308
rect 67234 36268 67276 36308
rect 67316 36268 67358 36308
rect 67398 36268 67440 36308
rect 67480 36268 71112 36308
rect 71152 36268 71194 36308
rect 71234 36268 71276 36308
rect 71316 36268 71358 36308
rect 71398 36268 71440 36308
rect 71480 36268 75112 36308
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75480 36268 79112 36308
rect 79152 36268 79194 36308
rect 79234 36268 79276 36308
rect 79316 36268 79358 36308
rect 79398 36268 79440 36308
rect 79480 36268 83112 36308
rect 83152 36268 83194 36308
rect 83234 36268 83276 36308
rect 83316 36268 83358 36308
rect 83398 36268 83440 36308
rect 83480 36268 87112 36308
rect 87152 36268 87194 36308
rect 87234 36268 87276 36308
rect 87316 36268 87358 36308
rect 87398 36268 87440 36308
rect 87480 36268 91112 36308
rect 91152 36268 91194 36308
rect 91234 36268 91276 36308
rect 91316 36268 91358 36308
rect 91398 36268 91440 36308
rect 91480 36268 95112 36308
rect 95152 36268 95194 36308
rect 95234 36268 95276 36308
rect 95316 36268 95358 36308
rect 95398 36268 95440 36308
rect 95480 36268 99112 36308
rect 99152 36268 99194 36308
rect 99234 36268 99276 36308
rect 99316 36268 99358 36308
rect 99398 36268 99440 36308
rect 99480 36268 99516 36308
rect 576 36244 99516 36268
rect 74851 35972 74909 35973
rect 74851 35932 74860 35972
rect 74900 35932 74909 35972
rect 74851 35931 74909 35932
rect 76579 35972 76637 35973
rect 76579 35932 76588 35972
rect 76628 35932 76637 35972
rect 76579 35931 76637 35932
rect 77443 35972 77501 35973
rect 77443 35932 77452 35972
rect 77492 35932 77501 35972
rect 77443 35931 77501 35932
rect 78595 35972 78653 35973
rect 78595 35932 78604 35972
rect 78644 35932 78653 35972
rect 78595 35931 78653 35932
rect 79363 35972 79421 35973
rect 79363 35932 79372 35972
rect 79412 35932 79421 35972
rect 79363 35931 79421 35932
rect 81379 35972 81437 35973
rect 81379 35932 81388 35972
rect 81428 35932 81437 35972
rect 81379 35931 81437 35932
rect 85027 35972 85085 35973
rect 85027 35932 85036 35972
rect 85076 35932 85085 35972
rect 85027 35931 85085 35932
rect 85411 35972 85469 35973
rect 85411 35932 85420 35972
rect 85460 35932 85469 35972
rect 85411 35931 85469 35932
rect 92227 35972 92285 35973
rect 92227 35932 92236 35972
rect 92276 35932 92285 35972
rect 92227 35931 92285 35932
rect 80227 35888 80285 35889
rect 80227 35848 80236 35888
rect 80276 35848 80285 35888
rect 80227 35847 80285 35848
rect 86563 35888 86621 35889
rect 86563 35848 86572 35888
rect 86612 35848 86621 35888
rect 86563 35847 86621 35848
rect 87811 35888 87869 35889
rect 87811 35848 87820 35888
rect 87860 35848 87869 35888
rect 87811 35847 87869 35848
rect 89827 35888 89885 35889
rect 89827 35848 89836 35888
rect 89876 35848 89885 35888
rect 89827 35847 89885 35848
rect 90211 35888 90269 35889
rect 90211 35848 90220 35888
rect 90260 35848 90269 35888
rect 90211 35847 90269 35848
rect 93955 35888 94013 35889
rect 93955 35848 93964 35888
rect 94004 35848 94013 35888
rect 93955 35847 94013 35848
rect 94915 35888 94973 35889
rect 94915 35848 94924 35888
rect 94964 35848 94973 35888
rect 94915 35847 94973 35848
rect 75051 35720 75093 35729
rect 75051 35680 75052 35720
rect 75092 35680 75093 35720
rect 75051 35671 75093 35680
rect 76779 35720 76821 35729
rect 76779 35680 76780 35720
rect 76820 35680 76821 35720
rect 76779 35671 76821 35680
rect 77643 35720 77685 35729
rect 77643 35680 77644 35720
rect 77684 35680 77685 35720
rect 77643 35671 77685 35680
rect 78795 35720 78837 35729
rect 78795 35680 78796 35720
rect 78836 35680 78837 35720
rect 78795 35671 78837 35680
rect 79179 35720 79221 35729
rect 79179 35680 79180 35720
rect 79220 35680 79221 35720
rect 79179 35671 79221 35680
rect 80331 35720 80373 35729
rect 80331 35680 80332 35720
rect 80372 35680 80373 35720
rect 80331 35671 80373 35680
rect 81579 35720 81621 35729
rect 81579 35680 81580 35720
rect 81620 35680 81621 35720
rect 81579 35671 81621 35680
rect 85227 35720 85269 35729
rect 85227 35680 85228 35720
rect 85268 35680 85269 35720
rect 85227 35671 85269 35680
rect 85611 35720 85653 35729
rect 85611 35680 85612 35720
rect 85652 35680 85653 35720
rect 85611 35671 85653 35680
rect 86667 35720 86709 35729
rect 86667 35680 86668 35720
rect 86708 35680 86709 35720
rect 86667 35671 86709 35680
rect 87915 35720 87957 35729
rect 87915 35680 87916 35720
rect 87956 35680 87957 35720
rect 87915 35671 87957 35680
rect 89931 35720 89973 35729
rect 89931 35680 89932 35720
rect 89972 35680 89973 35720
rect 89931 35671 89973 35680
rect 90315 35720 90357 35729
rect 90315 35680 90316 35720
rect 90356 35680 90357 35720
rect 90315 35671 90357 35680
rect 92427 35720 92469 35729
rect 92427 35680 92428 35720
rect 92468 35680 92469 35720
rect 92427 35671 92469 35680
rect 93867 35720 93909 35729
rect 93867 35680 93868 35720
rect 93908 35680 93909 35720
rect 93867 35671 93909 35680
rect 95019 35720 95061 35729
rect 95019 35680 95020 35720
rect 95060 35680 95061 35720
rect 95019 35671 95061 35680
rect 576 35552 99360 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 8352 35552
rect 8392 35512 8434 35552
rect 8474 35512 8516 35552
rect 8556 35512 8598 35552
rect 8638 35512 8680 35552
rect 8720 35512 12352 35552
rect 12392 35512 12434 35552
rect 12474 35512 12516 35552
rect 12556 35512 12598 35552
rect 12638 35512 12680 35552
rect 12720 35512 16352 35552
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16720 35512 20352 35552
rect 20392 35512 20434 35552
rect 20474 35512 20516 35552
rect 20556 35512 20598 35552
rect 20638 35512 20680 35552
rect 20720 35512 24352 35552
rect 24392 35512 24434 35552
rect 24474 35512 24516 35552
rect 24556 35512 24598 35552
rect 24638 35512 24680 35552
rect 24720 35512 28352 35552
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28720 35512 32352 35552
rect 32392 35512 32434 35552
rect 32474 35512 32516 35552
rect 32556 35512 32598 35552
rect 32638 35512 32680 35552
rect 32720 35512 36352 35552
rect 36392 35512 36434 35552
rect 36474 35512 36516 35552
rect 36556 35512 36598 35552
rect 36638 35512 36680 35552
rect 36720 35512 40352 35552
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40720 35512 44352 35552
rect 44392 35512 44434 35552
rect 44474 35512 44516 35552
rect 44556 35512 44598 35552
rect 44638 35512 44680 35552
rect 44720 35512 48352 35552
rect 48392 35512 48434 35552
rect 48474 35512 48516 35552
rect 48556 35512 48598 35552
rect 48638 35512 48680 35552
rect 48720 35512 52352 35552
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52720 35512 56352 35552
rect 56392 35512 56434 35552
rect 56474 35512 56516 35552
rect 56556 35512 56598 35552
rect 56638 35512 56680 35552
rect 56720 35512 60352 35552
rect 60392 35512 60434 35552
rect 60474 35512 60516 35552
rect 60556 35512 60598 35552
rect 60638 35512 60680 35552
rect 60720 35512 64352 35552
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64720 35512 68352 35552
rect 68392 35512 68434 35552
rect 68474 35512 68516 35552
rect 68556 35512 68598 35552
rect 68638 35512 68680 35552
rect 68720 35512 72352 35552
rect 72392 35512 72434 35552
rect 72474 35512 72516 35552
rect 72556 35512 72598 35552
rect 72638 35512 72680 35552
rect 72720 35512 76352 35552
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76720 35512 80352 35552
rect 80392 35512 80434 35552
rect 80474 35512 80516 35552
rect 80556 35512 80598 35552
rect 80638 35512 80680 35552
rect 80720 35512 84352 35552
rect 84392 35512 84434 35552
rect 84474 35512 84516 35552
rect 84556 35512 84598 35552
rect 84638 35512 84680 35552
rect 84720 35512 88352 35552
rect 88392 35512 88434 35552
rect 88474 35512 88516 35552
rect 88556 35512 88598 35552
rect 88638 35512 88680 35552
rect 88720 35512 92352 35552
rect 92392 35512 92434 35552
rect 92474 35512 92516 35552
rect 92556 35512 92598 35552
rect 92638 35512 92680 35552
rect 92720 35512 96352 35552
rect 96392 35512 96434 35552
rect 96474 35512 96516 35552
rect 96556 35512 96598 35552
rect 96638 35512 96680 35552
rect 96720 35512 99360 35552
rect 576 35488 99360 35512
rect 79179 35384 79221 35393
rect 79179 35344 79180 35384
rect 79220 35344 79221 35384
rect 79179 35335 79221 35344
rect 88107 35384 88149 35393
rect 88107 35344 88108 35384
rect 88148 35344 88149 35384
rect 88107 35335 88149 35344
rect 93963 35384 94005 35393
rect 93963 35344 93964 35384
rect 94004 35344 94005 35384
rect 93963 35335 94005 35344
rect 76099 35216 76157 35217
rect 76099 35176 76108 35216
rect 76148 35176 76157 35216
rect 76099 35175 76157 35176
rect 76675 35216 76733 35217
rect 76675 35176 76684 35216
rect 76724 35176 76733 35216
rect 76675 35175 76733 35176
rect 77539 35216 77597 35217
rect 77539 35176 77548 35216
rect 77588 35176 77597 35216
rect 77539 35175 77597 35176
rect 78499 35216 78557 35217
rect 78499 35176 78508 35216
rect 78548 35176 78557 35216
rect 78499 35175 78557 35176
rect 79747 35216 79805 35217
rect 79747 35176 79756 35216
rect 79796 35176 79805 35216
rect 79747 35175 79805 35176
rect 80611 35216 80669 35217
rect 80611 35176 80620 35216
rect 80660 35176 80669 35216
rect 80611 35175 80669 35176
rect 81571 35216 81629 35217
rect 81571 35176 81580 35216
rect 81620 35176 81629 35216
rect 81571 35175 81629 35176
rect 82339 35216 82397 35217
rect 82339 35176 82348 35216
rect 82388 35176 82397 35216
rect 82339 35175 82397 35176
rect 84643 35216 84701 35217
rect 84643 35176 84652 35216
rect 84692 35176 84701 35216
rect 84643 35175 84701 35176
rect 85027 35216 85085 35217
rect 85027 35176 85036 35216
rect 85076 35176 85085 35216
rect 85027 35175 85085 35176
rect 85795 35216 85853 35217
rect 85795 35176 85804 35216
rect 85844 35176 85853 35216
rect 85795 35175 85853 35176
rect 87715 35216 87773 35217
rect 87715 35176 87724 35216
rect 87764 35176 87773 35216
rect 87715 35175 87773 35176
rect 91459 35216 91517 35217
rect 91459 35176 91468 35216
rect 91508 35176 91517 35216
rect 91459 35175 91517 35176
rect 92227 35216 92285 35217
rect 92227 35176 92236 35216
rect 92276 35176 92285 35216
rect 92227 35175 92285 35176
rect 93091 35216 93149 35217
rect 93091 35176 93100 35216
rect 93140 35176 93149 35216
rect 93091 35175 93149 35176
rect 94819 35216 94877 35217
rect 94819 35176 94828 35216
rect 94868 35176 94877 35216
rect 94819 35175 94877 35176
rect 95203 35216 95261 35217
rect 95203 35176 95212 35216
rect 95252 35176 95261 35216
rect 95203 35175 95261 35176
rect 97027 35216 97085 35217
rect 97027 35176 97036 35216
rect 97076 35176 97085 35216
rect 97027 35175 97085 35176
rect 73699 35132 73757 35133
rect 73699 35092 73708 35132
rect 73748 35092 73757 35132
rect 73699 35091 73757 35092
rect 74083 35132 74141 35133
rect 74083 35092 74092 35132
rect 74132 35092 74141 35132
rect 74083 35091 74141 35092
rect 74659 35132 74717 35133
rect 74659 35092 74668 35132
rect 74708 35092 74717 35132
rect 74659 35091 74717 35092
rect 75619 35132 75677 35133
rect 75619 35092 75628 35132
rect 75668 35092 75677 35132
rect 75619 35091 75677 35092
rect 77059 35132 77117 35133
rect 77059 35092 77068 35132
rect 77108 35092 77117 35132
rect 77059 35091 77117 35092
rect 78979 35132 79037 35133
rect 78979 35092 78988 35132
rect 79028 35092 79037 35132
rect 78979 35091 79037 35092
rect 79363 35132 79421 35133
rect 79363 35092 79372 35132
rect 79412 35092 79421 35132
rect 79363 35091 79421 35092
rect 80131 35132 80189 35133
rect 80131 35092 80140 35132
rect 80180 35092 80189 35132
rect 80131 35091 80189 35092
rect 80899 35132 80957 35133
rect 80899 35092 80908 35132
rect 80948 35092 80957 35132
rect 80899 35091 80957 35092
rect 81763 35132 81821 35133
rect 81763 35092 81772 35132
rect 81812 35092 81821 35132
rect 81763 35091 81821 35092
rect 82627 35132 82685 35133
rect 82627 35092 82636 35132
rect 82676 35092 82685 35132
rect 82627 35091 82685 35092
rect 83299 35132 83357 35133
rect 83299 35092 83308 35132
rect 83348 35092 83357 35132
rect 83299 35091 83357 35092
rect 83491 35132 83549 35133
rect 83491 35092 83500 35132
rect 83540 35092 83549 35132
rect 83491 35091 83549 35092
rect 83875 35132 83933 35133
rect 83875 35092 83884 35132
rect 83924 35092 83933 35132
rect 83875 35091 83933 35092
rect 84259 35132 84317 35133
rect 84259 35092 84268 35132
rect 84308 35092 84317 35132
rect 84259 35091 84317 35092
rect 86083 35132 86141 35133
rect 86083 35092 86092 35132
rect 86132 35092 86141 35132
rect 86083 35091 86141 35092
rect 86659 35132 86717 35133
rect 86659 35092 86668 35132
rect 86708 35092 86717 35132
rect 86659 35091 86717 35092
rect 87043 35132 87101 35133
rect 87043 35092 87052 35132
rect 87092 35092 87101 35132
rect 87043 35091 87101 35092
rect 87427 35132 87485 35133
rect 87427 35092 87436 35132
rect 87476 35092 87485 35132
rect 87427 35091 87485 35092
rect 87907 35132 87965 35133
rect 87907 35092 87916 35132
rect 87956 35092 87965 35132
rect 87907 35091 87965 35092
rect 88483 35132 88541 35133
rect 88483 35092 88492 35132
rect 88532 35092 88541 35132
rect 88483 35091 88541 35092
rect 88675 35132 88733 35133
rect 88675 35092 88684 35132
rect 88724 35092 88733 35132
rect 88675 35091 88733 35092
rect 89059 35132 89117 35133
rect 89059 35092 89068 35132
rect 89108 35092 89117 35132
rect 89059 35091 89117 35092
rect 89443 35132 89501 35133
rect 89443 35092 89452 35132
rect 89492 35092 89501 35132
rect 89443 35091 89501 35092
rect 89827 35132 89885 35133
rect 89827 35092 89836 35132
rect 89876 35092 89885 35132
rect 89827 35091 89885 35092
rect 90211 35132 90269 35133
rect 90211 35092 90220 35132
rect 90260 35092 90269 35132
rect 90211 35091 90269 35092
rect 90681 35129 90723 35138
rect 90681 35089 90682 35129
rect 90722 35089 90723 35129
rect 91075 35132 91133 35133
rect 91075 35092 91084 35132
rect 91124 35092 91133 35132
rect 91075 35091 91133 35092
rect 91747 35132 91805 35133
rect 91747 35092 91756 35132
rect 91796 35092 91805 35132
rect 91747 35091 91805 35092
rect 92611 35132 92669 35133
rect 92611 35092 92620 35132
rect 92660 35092 92669 35132
rect 92611 35091 92669 35092
rect 93379 35132 93437 35133
rect 93379 35092 93388 35132
rect 93428 35092 93437 35132
rect 93379 35091 93437 35092
rect 94147 35132 94205 35133
rect 94147 35092 94156 35132
rect 94196 35092 94205 35132
rect 94147 35091 94205 35092
rect 94531 35132 94589 35133
rect 94531 35092 94540 35132
rect 94580 35092 94589 35132
rect 94531 35091 94589 35092
rect 95395 35132 95453 35133
rect 95395 35092 95404 35132
rect 95444 35092 95453 35132
rect 95395 35091 95453 35092
rect 95779 35132 95837 35133
rect 95779 35092 95788 35132
rect 95828 35092 95837 35132
rect 95779 35091 95837 35092
rect 96163 35132 96221 35133
rect 96163 35092 96172 35132
rect 96212 35092 96221 35132
rect 96163 35091 96221 35092
rect 96547 35132 96605 35133
rect 96547 35092 96556 35132
rect 96596 35092 96605 35132
rect 96547 35091 96605 35092
rect 97795 35132 97853 35133
rect 97795 35092 97804 35132
rect 97844 35092 97853 35132
rect 97795 35091 97853 35092
rect 90681 35080 90723 35089
rect 74475 35048 74517 35057
rect 74475 35008 74476 35048
rect 74516 35008 74517 35048
rect 74475 34999 74517 35008
rect 77259 35048 77301 35057
rect 77259 35008 77260 35048
rect 77300 35008 77301 35048
rect 77259 34999 77301 35008
rect 86475 35048 86517 35057
rect 86475 35008 86476 35048
rect 86516 35008 86517 35048
rect 86475 34999 86517 35008
rect 73899 34964 73941 34973
rect 73899 34924 73900 34964
rect 73940 34924 73941 34964
rect 73899 34915 73941 34924
rect 74283 34964 74325 34973
rect 74283 34924 74284 34964
rect 74324 34924 74325 34964
rect 74283 34915 74325 34924
rect 75819 34964 75861 34973
rect 75819 34924 75820 34964
rect 75860 34924 75861 34964
rect 75819 34915 75861 34924
rect 76011 34964 76053 34973
rect 76011 34924 76012 34964
rect 76052 34924 76053 34964
rect 76011 34915 76053 34924
rect 76779 34964 76821 34973
rect 76779 34924 76780 34964
rect 76820 34924 76821 34964
rect 76779 34915 76821 34924
rect 77451 34964 77493 34973
rect 77451 34924 77452 34964
rect 77492 34924 77493 34964
rect 77451 34915 77493 34924
rect 78603 34964 78645 34973
rect 78603 34924 78604 34964
rect 78644 34924 78645 34964
rect 78603 34915 78645 34924
rect 79563 34964 79605 34973
rect 79563 34924 79564 34964
rect 79604 34924 79605 34964
rect 79563 34915 79605 34924
rect 79851 34964 79893 34973
rect 79851 34924 79852 34964
rect 79892 34924 79893 34964
rect 79851 34915 79893 34924
rect 80331 34964 80373 34973
rect 80331 34924 80332 34964
rect 80372 34924 80373 34964
rect 80331 34915 80373 34924
rect 80715 34964 80757 34973
rect 80715 34924 80716 34964
rect 80756 34924 80757 34964
rect 80715 34915 80757 34924
rect 81099 34964 81141 34973
rect 81099 34924 81100 34964
rect 81140 34924 81141 34964
rect 81099 34915 81141 34924
rect 81483 34964 81525 34973
rect 81483 34924 81484 34964
rect 81524 34924 81525 34964
rect 81483 34915 81525 34924
rect 81963 34964 82005 34973
rect 81963 34924 81964 34964
rect 82004 34924 82005 34964
rect 81963 34915 82005 34924
rect 82443 34964 82485 34973
rect 82443 34924 82444 34964
rect 82484 34924 82485 34964
rect 82443 34915 82485 34924
rect 82827 34964 82869 34973
rect 82827 34924 82828 34964
rect 82868 34924 82869 34964
rect 82827 34915 82869 34924
rect 83115 34964 83157 34973
rect 83115 34924 83116 34964
rect 83156 34924 83157 34964
rect 83115 34915 83157 34924
rect 83691 34964 83733 34973
rect 83691 34924 83692 34964
rect 83732 34924 83733 34964
rect 83691 34915 83733 34924
rect 84075 34964 84117 34973
rect 84075 34924 84076 34964
rect 84116 34924 84117 34964
rect 84075 34915 84117 34924
rect 84459 34964 84501 34973
rect 84459 34924 84460 34964
rect 84500 34924 84501 34964
rect 84459 34915 84501 34924
rect 84747 34964 84789 34973
rect 84747 34924 84748 34964
rect 84788 34924 84789 34964
rect 84747 34915 84789 34924
rect 85131 34964 85173 34973
rect 85131 34924 85132 34964
rect 85172 34924 85173 34964
rect 85131 34915 85173 34924
rect 85899 34964 85941 34973
rect 85899 34924 85900 34964
rect 85940 34924 85941 34964
rect 85899 34915 85941 34924
rect 86283 34964 86325 34973
rect 86283 34924 86284 34964
rect 86324 34924 86325 34964
rect 86283 34915 86325 34924
rect 86859 34964 86901 34973
rect 86859 34924 86860 34964
rect 86900 34924 86901 34964
rect 86859 34915 86901 34924
rect 87243 34964 87285 34973
rect 87243 34924 87244 34964
rect 87284 34924 87285 34964
rect 87243 34915 87285 34924
rect 87627 34964 87669 34973
rect 87627 34924 87628 34964
rect 87668 34924 87669 34964
rect 87627 34915 87669 34924
rect 88299 34964 88341 34973
rect 88299 34924 88300 34964
rect 88340 34924 88341 34964
rect 88299 34915 88341 34924
rect 88875 34964 88917 34973
rect 88875 34924 88876 34964
rect 88916 34924 88917 34964
rect 88875 34915 88917 34924
rect 89259 34964 89301 34973
rect 89259 34924 89260 34964
rect 89300 34924 89301 34964
rect 89259 34915 89301 34924
rect 89643 34964 89685 34973
rect 89643 34924 89644 34964
rect 89684 34924 89685 34964
rect 89643 34915 89685 34924
rect 90027 34964 90069 34973
rect 90027 34924 90028 34964
rect 90068 34924 90069 34964
rect 90027 34915 90069 34924
rect 90411 34964 90453 34973
rect 90411 34924 90412 34964
rect 90452 34924 90453 34964
rect 90411 34915 90453 34924
rect 90891 34964 90933 34973
rect 90891 34924 90892 34964
rect 90932 34924 90933 34964
rect 90891 34915 90933 34924
rect 91275 34964 91317 34973
rect 91275 34924 91276 34964
rect 91316 34924 91317 34964
rect 91275 34915 91317 34924
rect 91563 34964 91605 34973
rect 91563 34924 91564 34964
rect 91604 34924 91605 34964
rect 91563 34915 91605 34924
rect 91947 34964 91989 34973
rect 91947 34924 91948 34964
rect 91988 34924 91989 34964
rect 91947 34915 91989 34924
rect 92331 34964 92373 34973
rect 92331 34924 92332 34964
rect 92372 34924 92373 34964
rect 92331 34915 92373 34924
rect 92811 34964 92853 34973
rect 92811 34924 92812 34964
rect 92852 34924 92853 34964
rect 92811 34915 92853 34924
rect 93195 34964 93237 34973
rect 93195 34924 93196 34964
rect 93236 34924 93237 34964
rect 93195 34915 93237 34924
rect 93579 34964 93621 34973
rect 93579 34924 93580 34964
rect 93620 34924 93621 34964
rect 93579 34915 93621 34924
rect 93963 34964 94005 34973
rect 93963 34924 93964 34964
rect 94004 34924 94005 34964
rect 93963 34915 94005 34924
rect 94347 34964 94389 34973
rect 94347 34924 94348 34964
rect 94388 34924 94389 34964
rect 94347 34915 94389 34924
rect 94731 34964 94773 34973
rect 94731 34924 94732 34964
rect 94772 34924 94773 34964
rect 94731 34915 94773 34924
rect 95115 34964 95157 34973
rect 95115 34924 95116 34964
rect 95156 34924 95157 34964
rect 95115 34915 95157 34924
rect 95595 34964 95637 34973
rect 95595 34924 95596 34964
rect 95636 34924 95637 34964
rect 95595 34915 95637 34924
rect 95979 34964 96021 34973
rect 95979 34924 95980 34964
rect 96020 34924 96021 34964
rect 95979 34915 96021 34924
rect 96363 34964 96405 34973
rect 96363 34924 96364 34964
rect 96404 34924 96405 34964
rect 96363 34915 96405 34924
rect 96747 34964 96789 34973
rect 96747 34924 96748 34964
rect 96788 34924 96789 34964
rect 96747 34915 96789 34924
rect 96939 34964 96981 34973
rect 96939 34924 96940 34964
rect 96980 34924 96981 34964
rect 96939 34915 96981 34924
rect 97995 34964 98037 34973
rect 97995 34924 97996 34964
rect 98036 34924 98037 34964
rect 97995 34915 98037 34924
rect 576 34796 99516 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 7112 34796
rect 7152 34756 7194 34796
rect 7234 34756 7276 34796
rect 7316 34756 7358 34796
rect 7398 34756 7440 34796
rect 7480 34756 11112 34796
rect 11152 34756 11194 34796
rect 11234 34756 11276 34796
rect 11316 34756 11358 34796
rect 11398 34756 11440 34796
rect 11480 34756 15112 34796
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15480 34756 19112 34796
rect 19152 34756 19194 34796
rect 19234 34756 19276 34796
rect 19316 34756 19358 34796
rect 19398 34756 19440 34796
rect 19480 34756 23112 34796
rect 23152 34756 23194 34796
rect 23234 34756 23276 34796
rect 23316 34756 23358 34796
rect 23398 34756 23440 34796
rect 23480 34756 27112 34796
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27480 34756 31112 34796
rect 31152 34756 31194 34796
rect 31234 34756 31276 34796
rect 31316 34756 31358 34796
rect 31398 34756 31440 34796
rect 31480 34756 35112 34796
rect 35152 34756 35194 34796
rect 35234 34756 35276 34796
rect 35316 34756 35358 34796
rect 35398 34756 35440 34796
rect 35480 34756 39112 34796
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39480 34756 43112 34796
rect 43152 34756 43194 34796
rect 43234 34756 43276 34796
rect 43316 34756 43358 34796
rect 43398 34756 43440 34796
rect 43480 34756 47112 34796
rect 47152 34756 47194 34796
rect 47234 34756 47276 34796
rect 47316 34756 47358 34796
rect 47398 34756 47440 34796
rect 47480 34756 51112 34796
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51480 34756 55112 34796
rect 55152 34756 55194 34796
rect 55234 34756 55276 34796
rect 55316 34756 55358 34796
rect 55398 34756 55440 34796
rect 55480 34756 59112 34796
rect 59152 34756 59194 34796
rect 59234 34756 59276 34796
rect 59316 34756 59358 34796
rect 59398 34756 59440 34796
rect 59480 34756 63112 34796
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63480 34756 67112 34796
rect 67152 34756 67194 34796
rect 67234 34756 67276 34796
rect 67316 34756 67358 34796
rect 67398 34756 67440 34796
rect 67480 34756 71112 34796
rect 71152 34756 71194 34796
rect 71234 34756 71276 34796
rect 71316 34756 71358 34796
rect 71398 34756 71440 34796
rect 71480 34756 75112 34796
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75480 34756 79112 34796
rect 79152 34756 79194 34796
rect 79234 34756 79276 34796
rect 79316 34756 79358 34796
rect 79398 34756 79440 34796
rect 79480 34756 83112 34796
rect 83152 34756 83194 34796
rect 83234 34756 83276 34796
rect 83316 34756 83358 34796
rect 83398 34756 83440 34796
rect 83480 34756 87112 34796
rect 87152 34756 87194 34796
rect 87234 34756 87276 34796
rect 87316 34756 87358 34796
rect 87398 34756 87440 34796
rect 87480 34756 91112 34796
rect 91152 34756 91194 34796
rect 91234 34756 91276 34796
rect 91316 34756 91358 34796
rect 91398 34756 91440 34796
rect 91480 34756 95112 34796
rect 95152 34756 95194 34796
rect 95234 34756 95276 34796
rect 95316 34756 95358 34796
rect 95398 34756 95440 34796
rect 95480 34756 99112 34796
rect 99152 34756 99194 34796
rect 99234 34756 99276 34796
rect 99316 34756 99358 34796
rect 99398 34756 99440 34796
rect 99480 34756 99516 34796
rect 576 34732 99516 34756
rect 83307 34628 83349 34637
rect 83307 34588 83308 34628
rect 83348 34588 83349 34628
rect 83307 34579 83349 34588
rect 86379 34628 86421 34637
rect 86379 34588 86380 34628
rect 86420 34588 86421 34628
rect 86379 34579 86421 34588
rect 92427 34628 92469 34637
rect 92427 34588 92428 34628
rect 92468 34588 92469 34628
rect 92427 34579 92469 34588
rect 95883 34628 95925 34637
rect 95883 34588 95884 34628
rect 95924 34588 95925 34628
rect 95883 34579 95925 34588
rect 80619 34544 80661 34553
rect 80619 34504 80620 34544
rect 80660 34504 80661 34544
rect 80619 34495 80661 34504
rect 81867 34544 81909 34553
rect 81867 34504 81868 34544
rect 81908 34504 81909 34544
rect 81867 34495 81909 34504
rect 85227 34544 85269 34553
rect 85227 34504 85228 34544
rect 85268 34504 85269 34544
rect 85227 34495 85269 34504
rect 89163 34544 89205 34553
rect 89163 34504 89164 34544
rect 89204 34504 89205 34544
rect 89163 34495 89205 34504
rect 91179 34544 91221 34553
rect 91179 34504 91180 34544
rect 91220 34504 91221 34544
rect 91179 34495 91221 34504
rect 96459 34544 96501 34553
rect 96459 34504 96460 34544
rect 96500 34504 96501 34544
rect 96459 34495 96501 34504
rect 96843 34544 96885 34553
rect 96843 34504 96844 34544
rect 96884 34504 96885 34544
rect 96843 34495 96885 34504
rect 82243 34471 82301 34472
rect 73411 34460 73469 34461
rect 73411 34420 73420 34460
rect 73460 34420 73469 34460
rect 73411 34419 73469 34420
rect 73891 34460 73949 34461
rect 73891 34420 73900 34460
rect 73940 34420 73949 34460
rect 73891 34419 73949 34420
rect 74659 34460 74717 34461
rect 74659 34420 74668 34460
rect 74708 34420 74717 34460
rect 74659 34419 74717 34420
rect 75139 34460 75197 34461
rect 75139 34420 75148 34460
rect 75188 34420 75197 34460
rect 75139 34419 75197 34420
rect 76195 34460 76253 34461
rect 76195 34420 76204 34460
rect 76244 34420 76253 34460
rect 76195 34419 76253 34420
rect 76963 34460 77021 34461
rect 76963 34420 76972 34460
rect 77012 34420 77021 34460
rect 76963 34419 77021 34420
rect 77827 34460 77885 34461
rect 77827 34420 77836 34460
rect 77876 34420 77885 34460
rect 77827 34419 77885 34420
rect 78211 34460 78269 34461
rect 78211 34420 78220 34460
rect 78260 34420 78269 34460
rect 78211 34419 78269 34420
rect 79747 34460 79805 34461
rect 79747 34420 79756 34460
rect 79796 34420 79805 34460
rect 79747 34419 79805 34420
rect 80419 34460 80477 34461
rect 80419 34420 80428 34460
rect 80468 34420 80477 34460
rect 80419 34419 80477 34420
rect 80995 34460 81053 34461
rect 80995 34420 81004 34460
rect 81044 34420 81053 34460
rect 80995 34419 81053 34420
rect 81475 34460 81533 34461
rect 81475 34420 81484 34460
rect 81524 34420 81533 34460
rect 81475 34419 81533 34420
rect 82051 34460 82109 34461
rect 82051 34420 82060 34460
rect 82100 34420 82109 34460
rect 82243 34431 82252 34471
rect 82292 34431 82301 34471
rect 82243 34430 82301 34431
rect 83107 34460 83165 34461
rect 82051 34419 82109 34420
rect 83107 34420 83116 34460
rect 83156 34420 83165 34460
rect 83107 34419 83165 34420
rect 84643 34460 84701 34461
rect 84643 34420 84652 34460
rect 84692 34420 84701 34460
rect 84643 34419 84701 34420
rect 85027 34460 85085 34461
rect 85027 34420 85036 34460
rect 85076 34420 85085 34460
rect 85027 34419 85085 34420
rect 85795 34460 85853 34461
rect 85795 34420 85804 34460
rect 85844 34420 85853 34460
rect 85795 34419 85853 34420
rect 86563 34460 86621 34461
rect 86563 34420 86572 34460
rect 86612 34420 86621 34460
rect 86563 34419 86621 34420
rect 87811 34460 87869 34461
rect 87811 34420 87820 34460
rect 87860 34420 87869 34460
rect 87811 34419 87869 34420
rect 88291 34460 88349 34461
rect 88291 34420 88300 34460
rect 88340 34420 88349 34460
rect 88291 34419 88349 34420
rect 89347 34460 89405 34461
rect 89347 34420 89356 34460
rect 89396 34420 89405 34460
rect 89347 34419 89405 34420
rect 90499 34460 90557 34461
rect 90499 34420 90508 34460
rect 90548 34420 90557 34460
rect 90499 34419 90557 34420
rect 90979 34460 91037 34461
rect 90979 34420 90988 34460
rect 91028 34420 91037 34460
rect 90979 34419 91037 34420
rect 92227 34460 92285 34461
rect 92227 34420 92236 34460
rect 92276 34420 92285 34460
rect 92227 34419 92285 34420
rect 93091 34460 93149 34461
rect 93091 34420 93100 34460
rect 93140 34420 93149 34460
rect 93091 34419 93149 34420
rect 93859 34460 93917 34461
rect 93859 34420 93868 34460
rect 93908 34420 93917 34460
rect 93859 34419 93917 34420
rect 94627 34460 94685 34461
rect 94627 34420 94636 34460
rect 94676 34420 94685 34460
rect 94627 34419 94685 34420
rect 95011 34460 95069 34461
rect 95011 34420 95020 34460
rect 95060 34420 95069 34460
rect 95011 34419 95069 34420
rect 96067 34460 96125 34461
rect 96067 34420 96076 34460
rect 96116 34420 96125 34460
rect 96067 34419 96125 34420
rect 96259 34460 96317 34461
rect 96259 34420 96268 34460
rect 96308 34420 96317 34460
rect 96259 34419 96317 34420
rect 97027 34460 97085 34461
rect 97027 34420 97036 34460
rect 97076 34420 97085 34460
rect 97027 34419 97085 34420
rect 97507 34460 97565 34461
rect 97507 34420 97516 34460
rect 97556 34420 97565 34460
rect 97507 34419 97565 34420
rect 98659 34460 98717 34461
rect 98659 34420 98668 34460
rect 98708 34420 98717 34460
rect 98659 34419 98717 34420
rect 75619 34376 75677 34377
rect 74848 34365 74906 34366
rect 74848 34325 74857 34365
rect 74897 34325 74906 34365
rect 75619 34336 75628 34376
rect 75668 34336 75677 34376
rect 75619 34335 75677 34336
rect 75907 34376 75965 34377
rect 75907 34336 75916 34376
rect 75956 34336 75965 34376
rect 75907 34335 75965 34336
rect 76675 34376 76733 34377
rect 76675 34336 76684 34376
rect 76724 34336 76733 34376
rect 76675 34335 76733 34336
rect 77539 34376 77597 34377
rect 77539 34336 77548 34376
rect 77588 34336 77597 34376
rect 77539 34335 77597 34336
rect 78691 34376 78749 34377
rect 78691 34336 78700 34376
rect 78740 34336 78749 34376
rect 78691 34335 78749 34336
rect 78883 34376 78941 34377
rect 78883 34336 78892 34376
rect 78932 34336 78941 34376
rect 78883 34335 78941 34336
rect 79363 34376 79421 34377
rect 79363 34336 79372 34376
rect 79412 34336 79421 34376
rect 79363 34335 79421 34336
rect 80126 34373 80168 34382
rect 89923 34377 89981 34378
rect 74848 34324 74906 34325
rect 80126 34333 80127 34373
rect 80167 34333 80168 34373
rect 81187 34376 81245 34377
rect 81187 34336 81196 34376
rect 81236 34336 81245 34376
rect 81187 34335 81245 34336
rect 82627 34376 82685 34377
rect 82627 34336 82636 34376
rect 82676 34336 82685 34376
rect 82627 34335 82685 34336
rect 83587 34376 83645 34377
rect 83587 34336 83596 34376
rect 83636 34336 83645 34376
rect 83587 34335 83645 34336
rect 83875 34376 83933 34377
rect 83875 34336 83884 34376
rect 83924 34336 83933 34376
rect 83875 34335 83933 34336
rect 84163 34376 84221 34377
rect 84163 34336 84172 34376
rect 84212 34336 84221 34376
rect 84163 34335 84221 34336
rect 84451 34376 84509 34377
rect 84451 34336 84460 34376
rect 84500 34336 84509 34376
rect 84451 34335 84509 34336
rect 85411 34376 85469 34377
rect 85411 34336 85420 34376
rect 85460 34336 85469 34376
rect 85411 34335 85469 34336
rect 86851 34376 86909 34377
rect 86851 34336 86860 34376
rect 86900 34336 86909 34376
rect 86851 34335 86909 34336
rect 87043 34376 87101 34377
rect 87043 34336 87052 34376
rect 87092 34336 87101 34376
rect 87043 34335 87101 34336
rect 87331 34376 87389 34377
rect 87331 34336 87340 34376
rect 87380 34336 87389 34376
rect 87331 34335 87389 34336
rect 88675 34376 88733 34377
rect 88675 34336 88684 34376
rect 88724 34336 88733 34376
rect 88675 34335 88733 34336
rect 89635 34376 89693 34377
rect 89635 34336 89644 34376
rect 89684 34336 89693 34376
rect 89923 34337 89932 34377
rect 89972 34337 89981 34377
rect 89923 34336 89981 34337
rect 90211 34376 90269 34377
rect 90211 34336 90220 34376
rect 90260 34336 90269 34376
rect 89635 34335 89693 34336
rect 90211 34335 90269 34336
rect 91459 34376 91517 34377
rect 91459 34336 91468 34376
rect 91508 34336 91517 34376
rect 91459 34335 91517 34336
rect 91747 34376 91805 34377
rect 91747 34336 91756 34376
rect 91796 34336 91805 34376
rect 91747 34335 91805 34336
rect 92035 34376 92093 34377
rect 92035 34336 92044 34376
rect 92084 34336 92093 34376
rect 92035 34335 92093 34336
rect 92611 34376 92669 34377
rect 92611 34336 92620 34376
rect 92660 34336 92669 34376
rect 92611 34335 92669 34336
rect 92803 34376 92861 34377
rect 92803 34336 92812 34376
rect 92852 34336 92861 34376
rect 92803 34335 92861 34336
rect 93571 34376 93629 34377
rect 93571 34336 93580 34376
rect 93620 34336 93629 34376
rect 93571 34335 93629 34336
rect 94243 34376 94301 34377
rect 94243 34336 94252 34376
rect 94292 34336 94301 34376
rect 94243 34335 94301 34336
rect 95587 34376 95645 34377
rect 95587 34336 95596 34376
rect 95636 34336 95645 34376
rect 95587 34335 95645 34336
rect 96739 34376 96797 34377
rect 96739 34336 96748 34376
rect 96788 34336 96797 34376
rect 96739 34335 96797 34336
rect 97891 34376 97949 34377
rect 97891 34336 97900 34376
rect 97940 34336 97949 34376
rect 97891 34335 97949 34336
rect 98275 34376 98333 34377
rect 98275 34336 98284 34376
rect 98324 34336 98333 34376
rect 98275 34335 98333 34336
rect 98851 34376 98909 34377
rect 98851 34336 98860 34376
rect 98900 34336 98909 34376
rect 98851 34335 98909 34336
rect 99139 34376 99197 34377
rect 99139 34336 99148 34376
rect 99188 34336 99197 34376
rect 99139 34335 99197 34336
rect 80126 34324 80168 34333
rect 80235 34292 80277 34301
rect 80235 34252 80236 34292
rect 80276 34252 80277 34292
rect 80235 34243 80277 34252
rect 73611 34208 73653 34217
rect 73611 34168 73612 34208
rect 73652 34168 73653 34208
rect 73611 34159 73653 34168
rect 74091 34208 74133 34217
rect 74091 34168 74092 34208
rect 74132 34168 74133 34208
rect 74091 34159 74133 34168
rect 74475 34208 74517 34217
rect 74475 34168 74476 34208
rect 74516 34168 74517 34208
rect 74475 34159 74517 34168
rect 74955 34208 74997 34217
rect 74955 34168 74956 34208
rect 74996 34168 74997 34208
rect 74955 34159 74997 34168
rect 75339 34208 75381 34217
rect 75339 34168 75340 34208
rect 75380 34168 75381 34208
rect 75339 34159 75381 34168
rect 75531 34208 75573 34217
rect 75531 34168 75532 34208
rect 75572 34168 75573 34208
rect 75531 34159 75573 34168
rect 76011 34208 76053 34217
rect 76011 34168 76012 34208
rect 76052 34168 76053 34208
rect 76011 34159 76053 34168
rect 76395 34208 76437 34217
rect 76395 34168 76396 34208
rect 76436 34168 76437 34208
rect 76395 34159 76437 34168
rect 76779 34208 76821 34217
rect 76779 34168 76780 34208
rect 76820 34168 76821 34208
rect 76779 34159 76821 34168
rect 77163 34208 77205 34217
rect 77163 34168 77164 34208
rect 77204 34168 77205 34208
rect 77163 34159 77205 34168
rect 77643 34208 77685 34217
rect 77643 34168 77644 34208
rect 77684 34168 77685 34208
rect 77643 34159 77685 34168
rect 78027 34208 78069 34217
rect 78027 34168 78028 34208
rect 78068 34168 78069 34208
rect 78027 34159 78069 34168
rect 78411 34208 78453 34217
rect 78411 34168 78412 34208
rect 78452 34168 78453 34208
rect 78411 34159 78453 34168
rect 78603 34208 78645 34217
rect 78603 34168 78604 34208
rect 78644 34168 78645 34208
rect 78603 34159 78645 34168
rect 78987 34208 79029 34217
rect 78987 34168 78988 34208
rect 79028 34168 79029 34208
rect 78987 34159 79029 34168
rect 79467 34208 79509 34217
rect 79467 34168 79468 34208
rect 79508 34168 79509 34208
rect 79467 34159 79509 34168
rect 79947 34208 79989 34217
rect 79947 34168 79948 34208
rect 79988 34168 79989 34208
rect 79947 34159 79989 34168
rect 80811 34208 80853 34217
rect 80811 34168 80812 34208
rect 80852 34168 80853 34208
rect 80811 34159 80853 34168
rect 81291 34208 81333 34217
rect 81291 34168 81292 34208
rect 81332 34168 81333 34208
rect 81291 34159 81333 34168
rect 81675 34208 81717 34217
rect 81675 34168 81676 34208
rect 81716 34168 81717 34208
rect 81675 34159 81717 34168
rect 82443 34208 82485 34217
rect 82443 34168 82444 34208
rect 82484 34168 82485 34208
rect 82443 34159 82485 34168
rect 82731 34208 82773 34217
rect 82731 34168 82732 34208
rect 82772 34168 82773 34208
rect 82731 34159 82773 34168
rect 83499 34208 83541 34217
rect 83499 34168 83500 34208
rect 83540 34168 83541 34208
rect 83499 34159 83541 34168
rect 83787 34208 83829 34217
rect 83787 34168 83788 34208
rect 83828 34168 83829 34208
rect 83787 34159 83829 34168
rect 84075 34208 84117 34217
rect 84075 34168 84076 34208
rect 84116 34168 84117 34208
rect 84075 34159 84117 34168
rect 84363 34208 84405 34217
rect 84363 34168 84364 34208
rect 84404 34168 84405 34208
rect 84363 34159 84405 34168
rect 84843 34208 84885 34217
rect 84843 34168 84844 34208
rect 84884 34168 84885 34208
rect 84843 34159 84885 34168
rect 85515 34208 85557 34217
rect 85515 34168 85516 34208
rect 85556 34168 85557 34208
rect 85515 34159 85557 34168
rect 85995 34208 86037 34217
rect 85995 34168 85996 34208
rect 86036 34168 86037 34208
rect 85995 34159 86037 34168
rect 86763 34208 86805 34217
rect 86763 34168 86764 34208
rect 86804 34168 86805 34208
rect 86763 34159 86805 34168
rect 87147 34208 87189 34217
rect 87147 34168 87148 34208
rect 87188 34168 87189 34208
rect 87147 34159 87189 34168
rect 87435 34208 87477 34217
rect 87435 34168 87436 34208
rect 87476 34168 87477 34208
rect 87435 34159 87477 34168
rect 88011 34208 88053 34217
rect 88011 34168 88012 34208
rect 88052 34168 88053 34208
rect 88011 34159 88053 34168
rect 88491 34208 88533 34217
rect 88491 34168 88492 34208
rect 88532 34168 88533 34208
rect 88491 34159 88533 34168
rect 88779 34208 88821 34217
rect 88779 34168 88780 34208
rect 88820 34168 88821 34208
rect 88779 34159 88821 34168
rect 89547 34208 89589 34217
rect 89547 34168 89548 34208
rect 89588 34168 89589 34208
rect 89547 34159 89589 34168
rect 89835 34208 89877 34217
rect 89835 34168 89836 34208
rect 89876 34168 89877 34208
rect 89835 34159 89877 34168
rect 90315 34208 90357 34217
rect 90315 34168 90316 34208
rect 90356 34168 90357 34208
rect 90315 34159 90357 34168
rect 90699 34208 90741 34217
rect 90699 34168 90700 34208
rect 90740 34168 90741 34208
rect 90699 34159 90741 34168
rect 91371 34208 91413 34217
rect 91371 34168 91372 34208
rect 91412 34168 91413 34208
rect 91371 34159 91413 34168
rect 91659 34208 91701 34217
rect 91659 34168 91660 34208
rect 91700 34168 91701 34208
rect 91659 34159 91701 34168
rect 91947 34208 91989 34217
rect 91947 34168 91948 34208
rect 91988 34168 91989 34208
rect 91947 34159 91989 34168
rect 93291 34208 93333 34217
rect 93291 34168 93292 34208
rect 93332 34168 93333 34208
rect 93291 34159 93333 34168
rect 93483 34208 93525 34217
rect 93483 34168 93484 34208
rect 93524 34168 93525 34208
rect 93483 34159 93525 34168
rect 94059 34208 94101 34217
rect 94059 34168 94060 34208
rect 94100 34168 94101 34208
rect 94059 34159 94101 34168
rect 94347 34208 94389 34217
rect 94347 34168 94348 34208
rect 94388 34168 94389 34208
rect 94347 34159 94389 34168
rect 94827 34208 94869 34217
rect 94827 34168 94828 34208
rect 94868 34168 94869 34208
rect 94827 34159 94869 34168
rect 95211 34208 95253 34217
rect 95211 34168 95212 34208
rect 95252 34168 95253 34208
rect 95211 34159 95253 34168
rect 95499 34208 95541 34217
rect 95499 34168 95500 34208
rect 95540 34168 95541 34208
rect 95499 34159 95541 34168
rect 97227 34208 97269 34217
rect 97227 34168 97228 34208
rect 97268 34168 97269 34208
rect 97227 34159 97269 34168
rect 97707 34208 97749 34217
rect 97707 34168 97708 34208
rect 97748 34168 97749 34208
rect 97707 34159 97749 34168
rect 97995 34208 98037 34217
rect 97995 34168 97996 34208
rect 98036 34168 98037 34208
rect 97995 34159 98037 34168
rect 98187 34208 98229 34217
rect 98187 34168 98188 34208
rect 98228 34168 98229 34208
rect 98187 34159 98229 34168
rect 98475 34208 98517 34217
rect 98475 34168 98476 34208
rect 98516 34168 98517 34208
rect 98475 34159 98517 34168
rect 98955 34208 98997 34217
rect 98955 34168 98956 34208
rect 98996 34168 98997 34208
rect 98955 34159 98997 34168
rect 99243 34208 99285 34217
rect 99243 34168 99244 34208
rect 99284 34168 99285 34208
rect 99243 34159 99285 34168
rect 576 34040 99360 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 8352 34040
rect 8392 34000 8434 34040
rect 8474 34000 8516 34040
rect 8556 34000 8598 34040
rect 8638 34000 8680 34040
rect 8720 34000 12352 34040
rect 12392 34000 12434 34040
rect 12474 34000 12516 34040
rect 12556 34000 12598 34040
rect 12638 34000 12680 34040
rect 12720 34000 16352 34040
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16720 34000 20352 34040
rect 20392 34000 20434 34040
rect 20474 34000 20516 34040
rect 20556 34000 20598 34040
rect 20638 34000 20680 34040
rect 20720 34000 24352 34040
rect 24392 34000 24434 34040
rect 24474 34000 24516 34040
rect 24556 34000 24598 34040
rect 24638 34000 24680 34040
rect 24720 34000 28352 34040
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28720 34000 32352 34040
rect 32392 34000 32434 34040
rect 32474 34000 32516 34040
rect 32556 34000 32598 34040
rect 32638 34000 32680 34040
rect 32720 34000 36352 34040
rect 36392 34000 36434 34040
rect 36474 34000 36516 34040
rect 36556 34000 36598 34040
rect 36638 34000 36680 34040
rect 36720 34000 40352 34040
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40720 34000 44352 34040
rect 44392 34000 44434 34040
rect 44474 34000 44516 34040
rect 44556 34000 44598 34040
rect 44638 34000 44680 34040
rect 44720 34000 48352 34040
rect 48392 34000 48434 34040
rect 48474 34000 48516 34040
rect 48556 34000 48598 34040
rect 48638 34000 48680 34040
rect 48720 34000 52352 34040
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52720 34000 56352 34040
rect 56392 34000 56434 34040
rect 56474 34000 56516 34040
rect 56556 34000 56598 34040
rect 56638 34000 56680 34040
rect 56720 34000 60352 34040
rect 60392 34000 60434 34040
rect 60474 34000 60516 34040
rect 60556 34000 60598 34040
rect 60638 34000 60680 34040
rect 60720 34000 64352 34040
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64720 34000 68352 34040
rect 68392 34000 68434 34040
rect 68474 34000 68516 34040
rect 68556 34000 68598 34040
rect 68638 34000 68680 34040
rect 68720 34000 72352 34040
rect 72392 34000 72434 34040
rect 72474 34000 72516 34040
rect 72556 34000 72598 34040
rect 72638 34000 72680 34040
rect 72720 34000 76352 34040
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76720 34000 80352 34040
rect 80392 34000 80434 34040
rect 80474 34000 80516 34040
rect 80556 34000 80598 34040
rect 80638 34000 80680 34040
rect 80720 34000 84352 34040
rect 84392 34000 84434 34040
rect 84474 34000 84516 34040
rect 84556 34000 84598 34040
rect 84638 34000 84680 34040
rect 84720 34000 88352 34040
rect 88392 34000 88434 34040
rect 88474 34000 88516 34040
rect 88556 34000 88598 34040
rect 88638 34000 88680 34040
rect 88720 34000 92352 34040
rect 92392 34000 92434 34040
rect 92474 34000 92516 34040
rect 92556 34000 92598 34040
rect 92638 34000 92680 34040
rect 92720 34000 96352 34040
rect 96392 34000 96434 34040
rect 96474 34000 96516 34040
rect 96556 34000 96598 34040
rect 96638 34000 96680 34040
rect 96720 34000 99360 34040
rect 576 33976 99360 34000
rect 576 33284 69984 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 7112 33284
rect 7152 33244 7194 33284
rect 7234 33244 7276 33284
rect 7316 33244 7358 33284
rect 7398 33244 7440 33284
rect 7480 33244 11112 33284
rect 11152 33244 11194 33284
rect 11234 33244 11276 33284
rect 11316 33244 11358 33284
rect 11398 33244 11440 33284
rect 11480 33244 15112 33284
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15480 33244 19112 33284
rect 19152 33244 19194 33284
rect 19234 33244 19276 33284
rect 19316 33244 19358 33284
rect 19398 33244 19440 33284
rect 19480 33244 23112 33284
rect 23152 33244 23194 33284
rect 23234 33244 23276 33284
rect 23316 33244 23358 33284
rect 23398 33244 23440 33284
rect 23480 33244 27112 33284
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27480 33244 31112 33284
rect 31152 33244 31194 33284
rect 31234 33244 31276 33284
rect 31316 33244 31358 33284
rect 31398 33244 31440 33284
rect 31480 33244 35112 33284
rect 35152 33244 35194 33284
rect 35234 33244 35276 33284
rect 35316 33244 35358 33284
rect 35398 33244 35440 33284
rect 35480 33244 39112 33284
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39480 33244 43112 33284
rect 43152 33244 43194 33284
rect 43234 33244 43276 33284
rect 43316 33244 43358 33284
rect 43398 33244 43440 33284
rect 43480 33244 47112 33284
rect 47152 33244 47194 33284
rect 47234 33244 47276 33284
rect 47316 33244 47358 33284
rect 47398 33244 47440 33284
rect 47480 33244 51112 33284
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51480 33244 55112 33284
rect 55152 33244 55194 33284
rect 55234 33244 55276 33284
rect 55316 33244 55358 33284
rect 55398 33244 55440 33284
rect 55480 33244 59112 33284
rect 59152 33244 59194 33284
rect 59234 33244 59276 33284
rect 59316 33244 59358 33284
rect 59398 33244 59440 33284
rect 59480 33244 63112 33284
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63480 33244 67112 33284
rect 67152 33244 67194 33284
rect 67234 33244 67276 33284
rect 67316 33244 67358 33284
rect 67398 33244 67440 33284
rect 67480 33244 69984 33284
rect 576 33220 69984 33244
rect 576 32528 69984 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 8352 32528
rect 8392 32488 8434 32528
rect 8474 32488 8516 32528
rect 8556 32488 8598 32528
rect 8638 32488 8680 32528
rect 8720 32488 12352 32528
rect 12392 32488 12434 32528
rect 12474 32488 12516 32528
rect 12556 32488 12598 32528
rect 12638 32488 12680 32528
rect 12720 32488 16352 32528
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16720 32488 20352 32528
rect 20392 32488 20434 32528
rect 20474 32488 20516 32528
rect 20556 32488 20598 32528
rect 20638 32488 20680 32528
rect 20720 32488 24352 32528
rect 24392 32488 24434 32528
rect 24474 32488 24516 32528
rect 24556 32488 24598 32528
rect 24638 32488 24680 32528
rect 24720 32488 28352 32528
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28720 32488 32352 32528
rect 32392 32488 32434 32528
rect 32474 32488 32516 32528
rect 32556 32488 32598 32528
rect 32638 32488 32680 32528
rect 32720 32488 36352 32528
rect 36392 32488 36434 32528
rect 36474 32488 36516 32528
rect 36556 32488 36598 32528
rect 36638 32488 36680 32528
rect 36720 32488 40352 32528
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40720 32488 44352 32528
rect 44392 32488 44434 32528
rect 44474 32488 44516 32528
rect 44556 32488 44598 32528
rect 44638 32488 44680 32528
rect 44720 32488 48352 32528
rect 48392 32488 48434 32528
rect 48474 32488 48516 32528
rect 48556 32488 48598 32528
rect 48638 32488 48680 32528
rect 48720 32488 52352 32528
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52720 32488 56352 32528
rect 56392 32488 56434 32528
rect 56474 32488 56516 32528
rect 56556 32488 56598 32528
rect 56638 32488 56680 32528
rect 56720 32488 60352 32528
rect 60392 32488 60434 32528
rect 60474 32488 60516 32528
rect 60556 32488 60598 32528
rect 60638 32488 60680 32528
rect 60720 32488 64352 32528
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64720 32488 68352 32528
rect 68392 32488 68434 32528
rect 68474 32488 68516 32528
rect 68556 32488 68598 32528
rect 68638 32488 68680 32528
rect 68720 32488 69984 32528
rect 576 32464 69984 32488
rect 69763 32192 69821 32193
rect 69763 32152 69772 32192
rect 69812 32152 69821 32192
rect 69763 32151 69821 32152
rect 69867 31940 69909 31949
rect 69867 31900 69868 31940
rect 69908 31900 69909 31940
rect 69867 31891 69909 31900
rect 576 31772 69984 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 7112 31772
rect 7152 31732 7194 31772
rect 7234 31732 7276 31772
rect 7316 31732 7358 31772
rect 7398 31732 7440 31772
rect 7480 31732 11112 31772
rect 11152 31732 11194 31772
rect 11234 31732 11276 31772
rect 11316 31732 11358 31772
rect 11398 31732 11440 31772
rect 11480 31732 15112 31772
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15480 31732 19112 31772
rect 19152 31732 19194 31772
rect 19234 31732 19276 31772
rect 19316 31732 19358 31772
rect 19398 31732 19440 31772
rect 19480 31732 23112 31772
rect 23152 31732 23194 31772
rect 23234 31732 23276 31772
rect 23316 31732 23358 31772
rect 23398 31732 23440 31772
rect 23480 31732 27112 31772
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27480 31732 31112 31772
rect 31152 31732 31194 31772
rect 31234 31732 31276 31772
rect 31316 31732 31358 31772
rect 31398 31732 31440 31772
rect 31480 31732 35112 31772
rect 35152 31732 35194 31772
rect 35234 31732 35276 31772
rect 35316 31732 35358 31772
rect 35398 31732 35440 31772
rect 35480 31732 39112 31772
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39480 31732 43112 31772
rect 43152 31732 43194 31772
rect 43234 31732 43276 31772
rect 43316 31732 43358 31772
rect 43398 31732 43440 31772
rect 43480 31732 47112 31772
rect 47152 31732 47194 31772
rect 47234 31732 47276 31772
rect 47316 31732 47358 31772
rect 47398 31732 47440 31772
rect 47480 31732 51112 31772
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51480 31732 55112 31772
rect 55152 31732 55194 31772
rect 55234 31732 55276 31772
rect 55316 31732 55358 31772
rect 55398 31732 55440 31772
rect 55480 31732 59112 31772
rect 59152 31732 59194 31772
rect 59234 31732 59276 31772
rect 59316 31732 59358 31772
rect 59398 31732 59440 31772
rect 59480 31732 63112 31772
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63480 31732 67112 31772
rect 67152 31732 67194 31772
rect 67234 31732 67276 31772
rect 67316 31732 67358 31772
rect 67398 31732 67440 31772
rect 67480 31732 69984 31772
rect 576 31708 69984 31732
rect 68811 31604 68853 31613
rect 68811 31564 68812 31604
rect 68852 31564 68853 31604
rect 68811 31555 68853 31564
rect 69867 31604 69909 31613
rect 69867 31564 69868 31604
rect 69908 31564 69909 31604
rect 69867 31555 69909 31564
rect 67179 31520 67221 31529
rect 67179 31480 67180 31520
rect 67220 31480 67221 31520
rect 67179 31471 67221 31480
rect 69195 31520 69237 31529
rect 69195 31480 69196 31520
rect 69236 31480 69237 31520
rect 69195 31471 69237 31480
rect 69579 31520 69621 31529
rect 69579 31480 69580 31520
rect 69620 31480 69621 31520
rect 69579 31471 69621 31480
rect 68611 31436 68669 31437
rect 68611 31396 68620 31436
rect 68660 31396 68669 31436
rect 68611 31395 68669 31396
rect 68995 31436 69053 31437
rect 68995 31396 69004 31436
rect 69044 31396 69053 31436
rect 68995 31395 69053 31396
rect 69379 31436 69437 31437
rect 69379 31396 69388 31436
rect 69428 31396 69437 31436
rect 69379 31395 69437 31396
rect 67267 31352 67325 31353
rect 67267 31312 67276 31352
rect 67316 31312 67325 31352
rect 67267 31311 67325 31312
rect 67555 31352 67613 31353
rect 67555 31312 67564 31352
rect 67604 31312 67613 31352
rect 67555 31311 67613 31312
rect 67747 31352 67805 31353
rect 67747 31312 67756 31352
rect 67796 31312 67805 31352
rect 67747 31311 67805 31312
rect 69763 31352 69821 31353
rect 69763 31312 69772 31352
rect 69812 31312 69821 31352
rect 69763 31311 69821 31312
rect 576 31016 69984 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 8352 31016
rect 8392 30976 8434 31016
rect 8474 30976 8516 31016
rect 8556 30976 8598 31016
rect 8638 30976 8680 31016
rect 8720 30976 12352 31016
rect 12392 30976 12434 31016
rect 12474 30976 12516 31016
rect 12556 30976 12598 31016
rect 12638 30976 12680 31016
rect 12720 30976 16352 31016
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16720 30976 20352 31016
rect 20392 30976 20434 31016
rect 20474 30976 20516 31016
rect 20556 30976 20598 31016
rect 20638 30976 20680 31016
rect 20720 30976 24352 31016
rect 24392 30976 24434 31016
rect 24474 30976 24516 31016
rect 24556 30976 24598 31016
rect 24638 30976 24680 31016
rect 24720 30976 28352 31016
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28720 30976 32352 31016
rect 32392 30976 32434 31016
rect 32474 30976 32516 31016
rect 32556 30976 32598 31016
rect 32638 30976 32680 31016
rect 32720 30976 36352 31016
rect 36392 30976 36434 31016
rect 36474 30976 36516 31016
rect 36556 30976 36598 31016
rect 36638 30976 36680 31016
rect 36720 30976 40352 31016
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40720 30976 44352 31016
rect 44392 30976 44434 31016
rect 44474 30976 44516 31016
rect 44556 30976 44598 31016
rect 44638 30976 44680 31016
rect 44720 30976 48352 31016
rect 48392 30976 48434 31016
rect 48474 30976 48516 31016
rect 48556 30976 48598 31016
rect 48638 30976 48680 31016
rect 48720 30976 52352 31016
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52720 30976 56352 31016
rect 56392 30976 56434 31016
rect 56474 30976 56516 31016
rect 56556 30976 56598 31016
rect 56638 30976 56680 31016
rect 56720 30976 60352 31016
rect 60392 30976 60434 31016
rect 60474 30976 60516 31016
rect 60556 30976 60598 31016
rect 60638 30976 60680 31016
rect 60720 30976 64352 31016
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64720 30976 68352 31016
rect 68392 30976 68434 31016
rect 68474 30976 68516 31016
rect 68556 30976 68598 31016
rect 68638 30976 68680 31016
rect 68720 30976 69984 31016
rect 576 30952 69984 30976
rect 67563 30848 67605 30857
rect 67563 30808 67564 30848
rect 67604 30808 67605 30848
rect 67563 30799 67605 30808
rect 68619 30848 68661 30857
rect 68619 30808 68620 30848
rect 68660 30808 68661 30848
rect 68619 30799 68661 30808
rect 69099 30848 69141 30857
rect 69099 30808 69100 30848
rect 69140 30808 69141 30848
rect 69099 30799 69141 30808
rect 69387 30848 69429 30857
rect 69387 30808 69388 30848
rect 69428 30808 69429 30848
rect 69387 30799 69429 30808
rect 69675 30848 69717 30857
rect 69675 30808 69676 30848
rect 69716 30808 69717 30848
rect 69675 30799 69717 30808
rect 68515 30680 68573 30681
rect 68515 30640 68524 30680
rect 68564 30640 68573 30680
rect 68515 30639 68573 30640
rect 68995 30680 69053 30681
rect 68995 30640 69004 30680
rect 69044 30640 69053 30680
rect 68995 30639 69053 30640
rect 69283 30680 69341 30681
rect 69283 30640 69292 30680
rect 69332 30640 69341 30680
rect 69283 30639 69341 30640
rect 69571 30680 69629 30681
rect 69571 30640 69580 30680
rect 69620 30640 69629 30680
rect 69571 30639 69629 30640
rect 67363 30596 67421 30597
rect 67363 30556 67372 30596
rect 67412 30556 67421 30596
rect 67363 30555 67421 30556
rect 576 30260 69984 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 7112 30260
rect 7152 30220 7194 30260
rect 7234 30220 7276 30260
rect 7316 30220 7358 30260
rect 7398 30220 7440 30260
rect 7480 30220 11112 30260
rect 11152 30220 11194 30260
rect 11234 30220 11276 30260
rect 11316 30220 11358 30260
rect 11398 30220 11440 30260
rect 11480 30220 15112 30260
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15480 30220 19112 30260
rect 19152 30220 19194 30260
rect 19234 30220 19276 30260
rect 19316 30220 19358 30260
rect 19398 30220 19440 30260
rect 19480 30220 23112 30260
rect 23152 30220 23194 30260
rect 23234 30220 23276 30260
rect 23316 30220 23358 30260
rect 23398 30220 23440 30260
rect 23480 30220 27112 30260
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27480 30220 31112 30260
rect 31152 30220 31194 30260
rect 31234 30220 31276 30260
rect 31316 30220 31358 30260
rect 31398 30220 31440 30260
rect 31480 30220 35112 30260
rect 35152 30220 35194 30260
rect 35234 30220 35276 30260
rect 35316 30220 35358 30260
rect 35398 30220 35440 30260
rect 35480 30220 39112 30260
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39480 30220 43112 30260
rect 43152 30220 43194 30260
rect 43234 30220 43276 30260
rect 43316 30220 43358 30260
rect 43398 30220 43440 30260
rect 43480 30220 47112 30260
rect 47152 30220 47194 30260
rect 47234 30220 47276 30260
rect 47316 30220 47358 30260
rect 47398 30220 47440 30260
rect 47480 30220 51112 30260
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51480 30220 55112 30260
rect 55152 30220 55194 30260
rect 55234 30220 55276 30260
rect 55316 30220 55358 30260
rect 55398 30220 55440 30260
rect 55480 30220 59112 30260
rect 59152 30220 59194 30260
rect 59234 30220 59276 30260
rect 59316 30220 59358 30260
rect 59398 30220 59440 30260
rect 59480 30220 63112 30260
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63480 30220 67112 30260
rect 67152 30220 67194 30260
rect 67234 30220 67276 30260
rect 67316 30220 67358 30260
rect 67398 30220 67440 30260
rect 67480 30220 69984 30260
rect 576 30196 69984 30220
rect 576 29504 69984 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 8352 29504
rect 8392 29464 8434 29504
rect 8474 29464 8516 29504
rect 8556 29464 8598 29504
rect 8638 29464 8680 29504
rect 8720 29464 12352 29504
rect 12392 29464 12434 29504
rect 12474 29464 12516 29504
rect 12556 29464 12598 29504
rect 12638 29464 12680 29504
rect 12720 29464 16352 29504
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16720 29464 20352 29504
rect 20392 29464 20434 29504
rect 20474 29464 20516 29504
rect 20556 29464 20598 29504
rect 20638 29464 20680 29504
rect 20720 29464 24352 29504
rect 24392 29464 24434 29504
rect 24474 29464 24516 29504
rect 24556 29464 24598 29504
rect 24638 29464 24680 29504
rect 24720 29464 28352 29504
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28720 29464 32352 29504
rect 32392 29464 32434 29504
rect 32474 29464 32516 29504
rect 32556 29464 32598 29504
rect 32638 29464 32680 29504
rect 32720 29464 36352 29504
rect 36392 29464 36434 29504
rect 36474 29464 36516 29504
rect 36556 29464 36598 29504
rect 36638 29464 36680 29504
rect 36720 29464 40352 29504
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40720 29464 44352 29504
rect 44392 29464 44434 29504
rect 44474 29464 44516 29504
rect 44556 29464 44598 29504
rect 44638 29464 44680 29504
rect 44720 29464 48352 29504
rect 48392 29464 48434 29504
rect 48474 29464 48516 29504
rect 48556 29464 48598 29504
rect 48638 29464 48680 29504
rect 48720 29464 52352 29504
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52720 29464 56352 29504
rect 56392 29464 56434 29504
rect 56474 29464 56516 29504
rect 56556 29464 56598 29504
rect 56638 29464 56680 29504
rect 56720 29464 60352 29504
rect 60392 29464 60434 29504
rect 60474 29464 60516 29504
rect 60556 29464 60598 29504
rect 60638 29464 60680 29504
rect 60720 29464 64352 29504
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64720 29464 68352 29504
rect 68392 29464 68434 29504
rect 68474 29464 68516 29504
rect 68556 29464 68598 29504
rect 68638 29464 68680 29504
rect 68720 29464 69984 29504
rect 576 29440 69984 29464
rect 576 28748 69984 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 7112 28748
rect 7152 28708 7194 28748
rect 7234 28708 7276 28748
rect 7316 28708 7358 28748
rect 7398 28708 7440 28748
rect 7480 28708 11112 28748
rect 11152 28708 11194 28748
rect 11234 28708 11276 28748
rect 11316 28708 11358 28748
rect 11398 28708 11440 28748
rect 11480 28708 15112 28748
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15480 28708 19112 28748
rect 19152 28708 19194 28748
rect 19234 28708 19276 28748
rect 19316 28708 19358 28748
rect 19398 28708 19440 28748
rect 19480 28708 23112 28748
rect 23152 28708 23194 28748
rect 23234 28708 23276 28748
rect 23316 28708 23358 28748
rect 23398 28708 23440 28748
rect 23480 28708 27112 28748
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27480 28708 31112 28748
rect 31152 28708 31194 28748
rect 31234 28708 31276 28748
rect 31316 28708 31358 28748
rect 31398 28708 31440 28748
rect 31480 28708 35112 28748
rect 35152 28708 35194 28748
rect 35234 28708 35276 28748
rect 35316 28708 35358 28748
rect 35398 28708 35440 28748
rect 35480 28708 39112 28748
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39480 28708 43112 28748
rect 43152 28708 43194 28748
rect 43234 28708 43276 28748
rect 43316 28708 43358 28748
rect 43398 28708 43440 28748
rect 43480 28708 47112 28748
rect 47152 28708 47194 28748
rect 47234 28708 47276 28748
rect 47316 28708 47358 28748
rect 47398 28708 47440 28748
rect 47480 28708 51112 28748
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51480 28708 55112 28748
rect 55152 28708 55194 28748
rect 55234 28708 55276 28748
rect 55316 28708 55358 28748
rect 55398 28708 55440 28748
rect 55480 28708 59112 28748
rect 59152 28708 59194 28748
rect 59234 28708 59276 28748
rect 59316 28708 59358 28748
rect 59398 28708 59440 28748
rect 59480 28708 63112 28748
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63480 28708 67112 28748
rect 67152 28708 67194 28748
rect 67234 28708 67276 28748
rect 67316 28708 67358 28748
rect 67398 28708 67440 28748
rect 67480 28708 69984 28748
rect 576 28684 69984 28708
rect 576 27992 69984 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 8352 27992
rect 8392 27952 8434 27992
rect 8474 27952 8516 27992
rect 8556 27952 8598 27992
rect 8638 27952 8680 27992
rect 8720 27952 12352 27992
rect 12392 27952 12434 27992
rect 12474 27952 12516 27992
rect 12556 27952 12598 27992
rect 12638 27952 12680 27992
rect 12720 27952 16352 27992
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16720 27952 20352 27992
rect 20392 27952 20434 27992
rect 20474 27952 20516 27992
rect 20556 27952 20598 27992
rect 20638 27952 20680 27992
rect 20720 27952 24352 27992
rect 24392 27952 24434 27992
rect 24474 27952 24516 27992
rect 24556 27952 24598 27992
rect 24638 27952 24680 27992
rect 24720 27952 28352 27992
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28720 27952 32352 27992
rect 32392 27952 32434 27992
rect 32474 27952 32516 27992
rect 32556 27952 32598 27992
rect 32638 27952 32680 27992
rect 32720 27952 36352 27992
rect 36392 27952 36434 27992
rect 36474 27952 36516 27992
rect 36556 27952 36598 27992
rect 36638 27952 36680 27992
rect 36720 27952 40352 27992
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40720 27952 44352 27992
rect 44392 27952 44434 27992
rect 44474 27952 44516 27992
rect 44556 27952 44598 27992
rect 44638 27952 44680 27992
rect 44720 27952 48352 27992
rect 48392 27952 48434 27992
rect 48474 27952 48516 27992
rect 48556 27952 48598 27992
rect 48638 27952 48680 27992
rect 48720 27952 52352 27992
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52720 27952 56352 27992
rect 56392 27952 56434 27992
rect 56474 27952 56516 27992
rect 56556 27952 56598 27992
rect 56638 27952 56680 27992
rect 56720 27952 60352 27992
rect 60392 27952 60434 27992
rect 60474 27952 60516 27992
rect 60556 27952 60598 27992
rect 60638 27952 60680 27992
rect 60720 27952 64352 27992
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64720 27952 68352 27992
rect 68392 27952 68434 27992
rect 68474 27952 68516 27992
rect 68556 27952 68598 27992
rect 68638 27952 68680 27992
rect 68720 27952 69984 27992
rect 576 27928 69984 27952
rect 68803 27572 68861 27573
rect 68803 27532 68812 27572
rect 68852 27532 68861 27572
rect 68803 27531 68861 27532
rect 69003 27404 69045 27413
rect 69003 27364 69004 27404
rect 69044 27364 69045 27404
rect 69003 27355 69045 27364
rect 576 27236 69984 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 7112 27236
rect 7152 27196 7194 27236
rect 7234 27196 7276 27236
rect 7316 27196 7358 27236
rect 7398 27196 7440 27236
rect 7480 27196 11112 27236
rect 11152 27196 11194 27236
rect 11234 27196 11276 27236
rect 11316 27196 11358 27236
rect 11398 27196 11440 27236
rect 11480 27196 15112 27236
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15480 27196 19112 27236
rect 19152 27196 19194 27236
rect 19234 27196 19276 27236
rect 19316 27196 19358 27236
rect 19398 27196 19440 27236
rect 19480 27196 23112 27236
rect 23152 27196 23194 27236
rect 23234 27196 23276 27236
rect 23316 27196 23358 27236
rect 23398 27196 23440 27236
rect 23480 27196 27112 27236
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27480 27196 31112 27236
rect 31152 27196 31194 27236
rect 31234 27196 31276 27236
rect 31316 27196 31358 27236
rect 31398 27196 31440 27236
rect 31480 27196 35112 27236
rect 35152 27196 35194 27236
rect 35234 27196 35276 27236
rect 35316 27196 35358 27236
rect 35398 27196 35440 27236
rect 35480 27196 39112 27236
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39480 27196 43112 27236
rect 43152 27196 43194 27236
rect 43234 27196 43276 27236
rect 43316 27196 43358 27236
rect 43398 27196 43440 27236
rect 43480 27196 47112 27236
rect 47152 27196 47194 27236
rect 47234 27196 47276 27236
rect 47316 27196 47358 27236
rect 47398 27196 47440 27236
rect 47480 27196 51112 27236
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51480 27196 55112 27236
rect 55152 27196 55194 27236
rect 55234 27196 55276 27236
rect 55316 27196 55358 27236
rect 55398 27196 55440 27236
rect 55480 27196 59112 27236
rect 59152 27196 59194 27236
rect 59234 27196 59276 27236
rect 59316 27196 59358 27236
rect 59398 27196 59440 27236
rect 59480 27196 63112 27236
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63480 27196 67112 27236
rect 67152 27196 67194 27236
rect 67234 27196 67276 27236
rect 67316 27196 67358 27236
rect 67398 27196 67440 27236
rect 67480 27196 69984 27236
rect 576 27172 69984 27196
rect 68139 26984 68181 26993
rect 68139 26944 68140 26984
rect 68180 26944 68181 26984
rect 68139 26935 68181 26944
rect 67939 26900 67997 26901
rect 67939 26860 67948 26900
rect 67988 26860 67997 26900
rect 67939 26859 67997 26860
rect 68323 26900 68381 26901
rect 68323 26860 68332 26900
rect 68372 26860 68381 26900
rect 68323 26859 68381 26860
rect 69475 26900 69533 26901
rect 69475 26860 69484 26900
rect 69524 26860 69533 26900
rect 69475 26859 69533 26860
rect 67755 26648 67797 26657
rect 67755 26608 67756 26648
rect 67796 26608 67797 26648
rect 67755 26599 67797 26608
rect 69675 26648 69717 26657
rect 69675 26608 69676 26648
rect 69716 26608 69717 26648
rect 69675 26599 69717 26608
rect 576 26480 69984 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 8352 26480
rect 8392 26440 8434 26480
rect 8474 26440 8516 26480
rect 8556 26440 8598 26480
rect 8638 26440 8680 26480
rect 8720 26440 12352 26480
rect 12392 26440 12434 26480
rect 12474 26440 12516 26480
rect 12556 26440 12598 26480
rect 12638 26440 12680 26480
rect 12720 26440 16352 26480
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16720 26440 20352 26480
rect 20392 26440 20434 26480
rect 20474 26440 20516 26480
rect 20556 26440 20598 26480
rect 20638 26440 20680 26480
rect 20720 26440 24352 26480
rect 24392 26440 24434 26480
rect 24474 26440 24516 26480
rect 24556 26440 24598 26480
rect 24638 26440 24680 26480
rect 24720 26440 28352 26480
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28720 26440 32352 26480
rect 32392 26440 32434 26480
rect 32474 26440 32516 26480
rect 32556 26440 32598 26480
rect 32638 26440 32680 26480
rect 32720 26440 36352 26480
rect 36392 26440 36434 26480
rect 36474 26440 36516 26480
rect 36556 26440 36598 26480
rect 36638 26440 36680 26480
rect 36720 26440 40352 26480
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40720 26440 44352 26480
rect 44392 26440 44434 26480
rect 44474 26440 44516 26480
rect 44556 26440 44598 26480
rect 44638 26440 44680 26480
rect 44720 26440 48352 26480
rect 48392 26440 48434 26480
rect 48474 26440 48516 26480
rect 48556 26440 48598 26480
rect 48638 26440 48680 26480
rect 48720 26440 52352 26480
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52720 26440 56352 26480
rect 56392 26440 56434 26480
rect 56474 26440 56516 26480
rect 56556 26440 56598 26480
rect 56638 26440 56680 26480
rect 56720 26440 60352 26480
rect 60392 26440 60434 26480
rect 60474 26440 60516 26480
rect 60556 26440 60598 26480
rect 60638 26440 60680 26480
rect 60720 26440 64352 26480
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64720 26440 68352 26480
rect 68392 26440 68434 26480
rect 68474 26440 68516 26480
rect 68556 26440 68598 26480
rect 68638 26440 68680 26480
rect 68720 26440 69984 26480
rect 576 26416 69984 26440
rect 67555 26144 67613 26145
rect 67555 26104 67564 26144
rect 67604 26104 67613 26144
rect 67555 26103 67613 26104
rect 68611 26144 68669 26145
rect 68611 26104 68620 26144
rect 68660 26104 68669 26144
rect 68611 26103 68669 26104
rect 68803 26144 68861 26145
rect 68803 26104 68812 26144
rect 68852 26104 68861 26144
rect 68803 26103 68861 26104
rect 69091 26144 69149 26145
rect 69091 26104 69100 26144
rect 69140 26104 69149 26144
rect 69091 26103 69149 26104
rect 69763 26144 69821 26145
rect 69763 26104 69772 26144
rect 69812 26104 69821 26144
rect 69763 26103 69821 26104
rect 67747 26060 67805 26061
rect 67747 26020 67756 26060
rect 67796 26020 67805 26060
rect 67747 26019 67805 26020
rect 69379 26060 69437 26061
rect 69379 26020 69388 26060
rect 69428 26020 69437 26060
rect 69379 26019 69437 26020
rect 67467 25892 67509 25901
rect 67467 25852 67468 25892
rect 67508 25852 67509 25892
rect 67467 25843 67509 25852
rect 67947 25892 67989 25901
rect 67947 25852 67948 25892
rect 67988 25852 67989 25892
rect 67947 25843 67989 25852
rect 68523 25892 68565 25901
rect 68523 25852 68524 25892
rect 68564 25852 68565 25892
rect 68523 25843 68565 25852
rect 68907 25892 68949 25901
rect 68907 25852 68908 25892
rect 68948 25852 68949 25892
rect 68907 25843 68949 25852
rect 69195 25892 69237 25901
rect 69195 25852 69196 25892
rect 69236 25852 69237 25892
rect 69195 25843 69237 25852
rect 69579 25892 69621 25901
rect 69579 25852 69580 25892
rect 69620 25852 69621 25892
rect 69579 25843 69621 25852
rect 69867 25892 69909 25901
rect 69867 25852 69868 25892
rect 69908 25852 69909 25892
rect 69867 25843 69909 25852
rect 576 25724 69984 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 7112 25724
rect 7152 25684 7194 25724
rect 7234 25684 7276 25724
rect 7316 25684 7358 25724
rect 7398 25684 7440 25724
rect 7480 25684 11112 25724
rect 11152 25684 11194 25724
rect 11234 25684 11276 25724
rect 11316 25684 11358 25724
rect 11398 25684 11440 25724
rect 11480 25684 15112 25724
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15480 25684 19112 25724
rect 19152 25684 19194 25724
rect 19234 25684 19276 25724
rect 19316 25684 19358 25724
rect 19398 25684 19440 25724
rect 19480 25684 23112 25724
rect 23152 25684 23194 25724
rect 23234 25684 23276 25724
rect 23316 25684 23358 25724
rect 23398 25684 23440 25724
rect 23480 25684 27112 25724
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27480 25684 31112 25724
rect 31152 25684 31194 25724
rect 31234 25684 31276 25724
rect 31316 25684 31358 25724
rect 31398 25684 31440 25724
rect 31480 25684 35112 25724
rect 35152 25684 35194 25724
rect 35234 25684 35276 25724
rect 35316 25684 35358 25724
rect 35398 25684 35440 25724
rect 35480 25684 39112 25724
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39480 25684 43112 25724
rect 43152 25684 43194 25724
rect 43234 25684 43276 25724
rect 43316 25684 43358 25724
rect 43398 25684 43440 25724
rect 43480 25684 47112 25724
rect 47152 25684 47194 25724
rect 47234 25684 47276 25724
rect 47316 25684 47358 25724
rect 47398 25684 47440 25724
rect 47480 25684 51112 25724
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51480 25684 55112 25724
rect 55152 25684 55194 25724
rect 55234 25684 55276 25724
rect 55316 25684 55358 25724
rect 55398 25684 55440 25724
rect 55480 25684 59112 25724
rect 59152 25684 59194 25724
rect 59234 25684 59276 25724
rect 59316 25684 59358 25724
rect 59398 25684 59440 25724
rect 59480 25684 63112 25724
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63480 25684 67112 25724
rect 67152 25684 67194 25724
rect 67234 25684 67276 25724
rect 67316 25684 67358 25724
rect 67398 25684 67440 25724
rect 67480 25684 69984 25724
rect 576 25660 69984 25684
rect 68811 25556 68853 25565
rect 68811 25516 68812 25556
rect 68852 25516 68853 25556
rect 68811 25507 68853 25516
rect 69867 25556 69909 25565
rect 69867 25516 69868 25556
rect 69908 25516 69909 25556
rect 69867 25507 69909 25516
rect 68611 25388 68669 25389
rect 68611 25348 68620 25388
rect 68660 25348 68669 25388
rect 68611 25347 68669 25348
rect 69667 25388 69725 25389
rect 69667 25348 69676 25388
rect 69716 25348 69725 25388
rect 69667 25347 69725 25348
rect 643 25304 701 25305
rect 643 25264 652 25304
rect 692 25264 701 25304
rect 643 25263 701 25264
rect 835 25304 893 25305
rect 835 25264 844 25304
rect 884 25264 893 25304
rect 835 25263 893 25264
rect 69283 25304 69341 25305
rect 69283 25264 69292 25304
rect 69332 25264 69341 25304
rect 69283 25263 69341 25264
rect 69475 25304 69533 25305
rect 69475 25264 69484 25304
rect 69524 25264 69533 25304
rect 69475 25263 69533 25264
rect 576 24968 69984 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 8352 24968
rect 8392 24928 8434 24968
rect 8474 24928 8516 24968
rect 8556 24928 8598 24968
rect 8638 24928 8680 24968
rect 8720 24928 12352 24968
rect 12392 24928 12434 24968
rect 12474 24928 12516 24968
rect 12556 24928 12598 24968
rect 12638 24928 12680 24968
rect 12720 24928 16352 24968
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16720 24928 20352 24968
rect 20392 24928 20434 24968
rect 20474 24928 20516 24968
rect 20556 24928 20598 24968
rect 20638 24928 20680 24968
rect 20720 24928 24352 24968
rect 24392 24928 24434 24968
rect 24474 24928 24516 24968
rect 24556 24928 24598 24968
rect 24638 24928 24680 24968
rect 24720 24928 28352 24968
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28720 24928 32352 24968
rect 32392 24928 32434 24968
rect 32474 24928 32516 24968
rect 32556 24928 32598 24968
rect 32638 24928 32680 24968
rect 32720 24928 36352 24968
rect 36392 24928 36434 24968
rect 36474 24928 36516 24968
rect 36556 24928 36598 24968
rect 36638 24928 36680 24968
rect 36720 24928 40352 24968
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40720 24928 44352 24968
rect 44392 24928 44434 24968
rect 44474 24928 44516 24968
rect 44556 24928 44598 24968
rect 44638 24928 44680 24968
rect 44720 24928 48352 24968
rect 48392 24928 48434 24968
rect 48474 24928 48516 24968
rect 48556 24928 48598 24968
rect 48638 24928 48680 24968
rect 48720 24928 52352 24968
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52720 24928 56352 24968
rect 56392 24928 56434 24968
rect 56474 24928 56516 24968
rect 56556 24928 56598 24968
rect 56638 24928 56680 24968
rect 56720 24928 60352 24968
rect 60392 24928 60434 24968
rect 60474 24928 60516 24968
rect 60556 24928 60598 24968
rect 60638 24928 60680 24968
rect 60720 24928 64352 24968
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64720 24928 68352 24968
rect 68392 24928 68434 24968
rect 68474 24928 68516 24968
rect 68556 24928 68598 24968
rect 68638 24928 68680 24968
rect 68720 24928 69984 24968
rect 576 24904 69984 24928
rect 643 24632 701 24633
rect 643 24592 652 24632
rect 692 24592 701 24632
rect 643 24591 701 24592
rect 835 24632 893 24633
rect 835 24592 844 24632
rect 884 24592 893 24632
rect 835 24591 893 24592
rect 576 24212 69984 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 7112 24212
rect 7152 24172 7194 24212
rect 7234 24172 7276 24212
rect 7316 24172 7358 24212
rect 7398 24172 7440 24212
rect 7480 24172 11112 24212
rect 11152 24172 11194 24212
rect 11234 24172 11276 24212
rect 11316 24172 11358 24212
rect 11398 24172 11440 24212
rect 11480 24172 15112 24212
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15480 24172 19112 24212
rect 19152 24172 19194 24212
rect 19234 24172 19276 24212
rect 19316 24172 19358 24212
rect 19398 24172 19440 24212
rect 19480 24172 23112 24212
rect 23152 24172 23194 24212
rect 23234 24172 23276 24212
rect 23316 24172 23358 24212
rect 23398 24172 23440 24212
rect 23480 24172 27112 24212
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27480 24172 31112 24212
rect 31152 24172 31194 24212
rect 31234 24172 31276 24212
rect 31316 24172 31358 24212
rect 31398 24172 31440 24212
rect 31480 24172 35112 24212
rect 35152 24172 35194 24212
rect 35234 24172 35276 24212
rect 35316 24172 35358 24212
rect 35398 24172 35440 24212
rect 35480 24172 39112 24212
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39480 24172 43112 24212
rect 43152 24172 43194 24212
rect 43234 24172 43276 24212
rect 43316 24172 43358 24212
rect 43398 24172 43440 24212
rect 43480 24172 47112 24212
rect 47152 24172 47194 24212
rect 47234 24172 47276 24212
rect 47316 24172 47358 24212
rect 47398 24172 47440 24212
rect 47480 24172 51112 24212
rect 51152 24172 51194 24212
rect 51234 24172 51276 24212
rect 51316 24172 51358 24212
rect 51398 24172 51440 24212
rect 51480 24172 55112 24212
rect 55152 24172 55194 24212
rect 55234 24172 55276 24212
rect 55316 24172 55358 24212
rect 55398 24172 55440 24212
rect 55480 24172 59112 24212
rect 59152 24172 59194 24212
rect 59234 24172 59276 24212
rect 59316 24172 59358 24212
rect 59398 24172 59440 24212
rect 59480 24172 63112 24212
rect 63152 24172 63194 24212
rect 63234 24172 63276 24212
rect 63316 24172 63358 24212
rect 63398 24172 63440 24212
rect 63480 24172 67112 24212
rect 67152 24172 67194 24212
rect 67234 24172 67276 24212
rect 67316 24172 67358 24212
rect 67398 24172 67440 24212
rect 67480 24172 69984 24212
rect 576 24148 69984 24172
rect 643 23792 701 23793
rect 643 23752 652 23792
rect 692 23752 701 23792
rect 643 23751 701 23752
rect 835 23792 893 23793
rect 835 23752 844 23792
rect 884 23752 893 23792
rect 835 23751 893 23752
rect 576 23456 99360 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 8352 23456
rect 8392 23416 8434 23456
rect 8474 23416 8516 23456
rect 8556 23416 8598 23456
rect 8638 23416 8680 23456
rect 8720 23416 12352 23456
rect 12392 23416 12434 23456
rect 12474 23416 12516 23456
rect 12556 23416 12598 23456
rect 12638 23416 12680 23456
rect 12720 23416 16352 23456
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16720 23416 20352 23456
rect 20392 23416 20434 23456
rect 20474 23416 20516 23456
rect 20556 23416 20598 23456
rect 20638 23416 20680 23456
rect 20720 23416 24352 23456
rect 24392 23416 24434 23456
rect 24474 23416 24516 23456
rect 24556 23416 24598 23456
rect 24638 23416 24680 23456
rect 24720 23416 28352 23456
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28720 23416 32352 23456
rect 32392 23416 32434 23456
rect 32474 23416 32516 23456
rect 32556 23416 32598 23456
rect 32638 23416 32680 23456
rect 32720 23416 36352 23456
rect 36392 23416 36434 23456
rect 36474 23416 36516 23456
rect 36556 23416 36598 23456
rect 36638 23416 36680 23456
rect 36720 23416 40352 23456
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40720 23416 44352 23456
rect 44392 23416 44434 23456
rect 44474 23416 44516 23456
rect 44556 23416 44598 23456
rect 44638 23416 44680 23456
rect 44720 23416 48352 23456
rect 48392 23416 48434 23456
rect 48474 23416 48516 23456
rect 48556 23416 48598 23456
rect 48638 23416 48680 23456
rect 48720 23416 52352 23456
rect 52392 23416 52434 23456
rect 52474 23416 52516 23456
rect 52556 23416 52598 23456
rect 52638 23416 52680 23456
rect 52720 23416 56352 23456
rect 56392 23416 56434 23456
rect 56474 23416 56516 23456
rect 56556 23416 56598 23456
rect 56638 23416 56680 23456
rect 56720 23416 60352 23456
rect 60392 23416 60434 23456
rect 60474 23416 60516 23456
rect 60556 23416 60598 23456
rect 60638 23416 60680 23456
rect 60720 23416 64352 23456
rect 64392 23416 64434 23456
rect 64474 23416 64516 23456
rect 64556 23416 64598 23456
rect 64638 23416 64680 23456
rect 64720 23416 68352 23456
rect 68392 23416 68434 23456
rect 68474 23416 68516 23456
rect 68556 23416 68598 23456
rect 68638 23416 68680 23456
rect 68720 23416 72352 23456
rect 72392 23416 72434 23456
rect 72474 23416 72516 23456
rect 72556 23416 72598 23456
rect 72638 23416 72680 23456
rect 72720 23416 76352 23456
rect 76392 23416 76434 23456
rect 76474 23416 76516 23456
rect 76556 23416 76598 23456
rect 76638 23416 76680 23456
rect 76720 23416 80352 23456
rect 80392 23416 80434 23456
rect 80474 23416 80516 23456
rect 80556 23416 80598 23456
rect 80638 23416 80680 23456
rect 80720 23416 84352 23456
rect 84392 23416 84434 23456
rect 84474 23416 84516 23456
rect 84556 23416 84598 23456
rect 84638 23416 84680 23456
rect 84720 23416 88352 23456
rect 88392 23416 88434 23456
rect 88474 23416 88516 23456
rect 88556 23416 88598 23456
rect 88638 23416 88680 23456
rect 88720 23416 92352 23456
rect 92392 23416 92434 23456
rect 92474 23416 92516 23456
rect 92556 23416 92598 23456
rect 92638 23416 92680 23456
rect 92720 23416 96352 23456
rect 96392 23416 96434 23456
rect 96474 23416 96516 23456
rect 96556 23416 96598 23456
rect 96638 23416 96680 23456
rect 96720 23416 99360 23456
rect 576 23392 99360 23416
rect 73131 23288 73173 23297
rect 73131 23248 73132 23288
rect 73172 23248 73173 23288
rect 73131 23239 73173 23248
rect 73419 23288 73461 23297
rect 73419 23248 73420 23288
rect 73460 23248 73461 23288
rect 73419 23239 73461 23248
rect 74091 23288 74133 23297
rect 74091 23248 74092 23288
rect 74132 23248 74133 23288
rect 74091 23239 74133 23248
rect 74955 23288 74997 23297
rect 74955 23248 74956 23288
rect 74996 23248 74997 23288
rect 74955 23239 74997 23248
rect 75531 23288 75573 23297
rect 75531 23248 75532 23288
rect 75572 23248 75573 23288
rect 75531 23239 75573 23248
rect 75915 23288 75957 23297
rect 75915 23248 75916 23288
rect 75956 23248 75957 23288
rect 75915 23239 75957 23248
rect 77067 23288 77109 23297
rect 77067 23248 77068 23288
rect 77108 23248 77109 23288
rect 77067 23239 77109 23248
rect 77451 23288 77493 23297
rect 77451 23248 77452 23288
rect 77492 23248 77493 23288
rect 77451 23239 77493 23248
rect 78027 23288 78069 23297
rect 78027 23248 78028 23288
rect 78068 23248 78069 23288
rect 78027 23239 78069 23248
rect 78603 23288 78645 23297
rect 78603 23248 78604 23288
rect 78644 23248 78645 23288
rect 78603 23239 78645 23248
rect 79179 23288 79221 23297
rect 79179 23248 79180 23288
rect 79220 23248 79221 23288
rect 79179 23239 79221 23248
rect 79467 23288 79509 23297
rect 79467 23248 79468 23288
rect 79508 23248 79509 23288
rect 79467 23239 79509 23248
rect 79851 23288 79893 23297
rect 79851 23248 79852 23288
rect 79892 23248 79893 23288
rect 79851 23239 79893 23248
rect 80907 23288 80949 23297
rect 80907 23248 80908 23288
rect 80948 23248 80949 23288
rect 80907 23239 80949 23248
rect 81195 23288 81237 23297
rect 81195 23248 81196 23288
rect 81236 23248 81237 23288
rect 81195 23239 81237 23248
rect 81483 23288 81525 23297
rect 81483 23248 81484 23288
rect 81524 23248 81525 23288
rect 81483 23239 81525 23248
rect 81771 23288 81813 23297
rect 81771 23248 81772 23288
rect 81812 23248 81813 23288
rect 81771 23239 81813 23248
rect 82059 23288 82101 23297
rect 82059 23248 82060 23288
rect 82100 23248 82101 23288
rect 82059 23239 82101 23248
rect 82635 23288 82677 23297
rect 82635 23248 82636 23288
rect 82676 23248 82677 23288
rect 82635 23239 82677 23248
rect 82923 23288 82965 23297
rect 82923 23248 82924 23288
rect 82964 23248 82965 23288
rect 82923 23239 82965 23248
rect 84459 23288 84501 23297
rect 84459 23248 84460 23288
rect 84500 23248 84501 23288
rect 84459 23239 84501 23248
rect 84843 23288 84885 23297
rect 84843 23248 84844 23288
rect 84884 23248 84885 23288
rect 84843 23239 84885 23248
rect 85227 23288 85269 23297
rect 85227 23248 85228 23288
rect 85268 23248 85269 23288
rect 85227 23239 85269 23248
rect 85515 23288 85557 23297
rect 85515 23248 85516 23288
rect 85556 23248 85557 23288
rect 85515 23239 85557 23248
rect 86283 23288 86325 23297
rect 86283 23248 86284 23288
rect 86324 23248 86325 23288
rect 86283 23239 86325 23248
rect 87147 23288 87189 23297
rect 87147 23248 87148 23288
rect 87188 23248 87189 23288
rect 87147 23239 87189 23248
rect 87723 23288 87765 23297
rect 87723 23248 87724 23288
rect 87764 23248 87765 23288
rect 87723 23239 87765 23248
rect 88011 23288 88053 23297
rect 88011 23248 88012 23288
rect 88052 23248 88053 23288
rect 88011 23239 88053 23248
rect 88395 23288 88437 23297
rect 88395 23248 88396 23288
rect 88436 23248 88437 23288
rect 88395 23239 88437 23248
rect 88875 23288 88917 23297
rect 88875 23248 88876 23288
rect 88916 23248 88917 23288
rect 88875 23239 88917 23248
rect 89355 23288 89397 23297
rect 89355 23248 89356 23288
rect 89396 23248 89397 23288
rect 89355 23239 89397 23248
rect 90507 23288 90549 23297
rect 90507 23248 90508 23288
rect 90548 23248 90549 23288
rect 90507 23239 90549 23248
rect 90795 23288 90837 23297
rect 90795 23248 90796 23288
rect 90836 23248 90837 23288
rect 90795 23239 90837 23248
rect 91083 23288 91125 23297
rect 91083 23248 91084 23288
rect 91124 23248 91125 23288
rect 91083 23239 91125 23248
rect 91467 23288 91509 23297
rect 91467 23248 91468 23288
rect 91508 23248 91509 23288
rect 91467 23239 91509 23248
rect 93099 23288 93141 23297
rect 93099 23248 93100 23288
rect 93140 23248 93141 23288
rect 93099 23239 93141 23248
rect 93483 23288 93525 23297
rect 93483 23248 93484 23288
rect 93524 23248 93525 23288
rect 93483 23239 93525 23248
rect 93963 23288 94005 23297
rect 93963 23248 93964 23288
rect 94004 23248 94005 23288
rect 93963 23239 94005 23248
rect 94635 23288 94677 23297
rect 94635 23248 94636 23288
rect 94676 23248 94677 23288
rect 94635 23239 94677 23248
rect 94827 23288 94869 23297
rect 94827 23248 94828 23288
rect 94868 23248 94869 23288
rect 94827 23239 94869 23248
rect 95403 23288 95445 23297
rect 95403 23248 95404 23288
rect 95444 23248 95445 23288
rect 95403 23239 95445 23248
rect 96459 23288 96501 23297
rect 96459 23248 96460 23288
rect 96500 23248 96501 23288
rect 96459 23239 96501 23248
rect 96747 23288 96789 23297
rect 96747 23248 96748 23288
rect 96788 23248 96789 23288
rect 96747 23239 96789 23248
rect 97035 23288 97077 23297
rect 97035 23248 97036 23288
rect 97076 23248 97077 23288
rect 97035 23239 97077 23248
rect 97323 23288 97365 23297
rect 97323 23248 97324 23288
rect 97364 23248 97365 23288
rect 97323 23239 97365 23248
rect 97707 23288 97749 23297
rect 97707 23248 97708 23288
rect 97748 23248 97749 23288
rect 97707 23239 97749 23248
rect 98091 23288 98133 23297
rect 98091 23248 98092 23288
rect 98132 23248 98133 23288
rect 98091 23239 98133 23248
rect 98475 23288 98517 23297
rect 98475 23248 98476 23288
rect 98516 23248 98517 23288
rect 98475 23239 98517 23248
rect 98859 23288 98901 23297
rect 98859 23248 98860 23288
rect 98900 23248 98901 23288
rect 98859 23239 98901 23248
rect 643 23120 701 23121
rect 643 23080 652 23120
rect 692 23080 701 23120
rect 643 23079 701 23080
rect 835 23120 893 23121
rect 835 23080 844 23120
rect 884 23080 893 23120
rect 835 23079 893 23080
rect 73027 23120 73085 23121
rect 73027 23080 73036 23120
rect 73076 23080 73085 23120
rect 73027 23079 73085 23080
rect 73315 23120 73373 23121
rect 73315 23080 73324 23120
rect 73364 23080 73373 23120
rect 73315 23079 73373 23080
rect 74179 23120 74237 23121
rect 74179 23080 74188 23120
rect 74228 23080 74237 23120
rect 74179 23079 74237 23080
rect 78115 23120 78173 23121
rect 78115 23080 78124 23120
rect 78164 23080 78173 23120
rect 78115 23079 78173 23080
rect 79267 23120 79325 23121
rect 79267 23080 79276 23120
rect 79316 23080 79325 23120
rect 79267 23079 79325 23080
rect 79555 23120 79613 23121
rect 79555 23080 79564 23120
rect 79604 23080 79613 23120
rect 79555 23079 79613 23080
rect 79747 23120 79805 23121
rect 79747 23080 79756 23120
rect 79796 23080 79805 23120
rect 79747 23079 79805 23080
rect 80035 23120 80093 23121
rect 80035 23080 80044 23120
rect 80084 23080 80093 23120
rect 80035 23079 80093 23080
rect 80227 23120 80285 23121
rect 80227 23080 80236 23120
rect 80276 23080 80285 23120
rect 80227 23079 80285 23080
rect 80995 23120 81053 23121
rect 80995 23080 81004 23120
rect 81044 23080 81053 23120
rect 80995 23079 81053 23080
rect 81283 23120 81341 23121
rect 81283 23080 81292 23120
rect 81332 23080 81341 23120
rect 81283 23079 81341 23080
rect 81571 23120 81629 23121
rect 81571 23080 81580 23120
rect 81620 23080 81629 23120
rect 81571 23079 81629 23080
rect 81859 23120 81917 23121
rect 81859 23080 81868 23120
rect 81908 23080 81917 23120
rect 81859 23079 81917 23080
rect 82147 23120 82205 23121
rect 82147 23080 82156 23120
rect 82196 23080 82205 23120
rect 82147 23079 82205 23080
rect 82819 23120 82877 23121
rect 82819 23080 82828 23120
rect 82868 23080 82877 23120
rect 82819 23079 82877 23080
rect 83203 23120 83261 23121
rect 83203 23080 83212 23120
rect 83252 23080 83261 23120
rect 83203 23079 83261 23080
rect 83395 23120 83453 23121
rect 83395 23080 83404 23120
rect 83444 23080 83453 23120
rect 83395 23079 83453 23080
rect 84067 23120 84125 23121
rect 84067 23080 84076 23120
rect 84116 23080 84125 23120
rect 84067 23079 84125 23080
rect 84355 23120 84413 23121
rect 84355 23080 84364 23120
rect 84404 23080 84413 23120
rect 84355 23079 84413 23080
rect 84739 23120 84797 23121
rect 84739 23080 84748 23120
rect 84788 23080 84797 23120
rect 84739 23079 84797 23080
rect 85123 23120 85181 23121
rect 85123 23080 85132 23120
rect 85172 23080 85181 23120
rect 85123 23079 85181 23080
rect 85411 23120 85469 23121
rect 85411 23080 85420 23120
rect 85460 23080 85469 23120
rect 85411 23079 85469 23080
rect 86467 23120 86525 23121
rect 86467 23080 86476 23120
rect 86516 23080 86525 23120
rect 86467 23079 86525 23080
rect 86659 23120 86717 23121
rect 86659 23080 86668 23120
rect 86708 23080 86717 23120
rect 86659 23079 86717 23080
rect 87811 23120 87869 23121
rect 87811 23080 87820 23120
rect 87860 23080 87869 23120
rect 87811 23079 87869 23080
rect 88099 23120 88157 23121
rect 88099 23080 88108 23120
rect 88148 23080 88157 23120
rect 88099 23079 88157 23080
rect 88483 23120 88541 23121
rect 88483 23080 88492 23120
rect 88532 23080 88541 23120
rect 88483 23079 88541 23080
rect 88771 23120 88829 23121
rect 88771 23080 88780 23120
rect 88820 23080 88829 23120
rect 88771 23079 88829 23080
rect 89443 23120 89501 23121
rect 89443 23080 89452 23120
rect 89492 23080 89501 23120
rect 89443 23079 89501 23080
rect 89635 23120 89693 23121
rect 89635 23080 89644 23120
rect 89684 23080 89693 23120
rect 89635 23079 89693 23080
rect 89827 23120 89885 23121
rect 89827 23080 89836 23120
rect 89876 23080 89885 23120
rect 89827 23079 89885 23080
rect 90595 23120 90653 23121
rect 90595 23080 90604 23120
rect 90644 23080 90653 23120
rect 90595 23079 90653 23080
rect 90883 23120 90941 23121
rect 90883 23080 90892 23120
rect 90932 23080 90941 23120
rect 90883 23079 90941 23080
rect 91171 23120 91229 23121
rect 91171 23080 91180 23120
rect 91220 23080 91229 23120
rect 91171 23079 91229 23080
rect 91363 23120 91421 23121
rect 91363 23080 91372 23120
rect 91412 23080 91421 23120
rect 91363 23079 91421 23080
rect 93675 23120 93717 23129
rect 93675 23080 93676 23120
rect 93716 23080 93717 23120
rect 93675 23071 93717 23080
rect 93763 23120 93821 23121
rect 93763 23080 93772 23120
rect 93812 23080 93821 23120
rect 93763 23079 93821 23080
rect 94051 23120 94109 23121
rect 94051 23080 94060 23120
rect 94100 23080 94109 23120
rect 94051 23079 94109 23080
rect 94915 23120 94973 23121
rect 94915 23080 94924 23120
rect 94964 23080 94973 23120
rect 94915 23079 94973 23080
rect 95299 23120 95357 23121
rect 95299 23080 95308 23120
rect 95348 23080 95357 23120
rect 95299 23079 95357 23080
rect 95683 23120 95741 23121
rect 95683 23080 95692 23120
rect 95732 23080 95741 23120
rect 95683 23079 95741 23080
rect 95875 23120 95933 23121
rect 95875 23080 95884 23120
rect 95924 23080 95933 23120
rect 95875 23079 95933 23080
rect 96547 23120 96605 23121
rect 96547 23080 96556 23120
rect 96596 23080 96605 23120
rect 96547 23079 96605 23080
rect 96835 23120 96893 23121
rect 96835 23080 96844 23120
rect 96884 23080 96893 23120
rect 96835 23079 96893 23080
rect 97123 23120 97181 23121
rect 97123 23080 97132 23120
rect 97172 23080 97181 23120
rect 97123 23079 97181 23080
rect 97411 23120 97469 23121
rect 97411 23080 97420 23120
rect 97460 23080 97469 23120
rect 97411 23079 97469 23080
rect 97795 23120 97853 23121
rect 97795 23080 97804 23120
rect 97844 23080 97853 23120
rect 97795 23079 97853 23080
rect 98179 23120 98237 23121
rect 98179 23080 98188 23120
rect 98228 23080 98237 23120
rect 98179 23079 98237 23080
rect 98947 23120 99005 23121
rect 98947 23080 98956 23120
rect 98996 23080 99005 23120
rect 98947 23079 99005 23080
rect 74371 23036 74429 23037
rect 74371 22996 74380 23036
rect 74420 22996 74429 23036
rect 74371 22995 74429 22996
rect 74755 23036 74813 23037
rect 74755 22996 74764 23036
rect 74804 22996 74813 23036
rect 74755 22995 74813 22996
rect 75331 23036 75389 23037
rect 75331 22996 75340 23036
rect 75380 22996 75389 23036
rect 75331 22995 75389 22996
rect 75715 23036 75773 23037
rect 75715 22996 75724 23036
rect 75764 22996 75773 23036
rect 75715 22995 75773 22996
rect 76099 23036 76157 23037
rect 76099 22996 76108 23036
rect 76148 22996 76157 23036
rect 76099 22995 76157 22996
rect 76291 23036 76349 23037
rect 76291 22996 76300 23036
rect 76340 22996 76349 23036
rect 76291 22995 76349 22996
rect 76867 23036 76925 23037
rect 76867 22996 76876 23036
rect 76916 22996 76925 23036
rect 76867 22995 76925 22996
rect 77251 23036 77309 23037
rect 77251 22996 77260 23036
rect 77300 22996 77309 23036
rect 77251 22995 77309 22996
rect 77827 23036 77885 23037
rect 77827 22996 77836 23036
rect 77876 22996 77885 23036
rect 77827 22995 77885 22996
rect 78403 23036 78461 23037
rect 78403 22996 78412 23036
rect 78452 22996 78461 23036
rect 78403 22995 78461 22996
rect 78787 23036 78845 23037
rect 78787 22996 78796 23036
rect 78836 22996 78845 23036
rect 78787 22995 78845 22996
rect 80707 23036 80765 23037
rect 80707 22996 80716 23036
rect 80756 22996 80765 23036
rect 80707 22995 80765 22996
rect 82435 23036 82493 23037
rect 82435 22996 82444 23036
rect 82484 22996 82493 23036
rect 82435 22995 82493 22996
rect 83779 23036 83837 23037
rect 83779 22996 83788 23036
rect 83828 22996 83837 23036
rect 83779 22995 83837 22996
rect 85699 23036 85757 23037
rect 85699 22996 85708 23036
rect 85748 22996 85757 23036
rect 85699 22995 85757 22996
rect 86083 23036 86141 23037
rect 86083 22996 86092 23036
rect 86132 22996 86141 23036
rect 86083 22995 86141 22996
rect 86947 23036 87005 23037
rect 86947 22996 86956 23036
rect 86996 22996 87005 23036
rect 86947 22995 87005 22996
rect 87523 23036 87581 23037
rect 87523 22996 87532 23036
rect 87572 22996 87581 23036
rect 87523 22995 87581 22996
rect 90307 23036 90365 23037
rect 90307 22996 90316 23036
rect 90356 22996 90365 23036
rect 90307 22995 90365 22996
rect 91651 23036 91709 23037
rect 91651 22996 91660 23036
rect 91700 22996 91709 23036
rect 91651 22995 91709 22996
rect 92035 23036 92093 23037
rect 92035 22996 92044 23036
rect 92084 22996 92093 23036
rect 92035 22995 92093 22996
rect 92419 23036 92477 23037
rect 92419 22996 92428 23036
rect 92468 22996 92477 23036
rect 92419 22995 92477 22996
rect 92899 23036 92957 23037
rect 92899 22996 92908 23036
rect 92948 22996 92957 23036
rect 92899 22995 92957 22996
rect 93283 23036 93341 23037
rect 93283 22996 93292 23036
rect 93332 22996 93341 23036
rect 93283 22995 93341 22996
rect 94435 23036 94493 23037
rect 94435 22996 94444 23036
rect 94484 22996 94493 23036
rect 94435 22995 94493 22996
rect 96067 23036 96125 23037
rect 96067 22996 96076 23036
rect 96116 22996 96125 23036
rect 96067 22995 96125 22996
rect 98659 23036 98717 23037
rect 98659 22996 98668 23036
rect 98708 22996 98717 23036
rect 98659 22995 98717 22996
rect 75147 22952 75189 22961
rect 75147 22912 75148 22952
rect 75188 22912 75189 22952
rect 75147 22903 75189 22912
rect 76491 22952 76533 22961
rect 76491 22912 76492 22952
rect 76532 22912 76533 22952
rect 76491 22903 76533 22912
rect 78987 22952 79029 22961
rect 78987 22912 78988 22952
rect 79028 22912 79029 22952
rect 78987 22903 79029 22912
rect 83595 22952 83637 22961
rect 83595 22912 83596 22952
rect 83636 22912 83637 22952
rect 83595 22903 83637 22912
rect 91851 22952 91893 22961
rect 91851 22912 91852 22952
rect 91892 22912 91893 22952
rect 91851 22903 91893 22912
rect 74571 22868 74613 22877
rect 74571 22828 74572 22868
rect 74612 22828 74613 22868
rect 74571 22819 74613 22828
rect 77643 22868 77685 22877
rect 77643 22828 77644 22868
rect 77684 22828 77685 22868
rect 77643 22819 77685 22828
rect 80523 22868 80565 22877
rect 80523 22828 80524 22868
rect 80564 22828 80565 22868
rect 80523 22819 80565 22828
rect 83979 22868 84021 22877
rect 83979 22828 83980 22868
rect 84020 22828 84021 22868
rect 83979 22819 84021 22828
rect 85899 22868 85941 22877
rect 85899 22828 85900 22868
rect 85940 22828 85941 22868
rect 85899 22819 85941 22828
rect 87339 22868 87381 22877
rect 87339 22828 87340 22868
rect 87380 22828 87381 22868
rect 87339 22819 87381 22828
rect 90123 22868 90165 22877
rect 90123 22828 90124 22868
rect 90164 22828 90165 22868
rect 90123 22819 90165 22828
rect 92235 22868 92277 22877
rect 92235 22828 92236 22868
rect 92276 22828 92277 22868
rect 92235 22819 92277 22828
rect 92619 22868 92661 22877
rect 92619 22828 92620 22868
rect 92660 22828 92661 22868
rect 92619 22819 92661 22828
rect 96267 22868 96309 22877
rect 96267 22828 96268 22868
rect 96308 22828 96309 22868
rect 96267 22819 96309 22828
rect 576 22700 99516 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 7112 22700
rect 7152 22660 7194 22700
rect 7234 22660 7276 22700
rect 7316 22660 7358 22700
rect 7398 22660 7440 22700
rect 7480 22660 11112 22700
rect 11152 22660 11194 22700
rect 11234 22660 11276 22700
rect 11316 22660 11358 22700
rect 11398 22660 11440 22700
rect 11480 22660 15112 22700
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15480 22660 19112 22700
rect 19152 22660 19194 22700
rect 19234 22660 19276 22700
rect 19316 22660 19358 22700
rect 19398 22660 19440 22700
rect 19480 22660 23112 22700
rect 23152 22660 23194 22700
rect 23234 22660 23276 22700
rect 23316 22660 23358 22700
rect 23398 22660 23440 22700
rect 23480 22660 27112 22700
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27480 22660 31112 22700
rect 31152 22660 31194 22700
rect 31234 22660 31276 22700
rect 31316 22660 31358 22700
rect 31398 22660 31440 22700
rect 31480 22660 35112 22700
rect 35152 22660 35194 22700
rect 35234 22660 35276 22700
rect 35316 22660 35358 22700
rect 35398 22660 35440 22700
rect 35480 22660 39112 22700
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39480 22660 43112 22700
rect 43152 22660 43194 22700
rect 43234 22660 43276 22700
rect 43316 22660 43358 22700
rect 43398 22660 43440 22700
rect 43480 22660 47112 22700
rect 47152 22660 47194 22700
rect 47234 22660 47276 22700
rect 47316 22660 47358 22700
rect 47398 22660 47440 22700
rect 47480 22660 51112 22700
rect 51152 22660 51194 22700
rect 51234 22660 51276 22700
rect 51316 22660 51358 22700
rect 51398 22660 51440 22700
rect 51480 22660 55112 22700
rect 55152 22660 55194 22700
rect 55234 22660 55276 22700
rect 55316 22660 55358 22700
rect 55398 22660 55440 22700
rect 55480 22660 59112 22700
rect 59152 22660 59194 22700
rect 59234 22660 59276 22700
rect 59316 22660 59358 22700
rect 59398 22660 59440 22700
rect 59480 22660 63112 22700
rect 63152 22660 63194 22700
rect 63234 22660 63276 22700
rect 63316 22660 63358 22700
rect 63398 22660 63440 22700
rect 63480 22660 67112 22700
rect 67152 22660 67194 22700
rect 67234 22660 67276 22700
rect 67316 22660 67358 22700
rect 67398 22660 67440 22700
rect 67480 22660 71112 22700
rect 71152 22660 71194 22700
rect 71234 22660 71276 22700
rect 71316 22660 71358 22700
rect 71398 22660 71440 22700
rect 71480 22660 75112 22700
rect 75152 22660 75194 22700
rect 75234 22660 75276 22700
rect 75316 22660 75358 22700
rect 75398 22660 75440 22700
rect 75480 22660 79112 22700
rect 79152 22660 79194 22700
rect 79234 22660 79276 22700
rect 79316 22660 79358 22700
rect 79398 22660 79440 22700
rect 79480 22660 83112 22700
rect 83152 22660 83194 22700
rect 83234 22660 83276 22700
rect 83316 22660 83358 22700
rect 83398 22660 83440 22700
rect 83480 22660 87112 22700
rect 87152 22660 87194 22700
rect 87234 22660 87276 22700
rect 87316 22660 87358 22700
rect 87398 22660 87440 22700
rect 87480 22660 91112 22700
rect 91152 22660 91194 22700
rect 91234 22660 91276 22700
rect 91316 22660 91358 22700
rect 91398 22660 91440 22700
rect 91480 22660 95112 22700
rect 95152 22660 95194 22700
rect 95234 22660 95276 22700
rect 95316 22660 95358 22700
rect 95398 22660 95440 22700
rect 95480 22660 99112 22700
rect 99152 22660 99194 22700
rect 99234 22660 99276 22700
rect 99316 22660 99358 22700
rect 99398 22660 99440 22700
rect 99480 22660 99516 22700
rect 576 22636 99516 22660
rect 73899 22532 73941 22541
rect 73899 22492 73900 22532
rect 73940 22492 73941 22532
rect 73899 22483 73941 22492
rect 74571 22532 74613 22541
rect 74571 22492 74572 22532
rect 74612 22492 74613 22532
rect 74571 22483 74613 22492
rect 75435 22532 75477 22541
rect 75435 22492 75436 22532
rect 75476 22492 75477 22532
rect 75435 22483 75477 22492
rect 75915 22532 75957 22541
rect 75915 22492 75916 22532
rect 75956 22492 75957 22532
rect 75915 22483 75957 22492
rect 76299 22532 76341 22541
rect 76299 22492 76300 22532
rect 76340 22492 76341 22532
rect 76299 22483 76341 22492
rect 76683 22532 76725 22541
rect 76683 22492 76684 22532
rect 76724 22492 76725 22532
rect 76683 22483 76725 22492
rect 77259 22532 77301 22541
rect 77259 22492 77260 22532
rect 77300 22492 77301 22532
rect 77259 22483 77301 22492
rect 77931 22532 77973 22541
rect 77931 22492 77932 22532
rect 77972 22492 77973 22532
rect 77931 22483 77973 22492
rect 78315 22532 78357 22541
rect 78315 22492 78316 22532
rect 78356 22492 78357 22532
rect 78315 22483 78357 22492
rect 79755 22532 79797 22541
rect 79755 22492 79756 22532
rect 79796 22492 79797 22532
rect 79755 22483 79797 22492
rect 80139 22532 80181 22541
rect 80139 22492 80140 22532
rect 80180 22492 80181 22532
rect 80139 22483 80181 22492
rect 80619 22532 80661 22541
rect 80619 22492 80620 22532
rect 80660 22492 80661 22532
rect 80619 22483 80661 22492
rect 80811 22532 80853 22541
rect 80811 22492 80812 22532
rect 80852 22492 80853 22532
rect 80811 22483 80853 22492
rect 81483 22532 81525 22541
rect 81483 22492 81484 22532
rect 81524 22492 81525 22532
rect 81483 22483 81525 22492
rect 81867 22532 81909 22541
rect 81867 22492 81868 22532
rect 81908 22492 81909 22532
rect 81867 22483 81909 22492
rect 83019 22532 83061 22541
rect 83019 22492 83020 22532
rect 83060 22492 83061 22532
rect 83019 22483 83061 22492
rect 83595 22532 83637 22541
rect 83595 22492 83596 22532
rect 83636 22492 83637 22532
rect 83595 22483 83637 22492
rect 83979 22532 84021 22541
rect 83979 22492 83980 22532
rect 84020 22492 84021 22532
rect 83979 22483 84021 22492
rect 84747 22532 84789 22541
rect 84747 22492 84748 22532
rect 84788 22492 84789 22532
rect 84747 22483 84789 22492
rect 85131 22532 85173 22541
rect 85131 22492 85132 22532
rect 85172 22492 85173 22532
rect 85131 22483 85173 22492
rect 85419 22532 85461 22541
rect 85419 22492 85420 22532
rect 85460 22492 85461 22532
rect 85419 22483 85461 22492
rect 85995 22532 86037 22541
rect 85995 22492 85996 22532
rect 86036 22492 86037 22532
rect 85995 22483 86037 22492
rect 86763 22532 86805 22541
rect 86763 22492 86764 22532
rect 86804 22492 86805 22532
rect 86763 22483 86805 22492
rect 87051 22532 87093 22541
rect 87051 22492 87052 22532
rect 87092 22492 87093 22532
rect 87051 22483 87093 22492
rect 87435 22532 87477 22541
rect 87435 22492 87436 22532
rect 87476 22492 87477 22532
rect 87435 22483 87477 22492
rect 87819 22532 87861 22541
rect 87819 22492 87820 22532
rect 87860 22492 87861 22532
rect 87819 22483 87861 22492
rect 88203 22532 88245 22541
rect 88203 22492 88204 22532
rect 88244 22492 88245 22532
rect 88203 22483 88245 22492
rect 88587 22532 88629 22541
rect 88587 22492 88588 22532
rect 88628 22492 88629 22532
rect 88587 22483 88629 22492
rect 89067 22532 89109 22541
rect 89067 22492 89068 22532
rect 89108 22492 89109 22532
rect 89067 22483 89109 22492
rect 89931 22532 89973 22541
rect 89931 22492 89932 22532
rect 89972 22492 89973 22532
rect 89931 22483 89973 22492
rect 90219 22532 90261 22541
rect 90219 22492 90220 22532
rect 90260 22492 90261 22532
rect 90219 22483 90261 22492
rect 90795 22532 90837 22541
rect 90795 22492 90796 22532
rect 90836 22492 90837 22532
rect 90795 22483 90837 22492
rect 91467 22532 91509 22541
rect 91467 22492 91468 22532
rect 91508 22492 91509 22532
rect 91467 22483 91509 22492
rect 91659 22532 91701 22541
rect 91659 22492 91660 22532
rect 91700 22492 91701 22532
rect 91659 22483 91701 22492
rect 92043 22532 92085 22541
rect 92043 22492 92044 22532
rect 92084 22492 92085 22532
rect 92043 22483 92085 22492
rect 92427 22532 92469 22541
rect 92427 22492 92428 22532
rect 92468 22492 92469 22532
rect 92427 22483 92469 22492
rect 92811 22532 92853 22541
rect 92811 22492 92812 22532
rect 92852 22492 92853 22532
rect 92811 22483 92853 22492
rect 93963 22532 94005 22541
rect 93963 22492 93964 22532
rect 94004 22492 94005 22532
rect 93963 22483 94005 22492
rect 94347 22532 94389 22541
rect 94347 22492 94348 22532
rect 94388 22492 94389 22532
rect 94347 22483 94389 22492
rect 94635 22532 94677 22541
rect 94635 22492 94636 22532
rect 94676 22492 94677 22532
rect 94635 22483 94677 22492
rect 95499 22532 95541 22541
rect 95499 22492 95500 22532
rect 95540 22492 95541 22532
rect 95499 22483 95541 22492
rect 95883 22532 95925 22541
rect 95883 22492 95884 22532
rect 95924 22492 95925 22532
rect 95883 22483 95925 22492
rect 96267 22532 96309 22541
rect 96267 22492 96268 22532
rect 96308 22492 96309 22532
rect 96267 22483 96309 22492
rect 96747 22532 96789 22541
rect 96747 22492 96748 22532
rect 96788 22492 96789 22532
rect 96747 22483 96789 22492
rect 97035 22532 97077 22541
rect 97035 22492 97036 22532
rect 97076 22492 97077 22532
rect 97035 22483 97077 22492
rect 97611 22532 97653 22541
rect 97611 22492 97612 22532
rect 97652 22492 97653 22532
rect 97611 22483 97653 22492
rect 97995 22532 98037 22541
rect 97995 22492 97996 22532
rect 98036 22492 98037 22532
rect 97995 22483 98037 22492
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 75051 22448 75093 22457
rect 75051 22408 75052 22448
rect 75092 22408 75093 22448
rect 75051 22399 75093 22408
rect 95115 22448 95157 22457
rect 95115 22408 95116 22448
rect 95156 22408 95157 22448
rect 95115 22399 95157 22408
rect 74755 22364 74813 22365
rect 74755 22324 74764 22364
rect 74804 22324 74813 22364
rect 74755 22323 74813 22324
rect 75235 22364 75293 22365
rect 75235 22324 75244 22364
rect 75284 22324 75293 22364
rect 75235 22323 75293 22324
rect 75619 22364 75677 22365
rect 75619 22324 75628 22364
rect 75668 22324 75677 22364
rect 75619 22323 75677 22324
rect 76099 22364 76157 22365
rect 76099 22324 76108 22364
rect 76148 22324 76157 22364
rect 76099 22323 76157 22324
rect 77731 22364 77789 22365
rect 77731 22324 77740 22364
rect 77780 22324 77789 22364
rect 77731 22323 77789 22324
rect 78115 22364 78173 22365
rect 78115 22324 78124 22364
rect 78164 22324 78173 22364
rect 78115 22323 78173 22324
rect 79555 22364 79613 22365
rect 79555 22324 79564 22364
rect 79604 22324 79613 22364
rect 79555 22323 79613 22324
rect 79939 22364 79997 22365
rect 79939 22324 79948 22364
rect 79988 22324 79997 22364
rect 79939 22323 79997 22324
rect 80419 22364 80477 22365
rect 80419 22324 80428 22364
rect 80468 22324 80477 22364
rect 80419 22323 80477 22324
rect 81283 22364 81341 22365
rect 81283 22324 81292 22364
rect 81332 22324 81341 22364
rect 81283 22323 81341 22324
rect 81667 22364 81725 22365
rect 81667 22324 81676 22364
rect 81716 22324 81725 22364
rect 81667 22323 81725 22324
rect 83203 22364 83261 22365
rect 83203 22324 83212 22364
rect 83252 22324 83261 22364
rect 83203 22323 83261 22324
rect 83779 22364 83837 22365
rect 83779 22324 83788 22364
rect 83828 22324 83837 22364
rect 83779 22323 83837 22324
rect 84547 22364 84605 22365
rect 84547 22324 84556 22364
rect 84596 22324 84605 22364
rect 84547 22323 84605 22324
rect 84931 22364 84989 22365
rect 84931 22324 84940 22364
rect 84980 22324 84989 22364
rect 84931 22323 84989 22324
rect 85603 22364 85661 22365
rect 85603 22324 85612 22364
rect 85652 22324 85661 22364
rect 85603 22323 85661 22324
rect 85795 22364 85853 22365
rect 85795 22324 85804 22364
rect 85844 22324 85853 22364
rect 85795 22323 85853 22324
rect 86371 22364 86429 22365
rect 86371 22324 86380 22364
rect 86420 22324 86429 22364
rect 86371 22323 86429 22324
rect 86563 22364 86621 22365
rect 86563 22324 86572 22364
rect 86612 22324 86621 22364
rect 86563 22323 86621 22324
rect 87235 22364 87293 22365
rect 87235 22324 87244 22364
rect 87284 22324 87293 22364
rect 87235 22323 87293 22324
rect 87619 22364 87677 22365
rect 87619 22324 87628 22364
rect 87668 22324 87677 22364
rect 87619 22323 87677 22324
rect 88003 22364 88061 22365
rect 88003 22324 88012 22364
rect 88052 22324 88061 22364
rect 88003 22323 88061 22324
rect 88387 22364 88445 22365
rect 88387 22324 88396 22364
rect 88436 22324 88445 22364
rect 88387 22323 88445 22324
rect 88867 22364 88925 22365
rect 88867 22324 88876 22364
rect 88916 22324 88925 22364
rect 88867 22323 88925 22324
rect 89731 22364 89789 22365
rect 89731 22324 89740 22364
rect 89780 22324 89789 22364
rect 89731 22323 89789 22324
rect 90403 22364 90461 22365
rect 90403 22324 90412 22364
rect 90452 22324 90461 22364
rect 90403 22323 90461 22324
rect 90595 22364 90653 22365
rect 90595 22324 90604 22364
rect 90644 22324 90653 22364
rect 90595 22323 90653 22324
rect 91267 22364 91325 22365
rect 91267 22324 91276 22364
rect 91316 22324 91325 22364
rect 91267 22323 91325 22324
rect 91843 22364 91901 22365
rect 91843 22324 91852 22364
rect 91892 22324 91901 22364
rect 91843 22323 91901 22324
rect 92227 22364 92285 22365
rect 92227 22324 92236 22364
rect 92276 22324 92285 22364
rect 92227 22323 92285 22324
rect 92611 22364 92669 22365
rect 92611 22324 92620 22364
rect 92660 22324 92669 22364
rect 92611 22323 92669 22324
rect 92995 22364 93053 22365
rect 92995 22324 93004 22364
rect 93044 22324 93053 22364
rect 92995 22323 93053 22324
rect 93763 22364 93821 22365
rect 93763 22324 93772 22364
rect 93812 22324 93821 22364
rect 93763 22323 93821 22324
rect 94147 22364 94205 22365
rect 94147 22324 94156 22364
rect 94196 22324 94205 22364
rect 94147 22323 94205 22324
rect 94915 22364 94973 22365
rect 94915 22324 94924 22364
rect 94964 22324 94973 22364
rect 94915 22323 94973 22324
rect 95299 22364 95357 22365
rect 95299 22324 95308 22364
rect 95348 22324 95357 22364
rect 95299 22323 95357 22324
rect 95683 22364 95741 22365
rect 95683 22324 95692 22364
rect 95732 22324 95741 22364
rect 95683 22323 95741 22324
rect 96067 22364 96125 22365
rect 96067 22324 96076 22364
rect 96116 22324 96125 22364
rect 96067 22323 96125 22324
rect 96547 22364 96605 22365
rect 96547 22324 96556 22364
rect 96596 22324 96605 22364
rect 96547 22323 96605 22324
rect 97219 22364 97277 22365
rect 97219 22324 97228 22364
rect 97268 22324 97277 22364
rect 97219 22323 97277 22324
rect 97795 22364 97853 22365
rect 97795 22324 97804 22364
rect 97844 22324 97853 22364
rect 97795 22323 97853 22324
rect 98179 22364 98237 22365
rect 98179 22324 98188 22364
rect 98228 22324 98237 22364
rect 98179 22323 98237 22324
rect 73795 22280 73853 22281
rect 73795 22240 73804 22280
rect 73844 22240 73853 22280
rect 73795 22239 73853 22240
rect 75811 22280 75869 22281
rect 75811 22240 75820 22280
rect 75860 22240 75869 22280
rect 75811 22239 75869 22240
rect 76579 22280 76637 22281
rect 76579 22240 76588 22280
rect 76628 22240 76637 22280
rect 76579 22239 76637 22240
rect 77155 22280 77213 22281
rect 77155 22240 77164 22280
rect 77204 22240 77213 22280
rect 77155 22239 77213 22240
rect 78787 22280 78845 22281
rect 78787 22240 78796 22280
rect 78836 22240 78845 22280
rect 78787 22239 78845 22240
rect 80899 22280 80957 22281
rect 80899 22240 80908 22280
rect 80948 22240 80957 22280
rect 80899 22239 80957 22240
rect 83491 22280 83549 22281
rect 83491 22240 83500 22280
rect 83540 22240 83549 22280
rect 83491 22239 83549 22240
rect 84259 22280 84317 22281
rect 84259 22240 84268 22280
rect 84308 22240 84317 22280
rect 84259 22239 84317 22240
rect 86947 22280 87005 22281
rect 86947 22240 86956 22280
rect 86996 22240 87005 22280
rect 86947 22239 87005 22240
rect 90979 22280 91037 22281
rect 90979 22240 90988 22280
rect 91028 22240 91037 22280
rect 90979 22239 91037 22240
rect 91083 22280 91125 22289
rect 91083 22240 91084 22280
rect 91124 22240 91125 22280
rect 91083 22231 91125 22240
rect 93475 22280 93533 22281
rect 93475 22240 93484 22280
rect 93524 22240 93533 22280
rect 93475 22239 93533 22240
rect 94531 22280 94589 22281
rect 94531 22240 94540 22280
rect 94580 22240 94589 22280
rect 94531 22239 94589 22240
rect 93579 22196 93621 22205
rect 93579 22156 93580 22196
rect 93620 22156 93621 22196
rect 93579 22147 93621 22156
rect 78891 22112 78933 22121
rect 78891 22072 78892 22112
rect 78932 22072 78933 22112
rect 78891 22063 78933 22072
rect 84171 22112 84213 22121
rect 84171 22072 84172 22112
rect 84212 22072 84213 22112
rect 84171 22063 84213 22072
rect 86187 22112 86229 22121
rect 86187 22072 86188 22112
rect 86228 22072 86229 22112
rect 86187 22063 86229 22072
rect 576 21944 99360 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 8352 21944
rect 8392 21904 8434 21944
rect 8474 21904 8516 21944
rect 8556 21904 8598 21944
rect 8638 21904 8680 21944
rect 8720 21904 12352 21944
rect 12392 21904 12434 21944
rect 12474 21904 12516 21944
rect 12556 21904 12598 21944
rect 12638 21904 12680 21944
rect 12720 21904 16352 21944
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16720 21904 20352 21944
rect 20392 21904 20434 21944
rect 20474 21904 20516 21944
rect 20556 21904 20598 21944
rect 20638 21904 20680 21944
rect 20720 21904 24352 21944
rect 24392 21904 24434 21944
rect 24474 21904 24516 21944
rect 24556 21904 24598 21944
rect 24638 21904 24680 21944
rect 24720 21904 28352 21944
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28720 21904 32352 21944
rect 32392 21904 32434 21944
rect 32474 21904 32516 21944
rect 32556 21904 32598 21944
rect 32638 21904 32680 21944
rect 32720 21904 36352 21944
rect 36392 21904 36434 21944
rect 36474 21904 36516 21944
rect 36556 21904 36598 21944
rect 36638 21904 36680 21944
rect 36720 21904 40352 21944
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40720 21904 44352 21944
rect 44392 21904 44434 21944
rect 44474 21904 44516 21944
rect 44556 21904 44598 21944
rect 44638 21904 44680 21944
rect 44720 21904 48352 21944
rect 48392 21904 48434 21944
rect 48474 21904 48516 21944
rect 48556 21904 48598 21944
rect 48638 21904 48680 21944
rect 48720 21904 52352 21944
rect 52392 21904 52434 21944
rect 52474 21904 52516 21944
rect 52556 21904 52598 21944
rect 52638 21904 52680 21944
rect 52720 21904 56352 21944
rect 56392 21904 56434 21944
rect 56474 21904 56516 21944
rect 56556 21904 56598 21944
rect 56638 21904 56680 21944
rect 56720 21904 60352 21944
rect 60392 21904 60434 21944
rect 60474 21904 60516 21944
rect 60556 21904 60598 21944
rect 60638 21904 60680 21944
rect 60720 21904 64352 21944
rect 64392 21904 64434 21944
rect 64474 21904 64516 21944
rect 64556 21904 64598 21944
rect 64638 21904 64680 21944
rect 64720 21904 68352 21944
rect 68392 21904 68434 21944
rect 68474 21904 68516 21944
rect 68556 21904 68598 21944
rect 68638 21904 68680 21944
rect 68720 21904 72352 21944
rect 72392 21904 72434 21944
rect 72474 21904 72516 21944
rect 72556 21904 72598 21944
rect 72638 21904 72680 21944
rect 72720 21904 76352 21944
rect 76392 21904 76434 21944
rect 76474 21904 76516 21944
rect 76556 21904 76598 21944
rect 76638 21904 76680 21944
rect 76720 21904 80352 21944
rect 80392 21904 80434 21944
rect 80474 21904 80516 21944
rect 80556 21904 80598 21944
rect 80638 21904 80680 21944
rect 80720 21904 84352 21944
rect 84392 21904 84434 21944
rect 84474 21904 84516 21944
rect 84556 21904 84598 21944
rect 84638 21904 84680 21944
rect 84720 21904 88352 21944
rect 88392 21904 88434 21944
rect 88474 21904 88516 21944
rect 88556 21904 88598 21944
rect 88638 21904 88680 21944
rect 88720 21904 92352 21944
rect 92392 21904 92434 21944
rect 92474 21904 92516 21944
rect 92556 21904 92598 21944
rect 92638 21904 92680 21944
rect 92720 21904 96352 21944
rect 96392 21904 96434 21944
rect 96474 21904 96516 21944
rect 96556 21904 96598 21944
rect 96638 21904 96680 21944
rect 96720 21904 99360 21944
rect 576 21880 99360 21904
rect 75819 21776 75861 21785
rect 75819 21736 75820 21776
rect 75860 21736 75861 21776
rect 75819 21727 75861 21736
rect 76779 21776 76821 21785
rect 76779 21736 76780 21776
rect 76820 21736 76821 21776
rect 76779 21727 76821 21736
rect 77643 21776 77685 21785
rect 77643 21736 77644 21776
rect 77684 21736 77685 21776
rect 77643 21727 77685 21736
rect 79083 21776 79125 21785
rect 79083 21736 79084 21776
rect 79124 21736 79125 21776
rect 79083 21727 79125 21736
rect 79467 21776 79509 21785
rect 79467 21736 79468 21776
rect 79508 21736 79509 21776
rect 79467 21727 79509 21736
rect 81003 21776 81045 21785
rect 81003 21736 81004 21776
rect 81044 21736 81045 21776
rect 81003 21727 81045 21736
rect 82347 21776 82389 21785
rect 82347 21736 82348 21776
rect 82388 21736 82389 21776
rect 82347 21727 82389 21736
rect 82539 21776 82581 21785
rect 82539 21736 82540 21776
rect 82580 21736 82581 21776
rect 82539 21727 82581 21736
rect 83595 21776 83637 21785
rect 83595 21736 83596 21776
rect 83636 21736 83637 21776
rect 83595 21727 83637 21736
rect 84363 21776 84405 21785
rect 84363 21736 84364 21776
rect 84404 21736 84405 21776
rect 84363 21727 84405 21736
rect 85995 21776 86037 21785
rect 85995 21736 85996 21776
rect 86036 21736 86037 21776
rect 85995 21727 86037 21736
rect 86379 21776 86421 21785
rect 86379 21736 86380 21776
rect 86420 21736 86421 21776
rect 86379 21727 86421 21736
rect 86859 21776 86901 21785
rect 86859 21736 86860 21776
rect 86900 21736 86901 21776
rect 86859 21727 86901 21736
rect 89067 21776 89109 21785
rect 89067 21736 89068 21776
rect 89108 21736 89109 21776
rect 89067 21727 89109 21736
rect 89547 21776 89589 21785
rect 89547 21736 89548 21776
rect 89588 21736 89589 21776
rect 89547 21727 89589 21736
rect 91179 21776 91221 21785
rect 91179 21736 91180 21776
rect 91220 21736 91221 21776
rect 91179 21727 91221 21736
rect 92811 21776 92853 21785
rect 92811 21736 92812 21776
rect 92852 21736 92853 21776
rect 92811 21727 92853 21736
rect 93291 21776 93333 21785
rect 93291 21736 93292 21776
rect 93332 21736 93333 21776
rect 93291 21727 93333 21736
rect 95211 21776 95253 21785
rect 95211 21736 95212 21776
rect 95252 21736 95253 21776
rect 95211 21727 95253 21736
rect 75715 21608 75773 21609
rect 75715 21568 75724 21608
rect 75764 21568 75773 21608
rect 75715 21567 75773 21568
rect 77539 21608 77597 21609
rect 77539 21568 77548 21608
rect 77588 21568 77597 21608
rect 77539 21567 77597 21568
rect 82627 21608 82685 21609
rect 82627 21568 82636 21608
rect 82676 21568 82685 21608
rect 82627 21567 82685 21568
rect 85891 21608 85949 21609
rect 85891 21568 85900 21608
rect 85940 21568 85949 21608
rect 85891 21567 85949 21568
rect 86467 21608 86525 21609
rect 86467 21568 86476 21608
rect 86516 21568 86525 21608
rect 86467 21567 86525 21568
rect 86755 21608 86813 21609
rect 86755 21568 86764 21608
rect 86804 21568 86813 21608
rect 86755 21567 86813 21568
rect 89155 21608 89213 21609
rect 89155 21568 89164 21608
rect 89204 21568 89213 21608
rect 89155 21567 89213 21568
rect 91075 21608 91133 21609
rect 91075 21568 91084 21608
rect 91124 21568 91133 21608
rect 91075 21567 91133 21568
rect 92707 21608 92765 21609
rect 92707 21568 92716 21608
rect 92756 21568 92765 21608
rect 92707 21567 92765 21568
rect 93379 21608 93437 21609
rect 93379 21568 93388 21608
rect 93428 21568 93437 21608
rect 93379 21567 93437 21568
rect 95299 21608 95357 21609
rect 95299 21568 95308 21608
rect 95348 21568 95357 21608
rect 95299 21567 95357 21568
rect 76579 21524 76637 21525
rect 76579 21484 76588 21524
rect 76628 21484 76637 21524
rect 76579 21483 76637 21484
rect 78883 21524 78941 21525
rect 78883 21484 78892 21524
rect 78932 21484 78941 21524
rect 78883 21483 78941 21484
rect 79267 21524 79325 21525
rect 79267 21484 79276 21524
rect 79316 21484 79325 21524
rect 79267 21483 79325 21484
rect 80803 21524 80861 21525
rect 80803 21484 80812 21524
rect 80852 21484 80861 21524
rect 80803 21483 80861 21484
rect 82147 21524 82205 21525
rect 82147 21484 82156 21524
rect 82196 21484 82205 21524
rect 82147 21483 82205 21484
rect 83395 21524 83453 21525
rect 83395 21484 83404 21524
rect 83444 21484 83453 21524
rect 83395 21483 83453 21484
rect 84163 21524 84221 21525
rect 84163 21484 84172 21524
rect 84212 21484 84221 21524
rect 84163 21483 84221 21484
rect 89347 21524 89405 21525
rect 89347 21484 89356 21524
rect 89396 21484 89405 21524
rect 89347 21483 89405 21484
rect 576 21188 99516 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 7112 21188
rect 7152 21148 7194 21188
rect 7234 21148 7276 21188
rect 7316 21148 7358 21188
rect 7398 21148 7440 21188
rect 7480 21148 11112 21188
rect 11152 21148 11194 21188
rect 11234 21148 11276 21188
rect 11316 21148 11358 21188
rect 11398 21148 11440 21188
rect 11480 21148 15112 21188
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15480 21148 19112 21188
rect 19152 21148 19194 21188
rect 19234 21148 19276 21188
rect 19316 21148 19358 21188
rect 19398 21148 19440 21188
rect 19480 21148 23112 21188
rect 23152 21148 23194 21188
rect 23234 21148 23276 21188
rect 23316 21148 23358 21188
rect 23398 21148 23440 21188
rect 23480 21148 27112 21188
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27480 21148 31112 21188
rect 31152 21148 31194 21188
rect 31234 21148 31276 21188
rect 31316 21148 31358 21188
rect 31398 21148 31440 21188
rect 31480 21148 35112 21188
rect 35152 21148 35194 21188
rect 35234 21148 35276 21188
rect 35316 21148 35358 21188
rect 35398 21148 35440 21188
rect 35480 21148 39112 21188
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39480 21148 43112 21188
rect 43152 21148 43194 21188
rect 43234 21148 43276 21188
rect 43316 21148 43358 21188
rect 43398 21148 43440 21188
rect 43480 21148 47112 21188
rect 47152 21148 47194 21188
rect 47234 21148 47276 21188
rect 47316 21148 47358 21188
rect 47398 21148 47440 21188
rect 47480 21148 51112 21188
rect 51152 21148 51194 21188
rect 51234 21148 51276 21188
rect 51316 21148 51358 21188
rect 51398 21148 51440 21188
rect 51480 21148 55112 21188
rect 55152 21148 55194 21188
rect 55234 21148 55276 21188
rect 55316 21148 55358 21188
rect 55398 21148 55440 21188
rect 55480 21148 59112 21188
rect 59152 21148 59194 21188
rect 59234 21148 59276 21188
rect 59316 21148 59358 21188
rect 59398 21148 59440 21188
rect 59480 21148 63112 21188
rect 63152 21148 63194 21188
rect 63234 21148 63276 21188
rect 63316 21148 63358 21188
rect 63398 21148 63440 21188
rect 63480 21148 67112 21188
rect 67152 21148 67194 21188
rect 67234 21148 67276 21188
rect 67316 21148 67358 21188
rect 67398 21148 67440 21188
rect 67480 21148 71112 21188
rect 71152 21148 71194 21188
rect 71234 21148 71276 21188
rect 71316 21148 71358 21188
rect 71398 21148 71440 21188
rect 71480 21148 75112 21188
rect 75152 21148 75194 21188
rect 75234 21148 75276 21188
rect 75316 21148 75358 21188
rect 75398 21148 75440 21188
rect 75480 21148 79112 21188
rect 79152 21148 79194 21188
rect 79234 21148 79276 21188
rect 79316 21148 79358 21188
rect 79398 21148 79440 21188
rect 79480 21148 83112 21188
rect 83152 21148 83194 21188
rect 83234 21148 83276 21188
rect 83316 21148 83358 21188
rect 83398 21148 83440 21188
rect 83480 21148 87112 21188
rect 87152 21148 87194 21188
rect 87234 21148 87276 21188
rect 87316 21148 87358 21188
rect 87398 21148 87440 21188
rect 87480 21148 91112 21188
rect 91152 21148 91194 21188
rect 91234 21148 91276 21188
rect 91316 21148 91358 21188
rect 91398 21148 91440 21188
rect 91480 21148 95112 21188
rect 95152 21148 95194 21188
rect 95234 21148 95276 21188
rect 95316 21148 95358 21188
rect 95398 21148 95440 21188
rect 95480 21148 99112 21188
rect 99152 21148 99194 21188
rect 99234 21148 99276 21188
rect 99316 21148 99358 21188
rect 99398 21148 99440 21188
rect 99480 21148 99516 21188
rect 576 21124 99516 21148
rect 651 20936 693 20945
rect 651 20896 652 20936
rect 692 20896 693 20936
rect 651 20887 693 20896
rect 576 20432 99360 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 8352 20432
rect 8392 20392 8434 20432
rect 8474 20392 8516 20432
rect 8556 20392 8598 20432
rect 8638 20392 8680 20432
rect 8720 20392 12352 20432
rect 12392 20392 12434 20432
rect 12474 20392 12516 20432
rect 12556 20392 12598 20432
rect 12638 20392 12680 20432
rect 12720 20392 16352 20432
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16720 20392 20352 20432
rect 20392 20392 20434 20432
rect 20474 20392 20516 20432
rect 20556 20392 20598 20432
rect 20638 20392 20680 20432
rect 20720 20392 24352 20432
rect 24392 20392 24434 20432
rect 24474 20392 24516 20432
rect 24556 20392 24598 20432
rect 24638 20392 24680 20432
rect 24720 20392 28352 20432
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28720 20392 32352 20432
rect 32392 20392 32434 20432
rect 32474 20392 32516 20432
rect 32556 20392 32598 20432
rect 32638 20392 32680 20432
rect 32720 20392 36352 20432
rect 36392 20392 36434 20432
rect 36474 20392 36516 20432
rect 36556 20392 36598 20432
rect 36638 20392 36680 20432
rect 36720 20392 40352 20432
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40720 20392 44352 20432
rect 44392 20392 44434 20432
rect 44474 20392 44516 20432
rect 44556 20392 44598 20432
rect 44638 20392 44680 20432
rect 44720 20392 48352 20432
rect 48392 20392 48434 20432
rect 48474 20392 48516 20432
rect 48556 20392 48598 20432
rect 48638 20392 48680 20432
rect 48720 20392 52352 20432
rect 52392 20392 52434 20432
rect 52474 20392 52516 20432
rect 52556 20392 52598 20432
rect 52638 20392 52680 20432
rect 52720 20392 56352 20432
rect 56392 20392 56434 20432
rect 56474 20392 56516 20432
rect 56556 20392 56598 20432
rect 56638 20392 56680 20432
rect 56720 20392 60352 20432
rect 60392 20392 60434 20432
rect 60474 20392 60516 20432
rect 60556 20392 60598 20432
rect 60638 20392 60680 20432
rect 60720 20392 64352 20432
rect 64392 20392 64434 20432
rect 64474 20392 64516 20432
rect 64556 20392 64598 20432
rect 64638 20392 64680 20432
rect 64720 20392 68352 20432
rect 68392 20392 68434 20432
rect 68474 20392 68516 20432
rect 68556 20392 68598 20432
rect 68638 20392 68680 20432
rect 68720 20392 72352 20432
rect 72392 20392 72434 20432
rect 72474 20392 72516 20432
rect 72556 20392 72598 20432
rect 72638 20392 72680 20432
rect 72720 20392 76352 20432
rect 76392 20392 76434 20432
rect 76474 20392 76516 20432
rect 76556 20392 76598 20432
rect 76638 20392 76680 20432
rect 76720 20392 80352 20432
rect 80392 20392 80434 20432
rect 80474 20392 80516 20432
rect 80556 20392 80598 20432
rect 80638 20392 80680 20432
rect 80720 20392 84352 20432
rect 84392 20392 84434 20432
rect 84474 20392 84516 20432
rect 84556 20392 84598 20432
rect 84638 20392 84680 20432
rect 84720 20392 88352 20432
rect 88392 20392 88434 20432
rect 88474 20392 88516 20432
rect 88556 20392 88598 20432
rect 88638 20392 88680 20432
rect 88720 20392 92352 20432
rect 92392 20392 92434 20432
rect 92474 20392 92516 20432
rect 92556 20392 92598 20432
rect 92638 20392 92680 20432
rect 92720 20392 96352 20432
rect 96392 20392 96434 20432
rect 96474 20392 96516 20432
rect 96556 20392 96598 20432
rect 96638 20392 96680 20432
rect 96720 20392 99360 20432
rect 576 20368 99360 20392
rect 75523 20012 75581 20013
rect 75523 19972 75532 20012
rect 75572 19972 75581 20012
rect 75523 19971 75581 19972
rect 80611 20012 80669 20013
rect 80611 19972 80620 20012
rect 80660 19972 80669 20012
rect 80611 19971 80669 19972
rect 86851 20012 86909 20013
rect 86851 19972 86860 20012
rect 86900 19972 86909 20012
rect 86851 19971 86909 19972
rect 93187 20012 93245 20013
rect 93187 19972 93196 20012
rect 93236 19972 93245 20012
rect 93187 19971 93245 19972
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 75723 19928 75765 19937
rect 75723 19888 75724 19928
rect 75764 19888 75765 19928
rect 75723 19879 75765 19888
rect 80427 19844 80469 19853
rect 80427 19804 80428 19844
rect 80468 19804 80469 19844
rect 80427 19795 80469 19804
rect 87051 19844 87093 19853
rect 87051 19804 87052 19844
rect 87092 19804 87093 19844
rect 87051 19795 87093 19804
rect 93003 19844 93045 19853
rect 93003 19804 93004 19844
rect 93044 19804 93045 19844
rect 93003 19795 93045 19804
rect 576 19676 99516 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 7112 19676
rect 7152 19636 7194 19676
rect 7234 19636 7276 19676
rect 7316 19636 7358 19676
rect 7398 19636 7440 19676
rect 7480 19636 11112 19676
rect 11152 19636 11194 19676
rect 11234 19636 11276 19676
rect 11316 19636 11358 19676
rect 11398 19636 11440 19676
rect 11480 19636 15112 19676
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15480 19636 19112 19676
rect 19152 19636 19194 19676
rect 19234 19636 19276 19676
rect 19316 19636 19358 19676
rect 19398 19636 19440 19676
rect 19480 19636 23112 19676
rect 23152 19636 23194 19676
rect 23234 19636 23276 19676
rect 23316 19636 23358 19676
rect 23398 19636 23440 19676
rect 23480 19636 27112 19676
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27480 19636 31112 19676
rect 31152 19636 31194 19676
rect 31234 19636 31276 19676
rect 31316 19636 31358 19676
rect 31398 19636 31440 19676
rect 31480 19636 35112 19676
rect 35152 19636 35194 19676
rect 35234 19636 35276 19676
rect 35316 19636 35358 19676
rect 35398 19636 35440 19676
rect 35480 19636 39112 19676
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39480 19636 43112 19676
rect 43152 19636 43194 19676
rect 43234 19636 43276 19676
rect 43316 19636 43358 19676
rect 43398 19636 43440 19676
rect 43480 19636 47112 19676
rect 47152 19636 47194 19676
rect 47234 19636 47276 19676
rect 47316 19636 47358 19676
rect 47398 19636 47440 19676
rect 47480 19636 51112 19676
rect 51152 19636 51194 19676
rect 51234 19636 51276 19676
rect 51316 19636 51358 19676
rect 51398 19636 51440 19676
rect 51480 19636 55112 19676
rect 55152 19636 55194 19676
rect 55234 19636 55276 19676
rect 55316 19636 55358 19676
rect 55398 19636 55440 19676
rect 55480 19636 59112 19676
rect 59152 19636 59194 19676
rect 59234 19636 59276 19676
rect 59316 19636 59358 19676
rect 59398 19636 59440 19676
rect 59480 19636 63112 19676
rect 63152 19636 63194 19676
rect 63234 19636 63276 19676
rect 63316 19636 63358 19676
rect 63398 19636 63440 19676
rect 63480 19636 67112 19676
rect 67152 19636 67194 19676
rect 67234 19636 67276 19676
rect 67316 19636 67358 19676
rect 67398 19636 67440 19676
rect 67480 19636 71112 19676
rect 71152 19636 71194 19676
rect 71234 19636 71276 19676
rect 71316 19636 71358 19676
rect 71398 19636 71440 19676
rect 71480 19636 75112 19676
rect 75152 19636 75194 19676
rect 75234 19636 75276 19676
rect 75316 19636 75358 19676
rect 75398 19636 75440 19676
rect 75480 19636 79112 19676
rect 79152 19636 79194 19676
rect 79234 19636 79276 19676
rect 79316 19636 79358 19676
rect 79398 19636 79440 19676
rect 79480 19636 83112 19676
rect 83152 19636 83194 19676
rect 83234 19636 83276 19676
rect 83316 19636 83358 19676
rect 83398 19636 83440 19676
rect 83480 19636 87112 19676
rect 87152 19636 87194 19676
rect 87234 19636 87276 19676
rect 87316 19636 87358 19676
rect 87398 19636 87440 19676
rect 87480 19636 91112 19676
rect 91152 19636 91194 19676
rect 91234 19636 91276 19676
rect 91316 19636 91358 19676
rect 91398 19636 91440 19676
rect 91480 19636 95112 19676
rect 95152 19636 95194 19676
rect 95234 19636 95276 19676
rect 95316 19636 95358 19676
rect 95398 19636 95440 19676
rect 95480 19636 99112 19676
rect 99152 19636 99194 19676
rect 99234 19636 99276 19676
rect 99316 19636 99358 19676
rect 99398 19636 99440 19676
rect 99480 19636 99516 19676
rect 576 19612 99516 19636
rect 90123 19508 90165 19517
rect 90123 19468 90124 19508
rect 90164 19468 90165 19508
rect 90123 19459 90165 19468
rect 651 19424 693 19433
rect 651 19384 652 19424
rect 692 19384 693 19424
rect 651 19375 693 19384
rect 92907 19424 92949 19433
rect 92907 19384 92908 19424
rect 92948 19384 92949 19424
rect 92907 19375 92949 19384
rect 74755 19340 74813 19341
rect 74755 19300 74764 19340
rect 74804 19300 74813 19340
rect 74755 19299 74813 19300
rect 77635 19340 77693 19341
rect 77635 19300 77644 19340
rect 77684 19300 77693 19340
rect 77635 19299 77693 19300
rect 78211 19340 78269 19341
rect 78211 19300 78220 19340
rect 78260 19300 78269 19340
rect 78211 19299 78269 19300
rect 80515 19340 80573 19341
rect 80515 19300 80524 19340
rect 80564 19300 80573 19340
rect 80515 19299 80573 19300
rect 82051 19340 82109 19341
rect 82051 19300 82060 19340
rect 82100 19300 82109 19340
rect 82051 19299 82109 19300
rect 84067 19340 84125 19341
rect 84067 19300 84076 19340
rect 84116 19300 84125 19340
rect 84067 19299 84125 19300
rect 85603 19340 85661 19341
rect 85603 19300 85612 19340
rect 85652 19300 85661 19340
rect 85603 19299 85661 19300
rect 86563 19340 86621 19341
rect 86563 19300 86572 19340
rect 86612 19300 86621 19340
rect 86563 19299 86621 19300
rect 86755 19340 86813 19341
rect 86755 19300 86764 19340
rect 86804 19300 86813 19340
rect 86755 19299 86813 19300
rect 87427 19340 87485 19341
rect 87427 19300 87436 19340
rect 87476 19300 87485 19340
rect 87427 19299 87485 19300
rect 88195 19340 88253 19341
rect 88195 19300 88204 19340
rect 88244 19300 88253 19340
rect 88195 19299 88253 19300
rect 89731 19340 89789 19341
rect 89731 19300 89740 19340
rect 89780 19300 89789 19340
rect 89731 19299 89789 19300
rect 89923 19340 89981 19341
rect 89923 19300 89932 19340
rect 89972 19300 89981 19340
rect 89923 19299 89981 19300
rect 91363 19340 91421 19341
rect 91363 19300 91372 19340
rect 91412 19300 91421 19340
rect 91363 19299 91421 19300
rect 92515 19340 92573 19341
rect 92515 19300 92524 19340
rect 92564 19300 92573 19340
rect 92515 19299 92573 19300
rect 93091 19340 93149 19341
rect 93091 19300 93100 19340
rect 93140 19300 93149 19340
rect 93091 19299 93149 19300
rect 94147 19340 94205 19341
rect 94147 19300 94156 19340
rect 94196 19300 94205 19340
rect 94147 19299 94205 19300
rect 95779 19340 95837 19341
rect 95779 19300 95788 19340
rect 95828 19300 95837 19340
rect 95779 19299 95837 19300
rect 75235 19256 75293 19257
rect 75235 19216 75244 19256
rect 75284 19216 75293 19256
rect 75235 19215 75293 19216
rect 75427 19256 75485 19257
rect 75427 19216 75436 19256
rect 75476 19216 75485 19256
rect 75427 19215 75485 19216
rect 75619 19256 75677 19257
rect 75619 19216 75628 19256
rect 75668 19216 75677 19256
rect 75619 19215 75677 19216
rect 76579 19256 76637 19257
rect 76579 19216 76588 19256
rect 76628 19216 76637 19256
rect 76579 19215 76637 19216
rect 77059 19256 77117 19257
rect 77059 19216 77068 19256
rect 77108 19216 77117 19256
rect 77059 19215 77117 19216
rect 78595 19256 78653 19257
rect 78595 19216 78604 19256
rect 78644 19216 78653 19256
rect 78595 19215 78653 19216
rect 80035 19256 80093 19257
rect 80035 19216 80044 19256
rect 80084 19216 80093 19256
rect 80035 19215 80093 19216
rect 82627 19256 82685 19257
rect 82627 19216 82636 19256
rect 82676 19216 82685 19256
rect 82627 19215 82685 19216
rect 88483 19256 88541 19257
rect 88483 19216 88492 19256
rect 88532 19216 88541 19256
rect 88483 19215 88541 19216
rect 74955 19088 74997 19097
rect 74955 19048 74956 19088
rect 74996 19048 74997 19088
rect 74955 19039 74997 19048
rect 75723 19088 75765 19097
rect 75723 19048 75724 19088
rect 75764 19048 75765 19088
rect 75723 19039 75765 19048
rect 76683 19088 76725 19097
rect 76683 19048 76684 19088
rect 76724 19048 76725 19088
rect 76683 19039 76725 19048
rect 77163 19088 77205 19097
rect 77163 19048 77164 19088
rect 77204 19048 77205 19088
rect 77163 19039 77205 19048
rect 77835 19088 77877 19097
rect 77835 19048 77836 19088
rect 77876 19048 77877 19088
rect 77835 19039 77877 19048
rect 78027 19088 78069 19097
rect 78027 19048 78028 19088
rect 78068 19048 78069 19088
rect 78027 19039 78069 19048
rect 78699 19088 78741 19097
rect 78699 19048 78700 19088
rect 78740 19048 78741 19088
rect 78699 19039 78741 19048
rect 80139 19088 80181 19097
rect 80139 19048 80140 19088
rect 80180 19048 80181 19088
rect 80139 19039 80181 19048
rect 80331 19088 80373 19097
rect 80331 19048 80332 19088
rect 80372 19048 80373 19088
rect 80331 19039 80373 19048
rect 81867 19088 81909 19097
rect 81867 19048 81868 19088
rect 81908 19048 81909 19088
rect 81867 19039 81909 19048
rect 82731 19088 82773 19097
rect 82731 19048 82732 19088
rect 82772 19048 82773 19088
rect 82731 19039 82773 19048
rect 83883 19088 83925 19097
rect 83883 19048 83884 19088
rect 83924 19048 83925 19088
rect 83883 19039 83925 19048
rect 85803 19088 85845 19097
rect 85803 19048 85804 19088
rect 85844 19048 85845 19088
rect 85803 19039 85845 19048
rect 86379 19088 86421 19097
rect 86379 19048 86380 19088
rect 86420 19048 86421 19088
rect 86379 19039 86421 19048
rect 86955 19088 86997 19097
rect 86955 19048 86956 19088
rect 86996 19048 86997 19088
rect 86955 19039 86997 19048
rect 87627 19088 87669 19097
rect 87627 19048 87628 19088
rect 87668 19048 87669 19088
rect 87627 19039 87669 19048
rect 88011 19088 88053 19097
rect 88011 19048 88012 19088
rect 88052 19048 88053 19088
rect 88011 19039 88053 19048
rect 88395 19088 88437 19097
rect 88395 19048 88396 19088
rect 88436 19048 88437 19088
rect 88395 19039 88437 19048
rect 89547 19088 89589 19097
rect 89547 19048 89548 19088
rect 89588 19048 89589 19088
rect 89547 19039 89589 19048
rect 90123 19088 90165 19097
rect 90123 19048 90124 19088
rect 90164 19048 90165 19088
rect 90123 19039 90165 19048
rect 91563 19088 91605 19097
rect 91563 19048 91564 19088
rect 91604 19048 91605 19088
rect 91563 19039 91605 19048
rect 92715 19088 92757 19097
rect 92715 19048 92716 19088
rect 92756 19048 92757 19088
rect 92715 19039 92757 19048
rect 93963 19088 94005 19097
rect 93963 19048 93964 19088
rect 94004 19048 94005 19088
rect 93963 19039 94005 19048
rect 95595 19088 95637 19097
rect 95595 19048 95596 19088
rect 95636 19048 95637 19088
rect 95595 19039 95637 19048
rect 576 18920 99360 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 8352 18920
rect 8392 18880 8434 18920
rect 8474 18880 8516 18920
rect 8556 18880 8598 18920
rect 8638 18880 8680 18920
rect 8720 18880 12352 18920
rect 12392 18880 12434 18920
rect 12474 18880 12516 18920
rect 12556 18880 12598 18920
rect 12638 18880 12680 18920
rect 12720 18880 16352 18920
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16720 18880 20352 18920
rect 20392 18880 20434 18920
rect 20474 18880 20516 18920
rect 20556 18880 20598 18920
rect 20638 18880 20680 18920
rect 20720 18880 24352 18920
rect 24392 18880 24434 18920
rect 24474 18880 24516 18920
rect 24556 18880 24598 18920
rect 24638 18880 24680 18920
rect 24720 18880 28352 18920
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28720 18880 32352 18920
rect 32392 18880 32434 18920
rect 32474 18880 32516 18920
rect 32556 18880 32598 18920
rect 32638 18880 32680 18920
rect 32720 18880 36352 18920
rect 36392 18880 36434 18920
rect 36474 18880 36516 18920
rect 36556 18880 36598 18920
rect 36638 18880 36680 18920
rect 36720 18880 40352 18920
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40720 18880 44352 18920
rect 44392 18880 44434 18920
rect 44474 18880 44516 18920
rect 44556 18880 44598 18920
rect 44638 18880 44680 18920
rect 44720 18880 48352 18920
rect 48392 18880 48434 18920
rect 48474 18880 48516 18920
rect 48556 18880 48598 18920
rect 48638 18880 48680 18920
rect 48720 18880 52352 18920
rect 52392 18880 52434 18920
rect 52474 18880 52516 18920
rect 52556 18880 52598 18920
rect 52638 18880 52680 18920
rect 52720 18880 56352 18920
rect 56392 18880 56434 18920
rect 56474 18880 56516 18920
rect 56556 18880 56598 18920
rect 56638 18880 56680 18920
rect 56720 18880 60352 18920
rect 60392 18880 60434 18920
rect 60474 18880 60516 18920
rect 60556 18880 60598 18920
rect 60638 18880 60680 18920
rect 60720 18880 64352 18920
rect 64392 18880 64434 18920
rect 64474 18880 64516 18920
rect 64556 18880 64598 18920
rect 64638 18880 64680 18920
rect 64720 18880 68352 18920
rect 68392 18880 68434 18920
rect 68474 18880 68516 18920
rect 68556 18880 68598 18920
rect 68638 18880 68680 18920
rect 68720 18880 72352 18920
rect 72392 18880 72434 18920
rect 72474 18880 72516 18920
rect 72556 18880 72598 18920
rect 72638 18880 72680 18920
rect 72720 18880 76352 18920
rect 76392 18880 76434 18920
rect 76474 18880 76516 18920
rect 76556 18880 76598 18920
rect 76638 18880 76680 18920
rect 76720 18880 80352 18920
rect 80392 18880 80434 18920
rect 80474 18880 80516 18920
rect 80556 18880 80598 18920
rect 80638 18880 80680 18920
rect 80720 18880 84352 18920
rect 84392 18880 84434 18920
rect 84474 18880 84516 18920
rect 84556 18880 84598 18920
rect 84638 18880 84680 18920
rect 84720 18880 88352 18920
rect 88392 18880 88434 18920
rect 88474 18880 88516 18920
rect 88556 18880 88598 18920
rect 88638 18880 88680 18920
rect 88720 18880 92352 18920
rect 92392 18880 92434 18920
rect 92474 18880 92516 18920
rect 92556 18880 92598 18920
rect 92638 18880 92680 18920
rect 92720 18880 96352 18920
rect 96392 18880 96434 18920
rect 96474 18880 96516 18920
rect 96556 18880 96598 18920
rect 96638 18880 96680 18920
rect 96720 18880 99360 18920
rect 576 18856 99360 18880
rect 74955 18752 74997 18761
rect 74955 18712 74956 18752
rect 74996 18712 74997 18752
rect 74955 18703 74997 18712
rect 89443 18595 89501 18596
rect 72931 18584 72989 18585
rect 72931 18544 72940 18584
rect 72980 18544 72989 18584
rect 72931 18543 72989 18544
rect 74275 18584 74333 18585
rect 74275 18544 74284 18584
rect 74324 18544 74333 18584
rect 74275 18543 74333 18544
rect 76483 18584 76541 18585
rect 76483 18544 76492 18584
rect 76532 18544 76541 18584
rect 76483 18543 76541 18544
rect 77443 18584 77501 18585
rect 77443 18544 77452 18584
rect 77492 18544 77501 18584
rect 77443 18543 77501 18544
rect 78115 18584 78173 18585
rect 78115 18544 78124 18584
rect 78164 18544 78173 18584
rect 78115 18543 78173 18544
rect 85027 18584 85085 18585
rect 85027 18544 85036 18584
rect 85076 18544 85085 18584
rect 85027 18543 85085 18544
rect 86275 18584 86333 18585
rect 86275 18544 86284 18584
rect 86324 18544 86333 18584
rect 89443 18555 89452 18595
rect 89492 18555 89501 18595
rect 89443 18554 89501 18555
rect 92899 18584 92957 18585
rect 86275 18543 86333 18544
rect 92899 18544 92908 18584
rect 92948 18544 92957 18584
rect 92899 18543 92957 18544
rect 95107 18584 95165 18585
rect 95107 18544 95116 18584
rect 95156 18544 95165 18584
rect 95107 18543 95165 18544
rect 95971 18584 96029 18585
rect 95971 18544 95980 18584
rect 96020 18544 96029 18584
rect 95971 18543 96029 18544
rect 96931 18584 96989 18585
rect 96931 18544 96940 18584
rect 96980 18544 96989 18584
rect 96931 18543 96989 18544
rect 97603 18584 97661 18585
rect 97603 18544 97612 18584
rect 97652 18544 97661 18584
rect 97603 18543 97661 18544
rect 74563 18500 74621 18501
rect 74563 18460 74572 18500
rect 74612 18460 74621 18500
rect 74563 18459 74621 18460
rect 75139 18500 75197 18501
rect 75139 18460 75148 18500
rect 75188 18460 75197 18500
rect 75139 18459 75197 18460
rect 75811 18500 75869 18501
rect 75811 18460 75820 18500
rect 75860 18460 75869 18500
rect 75811 18459 75869 18460
rect 78403 18500 78461 18501
rect 78403 18460 78412 18500
rect 78452 18460 78461 18500
rect 78403 18459 78461 18460
rect 78979 18500 79037 18501
rect 78979 18460 78988 18500
rect 79028 18460 79037 18500
rect 78979 18459 79037 18460
rect 79363 18500 79421 18501
rect 79363 18460 79372 18500
rect 79412 18460 79421 18500
rect 79363 18459 79421 18460
rect 79843 18500 79901 18501
rect 79843 18460 79852 18500
rect 79892 18460 79901 18500
rect 79843 18459 79901 18460
rect 80995 18500 81053 18501
rect 80995 18460 81004 18500
rect 81044 18460 81053 18500
rect 80995 18459 81053 18460
rect 81379 18500 81437 18501
rect 81379 18460 81388 18500
rect 81428 18460 81437 18500
rect 81379 18459 81437 18460
rect 81763 18500 81821 18501
rect 81763 18460 81772 18500
rect 81812 18460 81821 18500
rect 81763 18459 81821 18460
rect 82243 18500 82301 18501
rect 82243 18460 82252 18500
rect 82292 18460 82301 18500
rect 82243 18459 82301 18460
rect 83011 18500 83069 18501
rect 83011 18460 83020 18500
rect 83060 18460 83069 18500
rect 83011 18459 83069 18460
rect 83395 18500 83453 18501
rect 83395 18460 83404 18500
rect 83444 18460 83453 18500
rect 83395 18459 83453 18460
rect 83779 18500 83837 18501
rect 83779 18460 83788 18500
rect 83828 18460 83837 18500
rect 83779 18459 83837 18460
rect 84259 18500 84317 18501
rect 84259 18460 84268 18500
rect 84308 18460 84317 18500
rect 84259 18459 84317 18460
rect 84643 18500 84701 18501
rect 84643 18460 84652 18500
rect 84692 18460 84701 18500
rect 84643 18459 84701 18460
rect 85507 18500 85565 18501
rect 85507 18460 85516 18500
rect 85556 18460 85565 18500
rect 85507 18459 85565 18460
rect 85891 18500 85949 18501
rect 85891 18460 85900 18500
rect 85940 18460 85949 18500
rect 85891 18459 85949 18460
rect 86563 18500 86621 18501
rect 86563 18460 86572 18500
rect 86612 18460 86621 18500
rect 86563 18459 86621 18460
rect 87043 18500 87101 18501
rect 87043 18460 87052 18500
rect 87092 18460 87101 18500
rect 87043 18459 87101 18460
rect 87715 18500 87773 18501
rect 87715 18460 87724 18500
rect 87764 18460 87773 18500
rect 87715 18459 87773 18460
rect 88195 18500 88253 18501
rect 88195 18460 88204 18500
rect 88244 18460 88253 18500
rect 88195 18459 88253 18460
rect 88579 18500 88637 18501
rect 88579 18460 88588 18500
rect 88628 18460 88637 18500
rect 88579 18459 88637 18460
rect 88963 18500 89021 18501
rect 88963 18460 88972 18500
rect 89012 18460 89021 18500
rect 88963 18459 89021 18460
rect 89731 18500 89789 18501
rect 89731 18460 89740 18500
rect 89780 18460 89789 18500
rect 89731 18459 89789 18460
rect 90115 18500 90173 18501
rect 90115 18460 90124 18500
rect 90164 18460 90173 18500
rect 90115 18459 90173 18460
rect 90595 18500 90653 18501
rect 90595 18460 90604 18500
rect 90644 18460 90653 18500
rect 90595 18459 90653 18460
rect 91267 18500 91325 18501
rect 91267 18460 91276 18500
rect 91316 18460 91325 18500
rect 91267 18459 91325 18460
rect 91843 18500 91901 18501
rect 91843 18460 91852 18500
rect 91892 18460 91901 18500
rect 91843 18459 91901 18460
rect 92227 18500 92285 18501
rect 92227 18460 92236 18500
rect 92276 18460 92285 18500
rect 92227 18459 92285 18460
rect 92611 18500 92669 18501
rect 92611 18460 92620 18500
rect 92660 18460 92669 18500
rect 92611 18459 92669 18460
rect 93091 18500 93149 18501
rect 93091 18460 93100 18500
rect 93140 18460 93149 18500
rect 93091 18459 93149 18460
rect 93859 18500 93917 18501
rect 93859 18460 93868 18500
rect 93908 18460 93917 18500
rect 93859 18459 93917 18460
rect 94243 18500 94301 18501
rect 94243 18460 94252 18500
rect 94292 18460 94301 18500
rect 94243 18459 94301 18460
rect 94915 18500 94973 18501
rect 94915 18460 94924 18500
rect 94964 18460 94973 18500
rect 94915 18459 94973 18460
rect 95491 18500 95549 18501
rect 95491 18460 95500 18500
rect 95540 18460 95549 18500
rect 95491 18459 95549 18460
rect 96259 18500 96317 18501
rect 96259 18460 96268 18500
rect 96308 18460 96317 18500
rect 96259 18459 96317 18460
rect 97123 18500 97181 18501
rect 97123 18460 97132 18500
rect 97172 18460 97181 18500
rect 97123 18459 97181 18460
rect 651 18416 693 18425
rect 651 18376 652 18416
rect 692 18376 693 18416
rect 651 18367 693 18376
rect 78795 18416 78837 18425
rect 78795 18376 78796 18416
rect 78836 18376 78837 18416
rect 78795 18367 78837 18376
rect 73035 18332 73077 18341
rect 73035 18292 73036 18332
rect 73076 18292 73077 18332
rect 73035 18283 73077 18292
rect 74187 18332 74229 18341
rect 74187 18292 74188 18332
rect 74228 18292 74229 18332
rect 74187 18283 74229 18292
rect 74763 18332 74805 18341
rect 74763 18292 74764 18332
rect 74804 18292 74805 18332
rect 74763 18283 74805 18292
rect 74955 18332 74997 18341
rect 74955 18292 74956 18332
rect 74996 18292 74997 18332
rect 74955 18283 74997 18292
rect 76011 18332 76053 18341
rect 76011 18292 76012 18332
rect 76052 18292 76053 18332
rect 76011 18283 76053 18292
rect 76587 18332 76629 18341
rect 76587 18292 76588 18332
rect 76628 18292 76629 18332
rect 76587 18283 76629 18292
rect 77547 18332 77589 18341
rect 77547 18292 77548 18332
rect 77588 18292 77589 18332
rect 77547 18283 77589 18292
rect 78219 18332 78261 18341
rect 78219 18292 78220 18332
rect 78260 18292 78261 18332
rect 78219 18283 78261 18292
rect 78603 18332 78645 18341
rect 78603 18292 78604 18332
rect 78644 18292 78645 18332
rect 78603 18283 78645 18292
rect 79563 18332 79605 18341
rect 79563 18292 79564 18332
rect 79604 18292 79605 18332
rect 79563 18283 79605 18292
rect 80043 18332 80085 18341
rect 80043 18292 80044 18332
rect 80084 18292 80085 18332
rect 80043 18283 80085 18292
rect 81195 18332 81237 18341
rect 81195 18292 81196 18332
rect 81236 18292 81237 18332
rect 81195 18283 81237 18292
rect 81579 18332 81621 18341
rect 81579 18292 81580 18332
rect 81620 18292 81621 18332
rect 81579 18283 81621 18292
rect 81963 18332 82005 18341
rect 81963 18292 81964 18332
rect 82004 18292 82005 18332
rect 81963 18283 82005 18292
rect 82443 18332 82485 18341
rect 82443 18292 82444 18332
rect 82484 18292 82485 18332
rect 82443 18283 82485 18292
rect 83211 18332 83253 18341
rect 83211 18292 83212 18332
rect 83252 18292 83253 18332
rect 83211 18283 83253 18292
rect 83595 18332 83637 18341
rect 83595 18292 83596 18332
rect 83636 18292 83637 18332
rect 83595 18283 83637 18292
rect 83979 18332 84021 18341
rect 83979 18292 83980 18332
rect 84020 18292 84021 18332
rect 83979 18283 84021 18292
rect 84459 18332 84501 18341
rect 84459 18292 84460 18332
rect 84500 18292 84501 18332
rect 84459 18283 84501 18292
rect 84843 18332 84885 18341
rect 84843 18292 84844 18332
rect 84884 18292 84885 18332
rect 84843 18283 84885 18292
rect 85131 18332 85173 18341
rect 85131 18292 85132 18332
rect 85172 18292 85173 18332
rect 85131 18283 85173 18292
rect 85707 18332 85749 18341
rect 85707 18292 85708 18332
rect 85748 18292 85749 18332
rect 85707 18283 85749 18292
rect 86091 18332 86133 18341
rect 86091 18292 86092 18332
rect 86132 18292 86133 18332
rect 86091 18283 86133 18292
rect 86379 18332 86421 18341
rect 86379 18292 86380 18332
rect 86420 18292 86421 18332
rect 86379 18283 86421 18292
rect 86763 18332 86805 18341
rect 86763 18292 86764 18332
rect 86804 18292 86805 18332
rect 86763 18283 86805 18292
rect 87243 18332 87285 18341
rect 87243 18292 87244 18332
rect 87284 18292 87285 18332
rect 87243 18283 87285 18292
rect 87915 18332 87957 18341
rect 87915 18292 87916 18332
rect 87956 18292 87957 18332
rect 87915 18283 87957 18292
rect 88395 18332 88437 18341
rect 88395 18292 88396 18332
rect 88436 18292 88437 18332
rect 88395 18283 88437 18292
rect 88779 18332 88821 18341
rect 88779 18292 88780 18332
rect 88820 18292 88821 18332
rect 88779 18283 88821 18292
rect 89163 18332 89205 18341
rect 89163 18292 89164 18332
rect 89204 18292 89205 18332
rect 89163 18283 89205 18292
rect 89547 18332 89589 18341
rect 89547 18292 89548 18332
rect 89588 18292 89589 18332
rect 89547 18283 89589 18292
rect 89931 18332 89973 18341
rect 89931 18292 89932 18332
rect 89972 18292 89973 18332
rect 89931 18283 89973 18292
rect 90315 18332 90357 18341
rect 90315 18292 90316 18332
rect 90356 18292 90357 18332
rect 90315 18283 90357 18292
rect 90795 18332 90837 18341
rect 90795 18292 90796 18332
rect 90836 18292 90837 18332
rect 90795 18283 90837 18292
rect 91467 18332 91509 18341
rect 91467 18292 91468 18332
rect 91508 18292 91509 18332
rect 91467 18283 91509 18292
rect 91659 18332 91701 18341
rect 91659 18292 91660 18332
rect 91700 18292 91701 18332
rect 91659 18283 91701 18292
rect 92043 18332 92085 18341
rect 92043 18292 92044 18332
rect 92084 18292 92085 18332
rect 92043 18283 92085 18292
rect 92427 18332 92469 18341
rect 92427 18292 92428 18332
rect 92468 18292 92469 18332
rect 92427 18283 92469 18292
rect 92811 18332 92853 18341
rect 92811 18292 92812 18332
rect 92852 18292 92853 18332
rect 92811 18283 92853 18292
rect 93291 18332 93333 18341
rect 93291 18292 93292 18332
rect 93332 18292 93333 18332
rect 93291 18283 93333 18292
rect 94059 18332 94101 18341
rect 94059 18292 94060 18332
rect 94100 18292 94101 18332
rect 94059 18283 94101 18292
rect 94443 18332 94485 18341
rect 94443 18292 94444 18332
rect 94484 18292 94485 18332
rect 94443 18283 94485 18292
rect 94731 18332 94773 18341
rect 94731 18292 94732 18332
rect 94772 18292 94773 18332
rect 94731 18283 94773 18292
rect 95211 18332 95253 18341
rect 95211 18292 95212 18332
rect 95252 18292 95253 18332
rect 95211 18283 95253 18292
rect 95691 18332 95733 18341
rect 95691 18292 95692 18332
rect 95732 18292 95733 18332
rect 95691 18283 95733 18292
rect 95883 18332 95925 18341
rect 95883 18292 95884 18332
rect 95924 18292 95925 18332
rect 95883 18283 95925 18292
rect 96459 18332 96501 18341
rect 96459 18292 96460 18332
rect 96500 18292 96501 18332
rect 96459 18283 96501 18292
rect 96843 18332 96885 18341
rect 96843 18292 96844 18332
rect 96884 18292 96885 18332
rect 96843 18283 96885 18292
rect 97323 18332 97365 18341
rect 97323 18292 97324 18332
rect 97364 18292 97365 18332
rect 97323 18283 97365 18292
rect 97515 18332 97557 18341
rect 97515 18292 97516 18332
rect 97556 18292 97557 18332
rect 97515 18283 97557 18292
rect 576 18164 99516 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 7112 18164
rect 7152 18124 7194 18164
rect 7234 18124 7276 18164
rect 7316 18124 7358 18164
rect 7398 18124 7440 18164
rect 7480 18124 11112 18164
rect 11152 18124 11194 18164
rect 11234 18124 11276 18164
rect 11316 18124 11358 18164
rect 11398 18124 11440 18164
rect 11480 18124 15112 18164
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15480 18124 19112 18164
rect 19152 18124 19194 18164
rect 19234 18124 19276 18164
rect 19316 18124 19358 18164
rect 19398 18124 19440 18164
rect 19480 18124 23112 18164
rect 23152 18124 23194 18164
rect 23234 18124 23276 18164
rect 23316 18124 23358 18164
rect 23398 18124 23440 18164
rect 23480 18124 27112 18164
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27480 18124 31112 18164
rect 31152 18124 31194 18164
rect 31234 18124 31276 18164
rect 31316 18124 31358 18164
rect 31398 18124 31440 18164
rect 31480 18124 35112 18164
rect 35152 18124 35194 18164
rect 35234 18124 35276 18164
rect 35316 18124 35358 18164
rect 35398 18124 35440 18164
rect 35480 18124 39112 18164
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39480 18124 43112 18164
rect 43152 18124 43194 18164
rect 43234 18124 43276 18164
rect 43316 18124 43358 18164
rect 43398 18124 43440 18164
rect 43480 18124 47112 18164
rect 47152 18124 47194 18164
rect 47234 18124 47276 18164
rect 47316 18124 47358 18164
rect 47398 18124 47440 18164
rect 47480 18124 51112 18164
rect 51152 18124 51194 18164
rect 51234 18124 51276 18164
rect 51316 18124 51358 18164
rect 51398 18124 51440 18164
rect 51480 18124 55112 18164
rect 55152 18124 55194 18164
rect 55234 18124 55276 18164
rect 55316 18124 55358 18164
rect 55398 18124 55440 18164
rect 55480 18124 59112 18164
rect 59152 18124 59194 18164
rect 59234 18124 59276 18164
rect 59316 18124 59358 18164
rect 59398 18124 59440 18164
rect 59480 18124 63112 18164
rect 63152 18124 63194 18164
rect 63234 18124 63276 18164
rect 63316 18124 63358 18164
rect 63398 18124 63440 18164
rect 63480 18124 67112 18164
rect 67152 18124 67194 18164
rect 67234 18124 67276 18164
rect 67316 18124 67358 18164
rect 67398 18124 67440 18164
rect 67480 18124 71112 18164
rect 71152 18124 71194 18164
rect 71234 18124 71276 18164
rect 71316 18124 71358 18164
rect 71398 18124 71440 18164
rect 71480 18124 75112 18164
rect 75152 18124 75194 18164
rect 75234 18124 75276 18164
rect 75316 18124 75358 18164
rect 75398 18124 75440 18164
rect 75480 18124 79112 18164
rect 79152 18124 79194 18164
rect 79234 18124 79276 18164
rect 79316 18124 79358 18164
rect 79398 18124 79440 18164
rect 79480 18124 83112 18164
rect 83152 18124 83194 18164
rect 83234 18124 83276 18164
rect 83316 18124 83358 18164
rect 83398 18124 83440 18164
rect 83480 18124 87112 18164
rect 87152 18124 87194 18164
rect 87234 18124 87276 18164
rect 87316 18124 87358 18164
rect 87398 18124 87440 18164
rect 87480 18124 91112 18164
rect 91152 18124 91194 18164
rect 91234 18124 91276 18164
rect 91316 18124 91358 18164
rect 91398 18124 91440 18164
rect 91480 18124 95112 18164
rect 95152 18124 95194 18164
rect 95234 18124 95276 18164
rect 95316 18124 95358 18164
rect 95398 18124 95440 18164
rect 95480 18124 99112 18164
rect 99152 18124 99194 18164
rect 99234 18124 99276 18164
rect 99316 18124 99358 18164
rect 99398 18124 99440 18164
rect 99480 18124 99516 18164
rect 576 18100 99516 18124
rect 651 17912 693 17921
rect 651 17872 652 17912
rect 692 17872 693 17912
rect 651 17863 693 17872
rect 98283 17912 98325 17921
rect 98283 17872 98284 17912
rect 98324 17872 98325 17912
rect 98283 17863 98325 17872
rect 73699 17828 73757 17829
rect 73699 17788 73708 17828
rect 73748 17788 73757 17828
rect 73699 17787 73757 17788
rect 74083 17828 74141 17829
rect 74083 17788 74092 17828
rect 74132 17788 74141 17828
rect 74083 17787 74141 17788
rect 74467 17828 74525 17829
rect 74467 17788 74476 17828
rect 74516 17788 74525 17828
rect 74467 17787 74525 17788
rect 75331 17828 75389 17829
rect 75331 17788 75340 17828
rect 75380 17788 75389 17828
rect 75331 17787 75389 17788
rect 76195 17828 76253 17829
rect 76195 17788 76204 17828
rect 76244 17788 76253 17828
rect 76195 17787 76253 17788
rect 76579 17828 76637 17829
rect 76579 17788 76588 17828
rect 76628 17788 76637 17828
rect 76579 17787 76637 17788
rect 76963 17828 77021 17829
rect 76963 17788 76972 17828
rect 77012 17788 77021 17828
rect 76963 17787 77021 17788
rect 77347 17828 77405 17829
rect 77347 17788 77356 17828
rect 77396 17788 77405 17828
rect 77347 17787 77405 17788
rect 78211 17828 78269 17829
rect 78211 17788 78220 17828
rect 78260 17788 78269 17828
rect 78211 17787 78269 17788
rect 78691 17828 78749 17829
rect 78691 17788 78700 17828
rect 78740 17788 78749 17828
rect 78691 17787 78749 17788
rect 80131 17828 80189 17829
rect 80131 17788 80140 17828
rect 80180 17788 80189 17828
rect 80131 17787 80189 17788
rect 80515 17828 80573 17829
rect 80515 17788 80524 17828
rect 80564 17788 80573 17828
rect 80515 17787 80573 17788
rect 82627 17828 82685 17829
rect 82627 17788 82636 17828
rect 82676 17788 82685 17828
rect 82627 17787 82685 17788
rect 84931 17828 84989 17829
rect 84931 17788 84940 17828
rect 84980 17788 84989 17828
rect 84931 17787 84989 17788
rect 86179 17828 86237 17829
rect 86179 17788 86188 17828
rect 86228 17788 86237 17828
rect 86179 17787 86237 17788
rect 89443 17828 89501 17829
rect 89443 17788 89452 17828
rect 89492 17788 89501 17828
rect 89443 17787 89501 17788
rect 93763 17828 93821 17829
rect 93763 17788 93772 17828
rect 93812 17788 93821 17828
rect 93763 17787 93821 17788
rect 95011 17828 95069 17829
rect 95011 17788 95020 17828
rect 95060 17788 95069 17828
rect 95011 17787 95069 17788
rect 95875 17828 95933 17829
rect 95875 17788 95884 17828
rect 95924 17788 95933 17828
rect 95875 17787 95933 17788
rect 96643 17828 96701 17829
rect 96643 17788 96652 17828
rect 96692 17788 96701 17828
rect 96643 17787 96701 17788
rect 97027 17828 97085 17829
rect 97027 17788 97036 17828
rect 97076 17788 97085 17828
rect 97027 17787 97085 17788
rect 97891 17828 97949 17829
rect 97891 17788 97900 17828
rect 97940 17788 97949 17828
rect 97891 17787 97949 17788
rect 98467 17828 98525 17829
rect 98467 17788 98476 17828
rect 98516 17788 98525 17828
rect 98467 17787 98525 17788
rect 93187 17749 93229 17758
rect 75043 17744 75101 17745
rect 75043 17704 75052 17744
rect 75092 17704 75101 17744
rect 75043 17703 75101 17704
rect 75811 17744 75869 17745
rect 75811 17704 75820 17744
rect 75860 17704 75869 17744
rect 75811 17703 75869 17704
rect 77731 17744 77789 17745
rect 77731 17704 77740 17744
rect 77780 17704 77789 17744
rect 77731 17703 77789 17704
rect 79171 17744 79229 17745
rect 79171 17704 79180 17744
rect 79220 17704 79229 17744
rect 79171 17703 79229 17704
rect 79459 17744 79517 17745
rect 79459 17704 79468 17744
rect 79508 17704 79517 17744
rect 79459 17703 79517 17704
rect 79843 17744 79901 17745
rect 79843 17704 79852 17744
rect 79892 17704 79901 17744
rect 79843 17703 79901 17704
rect 80995 17744 81053 17745
rect 80995 17704 81004 17744
rect 81044 17704 81053 17744
rect 80995 17703 81053 17704
rect 81283 17744 81341 17745
rect 81283 17704 81292 17744
rect 81332 17704 81341 17744
rect 81283 17703 81341 17704
rect 81475 17744 81533 17745
rect 81475 17704 81484 17744
rect 81524 17704 81533 17744
rect 81475 17703 81533 17704
rect 81955 17744 82013 17745
rect 81955 17704 81964 17744
rect 82004 17704 82013 17744
rect 81955 17703 82013 17704
rect 82243 17744 82301 17745
rect 82243 17704 82252 17744
rect 82292 17704 82301 17744
rect 82243 17703 82301 17704
rect 83011 17744 83069 17745
rect 83011 17704 83020 17744
rect 83060 17704 83069 17744
rect 83011 17703 83069 17704
rect 83395 17744 83453 17745
rect 83395 17704 83404 17744
rect 83444 17704 83453 17744
rect 83395 17703 83453 17704
rect 83779 17744 83837 17745
rect 83779 17704 83788 17744
rect 83828 17704 83837 17744
rect 83779 17703 83837 17704
rect 84163 17744 84221 17745
rect 84163 17704 84172 17744
rect 84212 17704 84221 17744
rect 84163 17703 84221 17704
rect 84739 17744 84797 17745
rect 84739 17704 84748 17744
rect 84788 17704 84797 17744
rect 84739 17703 84797 17704
rect 85411 17744 85469 17745
rect 85411 17704 85420 17744
rect 85460 17704 85469 17744
rect 85411 17703 85469 17704
rect 85795 17744 85853 17745
rect 85795 17704 85804 17744
rect 85844 17704 85853 17744
rect 85795 17703 85853 17704
rect 86563 17744 86621 17745
rect 86563 17704 86572 17744
rect 86612 17704 86621 17744
rect 86563 17703 86621 17704
rect 87043 17744 87101 17745
rect 87043 17704 87052 17744
rect 87092 17704 87101 17744
rect 87043 17703 87101 17704
rect 87427 17744 87485 17745
rect 87427 17704 87436 17744
rect 87476 17704 87485 17744
rect 87427 17703 87485 17704
rect 88195 17744 88253 17745
rect 88195 17704 88204 17744
rect 88244 17704 88253 17744
rect 88195 17703 88253 17704
rect 88579 17744 88637 17745
rect 88579 17704 88588 17744
rect 88628 17704 88637 17744
rect 88579 17703 88637 17704
rect 89059 17744 89117 17745
rect 89059 17704 89068 17744
rect 89108 17704 89117 17744
rect 89059 17703 89117 17704
rect 89923 17744 89981 17745
rect 89923 17704 89932 17744
rect 89972 17704 89981 17744
rect 89923 17703 89981 17704
rect 90211 17744 90269 17745
rect 90211 17704 90220 17744
rect 90260 17704 90269 17744
rect 90211 17703 90269 17704
rect 90595 17744 90653 17745
rect 90595 17704 90604 17744
rect 90644 17704 90653 17744
rect 90595 17703 90653 17704
rect 90979 17744 91037 17745
rect 90979 17704 90988 17744
rect 91028 17704 91037 17744
rect 90979 17703 91037 17704
rect 91363 17744 91421 17745
rect 91363 17704 91372 17744
rect 91412 17704 91421 17744
rect 91363 17703 91421 17704
rect 91843 17744 91901 17745
rect 91843 17704 91852 17744
rect 91892 17704 91901 17744
rect 91843 17703 91901 17704
rect 92227 17744 92285 17745
rect 92227 17704 92236 17744
rect 92276 17704 92285 17744
rect 92227 17703 92285 17704
rect 92803 17744 92861 17745
rect 92803 17704 92812 17744
rect 92852 17704 92861 17744
rect 92803 17703 92861 17704
rect 93187 17709 93188 17749
rect 93228 17709 93229 17749
rect 93187 17700 93229 17709
rect 94051 17744 94109 17745
rect 94051 17704 94060 17744
rect 94100 17704 94109 17744
rect 94051 17703 94109 17704
rect 94243 17744 94301 17745
rect 94243 17704 94252 17744
rect 94292 17704 94301 17744
rect 94243 17703 94301 17704
rect 94723 17744 94781 17745
rect 94723 17704 94732 17744
rect 94772 17704 94781 17744
rect 94723 17703 94781 17704
rect 95395 17744 95453 17745
rect 95395 17704 95404 17744
rect 95444 17704 95453 17744
rect 95395 17703 95453 17704
rect 96355 17744 96413 17745
rect 96355 17704 96364 17744
rect 96404 17704 96413 17744
rect 96355 17703 96413 17704
rect 97411 17744 97469 17745
rect 97411 17704 97420 17744
rect 97460 17704 97469 17744
rect 97411 17703 97469 17704
rect 98659 17744 98717 17745
rect 98659 17704 98668 17744
rect 98708 17704 98717 17744
rect 98659 17703 98717 17704
rect 81867 17660 81909 17669
rect 81867 17620 81868 17660
rect 81908 17620 81909 17660
rect 81867 17611 81909 17620
rect 84651 17660 84693 17669
rect 84651 17620 84652 17660
rect 84692 17620 84693 17660
rect 84651 17611 84693 17620
rect 92907 17660 92949 17669
rect 92907 17620 92908 17660
rect 92948 17620 92949 17660
rect 92907 17611 92949 17620
rect 98763 17660 98805 17669
rect 98763 17620 98764 17660
rect 98804 17620 98805 17660
rect 98763 17611 98805 17620
rect 73899 17576 73941 17585
rect 73899 17536 73900 17576
rect 73940 17536 73941 17576
rect 73899 17527 73941 17536
rect 74283 17576 74325 17585
rect 74283 17536 74284 17576
rect 74324 17536 74325 17576
rect 74283 17527 74325 17536
rect 74667 17576 74709 17585
rect 74667 17536 74668 17576
rect 74708 17536 74709 17576
rect 74667 17527 74709 17536
rect 75147 17576 75189 17585
rect 75147 17536 75148 17576
rect 75188 17536 75189 17576
rect 75147 17527 75189 17536
rect 75531 17576 75573 17585
rect 75531 17536 75532 17576
rect 75572 17536 75573 17576
rect 75531 17527 75573 17536
rect 75723 17576 75765 17585
rect 75723 17536 75724 17576
rect 75764 17536 75765 17576
rect 75723 17527 75765 17536
rect 76395 17576 76437 17585
rect 76395 17536 76396 17576
rect 76436 17536 76437 17576
rect 76395 17527 76437 17536
rect 76779 17576 76821 17585
rect 76779 17536 76780 17576
rect 76820 17536 76821 17576
rect 76779 17527 76821 17536
rect 77163 17576 77205 17585
rect 77163 17536 77164 17576
rect 77204 17536 77205 17576
rect 77163 17527 77205 17536
rect 77547 17576 77589 17585
rect 77547 17536 77548 17576
rect 77588 17536 77589 17576
rect 77547 17527 77589 17536
rect 77835 17576 77877 17585
rect 77835 17536 77836 17576
rect 77876 17536 77877 17576
rect 77835 17527 77877 17536
rect 78411 17576 78453 17585
rect 78411 17536 78412 17576
rect 78452 17536 78453 17576
rect 78411 17527 78453 17536
rect 78891 17576 78933 17585
rect 78891 17536 78892 17576
rect 78932 17536 78933 17576
rect 78891 17527 78933 17536
rect 79083 17576 79125 17585
rect 79083 17536 79084 17576
rect 79124 17536 79125 17576
rect 79083 17527 79125 17536
rect 79563 17576 79605 17585
rect 79563 17536 79564 17576
rect 79604 17536 79605 17576
rect 79563 17527 79605 17536
rect 79947 17576 79989 17585
rect 79947 17536 79948 17576
rect 79988 17536 79989 17576
rect 79947 17527 79989 17536
rect 80331 17576 80373 17585
rect 80331 17536 80332 17576
rect 80372 17536 80373 17576
rect 80331 17527 80373 17536
rect 80715 17576 80757 17585
rect 80715 17536 80716 17576
rect 80756 17536 80757 17576
rect 80715 17527 80757 17536
rect 80907 17576 80949 17585
rect 80907 17536 80908 17576
rect 80948 17536 80949 17576
rect 80907 17527 80949 17536
rect 81195 17576 81237 17585
rect 81195 17536 81196 17576
rect 81236 17536 81237 17576
rect 81195 17527 81237 17536
rect 81579 17576 81621 17585
rect 81579 17536 81580 17576
rect 81620 17536 81621 17576
rect 81579 17527 81621 17536
rect 82347 17576 82389 17585
rect 82347 17536 82348 17576
rect 82388 17536 82389 17576
rect 82347 17527 82389 17536
rect 82827 17576 82869 17585
rect 82827 17536 82828 17576
rect 82868 17536 82869 17576
rect 82827 17527 82869 17536
rect 83115 17576 83157 17585
rect 83115 17536 83116 17576
rect 83156 17536 83157 17576
rect 83115 17527 83157 17536
rect 83499 17576 83541 17585
rect 83499 17536 83500 17576
rect 83540 17536 83541 17576
rect 83499 17527 83541 17536
rect 83883 17576 83925 17585
rect 83883 17536 83884 17576
rect 83924 17536 83925 17576
rect 83883 17527 83925 17536
rect 84267 17576 84309 17585
rect 84267 17536 84268 17576
rect 84308 17536 84309 17576
rect 84267 17527 84309 17536
rect 85131 17576 85173 17585
rect 85131 17536 85132 17576
rect 85172 17536 85173 17576
rect 85131 17527 85173 17536
rect 85515 17576 85557 17585
rect 85515 17536 85516 17576
rect 85556 17536 85557 17576
rect 85515 17527 85557 17536
rect 85899 17576 85941 17585
rect 85899 17536 85900 17576
rect 85940 17536 85941 17576
rect 85899 17527 85941 17536
rect 86379 17576 86421 17585
rect 86379 17536 86380 17576
rect 86420 17536 86421 17576
rect 86379 17527 86421 17536
rect 86667 17576 86709 17585
rect 86667 17536 86668 17576
rect 86708 17536 86709 17576
rect 86667 17527 86709 17536
rect 87147 17576 87189 17585
rect 87147 17536 87148 17576
rect 87188 17536 87189 17576
rect 87147 17527 87189 17536
rect 87531 17576 87573 17585
rect 87531 17536 87532 17576
rect 87572 17536 87573 17576
rect 87531 17527 87573 17536
rect 88299 17576 88341 17585
rect 88299 17536 88300 17576
rect 88340 17536 88341 17576
rect 88299 17527 88341 17536
rect 88683 17576 88725 17585
rect 88683 17536 88684 17576
rect 88724 17536 88725 17576
rect 88683 17527 88725 17536
rect 89163 17576 89205 17585
rect 89163 17536 89164 17576
rect 89204 17536 89205 17576
rect 89163 17527 89205 17536
rect 89643 17576 89685 17585
rect 89643 17536 89644 17576
rect 89684 17536 89685 17576
rect 89643 17527 89685 17536
rect 89835 17576 89877 17585
rect 89835 17536 89836 17576
rect 89876 17536 89877 17576
rect 89835 17527 89877 17536
rect 90315 17576 90357 17585
rect 90315 17536 90316 17576
rect 90356 17536 90357 17576
rect 90315 17527 90357 17536
rect 90699 17576 90741 17585
rect 90699 17536 90700 17576
rect 90740 17536 90741 17576
rect 90699 17527 90741 17536
rect 91083 17576 91125 17585
rect 91083 17536 91084 17576
rect 91124 17536 91125 17576
rect 91083 17527 91125 17536
rect 91467 17576 91509 17585
rect 91467 17536 91468 17576
rect 91508 17536 91509 17576
rect 91467 17527 91509 17536
rect 91947 17576 91989 17585
rect 91947 17536 91948 17576
rect 91988 17536 91989 17576
rect 91947 17527 91989 17536
rect 92331 17576 92373 17585
rect 92331 17536 92332 17576
rect 92372 17536 92373 17576
rect 92331 17527 92373 17536
rect 93099 17576 93141 17585
rect 93099 17536 93100 17576
rect 93140 17536 93141 17576
rect 93099 17527 93141 17536
rect 93579 17576 93621 17585
rect 93579 17536 93580 17576
rect 93620 17536 93621 17576
rect 93579 17527 93621 17536
rect 93963 17576 94005 17585
rect 93963 17536 93964 17576
rect 94004 17536 94005 17576
rect 93963 17527 94005 17536
rect 94347 17576 94389 17585
rect 94347 17536 94348 17576
rect 94388 17536 94389 17576
rect 94347 17527 94389 17536
rect 94827 17576 94869 17585
rect 94827 17536 94828 17576
rect 94868 17536 94869 17576
rect 94827 17527 94869 17536
rect 95211 17576 95253 17585
rect 95211 17536 95212 17576
rect 95252 17536 95253 17576
rect 95211 17527 95253 17536
rect 95499 17576 95541 17585
rect 95499 17536 95500 17576
rect 95540 17536 95541 17576
rect 95499 17527 95541 17536
rect 96075 17576 96117 17585
rect 96075 17536 96076 17576
rect 96116 17536 96117 17576
rect 96075 17527 96117 17536
rect 96267 17576 96309 17585
rect 96267 17536 96268 17576
rect 96308 17536 96309 17576
rect 96267 17527 96309 17536
rect 96843 17576 96885 17585
rect 96843 17536 96844 17576
rect 96884 17536 96885 17576
rect 96843 17527 96885 17536
rect 97227 17576 97269 17585
rect 97227 17536 97228 17576
rect 97268 17536 97269 17576
rect 97227 17527 97269 17536
rect 97515 17576 97557 17585
rect 97515 17536 97516 17576
rect 97556 17536 97557 17576
rect 97515 17527 97557 17536
rect 97707 17576 97749 17585
rect 97707 17536 97708 17576
rect 97748 17536 97749 17576
rect 97707 17527 97749 17536
rect 576 17408 99360 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 8352 17408
rect 8392 17368 8434 17408
rect 8474 17368 8516 17408
rect 8556 17368 8598 17408
rect 8638 17368 8680 17408
rect 8720 17368 12352 17408
rect 12392 17368 12434 17408
rect 12474 17368 12516 17408
rect 12556 17368 12598 17408
rect 12638 17368 12680 17408
rect 12720 17368 16352 17408
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16720 17368 20352 17408
rect 20392 17368 20434 17408
rect 20474 17368 20516 17408
rect 20556 17368 20598 17408
rect 20638 17368 20680 17408
rect 20720 17368 24352 17408
rect 24392 17368 24434 17408
rect 24474 17368 24516 17408
rect 24556 17368 24598 17408
rect 24638 17368 24680 17408
rect 24720 17368 28352 17408
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28720 17368 32352 17408
rect 32392 17368 32434 17408
rect 32474 17368 32516 17408
rect 32556 17368 32598 17408
rect 32638 17368 32680 17408
rect 32720 17368 36352 17408
rect 36392 17368 36434 17408
rect 36474 17368 36516 17408
rect 36556 17368 36598 17408
rect 36638 17368 36680 17408
rect 36720 17368 40352 17408
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40720 17368 44352 17408
rect 44392 17368 44434 17408
rect 44474 17368 44516 17408
rect 44556 17368 44598 17408
rect 44638 17368 44680 17408
rect 44720 17368 48352 17408
rect 48392 17368 48434 17408
rect 48474 17368 48516 17408
rect 48556 17368 48598 17408
rect 48638 17368 48680 17408
rect 48720 17368 52352 17408
rect 52392 17368 52434 17408
rect 52474 17368 52516 17408
rect 52556 17368 52598 17408
rect 52638 17368 52680 17408
rect 52720 17368 56352 17408
rect 56392 17368 56434 17408
rect 56474 17368 56516 17408
rect 56556 17368 56598 17408
rect 56638 17368 56680 17408
rect 56720 17368 60352 17408
rect 60392 17368 60434 17408
rect 60474 17368 60516 17408
rect 60556 17368 60598 17408
rect 60638 17368 60680 17408
rect 60720 17368 64352 17408
rect 64392 17368 64434 17408
rect 64474 17368 64516 17408
rect 64556 17368 64598 17408
rect 64638 17368 64680 17408
rect 64720 17368 68352 17408
rect 68392 17368 68434 17408
rect 68474 17368 68516 17408
rect 68556 17368 68598 17408
rect 68638 17368 68680 17408
rect 68720 17368 72352 17408
rect 72392 17368 72434 17408
rect 72474 17368 72516 17408
rect 72556 17368 72598 17408
rect 72638 17368 72680 17408
rect 72720 17368 76352 17408
rect 76392 17368 76434 17408
rect 76474 17368 76516 17408
rect 76556 17368 76598 17408
rect 76638 17368 76680 17408
rect 76720 17368 80352 17408
rect 80392 17368 80434 17408
rect 80474 17368 80516 17408
rect 80556 17368 80598 17408
rect 80638 17368 80680 17408
rect 80720 17368 84352 17408
rect 84392 17368 84434 17408
rect 84474 17368 84516 17408
rect 84556 17368 84598 17408
rect 84638 17368 84680 17408
rect 84720 17368 88352 17408
rect 88392 17368 88434 17408
rect 88474 17368 88516 17408
rect 88556 17368 88598 17408
rect 88638 17368 88680 17408
rect 88720 17368 92352 17408
rect 92392 17368 92434 17408
rect 92474 17368 92516 17408
rect 92556 17368 92598 17408
rect 92638 17368 92680 17408
rect 92720 17368 96352 17408
rect 96392 17368 96434 17408
rect 96474 17368 96516 17408
rect 96556 17368 96598 17408
rect 96638 17368 96680 17408
rect 96720 17368 99360 17408
rect 576 17344 99360 17368
rect 651 16904 693 16913
rect 651 16864 652 16904
rect 692 16864 693 16904
rect 651 16855 693 16864
rect 576 16652 69984 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 7112 16652
rect 7152 16612 7194 16652
rect 7234 16612 7276 16652
rect 7316 16612 7358 16652
rect 7398 16612 7440 16652
rect 7480 16612 11112 16652
rect 11152 16612 11194 16652
rect 11234 16612 11276 16652
rect 11316 16612 11358 16652
rect 11398 16612 11440 16652
rect 11480 16612 15112 16652
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15480 16612 19112 16652
rect 19152 16612 19194 16652
rect 19234 16612 19276 16652
rect 19316 16612 19358 16652
rect 19398 16612 19440 16652
rect 19480 16612 23112 16652
rect 23152 16612 23194 16652
rect 23234 16612 23276 16652
rect 23316 16612 23358 16652
rect 23398 16612 23440 16652
rect 23480 16612 27112 16652
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27480 16612 31112 16652
rect 31152 16612 31194 16652
rect 31234 16612 31276 16652
rect 31316 16612 31358 16652
rect 31398 16612 31440 16652
rect 31480 16612 35112 16652
rect 35152 16612 35194 16652
rect 35234 16612 35276 16652
rect 35316 16612 35358 16652
rect 35398 16612 35440 16652
rect 35480 16612 39112 16652
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39480 16612 43112 16652
rect 43152 16612 43194 16652
rect 43234 16612 43276 16652
rect 43316 16612 43358 16652
rect 43398 16612 43440 16652
rect 43480 16612 47112 16652
rect 47152 16612 47194 16652
rect 47234 16612 47276 16652
rect 47316 16612 47358 16652
rect 47398 16612 47440 16652
rect 47480 16612 51112 16652
rect 51152 16612 51194 16652
rect 51234 16612 51276 16652
rect 51316 16612 51358 16652
rect 51398 16612 51440 16652
rect 51480 16612 55112 16652
rect 55152 16612 55194 16652
rect 55234 16612 55276 16652
rect 55316 16612 55358 16652
rect 55398 16612 55440 16652
rect 55480 16612 59112 16652
rect 59152 16612 59194 16652
rect 59234 16612 59276 16652
rect 59316 16612 59358 16652
rect 59398 16612 59440 16652
rect 59480 16612 63112 16652
rect 63152 16612 63194 16652
rect 63234 16612 63276 16652
rect 63316 16612 63358 16652
rect 63398 16612 63440 16652
rect 63480 16612 67112 16652
rect 67152 16612 67194 16652
rect 67234 16612 67276 16652
rect 67316 16612 67358 16652
rect 67398 16612 67440 16652
rect 67480 16612 69984 16652
rect 576 16588 69984 16612
rect 651 16400 693 16409
rect 651 16360 652 16400
rect 692 16360 693 16400
rect 651 16351 693 16360
rect 69091 16316 69149 16317
rect 69091 16276 69100 16316
rect 69140 16276 69149 16316
rect 69091 16275 69149 16276
rect 69291 16064 69333 16073
rect 69291 16024 69292 16064
rect 69332 16024 69333 16064
rect 69291 16015 69333 16024
rect 576 15896 69984 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 8352 15896
rect 8392 15856 8434 15896
rect 8474 15856 8516 15896
rect 8556 15856 8598 15896
rect 8638 15856 8680 15896
rect 8720 15856 12352 15896
rect 12392 15856 12434 15896
rect 12474 15856 12516 15896
rect 12556 15856 12598 15896
rect 12638 15856 12680 15896
rect 12720 15856 16352 15896
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16720 15856 20352 15896
rect 20392 15856 20434 15896
rect 20474 15856 20516 15896
rect 20556 15856 20598 15896
rect 20638 15856 20680 15896
rect 20720 15856 24352 15896
rect 24392 15856 24434 15896
rect 24474 15856 24516 15896
rect 24556 15856 24598 15896
rect 24638 15856 24680 15896
rect 24720 15856 28352 15896
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28720 15856 32352 15896
rect 32392 15856 32434 15896
rect 32474 15856 32516 15896
rect 32556 15856 32598 15896
rect 32638 15856 32680 15896
rect 32720 15856 36352 15896
rect 36392 15856 36434 15896
rect 36474 15856 36516 15896
rect 36556 15856 36598 15896
rect 36638 15856 36680 15896
rect 36720 15856 40352 15896
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40720 15856 44352 15896
rect 44392 15856 44434 15896
rect 44474 15856 44516 15896
rect 44556 15856 44598 15896
rect 44638 15856 44680 15896
rect 44720 15856 48352 15896
rect 48392 15856 48434 15896
rect 48474 15856 48516 15896
rect 48556 15856 48598 15896
rect 48638 15856 48680 15896
rect 48720 15856 52352 15896
rect 52392 15856 52434 15896
rect 52474 15856 52516 15896
rect 52556 15856 52598 15896
rect 52638 15856 52680 15896
rect 52720 15856 56352 15896
rect 56392 15856 56434 15896
rect 56474 15856 56516 15896
rect 56556 15856 56598 15896
rect 56638 15856 56680 15896
rect 56720 15856 60352 15896
rect 60392 15856 60434 15896
rect 60474 15856 60516 15896
rect 60556 15856 60598 15896
rect 60638 15856 60680 15896
rect 60720 15856 64352 15896
rect 64392 15856 64434 15896
rect 64474 15856 64516 15896
rect 64556 15856 64598 15896
rect 64638 15856 64680 15896
rect 64720 15856 68352 15896
rect 68392 15856 68434 15896
rect 68474 15856 68516 15896
rect 68556 15856 68598 15896
rect 68638 15856 68680 15896
rect 68720 15856 69984 15896
rect 576 15832 69984 15856
rect 67371 15728 67413 15737
rect 67371 15688 67372 15728
rect 67412 15688 67413 15728
rect 67371 15679 67413 15688
rect 68227 15560 68285 15561
rect 68227 15520 68236 15560
rect 68276 15520 68285 15560
rect 68227 15519 68285 15520
rect 68419 15560 68477 15561
rect 68419 15520 68428 15560
rect 68468 15520 68477 15560
rect 68419 15519 68477 15520
rect 835 15476 893 15477
rect 835 15436 844 15476
rect 884 15436 893 15476
rect 835 15435 893 15436
rect 1987 15476 2045 15477
rect 1987 15436 1996 15476
rect 2036 15436 2045 15476
rect 1987 15435 2045 15436
rect 67171 15476 67229 15477
rect 67171 15436 67180 15476
rect 67220 15436 67229 15476
rect 67171 15435 67229 15436
rect 67747 15476 67805 15477
rect 67747 15436 67756 15476
rect 67796 15436 67805 15476
rect 67747 15435 67805 15436
rect 67563 15392 67605 15401
rect 67563 15352 67564 15392
rect 67604 15352 67605 15392
rect 67563 15343 67605 15352
rect 651 15308 693 15317
rect 651 15268 652 15308
rect 692 15268 693 15308
rect 651 15259 693 15268
rect 1803 15308 1845 15317
rect 1803 15268 1804 15308
rect 1844 15268 1845 15308
rect 1803 15259 1845 15268
rect 576 15140 69984 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 7112 15140
rect 7152 15100 7194 15140
rect 7234 15100 7276 15140
rect 7316 15100 7358 15140
rect 7398 15100 7440 15140
rect 7480 15100 11112 15140
rect 11152 15100 11194 15140
rect 11234 15100 11276 15140
rect 11316 15100 11358 15140
rect 11398 15100 11440 15140
rect 11480 15100 15112 15140
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15480 15100 19112 15140
rect 19152 15100 19194 15140
rect 19234 15100 19276 15140
rect 19316 15100 19358 15140
rect 19398 15100 19440 15140
rect 19480 15100 23112 15140
rect 23152 15100 23194 15140
rect 23234 15100 23276 15140
rect 23316 15100 23358 15140
rect 23398 15100 23440 15140
rect 23480 15100 27112 15140
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27480 15100 31112 15140
rect 31152 15100 31194 15140
rect 31234 15100 31276 15140
rect 31316 15100 31358 15140
rect 31398 15100 31440 15140
rect 31480 15100 35112 15140
rect 35152 15100 35194 15140
rect 35234 15100 35276 15140
rect 35316 15100 35358 15140
rect 35398 15100 35440 15140
rect 35480 15100 39112 15140
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39480 15100 43112 15140
rect 43152 15100 43194 15140
rect 43234 15100 43276 15140
rect 43316 15100 43358 15140
rect 43398 15100 43440 15140
rect 43480 15100 47112 15140
rect 47152 15100 47194 15140
rect 47234 15100 47276 15140
rect 47316 15100 47358 15140
rect 47398 15100 47440 15140
rect 47480 15100 51112 15140
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51480 15100 55112 15140
rect 55152 15100 55194 15140
rect 55234 15100 55276 15140
rect 55316 15100 55358 15140
rect 55398 15100 55440 15140
rect 55480 15100 59112 15140
rect 59152 15100 59194 15140
rect 59234 15100 59276 15140
rect 59316 15100 59358 15140
rect 59398 15100 59440 15140
rect 59480 15100 63112 15140
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63480 15100 67112 15140
rect 67152 15100 67194 15140
rect 67234 15100 67276 15140
rect 67316 15100 67358 15140
rect 67398 15100 67440 15140
rect 67480 15100 69984 15140
rect 576 15076 69984 15100
rect 1707 14972 1749 14981
rect 1707 14932 1708 14972
rect 1748 14932 1749 14972
rect 1707 14923 1749 14932
rect 68715 14972 68757 14981
rect 68715 14932 68716 14972
rect 68756 14932 68757 14972
rect 68715 14923 68757 14932
rect 69099 14972 69141 14981
rect 69099 14932 69100 14972
rect 69140 14932 69141 14972
rect 69099 14923 69141 14932
rect 69483 14972 69525 14981
rect 69483 14932 69484 14972
rect 69524 14932 69525 14972
rect 69483 14923 69525 14932
rect 69867 14972 69909 14981
rect 69867 14932 69868 14972
rect 69908 14932 69909 14972
rect 69867 14923 69909 14932
rect 835 14804 893 14805
rect 835 14764 844 14804
rect 884 14764 893 14804
rect 835 14763 893 14764
rect 1891 14804 1949 14805
rect 1891 14764 1900 14804
rect 1940 14764 1949 14804
rect 1891 14763 1949 14764
rect 68043 14804 68085 14813
rect 68043 14764 68044 14804
rect 68084 14764 68085 14804
rect 68043 14755 68085 14764
rect 69667 14804 69725 14805
rect 69667 14764 69676 14804
rect 69716 14764 69725 14804
rect 69667 14763 69725 14764
rect 68131 14720 68189 14721
rect 68131 14680 68140 14720
rect 68180 14680 68189 14720
rect 68131 14679 68189 14680
rect 68611 14720 68669 14721
rect 68611 14680 68620 14720
rect 68660 14680 68669 14720
rect 68611 14679 68669 14680
rect 68995 14720 69053 14721
rect 68995 14680 69004 14720
rect 69044 14680 69053 14720
rect 68995 14679 69053 14680
rect 69379 14720 69437 14721
rect 69379 14680 69388 14720
rect 69428 14680 69437 14720
rect 69379 14679 69437 14680
rect 651 14552 693 14561
rect 651 14512 652 14552
rect 692 14512 693 14552
rect 651 14503 693 14512
rect 576 14384 69984 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 8352 14384
rect 8392 14344 8434 14384
rect 8474 14344 8516 14384
rect 8556 14344 8598 14384
rect 8638 14344 8680 14384
rect 8720 14344 12352 14384
rect 12392 14344 12434 14384
rect 12474 14344 12516 14384
rect 12556 14344 12598 14384
rect 12638 14344 12680 14384
rect 12720 14344 16352 14384
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16720 14344 20352 14384
rect 20392 14344 20434 14384
rect 20474 14344 20516 14384
rect 20556 14344 20598 14384
rect 20638 14344 20680 14384
rect 20720 14344 24352 14384
rect 24392 14344 24434 14384
rect 24474 14344 24516 14384
rect 24556 14344 24598 14384
rect 24638 14344 24680 14384
rect 24720 14344 28352 14384
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28720 14344 32352 14384
rect 32392 14344 32434 14384
rect 32474 14344 32516 14384
rect 32556 14344 32598 14384
rect 32638 14344 32680 14384
rect 32720 14344 36352 14384
rect 36392 14344 36434 14384
rect 36474 14344 36516 14384
rect 36556 14344 36598 14384
rect 36638 14344 36680 14384
rect 36720 14344 40352 14384
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40720 14344 44352 14384
rect 44392 14344 44434 14384
rect 44474 14344 44516 14384
rect 44556 14344 44598 14384
rect 44638 14344 44680 14384
rect 44720 14344 48352 14384
rect 48392 14344 48434 14384
rect 48474 14344 48516 14384
rect 48556 14344 48598 14384
rect 48638 14344 48680 14384
rect 48720 14344 52352 14384
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52720 14344 56352 14384
rect 56392 14344 56434 14384
rect 56474 14344 56516 14384
rect 56556 14344 56598 14384
rect 56638 14344 56680 14384
rect 56720 14344 60352 14384
rect 60392 14344 60434 14384
rect 60474 14344 60516 14384
rect 60556 14344 60598 14384
rect 60638 14344 60680 14384
rect 60720 14344 64352 14384
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64720 14344 68352 14384
rect 68392 14344 68434 14384
rect 68474 14344 68516 14384
rect 68556 14344 68598 14384
rect 68638 14344 68680 14384
rect 68720 14344 69984 14384
rect 576 14320 69984 14344
rect 1323 14216 1365 14225
rect 1323 14176 1324 14216
rect 1364 14176 1365 14216
rect 1323 14167 1365 14176
rect 69387 14216 69429 14225
rect 69387 14176 69388 14216
rect 69428 14176 69429 14216
rect 69387 14167 69429 14176
rect 69867 14216 69909 14225
rect 69867 14176 69868 14216
rect 69908 14176 69909 14216
rect 69867 14167 69909 14176
rect 69763 14048 69821 14049
rect 69763 14008 69772 14048
rect 69812 14008 69821 14048
rect 69763 14007 69821 14008
rect 1507 13964 1565 13965
rect 1507 13924 1516 13964
rect 1556 13924 1565 13964
rect 1507 13923 1565 13924
rect 69187 13964 69245 13965
rect 69187 13924 69196 13964
rect 69236 13924 69245 13964
rect 69187 13923 69245 13924
rect 576 13628 69984 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 7112 13628
rect 7152 13588 7194 13628
rect 7234 13588 7276 13628
rect 7316 13588 7358 13628
rect 7398 13588 7440 13628
rect 7480 13588 11112 13628
rect 11152 13588 11194 13628
rect 11234 13588 11276 13628
rect 11316 13588 11358 13628
rect 11398 13588 11440 13628
rect 11480 13588 15112 13628
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15480 13588 19112 13628
rect 19152 13588 19194 13628
rect 19234 13588 19276 13628
rect 19316 13588 19358 13628
rect 19398 13588 19440 13628
rect 19480 13588 23112 13628
rect 23152 13588 23194 13628
rect 23234 13588 23276 13628
rect 23316 13588 23358 13628
rect 23398 13588 23440 13628
rect 23480 13588 27112 13628
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27480 13588 31112 13628
rect 31152 13588 31194 13628
rect 31234 13588 31276 13628
rect 31316 13588 31358 13628
rect 31398 13588 31440 13628
rect 31480 13588 35112 13628
rect 35152 13588 35194 13628
rect 35234 13588 35276 13628
rect 35316 13588 35358 13628
rect 35398 13588 35440 13628
rect 35480 13588 39112 13628
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39480 13588 43112 13628
rect 43152 13588 43194 13628
rect 43234 13588 43276 13628
rect 43316 13588 43358 13628
rect 43398 13588 43440 13628
rect 43480 13588 47112 13628
rect 47152 13588 47194 13628
rect 47234 13588 47276 13628
rect 47316 13588 47358 13628
rect 47398 13588 47440 13628
rect 47480 13588 51112 13628
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51480 13588 55112 13628
rect 55152 13588 55194 13628
rect 55234 13588 55276 13628
rect 55316 13588 55358 13628
rect 55398 13588 55440 13628
rect 55480 13588 59112 13628
rect 59152 13588 59194 13628
rect 59234 13588 59276 13628
rect 59316 13588 59358 13628
rect 59398 13588 59440 13628
rect 59480 13588 63112 13628
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63480 13588 67112 13628
rect 67152 13588 67194 13628
rect 67234 13588 67276 13628
rect 67316 13588 67358 13628
rect 67398 13588 67440 13628
rect 67480 13588 69984 13628
rect 576 13564 69984 13588
rect 1707 13376 1749 13385
rect 1707 13336 1708 13376
rect 1748 13336 1749 13376
rect 1707 13327 1749 13336
rect 835 13292 893 13293
rect 835 13252 844 13292
rect 884 13252 893 13292
rect 835 13251 893 13252
rect 1891 13292 1949 13293
rect 1891 13252 1900 13292
rect 1940 13252 1949 13292
rect 1891 13251 1949 13252
rect 651 13040 693 13049
rect 651 13000 652 13040
rect 692 13000 693 13040
rect 651 12991 693 13000
rect 576 12872 69984 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 8352 12872
rect 8392 12832 8434 12872
rect 8474 12832 8516 12872
rect 8556 12832 8598 12872
rect 8638 12832 8680 12872
rect 8720 12832 12352 12872
rect 12392 12832 12434 12872
rect 12474 12832 12516 12872
rect 12556 12832 12598 12872
rect 12638 12832 12680 12872
rect 12720 12832 16352 12872
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16720 12832 20352 12872
rect 20392 12832 20434 12872
rect 20474 12832 20516 12872
rect 20556 12832 20598 12872
rect 20638 12832 20680 12872
rect 20720 12832 24352 12872
rect 24392 12832 24434 12872
rect 24474 12832 24516 12872
rect 24556 12832 24598 12872
rect 24638 12832 24680 12872
rect 24720 12832 28352 12872
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28720 12832 32352 12872
rect 32392 12832 32434 12872
rect 32474 12832 32516 12872
rect 32556 12832 32598 12872
rect 32638 12832 32680 12872
rect 32720 12832 36352 12872
rect 36392 12832 36434 12872
rect 36474 12832 36516 12872
rect 36556 12832 36598 12872
rect 36638 12832 36680 12872
rect 36720 12832 40352 12872
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40720 12832 44352 12872
rect 44392 12832 44434 12872
rect 44474 12832 44516 12872
rect 44556 12832 44598 12872
rect 44638 12832 44680 12872
rect 44720 12832 48352 12872
rect 48392 12832 48434 12872
rect 48474 12832 48516 12872
rect 48556 12832 48598 12872
rect 48638 12832 48680 12872
rect 48720 12832 52352 12872
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52720 12832 56352 12872
rect 56392 12832 56434 12872
rect 56474 12832 56516 12872
rect 56556 12832 56598 12872
rect 56638 12832 56680 12872
rect 56720 12832 60352 12872
rect 60392 12832 60434 12872
rect 60474 12832 60516 12872
rect 60556 12832 60598 12872
rect 60638 12832 60680 12872
rect 60720 12832 64352 12872
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64720 12832 68352 12872
rect 68392 12832 68434 12872
rect 68474 12832 68516 12872
rect 68556 12832 68598 12872
rect 68638 12832 68680 12872
rect 68720 12832 69984 12872
rect 576 12808 69984 12832
rect 835 12452 893 12453
rect 835 12412 844 12452
rect 884 12412 893 12452
rect 835 12411 893 12412
rect 1795 12452 1853 12453
rect 1795 12412 1804 12452
rect 1844 12412 1853 12452
rect 1795 12411 1853 12412
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 1611 12284 1653 12293
rect 1611 12244 1612 12284
rect 1652 12244 1653 12284
rect 1611 12235 1653 12244
rect 576 12116 69984 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 7112 12116
rect 7152 12076 7194 12116
rect 7234 12076 7276 12116
rect 7316 12076 7358 12116
rect 7398 12076 7440 12116
rect 7480 12076 11112 12116
rect 11152 12076 11194 12116
rect 11234 12076 11276 12116
rect 11316 12076 11358 12116
rect 11398 12076 11440 12116
rect 11480 12076 15112 12116
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15480 12076 19112 12116
rect 19152 12076 19194 12116
rect 19234 12076 19276 12116
rect 19316 12076 19358 12116
rect 19398 12076 19440 12116
rect 19480 12076 23112 12116
rect 23152 12076 23194 12116
rect 23234 12076 23276 12116
rect 23316 12076 23358 12116
rect 23398 12076 23440 12116
rect 23480 12076 27112 12116
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27480 12076 31112 12116
rect 31152 12076 31194 12116
rect 31234 12076 31276 12116
rect 31316 12076 31358 12116
rect 31398 12076 31440 12116
rect 31480 12076 35112 12116
rect 35152 12076 35194 12116
rect 35234 12076 35276 12116
rect 35316 12076 35358 12116
rect 35398 12076 35440 12116
rect 35480 12076 39112 12116
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39480 12076 43112 12116
rect 43152 12076 43194 12116
rect 43234 12076 43276 12116
rect 43316 12076 43358 12116
rect 43398 12076 43440 12116
rect 43480 12076 47112 12116
rect 47152 12076 47194 12116
rect 47234 12076 47276 12116
rect 47316 12076 47358 12116
rect 47398 12076 47440 12116
rect 47480 12076 51112 12116
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51480 12076 55112 12116
rect 55152 12076 55194 12116
rect 55234 12076 55276 12116
rect 55316 12076 55358 12116
rect 55398 12076 55440 12116
rect 55480 12076 59112 12116
rect 59152 12076 59194 12116
rect 59234 12076 59276 12116
rect 59316 12076 59358 12116
rect 59398 12076 59440 12116
rect 59480 12076 63112 12116
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63480 12076 67112 12116
rect 67152 12076 67194 12116
rect 67234 12076 67276 12116
rect 67316 12076 67358 12116
rect 67398 12076 67440 12116
rect 67480 12076 69984 12116
rect 576 12052 69984 12076
rect 1995 11948 2037 11957
rect 1995 11908 1996 11948
rect 2036 11908 2037 11948
rect 1995 11899 2037 11908
rect 835 11780 893 11781
rect 835 11740 844 11780
rect 884 11740 893 11780
rect 835 11739 893 11740
rect 2179 11780 2237 11781
rect 2179 11740 2188 11780
rect 2228 11740 2237 11780
rect 2179 11739 2237 11740
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 576 11360 69984 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 8352 11360
rect 8392 11320 8434 11360
rect 8474 11320 8516 11360
rect 8556 11320 8598 11360
rect 8638 11320 8680 11360
rect 8720 11320 12352 11360
rect 12392 11320 12434 11360
rect 12474 11320 12516 11360
rect 12556 11320 12598 11360
rect 12638 11320 12680 11360
rect 12720 11320 16352 11360
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16720 11320 20352 11360
rect 20392 11320 20434 11360
rect 20474 11320 20516 11360
rect 20556 11320 20598 11360
rect 20638 11320 20680 11360
rect 20720 11320 24352 11360
rect 24392 11320 24434 11360
rect 24474 11320 24516 11360
rect 24556 11320 24598 11360
rect 24638 11320 24680 11360
rect 24720 11320 28352 11360
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28720 11320 32352 11360
rect 32392 11320 32434 11360
rect 32474 11320 32516 11360
rect 32556 11320 32598 11360
rect 32638 11320 32680 11360
rect 32720 11320 36352 11360
rect 36392 11320 36434 11360
rect 36474 11320 36516 11360
rect 36556 11320 36598 11360
rect 36638 11320 36680 11360
rect 36720 11320 40352 11360
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40720 11320 44352 11360
rect 44392 11320 44434 11360
rect 44474 11320 44516 11360
rect 44556 11320 44598 11360
rect 44638 11320 44680 11360
rect 44720 11320 48352 11360
rect 48392 11320 48434 11360
rect 48474 11320 48516 11360
rect 48556 11320 48598 11360
rect 48638 11320 48680 11360
rect 48720 11320 52352 11360
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52720 11320 56352 11360
rect 56392 11320 56434 11360
rect 56474 11320 56516 11360
rect 56556 11320 56598 11360
rect 56638 11320 56680 11360
rect 56720 11320 60352 11360
rect 60392 11320 60434 11360
rect 60474 11320 60516 11360
rect 60556 11320 60598 11360
rect 60638 11320 60680 11360
rect 60720 11320 64352 11360
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64720 11320 68352 11360
rect 68392 11320 68434 11360
rect 68474 11320 68516 11360
rect 68556 11320 68598 11360
rect 68638 11320 68680 11360
rect 68720 11320 69984 11360
rect 576 11296 69984 11320
rect 69763 11024 69821 11025
rect 69763 10984 69772 11024
rect 69812 10984 69821 11024
rect 69763 10983 69821 10984
rect 835 10940 893 10941
rect 835 10900 844 10940
rect 884 10900 893 10940
rect 835 10899 893 10900
rect 1603 10940 1661 10941
rect 1603 10900 1612 10940
rect 1652 10900 1661 10940
rect 1603 10899 1661 10900
rect 69283 10940 69341 10941
rect 69283 10900 69292 10940
rect 69332 10900 69341 10940
rect 69283 10899 69341 10900
rect 1419 10856 1461 10865
rect 1419 10816 1420 10856
rect 1460 10816 1461 10856
rect 1419 10807 1461 10816
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 69483 10772 69525 10781
rect 69483 10732 69484 10772
rect 69524 10732 69525 10772
rect 69483 10723 69525 10732
rect 69867 10772 69909 10781
rect 69867 10732 69868 10772
rect 69908 10732 69909 10772
rect 69867 10723 69909 10732
rect 576 10604 69984 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 7112 10604
rect 7152 10564 7194 10604
rect 7234 10564 7276 10604
rect 7316 10564 7358 10604
rect 7398 10564 7440 10604
rect 7480 10564 11112 10604
rect 11152 10564 11194 10604
rect 11234 10564 11276 10604
rect 11316 10564 11358 10604
rect 11398 10564 11440 10604
rect 11480 10564 15112 10604
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15480 10564 19112 10604
rect 19152 10564 19194 10604
rect 19234 10564 19276 10604
rect 19316 10564 19358 10604
rect 19398 10564 19440 10604
rect 19480 10564 23112 10604
rect 23152 10564 23194 10604
rect 23234 10564 23276 10604
rect 23316 10564 23358 10604
rect 23398 10564 23440 10604
rect 23480 10564 27112 10604
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27480 10564 31112 10604
rect 31152 10564 31194 10604
rect 31234 10564 31276 10604
rect 31316 10564 31358 10604
rect 31398 10564 31440 10604
rect 31480 10564 35112 10604
rect 35152 10564 35194 10604
rect 35234 10564 35276 10604
rect 35316 10564 35358 10604
rect 35398 10564 35440 10604
rect 35480 10564 39112 10604
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39480 10564 43112 10604
rect 43152 10564 43194 10604
rect 43234 10564 43276 10604
rect 43316 10564 43358 10604
rect 43398 10564 43440 10604
rect 43480 10564 47112 10604
rect 47152 10564 47194 10604
rect 47234 10564 47276 10604
rect 47316 10564 47358 10604
rect 47398 10564 47440 10604
rect 47480 10564 51112 10604
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51480 10564 55112 10604
rect 55152 10564 55194 10604
rect 55234 10564 55276 10604
rect 55316 10564 55358 10604
rect 55398 10564 55440 10604
rect 55480 10564 59112 10604
rect 59152 10564 59194 10604
rect 59234 10564 59276 10604
rect 59316 10564 59358 10604
rect 59398 10564 59440 10604
rect 59480 10564 63112 10604
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63480 10564 67112 10604
rect 67152 10564 67194 10604
rect 67234 10564 67276 10604
rect 67316 10564 67358 10604
rect 67398 10564 67440 10604
rect 67480 10564 69984 10604
rect 576 10540 69984 10564
rect 1323 10352 1365 10361
rect 1323 10312 1324 10352
rect 1364 10312 1365 10352
rect 1323 10303 1365 10312
rect 67659 10352 67701 10361
rect 67659 10312 67660 10352
rect 67700 10312 67701 10352
rect 67659 10303 67701 10312
rect 69195 10352 69237 10361
rect 69195 10312 69196 10352
rect 69236 10312 69237 10352
rect 69195 10303 69237 10312
rect 835 10268 893 10269
rect 835 10228 844 10268
rect 884 10228 893 10268
rect 835 10227 893 10228
rect 1507 10268 1565 10269
rect 1507 10228 1516 10268
rect 1556 10228 1565 10268
rect 1507 10227 1565 10228
rect 67459 10268 67517 10269
rect 67459 10228 67468 10268
rect 67508 10228 67517 10268
rect 67459 10227 67517 10228
rect 68995 10268 69053 10269
rect 68995 10228 69004 10268
rect 69044 10228 69053 10268
rect 68995 10227 69053 10228
rect 68323 10184 68381 10185
rect 68323 10144 68332 10184
rect 68372 10144 68381 10184
rect 68323 10143 68381 10144
rect 68515 10184 68573 10185
rect 68515 10144 68524 10184
rect 68564 10144 68573 10184
rect 68515 10143 68573 10144
rect 68707 10184 68765 10185
rect 68707 10144 68716 10184
rect 68756 10144 68765 10184
rect 68707 10143 68765 10144
rect 69379 10184 69437 10185
rect 69379 10144 69388 10184
rect 69428 10144 69437 10184
rect 69379 10143 69437 10144
rect 69667 10184 69725 10185
rect 69667 10144 69676 10184
rect 69716 10144 69725 10184
rect 69667 10143 69725 10144
rect 68235 10100 68277 10109
rect 68235 10060 68236 10100
rect 68276 10060 68277 10100
rect 68235 10051 68277 10060
rect 69483 10100 69525 10109
rect 69483 10060 69484 10100
rect 69524 10060 69525 10100
rect 69483 10051 69525 10060
rect 69771 10100 69813 10109
rect 69771 10060 69772 10100
rect 69812 10060 69813 10100
rect 69771 10051 69813 10060
rect 651 10016 693 10025
rect 651 9976 652 10016
rect 692 9976 693 10016
rect 651 9967 693 9976
rect 576 9848 69984 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 8352 9848
rect 8392 9808 8434 9848
rect 8474 9808 8516 9848
rect 8556 9808 8598 9848
rect 8638 9808 8680 9848
rect 8720 9808 12352 9848
rect 12392 9808 12434 9848
rect 12474 9808 12516 9848
rect 12556 9808 12598 9848
rect 12638 9808 12680 9848
rect 12720 9808 16352 9848
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16720 9808 20352 9848
rect 20392 9808 20434 9848
rect 20474 9808 20516 9848
rect 20556 9808 20598 9848
rect 20638 9808 20680 9848
rect 20720 9808 24352 9848
rect 24392 9808 24434 9848
rect 24474 9808 24516 9848
rect 24556 9808 24598 9848
rect 24638 9808 24680 9848
rect 24720 9808 28352 9848
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28720 9808 32352 9848
rect 32392 9808 32434 9848
rect 32474 9808 32516 9848
rect 32556 9808 32598 9848
rect 32638 9808 32680 9848
rect 32720 9808 36352 9848
rect 36392 9808 36434 9848
rect 36474 9808 36516 9848
rect 36556 9808 36598 9848
rect 36638 9808 36680 9848
rect 36720 9808 40352 9848
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40720 9808 44352 9848
rect 44392 9808 44434 9848
rect 44474 9808 44516 9848
rect 44556 9808 44598 9848
rect 44638 9808 44680 9848
rect 44720 9808 48352 9848
rect 48392 9808 48434 9848
rect 48474 9808 48516 9848
rect 48556 9808 48598 9848
rect 48638 9808 48680 9848
rect 48720 9808 52352 9848
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52720 9808 56352 9848
rect 56392 9808 56434 9848
rect 56474 9808 56516 9848
rect 56556 9808 56598 9848
rect 56638 9808 56680 9848
rect 56720 9808 60352 9848
rect 60392 9808 60434 9848
rect 60474 9808 60516 9848
rect 60556 9808 60598 9848
rect 60638 9808 60680 9848
rect 60720 9808 64352 9848
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64720 9808 68352 9848
rect 68392 9808 68434 9848
rect 68474 9808 68516 9848
rect 68556 9808 68598 9848
rect 68638 9808 68680 9848
rect 68720 9808 69984 9848
rect 576 9784 69984 9808
rect 69579 9680 69621 9689
rect 69579 9640 69580 9680
rect 69620 9640 69621 9680
rect 69579 9631 69621 9640
rect 69867 9680 69909 9689
rect 69867 9640 69868 9680
rect 69908 9640 69909 9680
rect 69867 9631 69909 9640
rect 69763 9512 69821 9513
rect 69763 9472 69772 9512
rect 69812 9472 69821 9512
rect 69763 9471 69821 9472
rect 835 9428 893 9429
rect 835 9388 844 9428
rect 884 9388 893 9428
rect 835 9387 893 9388
rect 1507 9428 1565 9429
rect 1507 9388 1516 9428
rect 1556 9388 1565 9428
rect 1507 9387 1565 9388
rect 68995 9428 69053 9429
rect 68995 9388 69004 9428
rect 69044 9388 69053 9428
rect 68995 9387 69053 9388
rect 69379 9428 69437 9429
rect 69379 9388 69388 9428
rect 69428 9388 69437 9428
rect 69379 9387 69437 9388
rect 1323 9344 1365 9353
rect 1323 9304 1324 9344
rect 1364 9304 1365 9344
rect 1323 9295 1365 9304
rect 69195 9344 69237 9353
rect 69195 9304 69196 9344
rect 69236 9304 69237 9344
rect 69195 9295 69237 9304
rect 651 9260 693 9269
rect 651 9220 652 9260
rect 692 9220 693 9260
rect 651 9211 693 9220
rect 576 9092 69984 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 7112 9092
rect 7152 9052 7194 9092
rect 7234 9052 7276 9092
rect 7316 9052 7358 9092
rect 7398 9052 7440 9092
rect 7480 9052 11112 9092
rect 11152 9052 11194 9092
rect 11234 9052 11276 9092
rect 11316 9052 11358 9092
rect 11398 9052 11440 9092
rect 11480 9052 15112 9092
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15480 9052 19112 9092
rect 19152 9052 19194 9092
rect 19234 9052 19276 9092
rect 19316 9052 19358 9092
rect 19398 9052 19440 9092
rect 19480 9052 23112 9092
rect 23152 9052 23194 9092
rect 23234 9052 23276 9092
rect 23316 9052 23358 9092
rect 23398 9052 23440 9092
rect 23480 9052 27112 9092
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27480 9052 31112 9092
rect 31152 9052 31194 9092
rect 31234 9052 31276 9092
rect 31316 9052 31358 9092
rect 31398 9052 31440 9092
rect 31480 9052 35112 9092
rect 35152 9052 35194 9092
rect 35234 9052 35276 9092
rect 35316 9052 35358 9092
rect 35398 9052 35440 9092
rect 35480 9052 39112 9092
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39480 9052 43112 9092
rect 43152 9052 43194 9092
rect 43234 9052 43276 9092
rect 43316 9052 43358 9092
rect 43398 9052 43440 9092
rect 43480 9052 47112 9092
rect 47152 9052 47194 9092
rect 47234 9052 47276 9092
rect 47316 9052 47358 9092
rect 47398 9052 47440 9092
rect 47480 9052 51112 9092
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51480 9052 55112 9092
rect 55152 9052 55194 9092
rect 55234 9052 55276 9092
rect 55316 9052 55358 9092
rect 55398 9052 55440 9092
rect 55480 9052 59112 9092
rect 59152 9052 59194 9092
rect 59234 9052 59276 9092
rect 59316 9052 59358 9092
rect 59398 9052 59440 9092
rect 59480 9052 63112 9092
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63480 9052 67112 9092
rect 67152 9052 67194 9092
rect 67234 9052 67276 9092
rect 67316 9052 67358 9092
rect 67398 9052 67440 9092
rect 67480 9052 69984 9092
rect 576 9028 69984 9052
rect 1419 8840 1461 8849
rect 1419 8800 1420 8840
rect 1460 8800 1461 8840
rect 1419 8791 1461 8800
rect 835 8756 893 8757
rect 835 8716 844 8756
rect 884 8716 893 8756
rect 835 8715 893 8716
rect 1603 8756 1661 8757
rect 1603 8716 1612 8756
rect 1652 8716 1661 8756
rect 1603 8715 1661 8716
rect 1987 8756 2045 8757
rect 1987 8716 1996 8756
rect 2036 8716 2045 8756
rect 1987 8715 2045 8716
rect 651 8504 693 8513
rect 651 8464 652 8504
rect 692 8464 693 8504
rect 651 8455 693 8464
rect 1803 8504 1845 8513
rect 1803 8464 1804 8504
rect 1844 8464 1845 8504
rect 1803 8455 1845 8464
rect 576 8336 69984 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 8352 8336
rect 8392 8296 8434 8336
rect 8474 8296 8516 8336
rect 8556 8296 8598 8336
rect 8638 8296 8680 8336
rect 8720 8296 12352 8336
rect 12392 8296 12434 8336
rect 12474 8296 12516 8336
rect 12556 8296 12598 8336
rect 12638 8296 12680 8336
rect 12720 8296 16352 8336
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16720 8296 20352 8336
rect 20392 8296 20434 8336
rect 20474 8296 20516 8336
rect 20556 8296 20598 8336
rect 20638 8296 20680 8336
rect 20720 8296 24352 8336
rect 24392 8296 24434 8336
rect 24474 8296 24516 8336
rect 24556 8296 24598 8336
rect 24638 8296 24680 8336
rect 24720 8296 28352 8336
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28720 8296 32352 8336
rect 32392 8296 32434 8336
rect 32474 8296 32516 8336
rect 32556 8296 32598 8336
rect 32638 8296 32680 8336
rect 32720 8296 36352 8336
rect 36392 8296 36434 8336
rect 36474 8296 36516 8336
rect 36556 8296 36598 8336
rect 36638 8296 36680 8336
rect 36720 8296 40352 8336
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40720 8296 44352 8336
rect 44392 8296 44434 8336
rect 44474 8296 44516 8336
rect 44556 8296 44598 8336
rect 44638 8296 44680 8336
rect 44720 8296 48352 8336
rect 48392 8296 48434 8336
rect 48474 8296 48516 8336
rect 48556 8296 48598 8336
rect 48638 8296 48680 8336
rect 48720 8296 52352 8336
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52720 8296 56352 8336
rect 56392 8296 56434 8336
rect 56474 8296 56516 8336
rect 56556 8296 56598 8336
rect 56638 8296 56680 8336
rect 56720 8296 60352 8336
rect 60392 8296 60434 8336
rect 60474 8296 60516 8336
rect 60556 8296 60598 8336
rect 60638 8296 60680 8336
rect 60720 8296 64352 8336
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64720 8296 68352 8336
rect 68392 8296 68434 8336
rect 68474 8296 68516 8336
rect 68556 8296 68598 8336
rect 68638 8296 68680 8336
rect 68720 8296 69984 8336
rect 576 8272 69984 8296
rect 835 7916 893 7917
rect 835 7876 844 7916
rect 884 7876 893 7916
rect 835 7875 893 7876
rect 1699 7916 1757 7917
rect 1699 7876 1708 7916
rect 1748 7876 1757 7916
rect 1699 7875 1757 7876
rect 1515 7832 1557 7841
rect 1515 7792 1516 7832
rect 1556 7792 1557 7832
rect 1515 7783 1557 7792
rect 651 7748 693 7757
rect 651 7708 652 7748
rect 692 7708 693 7748
rect 651 7699 693 7708
rect 576 7580 99516 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 7112 7580
rect 7152 7540 7194 7580
rect 7234 7540 7276 7580
rect 7316 7540 7358 7580
rect 7398 7540 7440 7580
rect 7480 7540 11112 7580
rect 11152 7540 11194 7580
rect 11234 7540 11276 7580
rect 11316 7540 11358 7580
rect 11398 7540 11440 7580
rect 11480 7540 15112 7580
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15480 7540 19112 7580
rect 19152 7540 19194 7580
rect 19234 7540 19276 7580
rect 19316 7540 19358 7580
rect 19398 7540 19440 7580
rect 19480 7540 23112 7580
rect 23152 7540 23194 7580
rect 23234 7540 23276 7580
rect 23316 7540 23358 7580
rect 23398 7540 23440 7580
rect 23480 7540 27112 7580
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27480 7540 31112 7580
rect 31152 7540 31194 7580
rect 31234 7540 31276 7580
rect 31316 7540 31358 7580
rect 31398 7540 31440 7580
rect 31480 7540 35112 7580
rect 35152 7540 35194 7580
rect 35234 7540 35276 7580
rect 35316 7540 35358 7580
rect 35398 7540 35440 7580
rect 35480 7540 39112 7580
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39480 7540 43112 7580
rect 43152 7540 43194 7580
rect 43234 7540 43276 7580
rect 43316 7540 43358 7580
rect 43398 7540 43440 7580
rect 43480 7540 47112 7580
rect 47152 7540 47194 7580
rect 47234 7540 47276 7580
rect 47316 7540 47358 7580
rect 47398 7540 47440 7580
rect 47480 7540 51112 7580
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51480 7540 55112 7580
rect 55152 7540 55194 7580
rect 55234 7540 55276 7580
rect 55316 7540 55358 7580
rect 55398 7540 55440 7580
rect 55480 7540 59112 7580
rect 59152 7540 59194 7580
rect 59234 7540 59276 7580
rect 59316 7540 59358 7580
rect 59398 7540 59440 7580
rect 59480 7540 63112 7580
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63480 7540 67112 7580
rect 67152 7540 67194 7580
rect 67234 7540 67276 7580
rect 67316 7540 67358 7580
rect 67398 7540 67440 7580
rect 67480 7540 71112 7580
rect 71152 7540 71194 7580
rect 71234 7540 71276 7580
rect 71316 7540 71358 7580
rect 71398 7540 71440 7580
rect 71480 7540 75112 7580
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75480 7540 79112 7580
rect 79152 7540 79194 7580
rect 79234 7540 79276 7580
rect 79316 7540 79358 7580
rect 79398 7540 79440 7580
rect 79480 7540 83112 7580
rect 83152 7540 83194 7580
rect 83234 7540 83276 7580
rect 83316 7540 83358 7580
rect 83398 7540 83440 7580
rect 83480 7540 87112 7580
rect 87152 7540 87194 7580
rect 87234 7540 87276 7580
rect 87316 7540 87358 7580
rect 87398 7540 87440 7580
rect 87480 7540 91112 7580
rect 91152 7540 91194 7580
rect 91234 7540 91276 7580
rect 91316 7540 91358 7580
rect 91398 7540 91440 7580
rect 91480 7540 95112 7580
rect 95152 7540 95194 7580
rect 95234 7540 95276 7580
rect 95316 7540 95358 7580
rect 95398 7540 95440 7580
rect 95480 7540 99112 7580
rect 99152 7540 99194 7580
rect 99234 7540 99276 7580
rect 99316 7540 99358 7580
rect 99398 7540 99440 7580
rect 99480 7540 99516 7580
rect 576 7516 99516 7540
rect 73419 7412 73461 7421
rect 73419 7372 73420 7412
rect 73460 7372 73461 7412
rect 73419 7363 73461 7372
rect 73803 7412 73845 7421
rect 73803 7372 73804 7412
rect 73844 7372 73845 7412
rect 73803 7363 73845 7372
rect 75243 7412 75285 7421
rect 75243 7372 75244 7412
rect 75284 7372 75285 7412
rect 75243 7363 75285 7372
rect 75915 7412 75957 7421
rect 75915 7372 75916 7412
rect 75956 7372 75957 7412
rect 75915 7363 75957 7372
rect 76299 7412 76341 7421
rect 76299 7372 76300 7412
rect 76340 7372 76341 7412
rect 76299 7363 76341 7372
rect 77067 7412 77109 7421
rect 77067 7372 77068 7412
rect 77108 7372 77109 7412
rect 77067 7363 77109 7372
rect 78027 7412 78069 7421
rect 78027 7372 78028 7412
rect 78068 7372 78069 7412
rect 78027 7363 78069 7372
rect 78315 7412 78357 7421
rect 78315 7372 78316 7412
rect 78356 7372 78357 7412
rect 78315 7363 78357 7372
rect 78795 7412 78837 7421
rect 78795 7372 78796 7412
rect 78836 7372 78837 7412
rect 78795 7363 78837 7372
rect 79179 7412 79221 7421
rect 79179 7372 79180 7412
rect 79220 7372 79221 7412
rect 79179 7363 79221 7372
rect 79467 7412 79509 7421
rect 79467 7372 79468 7412
rect 79508 7372 79509 7412
rect 79467 7363 79509 7372
rect 79851 7412 79893 7421
rect 79851 7372 79852 7412
rect 79892 7372 79893 7412
rect 79851 7363 79893 7372
rect 81483 7412 81525 7421
rect 81483 7372 81484 7412
rect 81524 7372 81525 7412
rect 81483 7363 81525 7372
rect 81675 7412 81717 7421
rect 81675 7372 81676 7412
rect 81716 7372 81717 7412
rect 81675 7363 81717 7372
rect 82347 7412 82389 7421
rect 82347 7372 82348 7412
rect 82388 7372 82389 7412
rect 82347 7363 82389 7372
rect 83403 7412 83445 7421
rect 83403 7372 83404 7412
rect 83444 7372 83445 7412
rect 83403 7363 83445 7372
rect 83883 7412 83925 7421
rect 83883 7372 83884 7412
rect 83924 7372 83925 7412
rect 83883 7363 83925 7372
rect 84651 7412 84693 7421
rect 84651 7372 84652 7412
rect 84692 7372 84693 7412
rect 84651 7363 84693 7372
rect 85035 7412 85077 7421
rect 85035 7372 85036 7412
rect 85076 7372 85077 7412
rect 85035 7363 85077 7372
rect 85707 7412 85749 7421
rect 85707 7372 85708 7412
rect 85748 7372 85749 7412
rect 85707 7363 85749 7372
rect 87147 7412 87189 7421
rect 87147 7372 87148 7412
rect 87188 7372 87189 7412
rect 87147 7363 87189 7372
rect 87723 7412 87765 7421
rect 87723 7372 87724 7412
rect 87764 7372 87765 7412
rect 87723 7363 87765 7372
rect 88779 7412 88821 7421
rect 88779 7372 88780 7412
rect 88820 7372 88821 7412
rect 88779 7363 88821 7372
rect 88971 7412 89013 7421
rect 88971 7372 88972 7412
rect 89012 7372 89013 7412
rect 88971 7363 89013 7372
rect 89643 7412 89685 7421
rect 89643 7372 89644 7412
rect 89684 7372 89685 7412
rect 89643 7363 89685 7372
rect 90411 7412 90453 7421
rect 90411 7372 90412 7412
rect 90452 7372 90453 7412
rect 90411 7363 90453 7372
rect 90603 7412 90645 7421
rect 90603 7372 90604 7412
rect 90644 7372 90645 7412
rect 90603 7363 90645 7372
rect 91851 7412 91893 7421
rect 91851 7372 91852 7412
rect 91892 7372 91893 7412
rect 91851 7363 91893 7372
rect 92907 7412 92949 7421
rect 92907 7372 92908 7412
rect 92948 7372 92949 7412
rect 92907 7363 92949 7372
rect 93291 7412 93333 7421
rect 93291 7372 93292 7412
rect 93332 7372 93333 7412
rect 93291 7363 93333 7372
rect 94731 7412 94773 7421
rect 94731 7372 94732 7412
rect 94772 7372 94773 7412
rect 94731 7363 94773 7372
rect 95115 7412 95157 7421
rect 95115 7372 95116 7412
rect 95156 7372 95157 7412
rect 95115 7363 95157 7372
rect 95883 7412 95925 7421
rect 95883 7372 95884 7412
rect 95924 7372 95925 7412
rect 95883 7363 95925 7372
rect 96843 7412 96885 7421
rect 96843 7372 96844 7412
rect 96884 7372 96885 7412
rect 96843 7363 96885 7372
rect 97131 7412 97173 7421
rect 97131 7372 97132 7412
rect 97172 7372 97173 7412
rect 97131 7363 97173 7372
rect 97419 7412 97461 7421
rect 97419 7372 97420 7412
rect 97460 7372 97461 7412
rect 97419 7363 97461 7372
rect 97995 7412 98037 7421
rect 97995 7372 97996 7412
rect 98036 7372 98037 7412
rect 97995 7363 98037 7372
rect 98475 7412 98517 7421
rect 98475 7372 98476 7412
rect 98516 7372 98517 7412
rect 98475 7363 98517 7372
rect 74475 7328 74517 7337
rect 74475 7288 74476 7328
rect 74516 7288 74517 7328
rect 74475 7279 74517 7288
rect 80043 7328 80085 7337
rect 80043 7288 80044 7328
rect 80084 7288 80085 7328
rect 80043 7279 80085 7288
rect 80715 7328 80757 7337
rect 80715 7288 80716 7328
rect 80756 7288 80757 7328
rect 80715 7279 80757 7288
rect 86283 7328 86325 7337
rect 86283 7288 86284 7328
rect 86324 7288 86325 7328
rect 86283 7279 86325 7288
rect 86475 7328 86517 7337
rect 86475 7288 86476 7328
rect 86516 7288 86517 7328
rect 86475 7279 86517 7288
rect 91179 7328 91221 7337
rect 91179 7288 91180 7328
rect 91220 7288 91221 7328
rect 91179 7279 91221 7288
rect 92331 7328 92373 7337
rect 92331 7288 92332 7328
rect 92372 7288 92373 7328
rect 92331 7279 92373 7288
rect 92523 7328 92565 7337
rect 92523 7288 92524 7328
rect 92564 7288 92565 7328
rect 92523 7279 92565 7288
rect 93963 7328 94005 7337
rect 93963 7288 93964 7328
rect 94004 7288 94005 7328
rect 93963 7279 94005 7288
rect 96651 7328 96693 7337
rect 96651 7288 96652 7328
rect 96692 7288 96693 7328
rect 96651 7279 96693 7288
rect 835 7244 893 7245
rect 835 7204 844 7244
rect 884 7204 893 7244
rect 835 7203 893 7204
rect 73603 7244 73661 7245
rect 73603 7204 73612 7244
rect 73652 7204 73661 7244
rect 73603 7203 73661 7204
rect 74275 7244 74333 7245
rect 74275 7204 74284 7244
rect 74324 7204 74333 7244
rect 74275 7203 74333 7204
rect 74659 7244 74717 7245
rect 74659 7204 74668 7244
rect 74708 7204 74717 7244
rect 74659 7203 74717 7204
rect 75043 7244 75101 7245
rect 75043 7204 75052 7244
rect 75092 7204 75101 7244
rect 75043 7203 75101 7204
rect 75427 7244 75485 7245
rect 75427 7204 75436 7244
rect 75476 7204 75485 7244
rect 75427 7203 75485 7204
rect 75715 7244 75773 7245
rect 75715 7204 75724 7244
rect 75764 7204 75773 7244
rect 75715 7203 75773 7204
rect 76099 7244 76157 7245
rect 76099 7204 76108 7244
rect 76148 7204 76157 7244
rect 76099 7203 76157 7204
rect 76867 7244 76925 7245
rect 76867 7204 76876 7244
rect 76916 7204 76925 7244
rect 76867 7203 76925 7204
rect 77443 7244 77501 7245
rect 77443 7204 77452 7244
rect 77492 7204 77501 7244
rect 77443 7203 77501 7204
rect 77827 7244 77885 7245
rect 77827 7204 77836 7244
rect 77876 7204 77885 7244
rect 77827 7203 77885 7204
rect 79651 7244 79709 7245
rect 79651 7204 79660 7244
rect 79700 7204 79709 7244
rect 79651 7203 79709 7204
rect 80227 7244 80285 7245
rect 80227 7204 80236 7244
rect 80276 7204 80285 7244
rect 80227 7203 80285 7204
rect 80515 7244 80573 7245
rect 80515 7204 80524 7244
rect 80564 7204 80573 7244
rect 80515 7203 80573 7204
rect 81091 7244 81149 7245
rect 81091 7204 81100 7244
rect 81140 7204 81149 7244
rect 81091 7203 81149 7204
rect 81283 7244 81341 7245
rect 81283 7204 81292 7244
rect 81332 7204 81341 7244
rect 81283 7203 81341 7204
rect 82819 7244 82877 7245
rect 82819 7204 82828 7244
rect 82868 7204 82877 7244
rect 82819 7203 82877 7204
rect 83019 7244 83061 7253
rect 83019 7204 83020 7244
rect 83060 7204 83061 7244
rect 83019 7195 83061 7204
rect 84259 7244 84317 7245
rect 84259 7204 84268 7244
rect 84308 7204 84317 7244
rect 84259 7203 84317 7204
rect 84835 7244 84893 7245
rect 84835 7204 84844 7244
rect 84884 7204 84893 7244
rect 84835 7203 84893 7204
rect 85219 7244 85277 7245
rect 85219 7204 85228 7244
rect 85268 7204 85277 7244
rect 85219 7203 85277 7204
rect 86083 7244 86141 7245
rect 86083 7204 86092 7244
rect 86132 7204 86141 7244
rect 86083 7203 86141 7204
rect 86659 7244 86717 7245
rect 86659 7204 86668 7244
rect 86708 7204 86717 7244
rect 86659 7203 86717 7204
rect 88003 7244 88061 7245
rect 88003 7204 88012 7244
rect 88052 7204 88061 7244
rect 88003 7203 88061 7204
rect 88579 7244 88637 7245
rect 88579 7204 88588 7244
rect 88628 7204 88637 7244
rect 88579 7203 88637 7204
rect 89443 7244 89501 7245
rect 89443 7204 89452 7244
rect 89492 7204 89501 7244
rect 89443 7203 89501 7204
rect 90019 7244 90077 7245
rect 90019 7204 90028 7244
rect 90068 7204 90077 7244
rect 90019 7203 90077 7204
rect 90979 7244 91037 7245
rect 90979 7204 90988 7244
rect 91028 7204 91037 7244
rect 90979 7203 91037 7204
rect 91363 7244 91421 7245
rect 91363 7204 91372 7244
rect 91412 7204 91421 7244
rect 91363 7203 91421 7204
rect 92131 7244 92189 7245
rect 92131 7204 92140 7244
rect 92180 7204 92189 7244
rect 92131 7203 92189 7204
rect 92707 7244 92765 7245
rect 92707 7204 92716 7244
rect 92756 7204 92765 7244
rect 92707 7203 92765 7204
rect 93091 7244 93149 7245
rect 93091 7204 93100 7244
rect 93140 7204 93149 7244
rect 93091 7203 93149 7204
rect 94147 7244 94205 7245
rect 94147 7204 94156 7244
rect 94196 7204 94205 7244
rect 94147 7203 94205 7204
rect 94339 7244 94397 7245
rect 94339 7204 94348 7244
rect 94388 7204 94397 7244
rect 94339 7203 94397 7204
rect 94915 7244 94973 7245
rect 94915 7204 94924 7244
rect 94964 7204 94973 7244
rect 94915 7203 94973 7204
rect 95299 7244 95357 7245
rect 95299 7204 95308 7244
rect 95348 7204 95357 7244
rect 95299 7203 95357 7204
rect 95683 7244 95741 7245
rect 95683 7204 95692 7244
rect 95732 7204 95741 7244
rect 95683 7203 95741 7204
rect 96259 7244 96317 7245
rect 96259 7204 96268 7244
rect 96308 7204 96317 7244
rect 96259 7203 96317 7204
rect 96451 7244 96509 7245
rect 96451 7204 96460 7244
rect 96500 7204 96509 7244
rect 96451 7203 96509 7204
rect 97603 7244 97661 7245
rect 97603 7204 97612 7244
rect 97652 7204 97661 7244
rect 97603 7203 97661 7204
rect 98179 7244 98237 7245
rect 98179 7204 98188 7244
rect 98228 7204 98237 7244
rect 98179 7203 98237 7204
rect 98659 7244 98717 7245
rect 98659 7204 98668 7244
rect 98708 7204 98717 7244
rect 98659 7203 98717 7204
rect 73315 7160 73373 7161
rect 73315 7120 73324 7160
rect 73364 7120 73373 7160
rect 73315 7119 73373 7120
rect 76675 7160 76733 7161
rect 76675 7120 76684 7160
rect 76724 7120 76733 7160
rect 76675 7119 76733 7120
rect 78115 7160 78173 7161
rect 78115 7120 78124 7160
rect 78164 7120 78173 7160
rect 78115 7119 78173 7120
rect 78403 7160 78461 7161
rect 78403 7120 78412 7160
rect 78452 7120 78461 7160
rect 79075 7160 79133 7161
rect 78403 7119 78461 7120
rect 78691 7149 78749 7150
rect 78691 7109 78700 7149
rect 78740 7109 78749 7149
rect 79075 7120 79084 7160
rect 79124 7120 79133 7160
rect 79075 7119 79133 7120
rect 79363 7160 79421 7161
rect 79363 7120 79372 7160
rect 79412 7120 79421 7160
rect 79363 7119 79421 7120
rect 81763 7160 81821 7161
rect 81763 7120 81772 7160
rect 81812 7120 81821 7160
rect 82059 7160 82101 7169
rect 81763 7119 81821 7120
rect 81955 7149 82013 7150
rect 78691 7108 78749 7109
rect 81955 7109 81964 7149
rect 82004 7109 82013 7149
rect 82059 7120 82060 7160
rect 82100 7120 82101 7160
rect 82059 7111 82101 7120
rect 82243 7160 82301 7161
rect 82243 7120 82252 7160
rect 82292 7120 82301 7160
rect 82243 7119 82301 7120
rect 83107 7160 83165 7161
rect 83107 7120 83116 7160
rect 83156 7120 83165 7160
rect 83107 7119 83165 7120
rect 83299 7160 83357 7161
rect 83299 7120 83308 7160
rect 83348 7120 83357 7160
rect 83299 7119 83357 7120
rect 83779 7160 83837 7161
rect 83779 7120 83788 7160
rect 83828 7120 83837 7160
rect 83779 7119 83837 7120
rect 84547 7160 84605 7161
rect 84547 7120 84556 7160
rect 84596 7120 84605 7160
rect 84547 7119 84605 7120
rect 85603 7160 85661 7161
rect 85603 7120 85612 7160
rect 85652 7120 85661 7160
rect 85603 7119 85661 7120
rect 86851 7160 86909 7161
rect 86851 7120 86860 7160
rect 86900 7120 86909 7160
rect 86851 7119 86909 7120
rect 87235 7160 87293 7161
rect 87235 7120 87244 7160
rect 87284 7120 87293 7160
rect 87235 7119 87293 7120
rect 87435 7160 87477 7169
rect 87435 7120 87436 7160
rect 87476 7120 87477 7160
rect 87435 7111 87477 7120
rect 87523 7160 87581 7161
rect 87523 7120 87532 7160
rect 87572 7120 87581 7160
rect 87523 7119 87581 7120
rect 87811 7160 87869 7161
rect 87811 7120 87820 7160
rect 87860 7120 87869 7160
rect 87811 7119 87869 7120
rect 89059 7160 89117 7161
rect 89059 7120 89068 7160
rect 89108 7120 89117 7160
rect 89059 7119 89117 7120
rect 90307 7160 90365 7161
rect 90307 7120 90316 7160
rect 90356 7120 90365 7160
rect 90307 7119 90365 7120
rect 90712 7160 90754 7169
rect 90712 7120 90713 7160
rect 90753 7120 90754 7160
rect 90712 7111 90754 7120
rect 91747 7160 91805 7161
rect 91747 7120 91756 7160
rect 91796 7120 91805 7160
rect 91747 7119 91805 7120
rect 93379 7160 93437 7161
rect 93379 7120 93388 7160
rect 93428 7120 93437 7160
rect 93379 7119 93437 7120
rect 93667 7160 93725 7161
rect 93667 7120 93676 7160
rect 93716 7120 93725 7160
rect 93667 7119 93725 7120
rect 96931 7160 96989 7161
rect 96931 7120 96940 7160
rect 96980 7120 96989 7160
rect 96931 7119 96989 7120
rect 97219 7160 97277 7161
rect 97219 7120 97228 7160
rect 97268 7120 97277 7160
rect 97219 7119 97277 7120
rect 81955 7108 82013 7109
rect 76587 7076 76629 7085
rect 76587 7036 76588 7076
rect 76628 7036 76629 7076
rect 76587 7027 76629 7036
rect 651 6992 693 7001
rect 651 6952 652 6992
rect 692 6952 693 6992
rect 651 6943 693 6952
rect 74091 6992 74133 7001
rect 74091 6952 74092 6992
rect 74132 6952 74133 6992
rect 74091 6943 74133 6952
rect 74859 6992 74901 7001
rect 74859 6952 74860 6992
rect 74900 6952 74901 6992
rect 74859 6943 74901 6952
rect 77259 6992 77301 7001
rect 77259 6952 77260 6992
rect 77300 6952 77301 6992
rect 77259 6943 77301 6952
rect 77643 6992 77685 7001
rect 77643 6952 77644 6992
rect 77684 6952 77685 6992
rect 77643 6943 77685 6952
rect 80907 6992 80949 7001
rect 80907 6952 80908 6992
rect 80948 6952 80949 6992
rect 80907 6943 80949 6952
rect 82635 6992 82677 7001
rect 82635 6952 82636 6992
rect 82676 6952 82677 6992
rect 82635 6943 82677 6952
rect 84075 6992 84117 7001
rect 84075 6952 84076 6992
rect 84116 6952 84117 6992
rect 84075 6943 84117 6952
rect 85419 6992 85461 7001
rect 85419 6952 85420 6992
rect 85460 6952 85461 6992
rect 85419 6943 85461 6952
rect 86955 6992 86997 7001
rect 86955 6952 86956 6992
rect 86996 6952 86997 6992
rect 86955 6943 86997 6952
rect 88203 6992 88245 7001
rect 88203 6952 88204 6992
rect 88244 6952 88245 6992
rect 88203 6943 88245 6952
rect 89835 6992 89877 7001
rect 89835 6952 89836 6992
rect 89876 6952 89877 6992
rect 89835 6943 89877 6952
rect 91563 6992 91605 7001
rect 91563 6952 91564 6992
rect 91604 6952 91605 6992
rect 91563 6943 91605 6952
rect 93771 6992 93813 7001
rect 93771 6952 93772 6992
rect 93812 6952 93813 6992
rect 93771 6943 93813 6952
rect 94539 6992 94581 7001
rect 94539 6952 94540 6992
rect 94580 6952 94581 6992
rect 94539 6943 94581 6952
rect 96075 6992 96117 7001
rect 96075 6952 96076 6992
rect 96116 6952 96117 6992
rect 96075 6943 96117 6952
rect 576 6824 99360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 8352 6824
rect 8392 6784 8434 6824
rect 8474 6784 8516 6824
rect 8556 6784 8598 6824
rect 8638 6784 8680 6824
rect 8720 6784 12352 6824
rect 12392 6784 12434 6824
rect 12474 6784 12516 6824
rect 12556 6784 12598 6824
rect 12638 6784 12680 6824
rect 12720 6784 16352 6824
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16720 6784 20352 6824
rect 20392 6784 20434 6824
rect 20474 6784 20516 6824
rect 20556 6784 20598 6824
rect 20638 6784 20680 6824
rect 20720 6784 24352 6824
rect 24392 6784 24434 6824
rect 24474 6784 24516 6824
rect 24556 6784 24598 6824
rect 24638 6784 24680 6824
rect 24720 6784 28352 6824
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28720 6784 32352 6824
rect 32392 6784 32434 6824
rect 32474 6784 32516 6824
rect 32556 6784 32598 6824
rect 32638 6784 32680 6824
rect 32720 6784 36352 6824
rect 36392 6784 36434 6824
rect 36474 6784 36516 6824
rect 36556 6784 36598 6824
rect 36638 6784 36680 6824
rect 36720 6784 40352 6824
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40720 6784 44352 6824
rect 44392 6784 44434 6824
rect 44474 6784 44516 6824
rect 44556 6784 44598 6824
rect 44638 6784 44680 6824
rect 44720 6784 48352 6824
rect 48392 6784 48434 6824
rect 48474 6784 48516 6824
rect 48556 6784 48598 6824
rect 48638 6784 48680 6824
rect 48720 6784 52352 6824
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52720 6784 56352 6824
rect 56392 6784 56434 6824
rect 56474 6784 56516 6824
rect 56556 6784 56598 6824
rect 56638 6784 56680 6824
rect 56720 6784 60352 6824
rect 60392 6784 60434 6824
rect 60474 6784 60516 6824
rect 60556 6784 60598 6824
rect 60638 6784 60680 6824
rect 60720 6784 64352 6824
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64720 6784 68352 6824
rect 68392 6784 68434 6824
rect 68474 6784 68516 6824
rect 68556 6784 68598 6824
rect 68638 6784 68680 6824
rect 68720 6784 72352 6824
rect 72392 6784 72434 6824
rect 72474 6784 72516 6824
rect 72556 6784 72598 6824
rect 72638 6784 72680 6824
rect 72720 6784 76352 6824
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76720 6784 80352 6824
rect 80392 6784 80434 6824
rect 80474 6784 80516 6824
rect 80556 6784 80598 6824
rect 80638 6784 80680 6824
rect 80720 6784 84352 6824
rect 84392 6784 84434 6824
rect 84474 6784 84516 6824
rect 84556 6784 84598 6824
rect 84638 6784 84680 6824
rect 84720 6784 88352 6824
rect 88392 6784 88434 6824
rect 88474 6784 88516 6824
rect 88556 6784 88598 6824
rect 88638 6784 88680 6824
rect 88720 6784 92352 6824
rect 92392 6784 92434 6824
rect 92474 6784 92516 6824
rect 92556 6784 92598 6824
rect 92638 6784 92680 6824
rect 92720 6784 96352 6824
rect 96392 6784 96434 6824
rect 96474 6784 96516 6824
rect 96556 6784 96598 6824
rect 96638 6784 96680 6824
rect 96720 6784 99360 6824
rect 576 6760 99360 6784
rect 1323 6656 1365 6665
rect 1323 6616 1324 6656
rect 1364 6616 1365 6656
rect 1323 6607 1365 6616
rect 74187 6656 74229 6665
rect 74187 6616 74188 6656
rect 74228 6616 74229 6656
rect 74187 6607 74229 6616
rect 75243 6656 75285 6665
rect 75243 6616 75244 6656
rect 75284 6616 75285 6656
rect 75243 6607 75285 6616
rect 75531 6656 75573 6665
rect 75531 6616 75532 6656
rect 75572 6616 75573 6656
rect 75531 6607 75573 6616
rect 75819 6656 75861 6665
rect 75819 6616 75820 6656
rect 75860 6616 75861 6656
rect 75819 6607 75861 6616
rect 76395 6656 76437 6665
rect 76395 6616 76396 6656
rect 76436 6616 76437 6656
rect 76395 6607 76437 6616
rect 76779 6656 76821 6665
rect 76779 6616 76780 6656
rect 76820 6616 76821 6656
rect 76779 6607 76821 6616
rect 77163 6656 77205 6665
rect 77163 6616 77164 6656
rect 77204 6616 77205 6656
rect 77163 6607 77205 6616
rect 77931 6656 77973 6665
rect 77931 6616 77932 6656
rect 77972 6616 77973 6656
rect 77931 6607 77973 6616
rect 78315 6656 78357 6665
rect 78315 6616 78316 6656
rect 78356 6616 78357 6656
rect 78315 6607 78357 6616
rect 79083 6656 79125 6665
rect 79083 6616 79084 6656
rect 79124 6616 79125 6656
rect 79083 6607 79125 6616
rect 80043 6656 80085 6665
rect 80043 6616 80044 6656
rect 80084 6616 80085 6656
rect 80043 6607 80085 6616
rect 80619 6656 80661 6665
rect 80619 6616 80620 6656
rect 80660 6616 80661 6656
rect 80619 6607 80661 6616
rect 81099 6656 81141 6665
rect 81099 6616 81100 6656
rect 81140 6616 81141 6656
rect 81099 6607 81141 6616
rect 81483 6656 81525 6665
rect 81483 6616 81484 6656
rect 81524 6616 81525 6656
rect 81483 6607 81525 6616
rect 81867 6656 81909 6665
rect 81867 6616 81868 6656
rect 81908 6616 81909 6656
rect 81867 6607 81909 6616
rect 82251 6656 82293 6665
rect 82251 6616 82252 6656
rect 82292 6616 82293 6656
rect 82251 6607 82293 6616
rect 82923 6656 82965 6665
rect 82923 6616 82924 6656
rect 82964 6616 82965 6656
rect 82923 6607 82965 6616
rect 83403 6656 83445 6665
rect 83403 6616 83404 6656
rect 83444 6616 83445 6656
rect 83403 6607 83445 6616
rect 83883 6656 83925 6665
rect 83883 6616 83884 6656
rect 83924 6616 83925 6656
rect 83883 6607 83925 6616
rect 84363 6656 84405 6665
rect 84363 6616 84364 6656
rect 84404 6616 84405 6656
rect 84363 6607 84405 6616
rect 84747 6656 84789 6665
rect 84747 6616 84748 6656
rect 84788 6616 84789 6656
rect 84747 6607 84789 6616
rect 84939 6656 84981 6665
rect 84939 6616 84940 6656
rect 84980 6616 84981 6656
rect 84939 6607 84981 6616
rect 85419 6656 85461 6665
rect 85419 6616 85420 6656
rect 85460 6616 85461 6656
rect 85419 6607 85461 6616
rect 85803 6656 85845 6665
rect 85803 6616 85804 6656
rect 85844 6616 85845 6656
rect 85803 6607 85845 6616
rect 86283 6656 86325 6665
rect 86283 6616 86284 6656
rect 86324 6616 86325 6656
rect 86283 6607 86325 6616
rect 87051 6656 87093 6665
rect 87051 6616 87052 6656
rect 87092 6616 87093 6656
rect 87051 6607 87093 6616
rect 87531 6656 87573 6665
rect 87531 6616 87532 6656
rect 87572 6616 87573 6656
rect 87531 6607 87573 6616
rect 87915 6656 87957 6665
rect 87915 6616 87916 6656
rect 87956 6616 87957 6656
rect 87915 6607 87957 6616
rect 88299 6656 88341 6665
rect 88299 6616 88300 6656
rect 88340 6616 88341 6656
rect 88299 6607 88341 6616
rect 88491 6656 88533 6665
rect 88491 6616 88492 6656
rect 88532 6616 88533 6656
rect 88491 6607 88533 6616
rect 89259 6656 89301 6665
rect 89259 6616 89260 6656
rect 89300 6616 89301 6656
rect 89259 6607 89301 6616
rect 90603 6656 90645 6665
rect 90603 6616 90604 6656
rect 90644 6616 90645 6656
rect 90603 6607 90645 6616
rect 91083 6656 91125 6665
rect 91083 6616 91084 6656
rect 91124 6616 91125 6656
rect 91083 6607 91125 6616
rect 91275 6656 91317 6665
rect 91275 6616 91276 6656
rect 91316 6616 91317 6656
rect 91275 6607 91317 6616
rect 91851 6656 91893 6665
rect 91851 6616 91852 6656
rect 91892 6616 91893 6656
rect 91851 6607 91893 6616
rect 92331 6656 92373 6665
rect 92331 6616 92332 6656
rect 92372 6616 92373 6656
rect 92331 6607 92373 6616
rect 92619 6656 92661 6665
rect 92619 6616 92620 6656
rect 92660 6616 92661 6656
rect 92619 6607 92661 6616
rect 93195 6656 93237 6665
rect 93195 6616 93196 6656
rect 93236 6616 93237 6656
rect 93195 6607 93237 6616
rect 93579 6656 93621 6665
rect 93579 6616 93580 6656
rect 93620 6616 93621 6656
rect 93579 6607 93621 6616
rect 94059 6656 94101 6665
rect 94059 6616 94060 6656
rect 94100 6616 94101 6656
rect 94059 6607 94101 6616
rect 94251 6656 94293 6665
rect 94251 6616 94252 6656
rect 94292 6616 94293 6656
rect 94251 6607 94293 6616
rect 94827 6656 94869 6665
rect 94827 6616 94828 6656
rect 94868 6616 94869 6656
rect 94827 6607 94869 6616
rect 95307 6656 95349 6665
rect 95307 6616 95308 6656
rect 95348 6616 95349 6656
rect 95307 6607 95349 6616
rect 95595 6656 95637 6665
rect 95595 6616 95596 6656
rect 95636 6616 95637 6656
rect 95595 6607 95637 6616
rect 96555 6656 96597 6665
rect 96555 6616 96556 6656
rect 96596 6616 96597 6656
rect 96555 6607 96597 6616
rect 97131 6656 97173 6665
rect 97131 6616 97132 6656
rect 97172 6616 97173 6656
rect 97131 6607 97173 6616
rect 97419 6656 97461 6665
rect 97419 6616 97420 6656
rect 97460 6616 97461 6656
rect 97419 6607 97461 6616
rect 97707 6656 97749 6665
rect 97707 6616 97708 6656
rect 97748 6616 97749 6656
rect 97707 6607 97749 6616
rect 98091 6656 98133 6665
rect 98091 6616 98092 6656
rect 98132 6616 98133 6656
rect 98091 6607 98133 6616
rect 74083 6488 74141 6489
rect 74083 6448 74092 6488
rect 74132 6448 74141 6488
rect 75427 6488 75485 6489
rect 74083 6447 74141 6448
rect 75136 6475 75194 6476
rect 75136 6435 75145 6475
rect 75185 6435 75194 6475
rect 75427 6448 75436 6488
rect 75476 6448 75485 6488
rect 75427 6447 75485 6448
rect 75715 6488 75773 6489
rect 75715 6448 75724 6488
rect 75764 6448 75773 6488
rect 75715 6447 75773 6448
rect 76291 6488 76349 6489
rect 76291 6448 76300 6488
rect 76340 6448 76349 6488
rect 76291 6447 76349 6448
rect 76675 6488 76733 6489
rect 76675 6448 76684 6488
rect 76724 6448 76733 6488
rect 76675 6447 76733 6448
rect 79939 6488 79997 6489
rect 79939 6448 79948 6488
rect 79988 6448 79997 6488
rect 79939 6447 79997 6448
rect 81379 6488 81437 6489
rect 81379 6448 81388 6488
rect 81428 6448 81437 6488
rect 81379 6447 81437 6448
rect 85027 6488 85085 6489
rect 85027 6448 85036 6488
rect 85076 6448 85085 6488
rect 85027 6447 85085 6448
rect 88579 6488 88637 6489
rect 88579 6448 88588 6488
rect 88628 6448 88637 6488
rect 88579 6447 88637 6448
rect 88779 6488 88821 6497
rect 88779 6448 88780 6488
rect 88820 6448 88821 6488
rect 88779 6439 88821 6448
rect 88867 6488 88925 6489
rect 88867 6448 88876 6488
rect 88916 6448 88925 6488
rect 88867 6447 88925 6448
rect 89155 6488 89213 6489
rect 89155 6448 89164 6488
rect 89204 6448 89213 6488
rect 89155 6447 89213 6448
rect 91363 6488 91421 6489
rect 91363 6448 91372 6488
rect 91412 6448 91421 6488
rect 91363 6447 91421 6448
rect 92515 6488 92573 6489
rect 92515 6448 92524 6488
rect 92564 6448 92573 6488
rect 92515 6447 92573 6448
rect 94723 6488 94781 6489
rect 94723 6448 94732 6488
rect 94772 6448 94781 6488
rect 94723 6447 94781 6448
rect 95683 6488 95741 6489
rect 95683 6448 95692 6488
rect 95732 6448 95741 6488
rect 95683 6447 95741 6448
rect 95875 6488 95933 6489
rect 95875 6448 95884 6488
rect 95924 6448 95933 6488
rect 95875 6447 95933 6448
rect 97315 6488 97373 6489
rect 97315 6448 97324 6488
rect 97364 6448 97373 6488
rect 97315 6447 97373 6448
rect 97795 6488 97853 6489
rect 97795 6448 97804 6488
rect 97844 6448 97853 6488
rect 97795 6447 97853 6448
rect 97987 6488 98045 6489
rect 97987 6448 97996 6488
rect 98036 6448 98045 6488
rect 97987 6447 98045 6448
rect 75136 6434 75194 6435
rect 1507 6404 1565 6405
rect 1507 6364 1516 6404
rect 1556 6364 1565 6404
rect 1507 6363 1565 6364
rect 74371 6404 74429 6405
rect 74371 6364 74380 6404
rect 74420 6364 74429 6404
rect 74371 6363 74429 6364
rect 74755 6404 74813 6405
rect 74755 6364 74764 6404
rect 74804 6364 74813 6404
rect 74755 6363 74813 6364
rect 76963 6404 77021 6405
rect 76963 6364 76972 6404
rect 77012 6364 77021 6404
rect 76963 6363 77021 6364
rect 77731 6404 77789 6405
rect 77731 6364 77740 6404
rect 77780 6364 77789 6404
rect 77731 6363 77789 6364
rect 78115 6404 78173 6405
rect 78115 6364 78124 6404
rect 78164 6364 78173 6404
rect 78115 6363 78173 6364
rect 78883 6404 78941 6405
rect 78883 6364 78892 6404
rect 78932 6364 78941 6404
rect 78883 6363 78941 6364
rect 79555 6404 79613 6405
rect 79555 6364 79564 6404
rect 79604 6364 79613 6404
rect 79555 6363 79613 6364
rect 80419 6404 80477 6405
rect 80419 6364 80428 6404
rect 80468 6364 80477 6404
rect 80419 6363 80477 6364
rect 80899 6404 80957 6405
rect 80899 6364 80908 6404
rect 80948 6364 80957 6404
rect 80899 6363 80957 6364
rect 81667 6404 81725 6405
rect 81667 6364 81676 6404
rect 81716 6364 81725 6404
rect 81667 6363 81725 6364
rect 82051 6404 82109 6405
rect 82051 6364 82060 6404
rect 82100 6364 82109 6404
rect 82051 6363 82109 6364
rect 82723 6404 82781 6405
rect 82723 6364 82732 6404
rect 82772 6364 82781 6404
rect 82723 6363 82781 6364
rect 83203 6404 83261 6405
rect 83203 6364 83212 6404
rect 83252 6364 83261 6404
rect 83203 6363 83261 6364
rect 83683 6404 83741 6405
rect 83683 6364 83692 6404
rect 83732 6364 83741 6404
rect 83683 6363 83741 6364
rect 84163 6404 84221 6405
rect 84163 6364 84172 6404
rect 84212 6364 84221 6404
rect 84163 6363 84221 6364
rect 84547 6404 84605 6405
rect 84547 6364 84556 6404
rect 84596 6364 84605 6404
rect 84547 6363 84605 6364
rect 85219 6404 85277 6405
rect 85219 6364 85228 6404
rect 85268 6364 85277 6404
rect 85219 6363 85277 6364
rect 85603 6404 85661 6405
rect 85603 6364 85612 6404
rect 85652 6364 85661 6404
rect 85603 6363 85661 6364
rect 86083 6404 86141 6405
rect 86083 6364 86092 6404
rect 86132 6364 86141 6404
rect 86083 6363 86141 6364
rect 86851 6404 86909 6405
rect 86851 6364 86860 6404
rect 86900 6364 86909 6404
rect 86851 6363 86909 6364
rect 87331 6404 87389 6405
rect 87331 6364 87340 6404
rect 87380 6364 87389 6404
rect 87331 6363 87389 6364
rect 87715 6404 87773 6405
rect 87715 6364 87724 6404
rect 87764 6364 87773 6404
rect 87715 6363 87773 6364
rect 88099 6404 88157 6405
rect 88099 6364 88108 6404
rect 88148 6364 88157 6404
rect 88099 6363 88157 6364
rect 89635 6404 89693 6405
rect 89635 6364 89644 6404
rect 89684 6364 89693 6404
rect 89635 6363 89693 6364
rect 90403 6404 90461 6405
rect 90403 6364 90412 6404
rect 90452 6364 90461 6404
rect 90403 6363 90461 6364
rect 90883 6404 90941 6405
rect 90883 6364 90892 6404
rect 90932 6364 90941 6404
rect 90883 6363 90941 6364
rect 91651 6404 91709 6405
rect 91651 6364 91660 6404
rect 91700 6364 91709 6404
rect 91651 6363 91709 6364
rect 92131 6404 92189 6405
rect 92131 6364 92140 6404
rect 92180 6364 92189 6404
rect 92131 6363 92189 6364
rect 92995 6404 93053 6405
rect 92995 6364 93004 6404
rect 93044 6364 93053 6404
rect 92995 6363 93053 6364
rect 93379 6404 93437 6405
rect 93379 6364 93388 6404
rect 93428 6364 93437 6404
rect 93379 6363 93437 6364
rect 93859 6404 93917 6405
rect 93859 6364 93868 6404
rect 93908 6364 93917 6404
rect 93859 6363 93917 6364
rect 94435 6404 94493 6405
rect 94435 6364 94444 6404
rect 94484 6364 94493 6404
rect 94435 6363 94493 6364
rect 95107 6404 95165 6405
rect 95107 6364 95116 6404
rect 95156 6364 95165 6404
rect 95107 6363 95165 6364
rect 96355 6404 96413 6405
rect 96355 6364 96364 6404
rect 96404 6364 96413 6404
rect 96355 6363 96413 6364
rect 96931 6404 96989 6405
rect 96931 6364 96940 6404
rect 96980 6364 96989 6404
rect 96931 6363 96989 6364
rect 74955 6320 74997 6329
rect 74955 6280 74956 6320
rect 74996 6280 74997 6320
rect 74955 6271 74997 6280
rect 79371 6320 79413 6329
rect 79371 6280 79372 6320
rect 79412 6280 79413 6320
rect 79371 6271 79413 6280
rect 89451 6320 89493 6329
rect 89451 6280 89452 6320
rect 89492 6280 89493 6320
rect 89451 6271 89493 6280
rect 74571 6236 74613 6245
rect 74571 6196 74572 6236
rect 74612 6196 74613 6236
rect 74571 6187 74613 6196
rect 95979 6236 96021 6245
rect 95979 6196 95980 6236
rect 96020 6196 96021 6236
rect 95979 6187 96021 6196
rect 576 6068 99516 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 7112 6068
rect 7152 6028 7194 6068
rect 7234 6028 7276 6068
rect 7316 6028 7358 6068
rect 7398 6028 7440 6068
rect 7480 6028 11112 6068
rect 11152 6028 11194 6068
rect 11234 6028 11276 6068
rect 11316 6028 11358 6068
rect 11398 6028 11440 6068
rect 11480 6028 15112 6068
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15480 6028 19112 6068
rect 19152 6028 19194 6068
rect 19234 6028 19276 6068
rect 19316 6028 19358 6068
rect 19398 6028 19440 6068
rect 19480 6028 23112 6068
rect 23152 6028 23194 6068
rect 23234 6028 23276 6068
rect 23316 6028 23358 6068
rect 23398 6028 23440 6068
rect 23480 6028 27112 6068
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27480 6028 31112 6068
rect 31152 6028 31194 6068
rect 31234 6028 31276 6068
rect 31316 6028 31358 6068
rect 31398 6028 31440 6068
rect 31480 6028 35112 6068
rect 35152 6028 35194 6068
rect 35234 6028 35276 6068
rect 35316 6028 35358 6068
rect 35398 6028 35440 6068
rect 35480 6028 39112 6068
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39480 6028 43112 6068
rect 43152 6028 43194 6068
rect 43234 6028 43276 6068
rect 43316 6028 43358 6068
rect 43398 6028 43440 6068
rect 43480 6028 47112 6068
rect 47152 6028 47194 6068
rect 47234 6028 47276 6068
rect 47316 6028 47358 6068
rect 47398 6028 47440 6068
rect 47480 6028 51112 6068
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51480 6028 55112 6068
rect 55152 6028 55194 6068
rect 55234 6028 55276 6068
rect 55316 6028 55358 6068
rect 55398 6028 55440 6068
rect 55480 6028 59112 6068
rect 59152 6028 59194 6068
rect 59234 6028 59276 6068
rect 59316 6028 59358 6068
rect 59398 6028 59440 6068
rect 59480 6028 63112 6068
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63480 6028 67112 6068
rect 67152 6028 67194 6068
rect 67234 6028 67276 6068
rect 67316 6028 67358 6068
rect 67398 6028 67440 6068
rect 67480 6028 71112 6068
rect 71152 6028 71194 6068
rect 71234 6028 71276 6068
rect 71316 6028 71358 6068
rect 71398 6028 71440 6068
rect 71480 6028 75112 6068
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75480 6028 79112 6068
rect 79152 6028 79194 6068
rect 79234 6028 79276 6068
rect 79316 6028 79358 6068
rect 79398 6028 79440 6068
rect 79480 6028 83112 6068
rect 83152 6028 83194 6068
rect 83234 6028 83276 6068
rect 83316 6028 83358 6068
rect 83398 6028 83440 6068
rect 83480 6028 87112 6068
rect 87152 6028 87194 6068
rect 87234 6028 87276 6068
rect 87316 6028 87358 6068
rect 87398 6028 87440 6068
rect 87480 6028 91112 6068
rect 91152 6028 91194 6068
rect 91234 6028 91276 6068
rect 91316 6028 91358 6068
rect 91398 6028 91440 6068
rect 91480 6028 95112 6068
rect 95152 6028 95194 6068
rect 95234 6028 95276 6068
rect 95316 6028 95358 6068
rect 95398 6028 95440 6068
rect 95480 6028 99112 6068
rect 99152 6028 99194 6068
rect 99234 6028 99276 6068
rect 99316 6028 99358 6068
rect 99398 6028 99440 6068
rect 99480 6028 99516 6068
rect 576 6004 99516 6028
rect 75339 5900 75381 5909
rect 75339 5860 75340 5900
rect 75380 5860 75381 5900
rect 75339 5851 75381 5860
rect 76683 5900 76725 5909
rect 76683 5860 76684 5900
rect 76724 5860 76725 5900
rect 76683 5851 76725 5860
rect 78315 5900 78357 5909
rect 78315 5860 78316 5900
rect 78356 5860 78357 5900
rect 78315 5851 78357 5860
rect 78795 5900 78837 5909
rect 78795 5860 78796 5900
rect 78836 5860 78837 5900
rect 78795 5851 78837 5860
rect 80139 5900 80181 5909
rect 80139 5860 80140 5900
rect 80180 5860 80181 5900
rect 80139 5851 80181 5860
rect 80331 5900 80373 5909
rect 80331 5860 80332 5900
rect 80372 5860 80373 5900
rect 80331 5851 80373 5860
rect 81195 5900 81237 5909
rect 81195 5860 81196 5900
rect 81236 5860 81237 5900
rect 81195 5851 81237 5860
rect 82635 5900 82677 5909
rect 82635 5860 82636 5900
rect 82676 5860 82677 5900
rect 82635 5851 82677 5860
rect 83595 5900 83637 5909
rect 83595 5860 83596 5900
rect 83636 5860 83637 5900
rect 83595 5851 83637 5860
rect 85515 5900 85557 5909
rect 85515 5860 85516 5900
rect 85556 5860 85557 5900
rect 85515 5851 85557 5860
rect 86763 5900 86805 5909
rect 86763 5860 86764 5900
rect 86804 5860 86805 5900
rect 86763 5851 86805 5860
rect 87627 5900 87669 5909
rect 87627 5860 87628 5900
rect 87668 5860 87669 5900
rect 87627 5851 87669 5860
rect 89067 5900 89109 5909
rect 89067 5860 89068 5900
rect 89108 5860 89109 5900
rect 89067 5851 89109 5860
rect 89643 5900 89685 5909
rect 89643 5860 89644 5900
rect 89684 5860 89685 5900
rect 89643 5851 89685 5860
rect 90219 5900 90261 5909
rect 90219 5860 90220 5900
rect 90260 5860 90261 5900
rect 90219 5851 90261 5860
rect 91659 5900 91701 5909
rect 91659 5860 91660 5900
rect 91700 5860 91701 5900
rect 91659 5851 91701 5860
rect 92811 5900 92853 5909
rect 92811 5860 92812 5900
rect 92852 5860 92853 5900
rect 92811 5851 92853 5860
rect 93195 5900 93237 5909
rect 93195 5860 93196 5900
rect 93236 5860 93237 5900
rect 93195 5851 93237 5860
rect 93579 5900 93621 5909
rect 93579 5860 93580 5900
rect 93620 5860 93621 5900
rect 93579 5851 93621 5860
rect 93963 5900 94005 5909
rect 93963 5860 93964 5900
rect 94004 5860 94005 5900
rect 93963 5851 94005 5860
rect 95691 5900 95733 5909
rect 95691 5860 95692 5900
rect 95732 5860 95733 5900
rect 95691 5851 95733 5860
rect 95979 5900 96021 5909
rect 95979 5860 95980 5900
rect 96020 5860 96021 5900
rect 95979 5851 96021 5860
rect 98763 5900 98805 5909
rect 98763 5860 98764 5900
rect 98804 5860 98805 5900
rect 98763 5851 98805 5860
rect 1803 5816 1845 5825
rect 1803 5776 1804 5816
rect 1844 5776 1845 5816
rect 1803 5767 1845 5776
rect 835 5732 893 5733
rect 835 5692 844 5732
rect 884 5692 893 5732
rect 835 5691 893 5692
rect 1603 5732 1661 5733
rect 1603 5692 1612 5732
rect 1652 5692 1661 5732
rect 1603 5691 1661 5692
rect 1987 5732 2045 5733
rect 1987 5692 1996 5732
rect 2036 5692 2045 5732
rect 1987 5691 2045 5692
rect 75139 5732 75197 5733
rect 75139 5692 75148 5732
rect 75188 5692 75197 5732
rect 75139 5691 75197 5692
rect 76483 5732 76541 5733
rect 76483 5692 76492 5732
rect 76532 5692 76541 5732
rect 76483 5691 76541 5692
rect 78595 5732 78653 5733
rect 78595 5692 78604 5732
rect 78644 5692 78653 5732
rect 78595 5691 78653 5692
rect 79939 5732 79997 5733
rect 79939 5692 79948 5732
rect 79988 5692 79997 5732
rect 79939 5691 79997 5692
rect 82435 5732 82493 5733
rect 82435 5692 82444 5732
rect 82484 5692 82493 5732
rect 82435 5691 82493 5692
rect 86563 5732 86621 5733
rect 86563 5692 86572 5732
rect 86612 5692 86621 5732
rect 86563 5691 86621 5692
rect 88867 5732 88925 5733
rect 88867 5692 88876 5732
rect 88916 5692 88925 5732
rect 88867 5691 88925 5692
rect 90403 5732 90461 5733
rect 90403 5692 90412 5732
rect 90452 5692 90461 5732
rect 90403 5691 90461 5692
rect 95491 5732 95549 5733
rect 95491 5692 95500 5732
rect 95540 5692 95549 5732
rect 95491 5691 95549 5692
rect 78211 5648 78269 5649
rect 78211 5608 78220 5648
rect 78260 5608 78269 5648
rect 78211 5607 78269 5608
rect 80419 5648 80477 5649
rect 80419 5608 80428 5648
rect 80468 5608 80477 5648
rect 80419 5607 80477 5608
rect 81091 5648 81149 5649
rect 81091 5608 81100 5648
rect 81140 5608 81149 5648
rect 81091 5607 81149 5608
rect 83491 5648 83549 5649
rect 83491 5608 83500 5648
rect 83540 5608 83549 5648
rect 83491 5607 83549 5608
rect 85411 5648 85469 5649
rect 85411 5608 85420 5648
rect 85460 5608 85469 5648
rect 85411 5607 85469 5608
rect 87523 5648 87581 5649
rect 87523 5608 87532 5648
rect 87572 5608 87581 5648
rect 87523 5607 87581 5608
rect 89539 5648 89597 5649
rect 89539 5608 89548 5648
rect 89588 5608 89597 5648
rect 89539 5607 89597 5608
rect 91555 5648 91613 5649
rect 91555 5608 91564 5648
rect 91604 5608 91613 5648
rect 91555 5607 91613 5608
rect 92899 5648 92957 5649
rect 92899 5608 92908 5648
rect 92948 5608 92957 5648
rect 92899 5607 92957 5608
rect 93283 5648 93341 5649
rect 93283 5608 93292 5648
rect 93332 5608 93341 5648
rect 93283 5607 93341 5608
rect 93667 5648 93725 5649
rect 93667 5608 93676 5648
rect 93716 5608 93725 5648
rect 93667 5607 93725 5608
rect 93859 5648 93917 5649
rect 93859 5608 93868 5648
rect 93908 5608 93917 5648
rect 93859 5607 93917 5608
rect 95875 5648 95933 5649
rect 95875 5608 95884 5648
rect 95924 5608 95933 5648
rect 95875 5607 95933 5608
rect 98371 5648 98429 5649
rect 98371 5608 98380 5648
rect 98420 5608 98429 5648
rect 98371 5607 98429 5608
rect 98659 5648 98717 5649
rect 98659 5608 98668 5648
rect 98708 5608 98717 5648
rect 98659 5607 98717 5608
rect 651 5480 693 5489
rect 651 5440 652 5480
rect 692 5440 693 5480
rect 651 5431 693 5440
rect 1419 5480 1461 5489
rect 1419 5440 1420 5480
rect 1460 5440 1461 5480
rect 1419 5431 1461 5440
rect 98283 5480 98325 5489
rect 98283 5440 98284 5480
rect 98324 5440 98325 5480
rect 98283 5431 98325 5440
rect 576 5312 99360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 8352 5312
rect 8392 5272 8434 5312
rect 8474 5272 8516 5312
rect 8556 5272 8598 5312
rect 8638 5272 8680 5312
rect 8720 5272 12352 5312
rect 12392 5272 12434 5312
rect 12474 5272 12516 5312
rect 12556 5272 12598 5312
rect 12638 5272 12680 5312
rect 12720 5272 16352 5312
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16720 5272 20352 5312
rect 20392 5272 20434 5312
rect 20474 5272 20516 5312
rect 20556 5272 20598 5312
rect 20638 5272 20680 5312
rect 20720 5272 24352 5312
rect 24392 5272 24434 5312
rect 24474 5272 24516 5312
rect 24556 5272 24598 5312
rect 24638 5272 24680 5312
rect 24720 5272 28352 5312
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28720 5272 32352 5312
rect 32392 5272 32434 5312
rect 32474 5272 32516 5312
rect 32556 5272 32598 5312
rect 32638 5272 32680 5312
rect 32720 5272 36352 5312
rect 36392 5272 36434 5312
rect 36474 5272 36516 5312
rect 36556 5272 36598 5312
rect 36638 5272 36680 5312
rect 36720 5272 40352 5312
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40720 5272 44352 5312
rect 44392 5272 44434 5312
rect 44474 5272 44516 5312
rect 44556 5272 44598 5312
rect 44638 5272 44680 5312
rect 44720 5272 48352 5312
rect 48392 5272 48434 5312
rect 48474 5272 48516 5312
rect 48556 5272 48598 5312
rect 48638 5272 48680 5312
rect 48720 5272 52352 5312
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52720 5272 56352 5312
rect 56392 5272 56434 5312
rect 56474 5272 56516 5312
rect 56556 5272 56598 5312
rect 56638 5272 56680 5312
rect 56720 5272 60352 5312
rect 60392 5272 60434 5312
rect 60474 5272 60516 5312
rect 60556 5272 60598 5312
rect 60638 5272 60680 5312
rect 60720 5272 64352 5312
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64720 5272 68352 5312
rect 68392 5272 68434 5312
rect 68474 5272 68516 5312
rect 68556 5272 68598 5312
rect 68638 5272 68680 5312
rect 68720 5272 72352 5312
rect 72392 5272 72434 5312
rect 72474 5272 72516 5312
rect 72556 5272 72598 5312
rect 72638 5272 72680 5312
rect 72720 5272 76352 5312
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76720 5272 80352 5312
rect 80392 5272 80434 5312
rect 80474 5272 80516 5312
rect 80556 5272 80598 5312
rect 80638 5272 80680 5312
rect 80720 5272 84352 5312
rect 84392 5272 84434 5312
rect 84474 5272 84516 5312
rect 84556 5272 84598 5312
rect 84638 5272 84680 5312
rect 84720 5272 88352 5312
rect 88392 5272 88434 5312
rect 88474 5272 88516 5312
rect 88556 5272 88598 5312
rect 88638 5272 88680 5312
rect 88720 5272 92352 5312
rect 92392 5272 92434 5312
rect 92474 5272 92516 5312
rect 92556 5272 92598 5312
rect 92638 5272 92680 5312
rect 92720 5272 96352 5312
rect 96392 5272 96434 5312
rect 96474 5272 96516 5312
rect 96556 5272 96598 5312
rect 96638 5272 96680 5312
rect 96720 5272 99360 5312
rect 576 5248 99360 5272
rect 835 4892 893 4893
rect 835 4852 844 4892
rect 884 4852 893 4892
rect 835 4851 893 4852
rect 1411 4892 1469 4893
rect 1411 4852 1420 4892
rect 1460 4852 1469 4892
rect 1411 4851 1469 4852
rect 1795 4892 1853 4893
rect 1795 4852 1804 4892
rect 1844 4852 1853 4892
rect 1795 4851 1853 4852
rect 2179 4892 2237 4893
rect 2179 4852 2188 4892
rect 2228 4852 2237 4892
rect 2179 4851 2237 4852
rect 96931 4892 96989 4893
rect 96931 4852 96940 4892
rect 96980 4852 96989 4892
rect 96931 4851 96989 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 97131 4808 97173 4817
rect 97131 4768 97132 4808
rect 97172 4768 97173 4808
rect 97131 4759 97173 4768
rect 1227 4724 1269 4733
rect 1227 4684 1228 4724
rect 1268 4684 1269 4724
rect 1227 4675 1269 4684
rect 1611 4724 1653 4733
rect 1611 4684 1612 4724
rect 1652 4684 1653 4724
rect 1611 4675 1653 4684
rect 1995 4724 2037 4733
rect 1995 4684 1996 4724
rect 2036 4684 2037 4724
rect 1995 4675 2037 4684
rect 576 4556 99516 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 7112 4556
rect 7152 4516 7194 4556
rect 7234 4516 7276 4556
rect 7316 4516 7358 4556
rect 7398 4516 7440 4556
rect 7480 4516 11112 4556
rect 11152 4516 11194 4556
rect 11234 4516 11276 4556
rect 11316 4516 11358 4556
rect 11398 4516 11440 4556
rect 11480 4516 15112 4556
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15480 4516 19112 4556
rect 19152 4516 19194 4556
rect 19234 4516 19276 4556
rect 19316 4516 19358 4556
rect 19398 4516 19440 4556
rect 19480 4516 23112 4556
rect 23152 4516 23194 4556
rect 23234 4516 23276 4556
rect 23316 4516 23358 4556
rect 23398 4516 23440 4556
rect 23480 4516 27112 4556
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27480 4516 31112 4556
rect 31152 4516 31194 4556
rect 31234 4516 31276 4556
rect 31316 4516 31358 4556
rect 31398 4516 31440 4556
rect 31480 4516 35112 4556
rect 35152 4516 35194 4556
rect 35234 4516 35276 4556
rect 35316 4516 35358 4556
rect 35398 4516 35440 4556
rect 35480 4516 39112 4556
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39480 4516 43112 4556
rect 43152 4516 43194 4556
rect 43234 4516 43276 4556
rect 43316 4516 43358 4556
rect 43398 4516 43440 4556
rect 43480 4516 47112 4556
rect 47152 4516 47194 4556
rect 47234 4516 47276 4556
rect 47316 4516 47358 4556
rect 47398 4516 47440 4556
rect 47480 4516 51112 4556
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51480 4516 55112 4556
rect 55152 4516 55194 4556
rect 55234 4516 55276 4556
rect 55316 4516 55358 4556
rect 55398 4516 55440 4556
rect 55480 4516 59112 4556
rect 59152 4516 59194 4556
rect 59234 4516 59276 4556
rect 59316 4516 59358 4556
rect 59398 4516 59440 4556
rect 59480 4516 63112 4556
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63480 4516 67112 4556
rect 67152 4516 67194 4556
rect 67234 4516 67276 4556
rect 67316 4516 67358 4556
rect 67398 4516 67440 4556
rect 67480 4516 71112 4556
rect 71152 4516 71194 4556
rect 71234 4516 71276 4556
rect 71316 4516 71358 4556
rect 71398 4516 71440 4556
rect 71480 4516 75112 4556
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75480 4516 79112 4556
rect 79152 4516 79194 4556
rect 79234 4516 79276 4556
rect 79316 4516 79358 4556
rect 79398 4516 79440 4556
rect 79480 4516 83112 4556
rect 83152 4516 83194 4556
rect 83234 4516 83276 4556
rect 83316 4516 83358 4556
rect 83398 4516 83440 4556
rect 83480 4516 87112 4556
rect 87152 4516 87194 4556
rect 87234 4516 87276 4556
rect 87316 4516 87358 4556
rect 87398 4516 87440 4556
rect 87480 4516 91112 4556
rect 91152 4516 91194 4556
rect 91234 4516 91276 4556
rect 91316 4516 91358 4556
rect 91398 4516 91440 4556
rect 91480 4516 95112 4556
rect 95152 4516 95194 4556
rect 95234 4516 95276 4556
rect 95316 4516 95358 4556
rect 95398 4516 95440 4556
rect 95480 4516 99112 4556
rect 99152 4516 99194 4556
rect 99234 4516 99276 4556
rect 99316 4516 99358 4556
rect 99398 4516 99440 4556
rect 99480 4516 99516 4556
rect 576 4492 99516 4516
rect 835 4220 893 4221
rect 835 4180 844 4220
rect 884 4180 893 4220
rect 835 4179 893 4180
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 576 3800 99360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 8352 3800
rect 8392 3760 8434 3800
rect 8474 3760 8516 3800
rect 8556 3760 8598 3800
rect 8638 3760 8680 3800
rect 8720 3760 12352 3800
rect 12392 3760 12434 3800
rect 12474 3760 12516 3800
rect 12556 3760 12598 3800
rect 12638 3760 12680 3800
rect 12720 3760 16352 3800
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16720 3760 20352 3800
rect 20392 3760 20434 3800
rect 20474 3760 20516 3800
rect 20556 3760 20598 3800
rect 20638 3760 20680 3800
rect 20720 3760 24352 3800
rect 24392 3760 24434 3800
rect 24474 3760 24516 3800
rect 24556 3760 24598 3800
rect 24638 3760 24680 3800
rect 24720 3760 28352 3800
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28720 3760 32352 3800
rect 32392 3760 32434 3800
rect 32474 3760 32516 3800
rect 32556 3760 32598 3800
rect 32638 3760 32680 3800
rect 32720 3760 36352 3800
rect 36392 3760 36434 3800
rect 36474 3760 36516 3800
rect 36556 3760 36598 3800
rect 36638 3760 36680 3800
rect 36720 3760 40352 3800
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40720 3760 44352 3800
rect 44392 3760 44434 3800
rect 44474 3760 44516 3800
rect 44556 3760 44598 3800
rect 44638 3760 44680 3800
rect 44720 3760 48352 3800
rect 48392 3760 48434 3800
rect 48474 3760 48516 3800
rect 48556 3760 48598 3800
rect 48638 3760 48680 3800
rect 48720 3760 52352 3800
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52720 3760 56352 3800
rect 56392 3760 56434 3800
rect 56474 3760 56516 3800
rect 56556 3760 56598 3800
rect 56638 3760 56680 3800
rect 56720 3760 60352 3800
rect 60392 3760 60434 3800
rect 60474 3760 60516 3800
rect 60556 3760 60598 3800
rect 60638 3760 60680 3800
rect 60720 3760 64352 3800
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64720 3760 68352 3800
rect 68392 3760 68434 3800
rect 68474 3760 68516 3800
rect 68556 3760 68598 3800
rect 68638 3760 68680 3800
rect 68720 3760 72352 3800
rect 72392 3760 72434 3800
rect 72474 3760 72516 3800
rect 72556 3760 72598 3800
rect 72638 3760 72680 3800
rect 72720 3760 76352 3800
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76720 3760 80352 3800
rect 80392 3760 80434 3800
rect 80474 3760 80516 3800
rect 80556 3760 80598 3800
rect 80638 3760 80680 3800
rect 80720 3760 84352 3800
rect 84392 3760 84434 3800
rect 84474 3760 84516 3800
rect 84556 3760 84598 3800
rect 84638 3760 84680 3800
rect 84720 3760 88352 3800
rect 88392 3760 88434 3800
rect 88474 3760 88516 3800
rect 88556 3760 88598 3800
rect 88638 3760 88680 3800
rect 88720 3760 92352 3800
rect 92392 3760 92434 3800
rect 92474 3760 92516 3800
rect 92556 3760 92598 3800
rect 92638 3760 92680 3800
rect 92720 3760 96352 3800
rect 96392 3760 96434 3800
rect 96474 3760 96516 3800
rect 96556 3760 96598 3800
rect 96638 3760 96680 3800
rect 96720 3760 99360 3800
rect 576 3736 99360 3760
rect 835 3380 893 3381
rect 835 3340 844 3380
rect 884 3340 893 3380
rect 835 3339 893 3340
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 576 3044 99516 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 7112 3044
rect 7152 3004 7194 3044
rect 7234 3004 7276 3044
rect 7316 3004 7358 3044
rect 7398 3004 7440 3044
rect 7480 3004 11112 3044
rect 11152 3004 11194 3044
rect 11234 3004 11276 3044
rect 11316 3004 11358 3044
rect 11398 3004 11440 3044
rect 11480 3004 15112 3044
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15480 3004 19112 3044
rect 19152 3004 19194 3044
rect 19234 3004 19276 3044
rect 19316 3004 19358 3044
rect 19398 3004 19440 3044
rect 19480 3004 23112 3044
rect 23152 3004 23194 3044
rect 23234 3004 23276 3044
rect 23316 3004 23358 3044
rect 23398 3004 23440 3044
rect 23480 3004 27112 3044
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27480 3004 31112 3044
rect 31152 3004 31194 3044
rect 31234 3004 31276 3044
rect 31316 3004 31358 3044
rect 31398 3004 31440 3044
rect 31480 3004 35112 3044
rect 35152 3004 35194 3044
rect 35234 3004 35276 3044
rect 35316 3004 35358 3044
rect 35398 3004 35440 3044
rect 35480 3004 39112 3044
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39480 3004 43112 3044
rect 43152 3004 43194 3044
rect 43234 3004 43276 3044
rect 43316 3004 43358 3044
rect 43398 3004 43440 3044
rect 43480 3004 47112 3044
rect 47152 3004 47194 3044
rect 47234 3004 47276 3044
rect 47316 3004 47358 3044
rect 47398 3004 47440 3044
rect 47480 3004 51112 3044
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51480 3004 55112 3044
rect 55152 3004 55194 3044
rect 55234 3004 55276 3044
rect 55316 3004 55358 3044
rect 55398 3004 55440 3044
rect 55480 3004 59112 3044
rect 59152 3004 59194 3044
rect 59234 3004 59276 3044
rect 59316 3004 59358 3044
rect 59398 3004 59440 3044
rect 59480 3004 63112 3044
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63480 3004 67112 3044
rect 67152 3004 67194 3044
rect 67234 3004 67276 3044
rect 67316 3004 67358 3044
rect 67398 3004 67440 3044
rect 67480 3004 71112 3044
rect 71152 3004 71194 3044
rect 71234 3004 71276 3044
rect 71316 3004 71358 3044
rect 71398 3004 71440 3044
rect 71480 3004 75112 3044
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75480 3004 79112 3044
rect 79152 3004 79194 3044
rect 79234 3004 79276 3044
rect 79316 3004 79358 3044
rect 79398 3004 79440 3044
rect 79480 3004 83112 3044
rect 83152 3004 83194 3044
rect 83234 3004 83276 3044
rect 83316 3004 83358 3044
rect 83398 3004 83440 3044
rect 83480 3004 87112 3044
rect 87152 3004 87194 3044
rect 87234 3004 87276 3044
rect 87316 3004 87358 3044
rect 87398 3004 87440 3044
rect 87480 3004 91112 3044
rect 91152 3004 91194 3044
rect 91234 3004 91276 3044
rect 91316 3004 91358 3044
rect 91398 3004 91440 3044
rect 91480 3004 95112 3044
rect 95152 3004 95194 3044
rect 95234 3004 95276 3044
rect 95316 3004 95358 3044
rect 95398 3004 95440 3044
rect 95480 3004 99112 3044
rect 99152 3004 99194 3044
rect 99234 3004 99276 3044
rect 99316 3004 99358 3044
rect 99398 3004 99440 3044
rect 99480 3004 99516 3044
rect 576 2980 99516 3004
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 576 2288 99360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 8352 2288
rect 8392 2248 8434 2288
rect 8474 2248 8516 2288
rect 8556 2248 8598 2288
rect 8638 2248 8680 2288
rect 8720 2248 12352 2288
rect 12392 2248 12434 2288
rect 12474 2248 12516 2288
rect 12556 2248 12598 2288
rect 12638 2248 12680 2288
rect 12720 2248 16352 2288
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16720 2248 20352 2288
rect 20392 2248 20434 2288
rect 20474 2248 20516 2288
rect 20556 2248 20598 2288
rect 20638 2248 20680 2288
rect 20720 2248 24352 2288
rect 24392 2248 24434 2288
rect 24474 2248 24516 2288
rect 24556 2248 24598 2288
rect 24638 2248 24680 2288
rect 24720 2248 28352 2288
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28720 2248 32352 2288
rect 32392 2248 32434 2288
rect 32474 2248 32516 2288
rect 32556 2248 32598 2288
rect 32638 2248 32680 2288
rect 32720 2248 36352 2288
rect 36392 2248 36434 2288
rect 36474 2248 36516 2288
rect 36556 2248 36598 2288
rect 36638 2248 36680 2288
rect 36720 2248 40352 2288
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40720 2248 44352 2288
rect 44392 2248 44434 2288
rect 44474 2248 44516 2288
rect 44556 2248 44598 2288
rect 44638 2248 44680 2288
rect 44720 2248 48352 2288
rect 48392 2248 48434 2288
rect 48474 2248 48516 2288
rect 48556 2248 48598 2288
rect 48638 2248 48680 2288
rect 48720 2248 52352 2288
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52720 2248 56352 2288
rect 56392 2248 56434 2288
rect 56474 2248 56516 2288
rect 56556 2248 56598 2288
rect 56638 2248 56680 2288
rect 56720 2248 60352 2288
rect 60392 2248 60434 2288
rect 60474 2248 60516 2288
rect 60556 2248 60598 2288
rect 60638 2248 60680 2288
rect 60720 2248 64352 2288
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64720 2248 68352 2288
rect 68392 2248 68434 2288
rect 68474 2248 68516 2288
rect 68556 2248 68598 2288
rect 68638 2248 68680 2288
rect 68720 2248 72352 2288
rect 72392 2248 72434 2288
rect 72474 2248 72516 2288
rect 72556 2248 72598 2288
rect 72638 2248 72680 2288
rect 72720 2248 76352 2288
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76720 2248 80352 2288
rect 80392 2248 80434 2288
rect 80474 2248 80516 2288
rect 80556 2248 80598 2288
rect 80638 2248 80680 2288
rect 80720 2248 84352 2288
rect 84392 2248 84434 2288
rect 84474 2248 84516 2288
rect 84556 2248 84598 2288
rect 84638 2248 84680 2288
rect 84720 2248 88352 2288
rect 88392 2248 88434 2288
rect 88474 2248 88516 2288
rect 88556 2248 88598 2288
rect 88638 2248 88680 2288
rect 88720 2248 92352 2288
rect 92392 2248 92434 2288
rect 92474 2248 92516 2288
rect 92556 2248 92598 2288
rect 92638 2248 92680 2288
rect 92720 2248 96352 2288
rect 96392 2248 96434 2288
rect 96474 2248 96516 2288
rect 96556 2248 96598 2288
rect 96638 2248 96680 2288
rect 96720 2248 99360 2288
rect 576 2224 99360 2248
rect 576 1532 99516 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 7112 1532
rect 7152 1492 7194 1532
rect 7234 1492 7276 1532
rect 7316 1492 7358 1532
rect 7398 1492 7440 1532
rect 7480 1492 11112 1532
rect 11152 1492 11194 1532
rect 11234 1492 11276 1532
rect 11316 1492 11358 1532
rect 11398 1492 11440 1532
rect 11480 1492 15112 1532
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15480 1492 19112 1532
rect 19152 1492 19194 1532
rect 19234 1492 19276 1532
rect 19316 1492 19358 1532
rect 19398 1492 19440 1532
rect 19480 1492 23112 1532
rect 23152 1492 23194 1532
rect 23234 1492 23276 1532
rect 23316 1492 23358 1532
rect 23398 1492 23440 1532
rect 23480 1492 27112 1532
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27480 1492 31112 1532
rect 31152 1492 31194 1532
rect 31234 1492 31276 1532
rect 31316 1492 31358 1532
rect 31398 1492 31440 1532
rect 31480 1492 35112 1532
rect 35152 1492 35194 1532
rect 35234 1492 35276 1532
rect 35316 1492 35358 1532
rect 35398 1492 35440 1532
rect 35480 1492 39112 1532
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39480 1492 43112 1532
rect 43152 1492 43194 1532
rect 43234 1492 43276 1532
rect 43316 1492 43358 1532
rect 43398 1492 43440 1532
rect 43480 1492 47112 1532
rect 47152 1492 47194 1532
rect 47234 1492 47276 1532
rect 47316 1492 47358 1532
rect 47398 1492 47440 1532
rect 47480 1492 51112 1532
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51480 1492 55112 1532
rect 55152 1492 55194 1532
rect 55234 1492 55276 1532
rect 55316 1492 55358 1532
rect 55398 1492 55440 1532
rect 55480 1492 59112 1532
rect 59152 1492 59194 1532
rect 59234 1492 59276 1532
rect 59316 1492 59358 1532
rect 59398 1492 59440 1532
rect 59480 1492 63112 1532
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63480 1492 67112 1532
rect 67152 1492 67194 1532
rect 67234 1492 67276 1532
rect 67316 1492 67358 1532
rect 67398 1492 67440 1532
rect 67480 1492 71112 1532
rect 71152 1492 71194 1532
rect 71234 1492 71276 1532
rect 71316 1492 71358 1532
rect 71398 1492 71440 1532
rect 71480 1492 75112 1532
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75480 1492 79112 1532
rect 79152 1492 79194 1532
rect 79234 1492 79276 1532
rect 79316 1492 79358 1532
rect 79398 1492 79440 1532
rect 79480 1492 83112 1532
rect 83152 1492 83194 1532
rect 83234 1492 83276 1532
rect 83316 1492 83358 1532
rect 83398 1492 83440 1532
rect 83480 1492 87112 1532
rect 87152 1492 87194 1532
rect 87234 1492 87276 1532
rect 87316 1492 87358 1532
rect 87398 1492 87440 1532
rect 87480 1492 91112 1532
rect 91152 1492 91194 1532
rect 91234 1492 91276 1532
rect 91316 1492 91358 1532
rect 91398 1492 91440 1532
rect 91480 1492 95112 1532
rect 95152 1492 95194 1532
rect 95234 1492 95276 1532
rect 95316 1492 95358 1532
rect 95398 1492 95440 1532
rect 95480 1492 99112 1532
rect 99152 1492 99194 1532
rect 99234 1492 99276 1532
rect 99316 1492 99358 1532
rect 99398 1492 99440 1532
rect 99480 1492 99516 1532
rect 576 1468 99516 1492
rect 576 776 99360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 8352 776
rect 8392 736 8434 776
rect 8474 736 8516 776
rect 8556 736 8598 776
rect 8638 736 8680 776
rect 8720 736 12352 776
rect 12392 736 12434 776
rect 12474 736 12516 776
rect 12556 736 12598 776
rect 12638 736 12680 776
rect 12720 736 16352 776
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16720 736 20352 776
rect 20392 736 20434 776
rect 20474 736 20516 776
rect 20556 736 20598 776
rect 20638 736 20680 776
rect 20720 736 24352 776
rect 24392 736 24434 776
rect 24474 736 24516 776
rect 24556 736 24598 776
rect 24638 736 24680 776
rect 24720 736 28352 776
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28720 736 32352 776
rect 32392 736 32434 776
rect 32474 736 32516 776
rect 32556 736 32598 776
rect 32638 736 32680 776
rect 32720 736 36352 776
rect 36392 736 36434 776
rect 36474 736 36516 776
rect 36556 736 36598 776
rect 36638 736 36680 776
rect 36720 736 40352 776
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40720 736 44352 776
rect 44392 736 44434 776
rect 44474 736 44516 776
rect 44556 736 44598 776
rect 44638 736 44680 776
rect 44720 736 48352 776
rect 48392 736 48434 776
rect 48474 736 48516 776
rect 48556 736 48598 776
rect 48638 736 48680 776
rect 48720 736 52352 776
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52720 736 56352 776
rect 56392 736 56434 776
rect 56474 736 56516 776
rect 56556 736 56598 776
rect 56638 736 56680 776
rect 56720 736 60352 776
rect 60392 736 60434 776
rect 60474 736 60516 776
rect 60556 736 60598 776
rect 60638 736 60680 776
rect 60720 736 64352 776
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64720 736 68352 776
rect 68392 736 68434 776
rect 68474 736 68516 776
rect 68556 736 68598 776
rect 68638 736 68680 776
rect 68720 736 72352 776
rect 72392 736 72434 776
rect 72474 736 72516 776
rect 72556 736 72598 776
rect 72638 736 72680 776
rect 72720 736 76352 776
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76720 736 80352 776
rect 80392 736 80434 776
rect 80474 736 80516 776
rect 80556 736 80598 776
rect 80638 736 80680 776
rect 80720 736 84352 776
rect 84392 736 84434 776
rect 84474 736 84516 776
rect 84556 736 84598 776
rect 84638 736 84680 776
rect 84720 736 88352 776
rect 88392 736 88434 776
rect 88474 736 88516 776
rect 88556 736 88598 776
rect 88638 736 88680 776
rect 88720 736 92352 776
rect 92392 736 92434 776
rect 92474 736 92516 776
rect 92556 736 92598 776
rect 92638 736 92680 776
rect 92720 736 96352 776
rect 96392 736 96434 776
rect 96474 736 96516 776
rect 96556 736 96598 776
rect 96638 736 96680 776
rect 96720 736 99360 776
rect 576 712 99360 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 8352 38536 8392 38576
rect 8434 38536 8474 38576
rect 8516 38536 8556 38576
rect 8598 38536 8638 38576
rect 8680 38536 8720 38576
rect 12352 38536 12392 38576
rect 12434 38536 12474 38576
rect 12516 38536 12556 38576
rect 12598 38536 12638 38576
rect 12680 38536 12720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 20352 38536 20392 38576
rect 20434 38536 20474 38576
rect 20516 38536 20556 38576
rect 20598 38536 20638 38576
rect 20680 38536 20720 38576
rect 24352 38536 24392 38576
rect 24434 38536 24474 38576
rect 24516 38536 24556 38576
rect 24598 38536 24638 38576
rect 24680 38536 24720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 32352 38536 32392 38576
rect 32434 38536 32474 38576
rect 32516 38536 32556 38576
rect 32598 38536 32638 38576
rect 32680 38536 32720 38576
rect 36352 38536 36392 38576
rect 36434 38536 36474 38576
rect 36516 38536 36556 38576
rect 36598 38536 36638 38576
rect 36680 38536 36720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 44352 38536 44392 38576
rect 44434 38536 44474 38576
rect 44516 38536 44556 38576
rect 44598 38536 44638 38576
rect 44680 38536 44720 38576
rect 48352 38536 48392 38576
rect 48434 38536 48474 38576
rect 48516 38536 48556 38576
rect 48598 38536 48638 38576
rect 48680 38536 48720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 56352 38536 56392 38576
rect 56434 38536 56474 38576
rect 56516 38536 56556 38576
rect 56598 38536 56638 38576
rect 56680 38536 56720 38576
rect 60352 38536 60392 38576
rect 60434 38536 60474 38576
rect 60516 38536 60556 38576
rect 60598 38536 60638 38576
rect 60680 38536 60720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 68352 38536 68392 38576
rect 68434 38536 68474 38576
rect 68516 38536 68556 38576
rect 68598 38536 68638 38576
rect 68680 38536 68720 38576
rect 72352 38536 72392 38576
rect 72434 38536 72474 38576
rect 72516 38536 72556 38576
rect 72598 38536 72638 38576
rect 72680 38536 72720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 80352 38536 80392 38576
rect 80434 38536 80474 38576
rect 80516 38536 80556 38576
rect 80598 38536 80638 38576
rect 80680 38536 80720 38576
rect 84352 38536 84392 38576
rect 84434 38536 84474 38576
rect 84516 38536 84556 38576
rect 84598 38536 84638 38576
rect 84680 38536 84720 38576
rect 88352 38536 88392 38576
rect 88434 38536 88474 38576
rect 88516 38536 88556 38576
rect 88598 38536 88638 38576
rect 88680 38536 88720 38576
rect 92352 38536 92392 38576
rect 92434 38536 92474 38576
rect 92516 38536 92556 38576
rect 92598 38536 92638 38576
rect 92680 38536 92720 38576
rect 96352 38536 96392 38576
rect 96434 38536 96474 38576
rect 96516 38536 96556 38576
rect 96598 38536 96638 38576
rect 96680 38536 96720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 7112 37780 7152 37820
rect 7194 37780 7234 37820
rect 7276 37780 7316 37820
rect 7358 37780 7398 37820
rect 7440 37780 7480 37820
rect 11112 37780 11152 37820
rect 11194 37780 11234 37820
rect 11276 37780 11316 37820
rect 11358 37780 11398 37820
rect 11440 37780 11480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 19112 37780 19152 37820
rect 19194 37780 19234 37820
rect 19276 37780 19316 37820
rect 19358 37780 19398 37820
rect 19440 37780 19480 37820
rect 23112 37780 23152 37820
rect 23194 37780 23234 37820
rect 23276 37780 23316 37820
rect 23358 37780 23398 37820
rect 23440 37780 23480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 31112 37780 31152 37820
rect 31194 37780 31234 37820
rect 31276 37780 31316 37820
rect 31358 37780 31398 37820
rect 31440 37780 31480 37820
rect 35112 37780 35152 37820
rect 35194 37780 35234 37820
rect 35276 37780 35316 37820
rect 35358 37780 35398 37820
rect 35440 37780 35480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 43112 37780 43152 37820
rect 43194 37780 43234 37820
rect 43276 37780 43316 37820
rect 43358 37780 43398 37820
rect 43440 37780 43480 37820
rect 47112 37780 47152 37820
rect 47194 37780 47234 37820
rect 47276 37780 47316 37820
rect 47358 37780 47398 37820
rect 47440 37780 47480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 55112 37780 55152 37820
rect 55194 37780 55234 37820
rect 55276 37780 55316 37820
rect 55358 37780 55398 37820
rect 55440 37780 55480 37820
rect 59112 37780 59152 37820
rect 59194 37780 59234 37820
rect 59276 37780 59316 37820
rect 59358 37780 59398 37820
rect 59440 37780 59480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 67112 37780 67152 37820
rect 67194 37780 67234 37820
rect 67276 37780 67316 37820
rect 67358 37780 67398 37820
rect 67440 37780 67480 37820
rect 71112 37780 71152 37820
rect 71194 37780 71234 37820
rect 71276 37780 71316 37820
rect 71358 37780 71398 37820
rect 71440 37780 71480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 79112 37780 79152 37820
rect 79194 37780 79234 37820
rect 79276 37780 79316 37820
rect 79358 37780 79398 37820
rect 79440 37780 79480 37820
rect 83112 37780 83152 37820
rect 83194 37780 83234 37820
rect 83276 37780 83316 37820
rect 83358 37780 83398 37820
rect 83440 37780 83480 37820
rect 87112 37780 87152 37820
rect 87194 37780 87234 37820
rect 87276 37780 87316 37820
rect 87358 37780 87398 37820
rect 87440 37780 87480 37820
rect 91112 37780 91152 37820
rect 91194 37780 91234 37820
rect 91276 37780 91316 37820
rect 91358 37780 91398 37820
rect 91440 37780 91480 37820
rect 95112 37780 95152 37820
rect 95194 37780 95234 37820
rect 95276 37780 95316 37820
rect 95358 37780 95398 37820
rect 95440 37780 95480 37820
rect 99112 37780 99152 37820
rect 99194 37780 99234 37820
rect 99276 37780 99316 37820
rect 99358 37780 99398 37820
rect 99440 37780 99480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 8352 37024 8392 37064
rect 8434 37024 8474 37064
rect 8516 37024 8556 37064
rect 8598 37024 8638 37064
rect 8680 37024 8720 37064
rect 12352 37024 12392 37064
rect 12434 37024 12474 37064
rect 12516 37024 12556 37064
rect 12598 37024 12638 37064
rect 12680 37024 12720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 20352 37024 20392 37064
rect 20434 37024 20474 37064
rect 20516 37024 20556 37064
rect 20598 37024 20638 37064
rect 20680 37024 20720 37064
rect 24352 37024 24392 37064
rect 24434 37024 24474 37064
rect 24516 37024 24556 37064
rect 24598 37024 24638 37064
rect 24680 37024 24720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 32352 37024 32392 37064
rect 32434 37024 32474 37064
rect 32516 37024 32556 37064
rect 32598 37024 32638 37064
rect 32680 37024 32720 37064
rect 36352 37024 36392 37064
rect 36434 37024 36474 37064
rect 36516 37024 36556 37064
rect 36598 37024 36638 37064
rect 36680 37024 36720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 44352 37024 44392 37064
rect 44434 37024 44474 37064
rect 44516 37024 44556 37064
rect 44598 37024 44638 37064
rect 44680 37024 44720 37064
rect 48352 37024 48392 37064
rect 48434 37024 48474 37064
rect 48516 37024 48556 37064
rect 48598 37024 48638 37064
rect 48680 37024 48720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 56352 37024 56392 37064
rect 56434 37024 56474 37064
rect 56516 37024 56556 37064
rect 56598 37024 56638 37064
rect 56680 37024 56720 37064
rect 60352 37024 60392 37064
rect 60434 37024 60474 37064
rect 60516 37024 60556 37064
rect 60598 37024 60638 37064
rect 60680 37024 60720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 68352 37024 68392 37064
rect 68434 37024 68474 37064
rect 68516 37024 68556 37064
rect 68598 37024 68638 37064
rect 68680 37024 68720 37064
rect 72352 37024 72392 37064
rect 72434 37024 72474 37064
rect 72516 37024 72556 37064
rect 72598 37024 72638 37064
rect 72680 37024 72720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 80352 37024 80392 37064
rect 80434 37024 80474 37064
rect 80516 37024 80556 37064
rect 80598 37024 80638 37064
rect 80680 37024 80720 37064
rect 84352 37024 84392 37064
rect 84434 37024 84474 37064
rect 84516 37024 84556 37064
rect 84598 37024 84638 37064
rect 84680 37024 84720 37064
rect 88352 37024 88392 37064
rect 88434 37024 88474 37064
rect 88516 37024 88556 37064
rect 88598 37024 88638 37064
rect 88680 37024 88720 37064
rect 92352 37024 92392 37064
rect 92434 37024 92474 37064
rect 92516 37024 92556 37064
rect 92598 37024 92638 37064
rect 92680 37024 92720 37064
rect 96352 37024 96392 37064
rect 96434 37024 96474 37064
rect 96516 37024 96556 37064
rect 96598 37024 96638 37064
rect 96680 37024 96720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 7112 36268 7152 36308
rect 7194 36268 7234 36308
rect 7276 36268 7316 36308
rect 7358 36268 7398 36308
rect 7440 36268 7480 36308
rect 11112 36268 11152 36308
rect 11194 36268 11234 36308
rect 11276 36268 11316 36308
rect 11358 36268 11398 36308
rect 11440 36268 11480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 19112 36268 19152 36308
rect 19194 36268 19234 36308
rect 19276 36268 19316 36308
rect 19358 36268 19398 36308
rect 19440 36268 19480 36308
rect 23112 36268 23152 36308
rect 23194 36268 23234 36308
rect 23276 36268 23316 36308
rect 23358 36268 23398 36308
rect 23440 36268 23480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 31112 36268 31152 36308
rect 31194 36268 31234 36308
rect 31276 36268 31316 36308
rect 31358 36268 31398 36308
rect 31440 36268 31480 36308
rect 35112 36268 35152 36308
rect 35194 36268 35234 36308
rect 35276 36268 35316 36308
rect 35358 36268 35398 36308
rect 35440 36268 35480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 43112 36268 43152 36308
rect 43194 36268 43234 36308
rect 43276 36268 43316 36308
rect 43358 36268 43398 36308
rect 43440 36268 43480 36308
rect 47112 36268 47152 36308
rect 47194 36268 47234 36308
rect 47276 36268 47316 36308
rect 47358 36268 47398 36308
rect 47440 36268 47480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 55112 36268 55152 36308
rect 55194 36268 55234 36308
rect 55276 36268 55316 36308
rect 55358 36268 55398 36308
rect 55440 36268 55480 36308
rect 59112 36268 59152 36308
rect 59194 36268 59234 36308
rect 59276 36268 59316 36308
rect 59358 36268 59398 36308
rect 59440 36268 59480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 67112 36268 67152 36308
rect 67194 36268 67234 36308
rect 67276 36268 67316 36308
rect 67358 36268 67398 36308
rect 67440 36268 67480 36308
rect 71112 36268 71152 36308
rect 71194 36268 71234 36308
rect 71276 36268 71316 36308
rect 71358 36268 71398 36308
rect 71440 36268 71480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 79112 36268 79152 36308
rect 79194 36268 79234 36308
rect 79276 36268 79316 36308
rect 79358 36268 79398 36308
rect 79440 36268 79480 36308
rect 83112 36268 83152 36308
rect 83194 36268 83234 36308
rect 83276 36268 83316 36308
rect 83358 36268 83398 36308
rect 83440 36268 83480 36308
rect 87112 36268 87152 36308
rect 87194 36268 87234 36308
rect 87276 36268 87316 36308
rect 87358 36268 87398 36308
rect 87440 36268 87480 36308
rect 91112 36268 91152 36308
rect 91194 36268 91234 36308
rect 91276 36268 91316 36308
rect 91358 36268 91398 36308
rect 91440 36268 91480 36308
rect 95112 36268 95152 36308
rect 95194 36268 95234 36308
rect 95276 36268 95316 36308
rect 95358 36268 95398 36308
rect 95440 36268 95480 36308
rect 99112 36268 99152 36308
rect 99194 36268 99234 36308
rect 99276 36268 99316 36308
rect 99358 36268 99398 36308
rect 99440 36268 99480 36308
rect 74860 35932 74900 35972
rect 76588 35932 76628 35972
rect 77452 35932 77492 35972
rect 78604 35932 78644 35972
rect 79372 35932 79412 35972
rect 81388 35932 81428 35972
rect 85036 35932 85076 35972
rect 85420 35932 85460 35972
rect 92236 35932 92276 35972
rect 80236 35848 80276 35888
rect 86572 35848 86612 35888
rect 87820 35848 87860 35888
rect 89836 35848 89876 35888
rect 90220 35848 90260 35888
rect 93964 35848 94004 35888
rect 94924 35848 94964 35888
rect 75052 35680 75092 35720
rect 76780 35680 76820 35720
rect 77644 35680 77684 35720
rect 78796 35680 78836 35720
rect 79180 35680 79220 35720
rect 80332 35680 80372 35720
rect 81580 35680 81620 35720
rect 85228 35680 85268 35720
rect 85612 35680 85652 35720
rect 86668 35680 86708 35720
rect 87916 35680 87956 35720
rect 89932 35680 89972 35720
rect 90316 35680 90356 35720
rect 92428 35680 92468 35720
rect 93868 35680 93908 35720
rect 95020 35680 95060 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 8352 35512 8392 35552
rect 8434 35512 8474 35552
rect 8516 35512 8556 35552
rect 8598 35512 8638 35552
rect 8680 35512 8720 35552
rect 12352 35512 12392 35552
rect 12434 35512 12474 35552
rect 12516 35512 12556 35552
rect 12598 35512 12638 35552
rect 12680 35512 12720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 20352 35512 20392 35552
rect 20434 35512 20474 35552
rect 20516 35512 20556 35552
rect 20598 35512 20638 35552
rect 20680 35512 20720 35552
rect 24352 35512 24392 35552
rect 24434 35512 24474 35552
rect 24516 35512 24556 35552
rect 24598 35512 24638 35552
rect 24680 35512 24720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 32352 35512 32392 35552
rect 32434 35512 32474 35552
rect 32516 35512 32556 35552
rect 32598 35512 32638 35552
rect 32680 35512 32720 35552
rect 36352 35512 36392 35552
rect 36434 35512 36474 35552
rect 36516 35512 36556 35552
rect 36598 35512 36638 35552
rect 36680 35512 36720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 44352 35512 44392 35552
rect 44434 35512 44474 35552
rect 44516 35512 44556 35552
rect 44598 35512 44638 35552
rect 44680 35512 44720 35552
rect 48352 35512 48392 35552
rect 48434 35512 48474 35552
rect 48516 35512 48556 35552
rect 48598 35512 48638 35552
rect 48680 35512 48720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 56352 35512 56392 35552
rect 56434 35512 56474 35552
rect 56516 35512 56556 35552
rect 56598 35512 56638 35552
rect 56680 35512 56720 35552
rect 60352 35512 60392 35552
rect 60434 35512 60474 35552
rect 60516 35512 60556 35552
rect 60598 35512 60638 35552
rect 60680 35512 60720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 68352 35512 68392 35552
rect 68434 35512 68474 35552
rect 68516 35512 68556 35552
rect 68598 35512 68638 35552
rect 68680 35512 68720 35552
rect 72352 35512 72392 35552
rect 72434 35512 72474 35552
rect 72516 35512 72556 35552
rect 72598 35512 72638 35552
rect 72680 35512 72720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 80352 35512 80392 35552
rect 80434 35512 80474 35552
rect 80516 35512 80556 35552
rect 80598 35512 80638 35552
rect 80680 35512 80720 35552
rect 84352 35512 84392 35552
rect 84434 35512 84474 35552
rect 84516 35512 84556 35552
rect 84598 35512 84638 35552
rect 84680 35512 84720 35552
rect 88352 35512 88392 35552
rect 88434 35512 88474 35552
rect 88516 35512 88556 35552
rect 88598 35512 88638 35552
rect 88680 35512 88720 35552
rect 92352 35512 92392 35552
rect 92434 35512 92474 35552
rect 92516 35512 92556 35552
rect 92598 35512 92638 35552
rect 92680 35512 92720 35552
rect 96352 35512 96392 35552
rect 96434 35512 96474 35552
rect 96516 35512 96556 35552
rect 96598 35512 96638 35552
rect 96680 35512 96720 35552
rect 79180 35344 79220 35384
rect 88108 35344 88148 35384
rect 93964 35344 94004 35384
rect 76108 35176 76148 35216
rect 76684 35176 76724 35216
rect 77548 35176 77588 35216
rect 78508 35176 78548 35216
rect 79756 35176 79796 35216
rect 80620 35176 80660 35216
rect 81580 35176 81620 35216
rect 82348 35176 82388 35216
rect 84652 35176 84692 35216
rect 85036 35176 85076 35216
rect 85804 35176 85844 35216
rect 87724 35176 87764 35216
rect 91468 35176 91508 35216
rect 92236 35176 92276 35216
rect 93100 35176 93140 35216
rect 94828 35176 94868 35216
rect 95212 35176 95252 35216
rect 97036 35176 97076 35216
rect 73708 35092 73748 35132
rect 74092 35092 74132 35132
rect 74668 35092 74708 35132
rect 75628 35092 75668 35132
rect 77068 35092 77108 35132
rect 78988 35092 79028 35132
rect 79372 35092 79412 35132
rect 80140 35092 80180 35132
rect 80908 35092 80948 35132
rect 81772 35092 81812 35132
rect 82636 35092 82676 35132
rect 83308 35092 83348 35132
rect 83500 35092 83540 35132
rect 83884 35092 83924 35132
rect 84268 35092 84308 35132
rect 86092 35092 86132 35132
rect 86668 35092 86708 35132
rect 87052 35092 87092 35132
rect 87436 35092 87476 35132
rect 87916 35092 87956 35132
rect 88492 35092 88532 35132
rect 88684 35092 88724 35132
rect 89068 35092 89108 35132
rect 89452 35092 89492 35132
rect 89836 35092 89876 35132
rect 90220 35092 90260 35132
rect 90682 35089 90722 35129
rect 91084 35092 91124 35132
rect 91756 35092 91796 35132
rect 92620 35092 92660 35132
rect 93388 35092 93428 35132
rect 94156 35092 94196 35132
rect 94540 35092 94580 35132
rect 95404 35092 95444 35132
rect 95788 35092 95828 35132
rect 96172 35092 96212 35132
rect 96556 35092 96596 35132
rect 97804 35092 97844 35132
rect 74476 35008 74516 35048
rect 77260 35008 77300 35048
rect 86476 35008 86516 35048
rect 73900 34924 73940 34964
rect 74284 34924 74324 34964
rect 75820 34924 75860 34964
rect 76012 34924 76052 34964
rect 76780 34924 76820 34964
rect 77452 34924 77492 34964
rect 78604 34924 78644 34964
rect 79564 34924 79604 34964
rect 79852 34924 79892 34964
rect 80332 34924 80372 34964
rect 80716 34924 80756 34964
rect 81100 34924 81140 34964
rect 81484 34924 81524 34964
rect 81964 34924 82004 34964
rect 82444 34924 82484 34964
rect 82828 34924 82868 34964
rect 83116 34924 83156 34964
rect 83692 34924 83732 34964
rect 84076 34924 84116 34964
rect 84460 34924 84500 34964
rect 84748 34924 84788 34964
rect 85132 34924 85172 34964
rect 85900 34924 85940 34964
rect 86284 34924 86324 34964
rect 86860 34924 86900 34964
rect 87244 34924 87284 34964
rect 87628 34924 87668 34964
rect 88300 34924 88340 34964
rect 88876 34924 88916 34964
rect 89260 34924 89300 34964
rect 89644 34924 89684 34964
rect 90028 34924 90068 34964
rect 90412 34924 90452 34964
rect 90892 34924 90932 34964
rect 91276 34924 91316 34964
rect 91564 34924 91604 34964
rect 91948 34924 91988 34964
rect 92332 34924 92372 34964
rect 92812 34924 92852 34964
rect 93196 34924 93236 34964
rect 93580 34924 93620 34964
rect 93964 34924 94004 34964
rect 94348 34924 94388 34964
rect 94732 34924 94772 34964
rect 95116 34924 95156 34964
rect 95596 34924 95636 34964
rect 95980 34924 96020 34964
rect 96364 34924 96404 34964
rect 96748 34924 96788 34964
rect 96940 34924 96980 34964
rect 97996 34924 98036 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 7112 34756 7152 34796
rect 7194 34756 7234 34796
rect 7276 34756 7316 34796
rect 7358 34756 7398 34796
rect 7440 34756 7480 34796
rect 11112 34756 11152 34796
rect 11194 34756 11234 34796
rect 11276 34756 11316 34796
rect 11358 34756 11398 34796
rect 11440 34756 11480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 19112 34756 19152 34796
rect 19194 34756 19234 34796
rect 19276 34756 19316 34796
rect 19358 34756 19398 34796
rect 19440 34756 19480 34796
rect 23112 34756 23152 34796
rect 23194 34756 23234 34796
rect 23276 34756 23316 34796
rect 23358 34756 23398 34796
rect 23440 34756 23480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 31112 34756 31152 34796
rect 31194 34756 31234 34796
rect 31276 34756 31316 34796
rect 31358 34756 31398 34796
rect 31440 34756 31480 34796
rect 35112 34756 35152 34796
rect 35194 34756 35234 34796
rect 35276 34756 35316 34796
rect 35358 34756 35398 34796
rect 35440 34756 35480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 43112 34756 43152 34796
rect 43194 34756 43234 34796
rect 43276 34756 43316 34796
rect 43358 34756 43398 34796
rect 43440 34756 43480 34796
rect 47112 34756 47152 34796
rect 47194 34756 47234 34796
rect 47276 34756 47316 34796
rect 47358 34756 47398 34796
rect 47440 34756 47480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 55112 34756 55152 34796
rect 55194 34756 55234 34796
rect 55276 34756 55316 34796
rect 55358 34756 55398 34796
rect 55440 34756 55480 34796
rect 59112 34756 59152 34796
rect 59194 34756 59234 34796
rect 59276 34756 59316 34796
rect 59358 34756 59398 34796
rect 59440 34756 59480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 67112 34756 67152 34796
rect 67194 34756 67234 34796
rect 67276 34756 67316 34796
rect 67358 34756 67398 34796
rect 67440 34756 67480 34796
rect 71112 34756 71152 34796
rect 71194 34756 71234 34796
rect 71276 34756 71316 34796
rect 71358 34756 71398 34796
rect 71440 34756 71480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 79112 34756 79152 34796
rect 79194 34756 79234 34796
rect 79276 34756 79316 34796
rect 79358 34756 79398 34796
rect 79440 34756 79480 34796
rect 83112 34756 83152 34796
rect 83194 34756 83234 34796
rect 83276 34756 83316 34796
rect 83358 34756 83398 34796
rect 83440 34756 83480 34796
rect 87112 34756 87152 34796
rect 87194 34756 87234 34796
rect 87276 34756 87316 34796
rect 87358 34756 87398 34796
rect 87440 34756 87480 34796
rect 91112 34756 91152 34796
rect 91194 34756 91234 34796
rect 91276 34756 91316 34796
rect 91358 34756 91398 34796
rect 91440 34756 91480 34796
rect 95112 34756 95152 34796
rect 95194 34756 95234 34796
rect 95276 34756 95316 34796
rect 95358 34756 95398 34796
rect 95440 34756 95480 34796
rect 99112 34756 99152 34796
rect 99194 34756 99234 34796
rect 99276 34756 99316 34796
rect 99358 34756 99398 34796
rect 99440 34756 99480 34796
rect 83308 34588 83348 34628
rect 86380 34588 86420 34628
rect 92428 34588 92468 34628
rect 95884 34588 95924 34628
rect 80620 34504 80660 34544
rect 81868 34504 81908 34544
rect 85228 34504 85268 34544
rect 89164 34504 89204 34544
rect 91180 34504 91220 34544
rect 96460 34504 96500 34544
rect 96844 34504 96884 34544
rect 73420 34420 73460 34460
rect 73900 34420 73940 34460
rect 74668 34420 74708 34460
rect 75148 34420 75188 34460
rect 76204 34420 76244 34460
rect 76972 34420 77012 34460
rect 77836 34420 77876 34460
rect 78220 34420 78260 34460
rect 79756 34420 79796 34460
rect 80428 34420 80468 34460
rect 81004 34420 81044 34460
rect 81484 34420 81524 34460
rect 82060 34420 82100 34460
rect 82252 34431 82292 34471
rect 83116 34420 83156 34460
rect 84652 34420 84692 34460
rect 85036 34420 85076 34460
rect 85804 34420 85844 34460
rect 86572 34420 86612 34460
rect 87820 34420 87860 34460
rect 88300 34420 88340 34460
rect 89356 34420 89396 34460
rect 90508 34420 90548 34460
rect 90988 34420 91028 34460
rect 92236 34420 92276 34460
rect 93100 34420 93140 34460
rect 93868 34420 93908 34460
rect 94636 34420 94676 34460
rect 95020 34420 95060 34460
rect 96076 34420 96116 34460
rect 96268 34420 96308 34460
rect 97036 34420 97076 34460
rect 97516 34420 97556 34460
rect 98668 34420 98708 34460
rect 74857 34325 74897 34365
rect 75628 34336 75668 34376
rect 75916 34336 75956 34376
rect 76684 34336 76724 34376
rect 77548 34336 77588 34376
rect 78700 34336 78740 34376
rect 78892 34336 78932 34376
rect 79372 34336 79412 34376
rect 80127 34333 80167 34373
rect 81196 34336 81236 34376
rect 82636 34336 82676 34376
rect 83596 34336 83636 34376
rect 83884 34336 83924 34376
rect 84172 34336 84212 34376
rect 84460 34336 84500 34376
rect 85420 34336 85460 34376
rect 86860 34336 86900 34376
rect 87052 34336 87092 34376
rect 87340 34336 87380 34376
rect 88684 34336 88724 34376
rect 89644 34336 89684 34376
rect 89932 34337 89972 34377
rect 90220 34336 90260 34376
rect 91468 34336 91508 34376
rect 91756 34336 91796 34376
rect 92044 34336 92084 34376
rect 92620 34336 92660 34376
rect 92812 34336 92852 34376
rect 93580 34336 93620 34376
rect 94252 34336 94292 34376
rect 95596 34336 95636 34376
rect 96748 34336 96788 34376
rect 97900 34336 97940 34376
rect 98284 34336 98324 34376
rect 98860 34336 98900 34376
rect 99148 34336 99188 34376
rect 80236 34252 80276 34292
rect 73612 34168 73652 34208
rect 74092 34168 74132 34208
rect 74476 34168 74516 34208
rect 74956 34168 74996 34208
rect 75340 34168 75380 34208
rect 75532 34168 75572 34208
rect 76012 34168 76052 34208
rect 76396 34168 76436 34208
rect 76780 34168 76820 34208
rect 77164 34168 77204 34208
rect 77644 34168 77684 34208
rect 78028 34168 78068 34208
rect 78412 34168 78452 34208
rect 78604 34168 78644 34208
rect 78988 34168 79028 34208
rect 79468 34168 79508 34208
rect 79948 34168 79988 34208
rect 80812 34168 80852 34208
rect 81292 34168 81332 34208
rect 81676 34168 81716 34208
rect 82444 34168 82484 34208
rect 82732 34168 82772 34208
rect 83500 34168 83540 34208
rect 83788 34168 83828 34208
rect 84076 34168 84116 34208
rect 84364 34168 84404 34208
rect 84844 34168 84884 34208
rect 85516 34168 85556 34208
rect 85996 34168 86036 34208
rect 86764 34168 86804 34208
rect 87148 34168 87188 34208
rect 87436 34168 87476 34208
rect 88012 34168 88052 34208
rect 88492 34168 88532 34208
rect 88780 34168 88820 34208
rect 89548 34168 89588 34208
rect 89836 34168 89876 34208
rect 90316 34168 90356 34208
rect 90700 34168 90740 34208
rect 91372 34168 91412 34208
rect 91660 34168 91700 34208
rect 91948 34168 91988 34208
rect 93292 34168 93332 34208
rect 93484 34168 93524 34208
rect 94060 34168 94100 34208
rect 94348 34168 94388 34208
rect 94828 34168 94868 34208
rect 95212 34168 95252 34208
rect 95500 34168 95540 34208
rect 97228 34168 97268 34208
rect 97708 34168 97748 34208
rect 97996 34168 98036 34208
rect 98188 34168 98228 34208
rect 98476 34168 98516 34208
rect 98956 34168 98996 34208
rect 99244 34168 99284 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 8352 34000 8392 34040
rect 8434 34000 8474 34040
rect 8516 34000 8556 34040
rect 8598 34000 8638 34040
rect 8680 34000 8720 34040
rect 12352 34000 12392 34040
rect 12434 34000 12474 34040
rect 12516 34000 12556 34040
rect 12598 34000 12638 34040
rect 12680 34000 12720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 20352 34000 20392 34040
rect 20434 34000 20474 34040
rect 20516 34000 20556 34040
rect 20598 34000 20638 34040
rect 20680 34000 20720 34040
rect 24352 34000 24392 34040
rect 24434 34000 24474 34040
rect 24516 34000 24556 34040
rect 24598 34000 24638 34040
rect 24680 34000 24720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 32352 34000 32392 34040
rect 32434 34000 32474 34040
rect 32516 34000 32556 34040
rect 32598 34000 32638 34040
rect 32680 34000 32720 34040
rect 36352 34000 36392 34040
rect 36434 34000 36474 34040
rect 36516 34000 36556 34040
rect 36598 34000 36638 34040
rect 36680 34000 36720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 44352 34000 44392 34040
rect 44434 34000 44474 34040
rect 44516 34000 44556 34040
rect 44598 34000 44638 34040
rect 44680 34000 44720 34040
rect 48352 34000 48392 34040
rect 48434 34000 48474 34040
rect 48516 34000 48556 34040
rect 48598 34000 48638 34040
rect 48680 34000 48720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 56352 34000 56392 34040
rect 56434 34000 56474 34040
rect 56516 34000 56556 34040
rect 56598 34000 56638 34040
rect 56680 34000 56720 34040
rect 60352 34000 60392 34040
rect 60434 34000 60474 34040
rect 60516 34000 60556 34040
rect 60598 34000 60638 34040
rect 60680 34000 60720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 68352 34000 68392 34040
rect 68434 34000 68474 34040
rect 68516 34000 68556 34040
rect 68598 34000 68638 34040
rect 68680 34000 68720 34040
rect 72352 34000 72392 34040
rect 72434 34000 72474 34040
rect 72516 34000 72556 34040
rect 72598 34000 72638 34040
rect 72680 34000 72720 34040
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 80352 34000 80392 34040
rect 80434 34000 80474 34040
rect 80516 34000 80556 34040
rect 80598 34000 80638 34040
rect 80680 34000 80720 34040
rect 84352 34000 84392 34040
rect 84434 34000 84474 34040
rect 84516 34000 84556 34040
rect 84598 34000 84638 34040
rect 84680 34000 84720 34040
rect 88352 34000 88392 34040
rect 88434 34000 88474 34040
rect 88516 34000 88556 34040
rect 88598 34000 88638 34040
rect 88680 34000 88720 34040
rect 92352 34000 92392 34040
rect 92434 34000 92474 34040
rect 92516 34000 92556 34040
rect 92598 34000 92638 34040
rect 92680 34000 92720 34040
rect 96352 34000 96392 34040
rect 96434 34000 96474 34040
rect 96516 34000 96556 34040
rect 96598 34000 96638 34040
rect 96680 34000 96720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 7112 33244 7152 33284
rect 7194 33244 7234 33284
rect 7276 33244 7316 33284
rect 7358 33244 7398 33284
rect 7440 33244 7480 33284
rect 11112 33244 11152 33284
rect 11194 33244 11234 33284
rect 11276 33244 11316 33284
rect 11358 33244 11398 33284
rect 11440 33244 11480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 19112 33244 19152 33284
rect 19194 33244 19234 33284
rect 19276 33244 19316 33284
rect 19358 33244 19398 33284
rect 19440 33244 19480 33284
rect 23112 33244 23152 33284
rect 23194 33244 23234 33284
rect 23276 33244 23316 33284
rect 23358 33244 23398 33284
rect 23440 33244 23480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 31112 33244 31152 33284
rect 31194 33244 31234 33284
rect 31276 33244 31316 33284
rect 31358 33244 31398 33284
rect 31440 33244 31480 33284
rect 35112 33244 35152 33284
rect 35194 33244 35234 33284
rect 35276 33244 35316 33284
rect 35358 33244 35398 33284
rect 35440 33244 35480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 43112 33244 43152 33284
rect 43194 33244 43234 33284
rect 43276 33244 43316 33284
rect 43358 33244 43398 33284
rect 43440 33244 43480 33284
rect 47112 33244 47152 33284
rect 47194 33244 47234 33284
rect 47276 33244 47316 33284
rect 47358 33244 47398 33284
rect 47440 33244 47480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 55112 33244 55152 33284
rect 55194 33244 55234 33284
rect 55276 33244 55316 33284
rect 55358 33244 55398 33284
rect 55440 33244 55480 33284
rect 59112 33244 59152 33284
rect 59194 33244 59234 33284
rect 59276 33244 59316 33284
rect 59358 33244 59398 33284
rect 59440 33244 59480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 67112 33244 67152 33284
rect 67194 33244 67234 33284
rect 67276 33244 67316 33284
rect 67358 33244 67398 33284
rect 67440 33244 67480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 8352 32488 8392 32528
rect 8434 32488 8474 32528
rect 8516 32488 8556 32528
rect 8598 32488 8638 32528
rect 8680 32488 8720 32528
rect 12352 32488 12392 32528
rect 12434 32488 12474 32528
rect 12516 32488 12556 32528
rect 12598 32488 12638 32528
rect 12680 32488 12720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 20352 32488 20392 32528
rect 20434 32488 20474 32528
rect 20516 32488 20556 32528
rect 20598 32488 20638 32528
rect 20680 32488 20720 32528
rect 24352 32488 24392 32528
rect 24434 32488 24474 32528
rect 24516 32488 24556 32528
rect 24598 32488 24638 32528
rect 24680 32488 24720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 32352 32488 32392 32528
rect 32434 32488 32474 32528
rect 32516 32488 32556 32528
rect 32598 32488 32638 32528
rect 32680 32488 32720 32528
rect 36352 32488 36392 32528
rect 36434 32488 36474 32528
rect 36516 32488 36556 32528
rect 36598 32488 36638 32528
rect 36680 32488 36720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 44352 32488 44392 32528
rect 44434 32488 44474 32528
rect 44516 32488 44556 32528
rect 44598 32488 44638 32528
rect 44680 32488 44720 32528
rect 48352 32488 48392 32528
rect 48434 32488 48474 32528
rect 48516 32488 48556 32528
rect 48598 32488 48638 32528
rect 48680 32488 48720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 56352 32488 56392 32528
rect 56434 32488 56474 32528
rect 56516 32488 56556 32528
rect 56598 32488 56638 32528
rect 56680 32488 56720 32528
rect 60352 32488 60392 32528
rect 60434 32488 60474 32528
rect 60516 32488 60556 32528
rect 60598 32488 60638 32528
rect 60680 32488 60720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 68352 32488 68392 32528
rect 68434 32488 68474 32528
rect 68516 32488 68556 32528
rect 68598 32488 68638 32528
rect 68680 32488 68720 32528
rect 69772 32152 69812 32192
rect 69868 31900 69908 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 7112 31732 7152 31772
rect 7194 31732 7234 31772
rect 7276 31732 7316 31772
rect 7358 31732 7398 31772
rect 7440 31732 7480 31772
rect 11112 31732 11152 31772
rect 11194 31732 11234 31772
rect 11276 31732 11316 31772
rect 11358 31732 11398 31772
rect 11440 31732 11480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 19112 31732 19152 31772
rect 19194 31732 19234 31772
rect 19276 31732 19316 31772
rect 19358 31732 19398 31772
rect 19440 31732 19480 31772
rect 23112 31732 23152 31772
rect 23194 31732 23234 31772
rect 23276 31732 23316 31772
rect 23358 31732 23398 31772
rect 23440 31732 23480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 31112 31732 31152 31772
rect 31194 31732 31234 31772
rect 31276 31732 31316 31772
rect 31358 31732 31398 31772
rect 31440 31732 31480 31772
rect 35112 31732 35152 31772
rect 35194 31732 35234 31772
rect 35276 31732 35316 31772
rect 35358 31732 35398 31772
rect 35440 31732 35480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 43112 31732 43152 31772
rect 43194 31732 43234 31772
rect 43276 31732 43316 31772
rect 43358 31732 43398 31772
rect 43440 31732 43480 31772
rect 47112 31732 47152 31772
rect 47194 31732 47234 31772
rect 47276 31732 47316 31772
rect 47358 31732 47398 31772
rect 47440 31732 47480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 55112 31732 55152 31772
rect 55194 31732 55234 31772
rect 55276 31732 55316 31772
rect 55358 31732 55398 31772
rect 55440 31732 55480 31772
rect 59112 31732 59152 31772
rect 59194 31732 59234 31772
rect 59276 31732 59316 31772
rect 59358 31732 59398 31772
rect 59440 31732 59480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 67112 31732 67152 31772
rect 67194 31732 67234 31772
rect 67276 31732 67316 31772
rect 67358 31732 67398 31772
rect 67440 31732 67480 31772
rect 68812 31564 68852 31604
rect 69868 31564 69908 31604
rect 67180 31480 67220 31520
rect 69196 31480 69236 31520
rect 69580 31480 69620 31520
rect 68620 31396 68660 31436
rect 69004 31396 69044 31436
rect 69388 31396 69428 31436
rect 67276 31312 67316 31352
rect 67564 31312 67604 31352
rect 67756 31312 67796 31352
rect 69772 31312 69812 31352
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 8352 30976 8392 31016
rect 8434 30976 8474 31016
rect 8516 30976 8556 31016
rect 8598 30976 8638 31016
rect 8680 30976 8720 31016
rect 12352 30976 12392 31016
rect 12434 30976 12474 31016
rect 12516 30976 12556 31016
rect 12598 30976 12638 31016
rect 12680 30976 12720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 20352 30976 20392 31016
rect 20434 30976 20474 31016
rect 20516 30976 20556 31016
rect 20598 30976 20638 31016
rect 20680 30976 20720 31016
rect 24352 30976 24392 31016
rect 24434 30976 24474 31016
rect 24516 30976 24556 31016
rect 24598 30976 24638 31016
rect 24680 30976 24720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 32352 30976 32392 31016
rect 32434 30976 32474 31016
rect 32516 30976 32556 31016
rect 32598 30976 32638 31016
rect 32680 30976 32720 31016
rect 36352 30976 36392 31016
rect 36434 30976 36474 31016
rect 36516 30976 36556 31016
rect 36598 30976 36638 31016
rect 36680 30976 36720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 44352 30976 44392 31016
rect 44434 30976 44474 31016
rect 44516 30976 44556 31016
rect 44598 30976 44638 31016
rect 44680 30976 44720 31016
rect 48352 30976 48392 31016
rect 48434 30976 48474 31016
rect 48516 30976 48556 31016
rect 48598 30976 48638 31016
rect 48680 30976 48720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 56352 30976 56392 31016
rect 56434 30976 56474 31016
rect 56516 30976 56556 31016
rect 56598 30976 56638 31016
rect 56680 30976 56720 31016
rect 60352 30976 60392 31016
rect 60434 30976 60474 31016
rect 60516 30976 60556 31016
rect 60598 30976 60638 31016
rect 60680 30976 60720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 68352 30976 68392 31016
rect 68434 30976 68474 31016
rect 68516 30976 68556 31016
rect 68598 30976 68638 31016
rect 68680 30976 68720 31016
rect 67564 30808 67604 30848
rect 68620 30808 68660 30848
rect 69100 30808 69140 30848
rect 69388 30808 69428 30848
rect 69676 30808 69716 30848
rect 68524 30640 68564 30680
rect 69004 30640 69044 30680
rect 69292 30640 69332 30680
rect 69580 30640 69620 30680
rect 67372 30556 67412 30596
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 7112 30220 7152 30260
rect 7194 30220 7234 30260
rect 7276 30220 7316 30260
rect 7358 30220 7398 30260
rect 7440 30220 7480 30260
rect 11112 30220 11152 30260
rect 11194 30220 11234 30260
rect 11276 30220 11316 30260
rect 11358 30220 11398 30260
rect 11440 30220 11480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 19112 30220 19152 30260
rect 19194 30220 19234 30260
rect 19276 30220 19316 30260
rect 19358 30220 19398 30260
rect 19440 30220 19480 30260
rect 23112 30220 23152 30260
rect 23194 30220 23234 30260
rect 23276 30220 23316 30260
rect 23358 30220 23398 30260
rect 23440 30220 23480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 31112 30220 31152 30260
rect 31194 30220 31234 30260
rect 31276 30220 31316 30260
rect 31358 30220 31398 30260
rect 31440 30220 31480 30260
rect 35112 30220 35152 30260
rect 35194 30220 35234 30260
rect 35276 30220 35316 30260
rect 35358 30220 35398 30260
rect 35440 30220 35480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 43112 30220 43152 30260
rect 43194 30220 43234 30260
rect 43276 30220 43316 30260
rect 43358 30220 43398 30260
rect 43440 30220 43480 30260
rect 47112 30220 47152 30260
rect 47194 30220 47234 30260
rect 47276 30220 47316 30260
rect 47358 30220 47398 30260
rect 47440 30220 47480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 55112 30220 55152 30260
rect 55194 30220 55234 30260
rect 55276 30220 55316 30260
rect 55358 30220 55398 30260
rect 55440 30220 55480 30260
rect 59112 30220 59152 30260
rect 59194 30220 59234 30260
rect 59276 30220 59316 30260
rect 59358 30220 59398 30260
rect 59440 30220 59480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 67112 30220 67152 30260
rect 67194 30220 67234 30260
rect 67276 30220 67316 30260
rect 67358 30220 67398 30260
rect 67440 30220 67480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 8352 29464 8392 29504
rect 8434 29464 8474 29504
rect 8516 29464 8556 29504
rect 8598 29464 8638 29504
rect 8680 29464 8720 29504
rect 12352 29464 12392 29504
rect 12434 29464 12474 29504
rect 12516 29464 12556 29504
rect 12598 29464 12638 29504
rect 12680 29464 12720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 20352 29464 20392 29504
rect 20434 29464 20474 29504
rect 20516 29464 20556 29504
rect 20598 29464 20638 29504
rect 20680 29464 20720 29504
rect 24352 29464 24392 29504
rect 24434 29464 24474 29504
rect 24516 29464 24556 29504
rect 24598 29464 24638 29504
rect 24680 29464 24720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 32352 29464 32392 29504
rect 32434 29464 32474 29504
rect 32516 29464 32556 29504
rect 32598 29464 32638 29504
rect 32680 29464 32720 29504
rect 36352 29464 36392 29504
rect 36434 29464 36474 29504
rect 36516 29464 36556 29504
rect 36598 29464 36638 29504
rect 36680 29464 36720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 44352 29464 44392 29504
rect 44434 29464 44474 29504
rect 44516 29464 44556 29504
rect 44598 29464 44638 29504
rect 44680 29464 44720 29504
rect 48352 29464 48392 29504
rect 48434 29464 48474 29504
rect 48516 29464 48556 29504
rect 48598 29464 48638 29504
rect 48680 29464 48720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 56352 29464 56392 29504
rect 56434 29464 56474 29504
rect 56516 29464 56556 29504
rect 56598 29464 56638 29504
rect 56680 29464 56720 29504
rect 60352 29464 60392 29504
rect 60434 29464 60474 29504
rect 60516 29464 60556 29504
rect 60598 29464 60638 29504
rect 60680 29464 60720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 68352 29464 68392 29504
rect 68434 29464 68474 29504
rect 68516 29464 68556 29504
rect 68598 29464 68638 29504
rect 68680 29464 68720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 7112 28708 7152 28748
rect 7194 28708 7234 28748
rect 7276 28708 7316 28748
rect 7358 28708 7398 28748
rect 7440 28708 7480 28748
rect 11112 28708 11152 28748
rect 11194 28708 11234 28748
rect 11276 28708 11316 28748
rect 11358 28708 11398 28748
rect 11440 28708 11480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 19112 28708 19152 28748
rect 19194 28708 19234 28748
rect 19276 28708 19316 28748
rect 19358 28708 19398 28748
rect 19440 28708 19480 28748
rect 23112 28708 23152 28748
rect 23194 28708 23234 28748
rect 23276 28708 23316 28748
rect 23358 28708 23398 28748
rect 23440 28708 23480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 31112 28708 31152 28748
rect 31194 28708 31234 28748
rect 31276 28708 31316 28748
rect 31358 28708 31398 28748
rect 31440 28708 31480 28748
rect 35112 28708 35152 28748
rect 35194 28708 35234 28748
rect 35276 28708 35316 28748
rect 35358 28708 35398 28748
rect 35440 28708 35480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 43112 28708 43152 28748
rect 43194 28708 43234 28748
rect 43276 28708 43316 28748
rect 43358 28708 43398 28748
rect 43440 28708 43480 28748
rect 47112 28708 47152 28748
rect 47194 28708 47234 28748
rect 47276 28708 47316 28748
rect 47358 28708 47398 28748
rect 47440 28708 47480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 55112 28708 55152 28748
rect 55194 28708 55234 28748
rect 55276 28708 55316 28748
rect 55358 28708 55398 28748
rect 55440 28708 55480 28748
rect 59112 28708 59152 28748
rect 59194 28708 59234 28748
rect 59276 28708 59316 28748
rect 59358 28708 59398 28748
rect 59440 28708 59480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 67112 28708 67152 28748
rect 67194 28708 67234 28748
rect 67276 28708 67316 28748
rect 67358 28708 67398 28748
rect 67440 28708 67480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 8352 27952 8392 27992
rect 8434 27952 8474 27992
rect 8516 27952 8556 27992
rect 8598 27952 8638 27992
rect 8680 27952 8720 27992
rect 12352 27952 12392 27992
rect 12434 27952 12474 27992
rect 12516 27952 12556 27992
rect 12598 27952 12638 27992
rect 12680 27952 12720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 20352 27952 20392 27992
rect 20434 27952 20474 27992
rect 20516 27952 20556 27992
rect 20598 27952 20638 27992
rect 20680 27952 20720 27992
rect 24352 27952 24392 27992
rect 24434 27952 24474 27992
rect 24516 27952 24556 27992
rect 24598 27952 24638 27992
rect 24680 27952 24720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 32352 27952 32392 27992
rect 32434 27952 32474 27992
rect 32516 27952 32556 27992
rect 32598 27952 32638 27992
rect 32680 27952 32720 27992
rect 36352 27952 36392 27992
rect 36434 27952 36474 27992
rect 36516 27952 36556 27992
rect 36598 27952 36638 27992
rect 36680 27952 36720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 44352 27952 44392 27992
rect 44434 27952 44474 27992
rect 44516 27952 44556 27992
rect 44598 27952 44638 27992
rect 44680 27952 44720 27992
rect 48352 27952 48392 27992
rect 48434 27952 48474 27992
rect 48516 27952 48556 27992
rect 48598 27952 48638 27992
rect 48680 27952 48720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 56352 27952 56392 27992
rect 56434 27952 56474 27992
rect 56516 27952 56556 27992
rect 56598 27952 56638 27992
rect 56680 27952 56720 27992
rect 60352 27952 60392 27992
rect 60434 27952 60474 27992
rect 60516 27952 60556 27992
rect 60598 27952 60638 27992
rect 60680 27952 60720 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 68352 27952 68392 27992
rect 68434 27952 68474 27992
rect 68516 27952 68556 27992
rect 68598 27952 68638 27992
rect 68680 27952 68720 27992
rect 68812 27532 68852 27572
rect 69004 27364 69044 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 7112 27196 7152 27236
rect 7194 27196 7234 27236
rect 7276 27196 7316 27236
rect 7358 27196 7398 27236
rect 7440 27196 7480 27236
rect 11112 27196 11152 27236
rect 11194 27196 11234 27236
rect 11276 27196 11316 27236
rect 11358 27196 11398 27236
rect 11440 27196 11480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 19112 27196 19152 27236
rect 19194 27196 19234 27236
rect 19276 27196 19316 27236
rect 19358 27196 19398 27236
rect 19440 27196 19480 27236
rect 23112 27196 23152 27236
rect 23194 27196 23234 27236
rect 23276 27196 23316 27236
rect 23358 27196 23398 27236
rect 23440 27196 23480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 31112 27196 31152 27236
rect 31194 27196 31234 27236
rect 31276 27196 31316 27236
rect 31358 27196 31398 27236
rect 31440 27196 31480 27236
rect 35112 27196 35152 27236
rect 35194 27196 35234 27236
rect 35276 27196 35316 27236
rect 35358 27196 35398 27236
rect 35440 27196 35480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 43112 27196 43152 27236
rect 43194 27196 43234 27236
rect 43276 27196 43316 27236
rect 43358 27196 43398 27236
rect 43440 27196 43480 27236
rect 47112 27196 47152 27236
rect 47194 27196 47234 27236
rect 47276 27196 47316 27236
rect 47358 27196 47398 27236
rect 47440 27196 47480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 55112 27196 55152 27236
rect 55194 27196 55234 27236
rect 55276 27196 55316 27236
rect 55358 27196 55398 27236
rect 55440 27196 55480 27236
rect 59112 27196 59152 27236
rect 59194 27196 59234 27236
rect 59276 27196 59316 27236
rect 59358 27196 59398 27236
rect 59440 27196 59480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 67112 27196 67152 27236
rect 67194 27196 67234 27236
rect 67276 27196 67316 27236
rect 67358 27196 67398 27236
rect 67440 27196 67480 27236
rect 68140 26944 68180 26984
rect 67948 26860 67988 26900
rect 68332 26860 68372 26900
rect 69484 26860 69524 26900
rect 67756 26608 67796 26648
rect 69676 26608 69716 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 8352 26440 8392 26480
rect 8434 26440 8474 26480
rect 8516 26440 8556 26480
rect 8598 26440 8638 26480
rect 8680 26440 8720 26480
rect 12352 26440 12392 26480
rect 12434 26440 12474 26480
rect 12516 26440 12556 26480
rect 12598 26440 12638 26480
rect 12680 26440 12720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 20352 26440 20392 26480
rect 20434 26440 20474 26480
rect 20516 26440 20556 26480
rect 20598 26440 20638 26480
rect 20680 26440 20720 26480
rect 24352 26440 24392 26480
rect 24434 26440 24474 26480
rect 24516 26440 24556 26480
rect 24598 26440 24638 26480
rect 24680 26440 24720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 32352 26440 32392 26480
rect 32434 26440 32474 26480
rect 32516 26440 32556 26480
rect 32598 26440 32638 26480
rect 32680 26440 32720 26480
rect 36352 26440 36392 26480
rect 36434 26440 36474 26480
rect 36516 26440 36556 26480
rect 36598 26440 36638 26480
rect 36680 26440 36720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 44352 26440 44392 26480
rect 44434 26440 44474 26480
rect 44516 26440 44556 26480
rect 44598 26440 44638 26480
rect 44680 26440 44720 26480
rect 48352 26440 48392 26480
rect 48434 26440 48474 26480
rect 48516 26440 48556 26480
rect 48598 26440 48638 26480
rect 48680 26440 48720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 56352 26440 56392 26480
rect 56434 26440 56474 26480
rect 56516 26440 56556 26480
rect 56598 26440 56638 26480
rect 56680 26440 56720 26480
rect 60352 26440 60392 26480
rect 60434 26440 60474 26480
rect 60516 26440 60556 26480
rect 60598 26440 60638 26480
rect 60680 26440 60720 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 68352 26440 68392 26480
rect 68434 26440 68474 26480
rect 68516 26440 68556 26480
rect 68598 26440 68638 26480
rect 68680 26440 68720 26480
rect 67564 26104 67604 26144
rect 68620 26104 68660 26144
rect 68812 26104 68852 26144
rect 69100 26104 69140 26144
rect 69772 26104 69812 26144
rect 67756 26020 67796 26060
rect 69388 26020 69428 26060
rect 67468 25852 67508 25892
rect 67948 25852 67988 25892
rect 68524 25852 68564 25892
rect 68908 25852 68948 25892
rect 69196 25852 69236 25892
rect 69580 25852 69620 25892
rect 69868 25852 69908 25892
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 7112 25684 7152 25724
rect 7194 25684 7234 25724
rect 7276 25684 7316 25724
rect 7358 25684 7398 25724
rect 7440 25684 7480 25724
rect 11112 25684 11152 25724
rect 11194 25684 11234 25724
rect 11276 25684 11316 25724
rect 11358 25684 11398 25724
rect 11440 25684 11480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 19112 25684 19152 25724
rect 19194 25684 19234 25724
rect 19276 25684 19316 25724
rect 19358 25684 19398 25724
rect 19440 25684 19480 25724
rect 23112 25684 23152 25724
rect 23194 25684 23234 25724
rect 23276 25684 23316 25724
rect 23358 25684 23398 25724
rect 23440 25684 23480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 31112 25684 31152 25724
rect 31194 25684 31234 25724
rect 31276 25684 31316 25724
rect 31358 25684 31398 25724
rect 31440 25684 31480 25724
rect 35112 25684 35152 25724
rect 35194 25684 35234 25724
rect 35276 25684 35316 25724
rect 35358 25684 35398 25724
rect 35440 25684 35480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 43112 25684 43152 25724
rect 43194 25684 43234 25724
rect 43276 25684 43316 25724
rect 43358 25684 43398 25724
rect 43440 25684 43480 25724
rect 47112 25684 47152 25724
rect 47194 25684 47234 25724
rect 47276 25684 47316 25724
rect 47358 25684 47398 25724
rect 47440 25684 47480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 55112 25684 55152 25724
rect 55194 25684 55234 25724
rect 55276 25684 55316 25724
rect 55358 25684 55398 25724
rect 55440 25684 55480 25724
rect 59112 25684 59152 25724
rect 59194 25684 59234 25724
rect 59276 25684 59316 25724
rect 59358 25684 59398 25724
rect 59440 25684 59480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 67112 25684 67152 25724
rect 67194 25684 67234 25724
rect 67276 25684 67316 25724
rect 67358 25684 67398 25724
rect 67440 25684 67480 25724
rect 68812 25516 68852 25556
rect 69868 25516 69908 25556
rect 68620 25348 68660 25388
rect 69676 25348 69716 25388
rect 652 25264 692 25304
rect 844 25264 884 25304
rect 69292 25264 69332 25304
rect 69484 25264 69524 25304
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 8352 24928 8392 24968
rect 8434 24928 8474 24968
rect 8516 24928 8556 24968
rect 8598 24928 8638 24968
rect 8680 24928 8720 24968
rect 12352 24928 12392 24968
rect 12434 24928 12474 24968
rect 12516 24928 12556 24968
rect 12598 24928 12638 24968
rect 12680 24928 12720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 20352 24928 20392 24968
rect 20434 24928 20474 24968
rect 20516 24928 20556 24968
rect 20598 24928 20638 24968
rect 20680 24928 20720 24968
rect 24352 24928 24392 24968
rect 24434 24928 24474 24968
rect 24516 24928 24556 24968
rect 24598 24928 24638 24968
rect 24680 24928 24720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 32352 24928 32392 24968
rect 32434 24928 32474 24968
rect 32516 24928 32556 24968
rect 32598 24928 32638 24968
rect 32680 24928 32720 24968
rect 36352 24928 36392 24968
rect 36434 24928 36474 24968
rect 36516 24928 36556 24968
rect 36598 24928 36638 24968
rect 36680 24928 36720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 44352 24928 44392 24968
rect 44434 24928 44474 24968
rect 44516 24928 44556 24968
rect 44598 24928 44638 24968
rect 44680 24928 44720 24968
rect 48352 24928 48392 24968
rect 48434 24928 48474 24968
rect 48516 24928 48556 24968
rect 48598 24928 48638 24968
rect 48680 24928 48720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 56352 24928 56392 24968
rect 56434 24928 56474 24968
rect 56516 24928 56556 24968
rect 56598 24928 56638 24968
rect 56680 24928 56720 24968
rect 60352 24928 60392 24968
rect 60434 24928 60474 24968
rect 60516 24928 60556 24968
rect 60598 24928 60638 24968
rect 60680 24928 60720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 68352 24928 68392 24968
rect 68434 24928 68474 24968
rect 68516 24928 68556 24968
rect 68598 24928 68638 24968
rect 68680 24928 68720 24968
rect 652 24592 692 24632
rect 844 24592 884 24632
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 7112 24172 7152 24212
rect 7194 24172 7234 24212
rect 7276 24172 7316 24212
rect 7358 24172 7398 24212
rect 7440 24172 7480 24212
rect 11112 24172 11152 24212
rect 11194 24172 11234 24212
rect 11276 24172 11316 24212
rect 11358 24172 11398 24212
rect 11440 24172 11480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 19112 24172 19152 24212
rect 19194 24172 19234 24212
rect 19276 24172 19316 24212
rect 19358 24172 19398 24212
rect 19440 24172 19480 24212
rect 23112 24172 23152 24212
rect 23194 24172 23234 24212
rect 23276 24172 23316 24212
rect 23358 24172 23398 24212
rect 23440 24172 23480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 31112 24172 31152 24212
rect 31194 24172 31234 24212
rect 31276 24172 31316 24212
rect 31358 24172 31398 24212
rect 31440 24172 31480 24212
rect 35112 24172 35152 24212
rect 35194 24172 35234 24212
rect 35276 24172 35316 24212
rect 35358 24172 35398 24212
rect 35440 24172 35480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 43112 24172 43152 24212
rect 43194 24172 43234 24212
rect 43276 24172 43316 24212
rect 43358 24172 43398 24212
rect 43440 24172 43480 24212
rect 47112 24172 47152 24212
rect 47194 24172 47234 24212
rect 47276 24172 47316 24212
rect 47358 24172 47398 24212
rect 47440 24172 47480 24212
rect 51112 24172 51152 24212
rect 51194 24172 51234 24212
rect 51276 24172 51316 24212
rect 51358 24172 51398 24212
rect 51440 24172 51480 24212
rect 55112 24172 55152 24212
rect 55194 24172 55234 24212
rect 55276 24172 55316 24212
rect 55358 24172 55398 24212
rect 55440 24172 55480 24212
rect 59112 24172 59152 24212
rect 59194 24172 59234 24212
rect 59276 24172 59316 24212
rect 59358 24172 59398 24212
rect 59440 24172 59480 24212
rect 63112 24172 63152 24212
rect 63194 24172 63234 24212
rect 63276 24172 63316 24212
rect 63358 24172 63398 24212
rect 63440 24172 63480 24212
rect 67112 24172 67152 24212
rect 67194 24172 67234 24212
rect 67276 24172 67316 24212
rect 67358 24172 67398 24212
rect 67440 24172 67480 24212
rect 652 23752 692 23792
rect 844 23752 884 23792
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 8352 23416 8392 23456
rect 8434 23416 8474 23456
rect 8516 23416 8556 23456
rect 8598 23416 8638 23456
rect 8680 23416 8720 23456
rect 12352 23416 12392 23456
rect 12434 23416 12474 23456
rect 12516 23416 12556 23456
rect 12598 23416 12638 23456
rect 12680 23416 12720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 20352 23416 20392 23456
rect 20434 23416 20474 23456
rect 20516 23416 20556 23456
rect 20598 23416 20638 23456
rect 20680 23416 20720 23456
rect 24352 23416 24392 23456
rect 24434 23416 24474 23456
rect 24516 23416 24556 23456
rect 24598 23416 24638 23456
rect 24680 23416 24720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 32352 23416 32392 23456
rect 32434 23416 32474 23456
rect 32516 23416 32556 23456
rect 32598 23416 32638 23456
rect 32680 23416 32720 23456
rect 36352 23416 36392 23456
rect 36434 23416 36474 23456
rect 36516 23416 36556 23456
rect 36598 23416 36638 23456
rect 36680 23416 36720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 44352 23416 44392 23456
rect 44434 23416 44474 23456
rect 44516 23416 44556 23456
rect 44598 23416 44638 23456
rect 44680 23416 44720 23456
rect 48352 23416 48392 23456
rect 48434 23416 48474 23456
rect 48516 23416 48556 23456
rect 48598 23416 48638 23456
rect 48680 23416 48720 23456
rect 52352 23416 52392 23456
rect 52434 23416 52474 23456
rect 52516 23416 52556 23456
rect 52598 23416 52638 23456
rect 52680 23416 52720 23456
rect 56352 23416 56392 23456
rect 56434 23416 56474 23456
rect 56516 23416 56556 23456
rect 56598 23416 56638 23456
rect 56680 23416 56720 23456
rect 60352 23416 60392 23456
rect 60434 23416 60474 23456
rect 60516 23416 60556 23456
rect 60598 23416 60638 23456
rect 60680 23416 60720 23456
rect 64352 23416 64392 23456
rect 64434 23416 64474 23456
rect 64516 23416 64556 23456
rect 64598 23416 64638 23456
rect 64680 23416 64720 23456
rect 68352 23416 68392 23456
rect 68434 23416 68474 23456
rect 68516 23416 68556 23456
rect 68598 23416 68638 23456
rect 68680 23416 68720 23456
rect 72352 23416 72392 23456
rect 72434 23416 72474 23456
rect 72516 23416 72556 23456
rect 72598 23416 72638 23456
rect 72680 23416 72720 23456
rect 76352 23416 76392 23456
rect 76434 23416 76474 23456
rect 76516 23416 76556 23456
rect 76598 23416 76638 23456
rect 76680 23416 76720 23456
rect 80352 23416 80392 23456
rect 80434 23416 80474 23456
rect 80516 23416 80556 23456
rect 80598 23416 80638 23456
rect 80680 23416 80720 23456
rect 84352 23416 84392 23456
rect 84434 23416 84474 23456
rect 84516 23416 84556 23456
rect 84598 23416 84638 23456
rect 84680 23416 84720 23456
rect 88352 23416 88392 23456
rect 88434 23416 88474 23456
rect 88516 23416 88556 23456
rect 88598 23416 88638 23456
rect 88680 23416 88720 23456
rect 92352 23416 92392 23456
rect 92434 23416 92474 23456
rect 92516 23416 92556 23456
rect 92598 23416 92638 23456
rect 92680 23416 92720 23456
rect 96352 23416 96392 23456
rect 96434 23416 96474 23456
rect 96516 23416 96556 23456
rect 96598 23416 96638 23456
rect 96680 23416 96720 23456
rect 73132 23248 73172 23288
rect 73420 23248 73460 23288
rect 74092 23248 74132 23288
rect 74956 23248 74996 23288
rect 75532 23248 75572 23288
rect 75916 23248 75956 23288
rect 77068 23248 77108 23288
rect 77452 23248 77492 23288
rect 78028 23248 78068 23288
rect 78604 23248 78644 23288
rect 79180 23248 79220 23288
rect 79468 23248 79508 23288
rect 79852 23248 79892 23288
rect 80908 23248 80948 23288
rect 81196 23248 81236 23288
rect 81484 23248 81524 23288
rect 81772 23248 81812 23288
rect 82060 23248 82100 23288
rect 82636 23248 82676 23288
rect 82924 23248 82964 23288
rect 84460 23248 84500 23288
rect 84844 23248 84884 23288
rect 85228 23248 85268 23288
rect 85516 23248 85556 23288
rect 86284 23248 86324 23288
rect 87148 23248 87188 23288
rect 87724 23248 87764 23288
rect 88012 23248 88052 23288
rect 88396 23248 88436 23288
rect 88876 23248 88916 23288
rect 89356 23248 89396 23288
rect 90508 23248 90548 23288
rect 90796 23248 90836 23288
rect 91084 23248 91124 23288
rect 91468 23248 91508 23288
rect 93100 23248 93140 23288
rect 93484 23248 93524 23288
rect 93964 23248 94004 23288
rect 94636 23248 94676 23288
rect 94828 23248 94868 23288
rect 95404 23248 95444 23288
rect 96460 23248 96500 23288
rect 96748 23248 96788 23288
rect 97036 23248 97076 23288
rect 97324 23248 97364 23288
rect 97708 23248 97748 23288
rect 98092 23248 98132 23288
rect 98476 23248 98516 23288
rect 98860 23248 98900 23288
rect 652 23080 692 23120
rect 844 23080 884 23120
rect 73036 23080 73076 23120
rect 73324 23080 73364 23120
rect 74188 23080 74228 23120
rect 78124 23080 78164 23120
rect 79276 23080 79316 23120
rect 79564 23080 79604 23120
rect 79756 23080 79796 23120
rect 80044 23080 80084 23120
rect 80236 23080 80276 23120
rect 81004 23080 81044 23120
rect 81292 23080 81332 23120
rect 81580 23080 81620 23120
rect 81868 23080 81908 23120
rect 82156 23080 82196 23120
rect 82828 23080 82868 23120
rect 83212 23080 83252 23120
rect 83404 23080 83444 23120
rect 84076 23080 84116 23120
rect 84364 23080 84404 23120
rect 84748 23080 84788 23120
rect 85132 23080 85172 23120
rect 85420 23080 85460 23120
rect 86476 23080 86516 23120
rect 86668 23080 86708 23120
rect 87820 23080 87860 23120
rect 88108 23080 88148 23120
rect 88492 23080 88532 23120
rect 88780 23080 88820 23120
rect 89452 23080 89492 23120
rect 89644 23080 89684 23120
rect 89836 23080 89876 23120
rect 90604 23080 90644 23120
rect 90892 23080 90932 23120
rect 91180 23080 91220 23120
rect 91372 23080 91412 23120
rect 93676 23080 93716 23120
rect 93772 23080 93812 23120
rect 94060 23080 94100 23120
rect 94924 23080 94964 23120
rect 95308 23080 95348 23120
rect 95692 23080 95732 23120
rect 95884 23080 95924 23120
rect 96556 23080 96596 23120
rect 96844 23080 96884 23120
rect 97132 23080 97172 23120
rect 97420 23080 97460 23120
rect 97804 23080 97844 23120
rect 98188 23080 98228 23120
rect 98956 23080 98996 23120
rect 74380 22996 74420 23036
rect 74764 22996 74804 23036
rect 75340 22996 75380 23036
rect 75724 22996 75764 23036
rect 76108 22996 76148 23036
rect 76300 22996 76340 23036
rect 76876 22996 76916 23036
rect 77260 22996 77300 23036
rect 77836 22996 77876 23036
rect 78412 22996 78452 23036
rect 78796 22996 78836 23036
rect 80716 22996 80756 23036
rect 82444 22996 82484 23036
rect 83788 22996 83828 23036
rect 85708 22996 85748 23036
rect 86092 22996 86132 23036
rect 86956 22996 86996 23036
rect 87532 22996 87572 23036
rect 90316 22996 90356 23036
rect 91660 22996 91700 23036
rect 92044 22996 92084 23036
rect 92428 22996 92468 23036
rect 92908 22996 92948 23036
rect 93292 22996 93332 23036
rect 94444 22996 94484 23036
rect 96076 22996 96116 23036
rect 98668 22996 98708 23036
rect 75148 22912 75188 22952
rect 76492 22912 76532 22952
rect 78988 22912 79028 22952
rect 83596 22912 83636 22952
rect 91852 22912 91892 22952
rect 74572 22828 74612 22868
rect 77644 22828 77684 22868
rect 80524 22828 80564 22868
rect 83980 22828 84020 22868
rect 85900 22828 85940 22868
rect 87340 22828 87380 22868
rect 90124 22828 90164 22868
rect 92236 22828 92276 22868
rect 92620 22828 92660 22868
rect 96268 22828 96308 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 7112 22660 7152 22700
rect 7194 22660 7234 22700
rect 7276 22660 7316 22700
rect 7358 22660 7398 22700
rect 7440 22660 7480 22700
rect 11112 22660 11152 22700
rect 11194 22660 11234 22700
rect 11276 22660 11316 22700
rect 11358 22660 11398 22700
rect 11440 22660 11480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 19112 22660 19152 22700
rect 19194 22660 19234 22700
rect 19276 22660 19316 22700
rect 19358 22660 19398 22700
rect 19440 22660 19480 22700
rect 23112 22660 23152 22700
rect 23194 22660 23234 22700
rect 23276 22660 23316 22700
rect 23358 22660 23398 22700
rect 23440 22660 23480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 31112 22660 31152 22700
rect 31194 22660 31234 22700
rect 31276 22660 31316 22700
rect 31358 22660 31398 22700
rect 31440 22660 31480 22700
rect 35112 22660 35152 22700
rect 35194 22660 35234 22700
rect 35276 22660 35316 22700
rect 35358 22660 35398 22700
rect 35440 22660 35480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 43112 22660 43152 22700
rect 43194 22660 43234 22700
rect 43276 22660 43316 22700
rect 43358 22660 43398 22700
rect 43440 22660 43480 22700
rect 47112 22660 47152 22700
rect 47194 22660 47234 22700
rect 47276 22660 47316 22700
rect 47358 22660 47398 22700
rect 47440 22660 47480 22700
rect 51112 22660 51152 22700
rect 51194 22660 51234 22700
rect 51276 22660 51316 22700
rect 51358 22660 51398 22700
rect 51440 22660 51480 22700
rect 55112 22660 55152 22700
rect 55194 22660 55234 22700
rect 55276 22660 55316 22700
rect 55358 22660 55398 22700
rect 55440 22660 55480 22700
rect 59112 22660 59152 22700
rect 59194 22660 59234 22700
rect 59276 22660 59316 22700
rect 59358 22660 59398 22700
rect 59440 22660 59480 22700
rect 63112 22660 63152 22700
rect 63194 22660 63234 22700
rect 63276 22660 63316 22700
rect 63358 22660 63398 22700
rect 63440 22660 63480 22700
rect 67112 22660 67152 22700
rect 67194 22660 67234 22700
rect 67276 22660 67316 22700
rect 67358 22660 67398 22700
rect 67440 22660 67480 22700
rect 71112 22660 71152 22700
rect 71194 22660 71234 22700
rect 71276 22660 71316 22700
rect 71358 22660 71398 22700
rect 71440 22660 71480 22700
rect 75112 22660 75152 22700
rect 75194 22660 75234 22700
rect 75276 22660 75316 22700
rect 75358 22660 75398 22700
rect 75440 22660 75480 22700
rect 79112 22660 79152 22700
rect 79194 22660 79234 22700
rect 79276 22660 79316 22700
rect 79358 22660 79398 22700
rect 79440 22660 79480 22700
rect 83112 22660 83152 22700
rect 83194 22660 83234 22700
rect 83276 22660 83316 22700
rect 83358 22660 83398 22700
rect 83440 22660 83480 22700
rect 87112 22660 87152 22700
rect 87194 22660 87234 22700
rect 87276 22660 87316 22700
rect 87358 22660 87398 22700
rect 87440 22660 87480 22700
rect 91112 22660 91152 22700
rect 91194 22660 91234 22700
rect 91276 22660 91316 22700
rect 91358 22660 91398 22700
rect 91440 22660 91480 22700
rect 95112 22660 95152 22700
rect 95194 22660 95234 22700
rect 95276 22660 95316 22700
rect 95358 22660 95398 22700
rect 95440 22660 95480 22700
rect 99112 22660 99152 22700
rect 99194 22660 99234 22700
rect 99276 22660 99316 22700
rect 99358 22660 99398 22700
rect 99440 22660 99480 22700
rect 73900 22492 73940 22532
rect 74572 22492 74612 22532
rect 75436 22492 75476 22532
rect 75916 22492 75956 22532
rect 76300 22492 76340 22532
rect 76684 22492 76724 22532
rect 77260 22492 77300 22532
rect 77932 22492 77972 22532
rect 78316 22492 78356 22532
rect 79756 22492 79796 22532
rect 80140 22492 80180 22532
rect 80620 22492 80660 22532
rect 80812 22492 80852 22532
rect 81484 22492 81524 22532
rect 81868 22492 81908 22532
rect 83020 22492 83060 22532
rect 83596 22492 83636 22532
rect 83980 22492 84020 22532
rect 84748 22492 84788 22532
rect 85132 22492 85172 22532
rect 85420 22492 85460 22532
rect 85996 22492 86036 22532
rect 86764 22492 86804 22532
rect 87052 22492 87092 22532
rect 87436 22492 87476 22532
rect 87820 22492 87860 22532
rect 88204 22492 88244 22532
rect 88588 22492 88628 22532
rect 89068 22492 89108 22532
rect 89932 22492 89972 22532
rect 90220 22492 90260 22532
rect 90796 22492 90836 22532
rect 91468 22492 91508 22532
rect 91660 22492 91700 22532
rect 92044 22492 92084 22532
rect 92428 22492 92468 22532
rect 92812 22492 92852 22532
rect 93964 22492 94004 22532
rect 94348 22492 94388 22532
rect 94636 22492 94676 22532
rect 95500 22492 95540 22532
rect 95884 22492 95924 22532
rect 96268 22492 96308 22532
rect 96748 22492 96788 22532
rect 97036 22492 97076 22532
rect 97612 22492 97652 22532
rect 97996 22492 98036 22532
rect 652 22408 692 22448
rect 75052 22408 75092 22448
rect 95116 22408 95156 22448
rect 74764 22324 74804 22364
rect 75244 22324 75284 22364
rect 75628 22324 75668 22364
rect 76108 22324 76148 22364
rect 77740 22324 77780 22364
rect 78124 22324 78164 22364
rect 79564 22324 79604 22364
rect 79948 22324 79988 22364
rect 80428 22324 80468 22364
rect 81292 22324 81332 22364
rect 81676 22324 81716 22364
rect 83212 22324 83252 22364
rect 83788 22324 83828 22364
rect 84556 22324 84596 22364
rect 84940 22324 84980 22364
rect 85612 22324 85652 22364
rect 85804 22324 85844 22364
rect 86380 22324 86420 22364
rect 86572 22324 86612 22364
rect 87244 22324 87284 22364
rect 87628 22324 87668 22364
rect 88012 22324 88052 22364
rect 88396 22324 88436 22364
rect 88876 22324 88916 22364
rect 89740 22324 89780 22364
rect 90412 22324 90452 22364
rect 90604 22324 90644 22364
rect 91276 22324 91316 22364
rect 91852 22324 91892 22364
rect 92236 22324 92276 22364
rect 92620 22324 92660 22364
rect 93004 22324 93044 22364
rect 93772 22324 93812 22364
rect 94156 22324 94196 22364
rect 94924 22324 94964 22364
rect 95308 22324 95348 22364
rect 95692 22324 95732 22364
rect 96076 22324 96116 22364
rect 96556 22324 96596 22364
rect 97228 22324 97268 22364
rect 97804 22324 97844 22364
rect 98188 22324 98228 22364
rect 73804 22240 73844 22280
rect 75820 22240 75860 22280
rect 76588 22240 76628 22280
rect 77164 22240 77204 22280
rect 78796 22240 78836 22280
rect 80908 22240 80948 22280
rect 83500 22240 83540 22280
rect 84268 22240 84308 22280
rect 86956 22240 86996 22280
rect 90988 22240 91028 22280
rect 91084 22240 91124 22280
rect 93484 22240 93524 22280
rect 94540 22240 94580 22280
rect 93580 22156 93620 22196
rect 78892 22072 78932 22112
rect 84172 22072 84212 22112
rect 86188 22072 86228 22112
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 8352 21904 8392 21944
rect 8434 21904 8474 21944
rect 8516 21904 8556 21944
rect 8598 21904 8638 21944
rect 8680 21904 8720 21944
rect 12352 21904 12392 21944
rect 12434 21904 12474 21944
rect 12516 21904 12556 21944
rect 12598 21904 12638 21944
rect 12680 21904 12720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 20352 21904 20392 21944
rect 20434 21904 20474 21944
rect 20516 21904 20556 21944
rect 20598 21904 20638 21944
rect 20680 21904 20720 21944
rect 24352 21904 24392 21944
rect 24434 21904 24474 21944
rect 24516 21904 24556 21944
rect 24598 21904 24638 21944
rect 24680 21904 24720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 32352 21904 32392 21944
rect 32434 21904 32474 21944
rect 32516 21904 32556 21944
rect 32598 21904 32638 21944
rect 32680 21904 32720 21944
rect 36352 21904 36392 21944
rect 36434 21904 36474 21944
rect 36516 21904 36556 21944
rect 36598 21904 36638 21944
rect 36680 21904 36720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 44352 21904 44392 21944
rect 44434 21904 44474 21944
rect 44516 21904 44556 21944
rect 44598 21904 44638 21944
rect 44680 21904 44720 21944
rect 48352 21904 48392 21944
rect 48434 21904 48474 21944
rect 48516 21904 48556 21944
rect 48598 21904 48638 21944
rect 48680 21904 48720 21944
rect 52352 21904 52392 21944
rect 52434 21904 52474 21944
rect 52516 21904 52556 21944
rect 52598 21904 52638 21944
rect 52680 21904 52720 21944
rect 56352 21904 56392 21944
rect 56434 21904 56474 21944
rect 56516 21904 56556 21944
rect 56598 21904 56638 21944
rect 56680 21904 56720 21944
rect 60352 21904 60392 21944
rect 60434 21904 60474 21944
rect 60516 21904 60556 21944
rect 60598 21904 60638 21944
rect 60680 21904 60720 21944
rect 64352 21904 64392 21944
rect 64434 21904 64474 21944
rect 64516 21904 64556 21944
rect 64598 21904 64638 21944
rect 64680 21904 64720 21944
rect 68352 21904 68392 21944
rect 68434 21904 68474 21944
rect 68516 21904 68556 21944
rect 68598 21904 68638 21944
rect 68680 21904 68720 21944
rect 72352 21904 72392 21944
rect 72434 21904 72474 21944
rect 72516 21904 72556 21944
rect 72598 21904 72638 21944
rect 72680 21904 72720 21944
rect 76352 21904 76392 21944
rect 76434 21904 76474 21944
rect 76516 21904 76556 21944
rect 76598 21904 76638 21944
rect 76680 21904 76720 21944
rect 80352 21904 80392 21944
rect 80434 21904 80474 21944
rect 80516 21904 80556 21944
rect 80598 21904 80638 21944
rect 80680 21904 80720 21944
rect 84352 21904 84392 21944
rect 84434 21904 84474 21944
rect 84516 21904 84556 21944
rect 84598 21904 84638 21944
rect 84680 21904 84720 21944
rect 88352 21904 88392 21944
rect 88434 21904 88474 21944
rect 88516 21904 88556 21944
rect 88598 21904 88638 21944
rect 88680 21904 88720 21944
rect 92352 21904 92392 21944
rect 92434 21904 92474 21944
rect 92516 21904 92556 21944
rect 92598 21904 92638 21944
rect 92680 21904 92720 21944
rect 96352 21904 96392 21944
rect 96434 21904 96474 21944
rect 96516 21904 96556 21944
rect 96598 21904 96638 21944
rect 96680 21904 96720 21944
rect 75820 21736 75860 21776
rect 76780 21736 76820 21776
rect 77644 21736 77684 21776
rect 79084 21736 79124 21776
rect 79468 21736 79508 21776
rect 81004 21736 81044 21776
rect 82348 21736 82388 21776
rect 82540 21736 82580 21776
rect 83596 21736 83636 21776
rect 84364 21736 84404 21776
rect 85996 21736 86036 21776
rect 86380 21736 86420 21776
rect 86860 21736 86900 21776
rect 89068 21736 89108 21776
rect 89548 21736 89588 21776
rect 91180 21736 91220 21776
rect 92812 21736 92852 21776
rect 93292 21736 93332 21776
rect 95212 21736 95252 21776
rect 75724 21568 75764 21608
rect 77548 21568 77588 21608
rect 82636 21568 82676 21608
rect 85900 21568 85940 21608
rect 86476 21568 86516 21608
rect 86764 21568 86804 21608
rect 89164 21568 89204 21608
rect 91084 21568 91124 21608
rect 92716 21568 92756 21608
rect 93388 21568 93428 21608
rect 95308 21568 95348 21608
rect 76588 21484 76628 21524
rect 78892 21484 78932 21524
rect 79276 21484 79316 21524
rect 80812 21484 80852 21524
rect 82156 21484 82196 21524
rect 83404 21484 83444 21524
rect 84172 21484 84212 21524
rect 89356 21484 89396 21524
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 7112 21148 7152 21188
rect 7194 21148 7234 21188
rect 7276 21148 7316 21188
rect 7358 21148 7398 21188
rect 7440 21148 7480 21188
rect 11112 21148 11152 21188
rect 11194 21148 11234 21188
rect 11276 21148 11316 21188
rect 11358 21148 11398 21188
rect 11440 21148 11480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 19112 21148 19152 21188
rect 19194 21148 19234 21188
rect 19276 21148 19316 21188
rect 19358 21148 19398 21188
rect 19440 21148 19480 21188
rect 23112 21148 23152 21188
rect 23194 21148 23234 21188
rect 23276 21148 23316 21188
rect 23358 21148 23398 21188
rect 23440 21148 23480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 31112 21148 31152 21188
rect 31194 21148 31234 21188
rect 31276 21148 31316 21188
rect 31358 21148 31398 21188
rect 31440 21148 31480 21188
rect 35112 21148 35152 21188
rect 35194 21148 35234 21188
rect 35276 21148 35316 21188
rect 35358 21148 35398 21188
rect 35440 21148 35480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 43112 21148 43152 21188
rect 43194 21148 43234 21188
rect 43276 21148 43316 21188
rect 43358 21148 43398 21188
rect 43440 21148 43480 21188
rect 47112 21148 47152 21188
rect 47194 21148 47234 21188
rect 47276 21148 47316 21188
rect 47358 21148 47398 21188
rect 47440 21148 47480 21188
rect 51112 21148 51152 21188
rect 51194 21148 51234 21188
rect 51276 21148 51316 21188
rect 51358 21148 51398 21188
rect 51440 21148 51480 21188
rect 55112 21148 55152 21188
rect 55194 21148 55234 21188
rect 55276 21148 55316 21188
rect 55358 21148 55398 21188
rect 55440 21148 55480 21188
rect 59112 21148 59152 21188
rect 59194 21148 59234 21188
rect 59276 21148 59316 21188
rect 59358 21148 59398 21188
rect 59440 21148 59480 21188
rect 63112 21148 63152 21188
rect 63194 21148 63234 21188
rect 63276 21148 63316 21188
rect 63358 21148 63398 21188
rect 63440 21148 63480 21188
rect 67112 21148 67152 21188
rect 67194 21148 67234 21188
rect 67276 21148 67316 21188
rect 67358 21148 67398 21188
rect 67440 21148 67480 21188
rect 71112 21148 71152 21188
rect 71194 21148 71234 21188
rect 71276 21148 71316 21188
rect 71358 21148 71398 21188
rect 71440 21148 71480 21188
rect 75112 21148 75152 21188
rect 75194 21148 75234 21188
rect 75276 21148 75316 21188
rect 75358 21148 75398 21188
rect 75440 21148 75480 21188
rect 79112 21148 79152 21188
rect 79194 21148 79234 21188
rect 79276 21148 79316 21188
rect 79358 21148 79398 21188
rect 79440 21148 79480 21188
rect 83112 21148 83152 21188
rect 83194 21148 83234 21188
rect 83276 21148 83316 21188
rect 83358 21148 83398 21188
rect 83440 21148 83480 21188
rect 87112 21148 87152 21188
rect 87194 21148 87234 21188
rect 87276 21148 87316 21188
rect 87358 21148 87398 21188
rect 87440 21148 87480 21188
rect 91112 21148 91152 21188
rect 91194 21148 91234 21188
rect 91276 21148 91316 21188
rect 91358 21148 91398 21188
rect 91440 21148 91480 21188
rect 95112 21148 95152 21188
rect 95194 21148 95234 21188
rect 95276 21148 95316 21188
rect 95358 21148 95398 21188
rect 95440 21148 95480 21188
rect 99112 21148 99152 21188
rect 99194 21148 99234 21188
rect 99276 21148 99316 21188
rect 99358 21148 99398 21188
rect 99440 21148 99480 21188
rect 652 20896 692 20936
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 8352 20392 8392 20432
rect 8434 20392 8474 20432
rect 8516 20392 8556 20432
rect 8598 20392 8638 20432
rect 8680 20392 8720 20432
rect 12352 20392 12392 20432
rect 12434 20392 12474 20432
rect 12516 20392 12556 20432
rect 12598 20392 12638 20432
rect 12680 20392 12720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 20352 20392 20392 20432
rect 20434 20392 20474 20432
rect 20516 20392 20556 20432
rect 20598 20392 20638 20432
rect 20680 20392 20720 20432
rect 24352 20392 24392 20432
rect 24434 20392 24474 20432
rect 24516 20392 24556 20432
rect 24598 20392 24638 20432
rect 24680 20392 24720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 32352 20392 32392 20432
rect 32434 20392 32474 20432
rect 32516 20392 32556 20432
rect 32598 20392 32638 20432
rect 32680 20392 32720 20432
rect 36352 20392 36392 20432
rect 36434 20392 36474 20432
rect 36516 20392 36556 20432
rect 36598 20392 36638 20432
rect 36680 20392 36720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 44352 20392 44392 20432
rect 44434 20392 44474 20432
rect 44516 20392 44556 20432
rect 44598 20392 44638 20432
rect 44680 20392 44720 20432
rect 48352 20392 48392 20432
rect 48434 20392 48474 20432
rect 48516 20392 48556 20432
rect 48598 20392 48638 20432
rect 48680 20392 48720 20432
rect 52352 20392 52392 20432
rect 52434 20392 52474 20432
rect 52516 20392 52556 20432
rect 52598 20392 52638 20432
rect 52680 20392 52720 20432
rect 56352 20392 56392 20432
rect 56434 20392 56474 20432
rect 56516 20392 56556 20432
rect 56598 20392 56638 20432
rect 56680 20392 56720 20432
rect 60352 20392 60392 20432
rect 60434 20392 60474 20432
rect 60516 20392 60556 20432
rect 60598 20392 60638 20432
rect 60680 20392 60720 20432
rect 64352 20392 64392 20432
rect 64434 20392 64474 20432
rect 64516 20392 64556 20432
rect 64598 20392 64638 20432
rect 64680 20392 64720 20432
rect 68352 20392 68392 20432
rect 68434 20392 68474 20432
rect 68516 20392 68556 20432
rect 68598 20392 68638 20432
rect 68680 20392 68720 20432
rect 72352 20392 72392 20432
rect 72434 20392 72474 20432
rect 72516 20392 72556 20432
rect 72598 20392 72638 20432
rect 72680 20392 72720 20432
rect 76352 20392 76392 20432
rect 76434 20392 76474 20432
rect 76516 20392 76556 20432
rect 76598 20392 76638 20432
rect 76680 20392 76720 20432
rect 80352 20392 80392 20432
rect 80434 20392 80474 20432
rect 80516 20392 80556 20432
rect 80598 20392 80638 20432
rect 80680 20392 80720 20432
rect 84352 20392 84392 20432
rect 84434 20392 84474 20432
rect 84516 20392 84556 20432
rect 84598 20392 84638 20432
rect 84680 20392 84720 20432
rect 88352 20392 88392 20432
rect 88434 20392 88474 20432
rect 88516 20392 88556 20432
rect 88598 20392 88638 20432
rect 88680 20392 88720 20432
rect 92352 20392 92392 20432
rect 92434 20392 92474 20432
rect 92516 20392 92556 20432
rect 92598 20392 92638 20432
rect 92680 20392 92720 20432
rect 96352 20392 96392 20432
rect 96434 20392 96474 20432
rect 96516 20392 96556 20432
rect 96598 20392 96638 20432
rect 96680 20392 96720 20432
rect 75532 19972 75572 20012
rect 80620 19972 80660 20012
rect 86860 19972 86900 20012
rect 93196 19972 93236 20012
rect 652 19888 692 19928
rect 75724 19888 75764 19928
rect 80428 19804 80468 19844
rect 87052 19804 87092 19844
rect 93004 19804 93044 19844
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 7112 19636 7152 19676
rect 7194 19636 7234 19676
rect 7276 19636 7316 19676
rect 7358 19636 7398 19676
rect 7440 19636 7480 19676
rect 11112 19636 11152 19676
rect 11194 19636 11234 19676
rect 11276 19636 11316 19676
rect 11358 19636 11398 19676
rect 11440 19636 11480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 19112 19636 19152 19676
rect 19194 19636 19234 19676
rect 19276 19636 19316 19676
rect 19358 19636 19398 19676
rect 19440 19636 19480 19676
rect 23112 19636 23152 19676
rect 23194 19636 23234 19676
rect 23276 19636 23316 19676
rect 23358 19636 23398 19676
rect 23440 19636 23480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 31112 19636 31152 19676
rect 31194 19636 31234 19676
rect 31276 19636 31316 19676
rect 31358 19636 31398 19676
rect 31440 19636 31480 19676
rect 35112 19636 35152 19676
rect 35194 19636 35234 19676
rect 35276 19636 35316 19676
rect 35358 19636 35398 19676
rect 35440 19636 35480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 43112 19636 43152 19676
rect 43194 19636 43234 19676
rect 43276 19636 43316 19676
rect 43358 19636 43398 19676
rect 43440 19636 43480 19676
rect 47112 19636 47152 19676
rect 47194 19636 47234 19676
rect 47276 19636 47316 19676
rect 47358 19636 47398 19676
rect 47440 19636 47480 19676
rect 51112 19636 51152 19676
rect 51194 19636 51234 19676
rect 51276 19636 51316 19676
rect 51358 19636 51398 19676
rect 51440 19636 51480 19676
rect 55112 19636 55152 19676
rect 55194 19636 55234 19676
rect 55276 19636 55316 19676
rect 55358 19636 55398 19676
rect 55440 19636 55480 19676
rect 59112 19636 59152 19676
rect 59194 19636 59234 19676
rect 59276 19636 59316 19676
rect 59358 19636 59398 19676
rect 59440 19636 59480 19676
rect 63112 19636 63152 19676
rect 63194 19636 63234 19676
rect 63276 19636 63316 19676
rect 63358 19636 63398 19676
rect 63440 19636 63480 19676
rect 67112 19636 67152 19676
rect 67194 19636 67234 19676
rect 67276 19636 67316 19676
rect 67358 19636 67398 19676
rect 67440 19636 67480 19676
rect 71112 19636 71152 19676
rect 71194 19636 71234 19676
rect 71276 19636 71316 19676
rect 71358 19636 71398 19676
rect 71440 19636 71480 19676
rect 75112 19636 75152 19676
rect 75194 19636 75234 19676
rect 75276 19636 75316 19676
rect 75358 19636 75398 19676
rect 75440 19636 75480 19676
rect 79112 19636 79152 19676
rect 79194 19636 79234 19676
rect 79276 19636 79316 19676
rect 79358 19636 79398 19676
rect 79440 19636 79480 19676
rect 83112 19636 83152 19676
rect 83194 19636 83234 19676
rect 83276 19636 83316 19676
rect 83358 19636 83398 19676
rect 83440 19636 83480 19676
rect 87112 19636 87152 19676
rect 87194 19636 87234 19676
rect 87276 19636 87316 19676
rect 87358 19636 87398 19676
rect 87440 19636 87480 19676
rect 91112 19636 91152 19676
rect 91194 19636 91234 19676
rect 91276 19636 91316 19676
rect 91358 19636 91398 19676
rect 91440 19636 91480 19676
rect 95112 19636 95152 19676
rect 95194 19636 95234 19676
rect 95276 19636 95316 19676
rect 95358 19636 95398 19676
rect 95440 19636 95480 19676
rect 99112 19636 99152 19676
rect 99194 19636 99234 19676
rect 99276 19636 99316 19676
rect 99358 19636 99398 19676
rect 99440 19636 99480 19676
rect 90124 19468 90164 19508
rect 652 19384 692 19424
rect 92908 19384 92948 19424
rect 74764 19300 74804 19340
rect 77644 19300 77684 19340
rect 78220 19300 78260 19340
rect 80524 19300 80564 19340
rect 82060 19300 82100 19340
rect 84076 19300 84116 19340
rect 85612 19300 85652 19340
rect 86572 19300 86612 19340
rect 86764 19300 86804 19340
rect 87436 19300 87476 19340
rect 88204 19300 88244 19340
rect 89740 19300 89780 19340
rect 89932 19300 89972 19340
rect 91372 19300 91412 19340
rect 92524 19300 92564 19340
rect 93100 19300 93140 19340
rect 94156 19300 94196 19340
rect 95788 19300 95828 19340
rect 75244 19216 75284 19256
rect 75436 19216 75476 19256
rect 75628 19216 75668 19256
rect 76588 19216 76628 19256
rect 77068 19216 77108 19256
rect 78604 19216 78644 19256
rect 80044 19216 80084 19256
rect 82636 19216 82676 19256
rect 88492 19216 88532 19256
rect 74956 19048 74996 19088
rect 75724 19048 75764 19088
rect 76684 19048 76724 19088
rect 77164 19048 77204 19088
rect 77836 19048 77876 19088
rect 78028 19048 78068 19088
rect 78700 19048 78740 19088
rect 80140 19048 80180 19088
rect 80332 19048 80372 19088
rect 81868 19048 81908 19088
rect 82732 19048 82772 19088
rect 83884 19048 83924 19088
rect 85804 19048 85844 19088
rect 86380 19048 86420 19088
rect 86956 19048 86996 19088
rect 87628 19048 87668 19088
rect 88012 19048 88052 19088
rect 88396 19048 88436 19088
rect 89548 19048 89588 19088
rect 90124 19048 90164 19088
rect 91564 19048 91604 19088
rect 92716 19048 92756 19088
rect 93964 19048 94004 19088
rect 95596 19048 95636 19088
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 8352 18880 8392 18920
rect 8434 18880 8474 18920
rect 8516 18880 8556 18920
rect 8598 18880 8638 18920
rect 8680 18880 8720 18920
rect 12352 18880 12392 18920
rect 12434 18880 12474 18920
rect 12516 18880 12556 18920
rect 12598 18880 12638 18920
rect 12680 18880 12720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 20352 18880 20392 18920
rect 20434 18880 20474 18920
rect 20516 18880 20556 18920
rect 20598 18880 20638 18920
rect 20680 18880 20720 18920
rect 24352 18880 24392 18920
rect 24434 18880 24474 18920
rect 24516 18880 24556 18920
rect 24598 18880 24638 18920
rect 24680 18880 24720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 32352 18880 32392 18920
rect 32434 18880 32474 18920
rect 32516 18880 32556 18920
rect 32598 18880 32638 18920
rect 32680 18880 32720 18920
rect 36352 18880 36392 18920
rect 36434 18880 36474 18920
rect 36516 18880 36556 18920
rect 36598 18880 36638 18920
rect 36680 18880 36720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 44352 18880 44392 18920
rect 44434 18880 44474 18920
rect 44516 18880 44556 18920
rect 44598 18880 44638 18920
rect 44680 18880 44720 18920
rect 48352 18880 48392 18920
rect 48434 18880 48474 18920
rect 48516 18880 48556 18920
rect 48598 18880 48638 18920
rect 48680 18880 48720 18920
rect 52352 18880 52392 18920
rect 52434 18880 52474 18920
rect 52516 18880 52556 18920
rect 52598 18880 52638 18920
rect 52680 18880 52720 18920
rect 56352 18880 56392 18920
rect 56434 18880 56474 18920
rect 56516 18880 56556 18920
rect 56598 18880 56638 18920
rect 56680 18880 56720 18920
rect 60352 18880 60392 18920
rect 60434 18880 60474 18920
rect 60516 18880 60556 18920
rect 60598 18880 60638 18920
rect 60680 18880 60720 18920
rect 64352 18880 64392 18920
rect 64434 18880 64474 18920
rect 64516 18880 64556 18920
rect 64598 18880 64638 18920
rect 64680 18880 64720 18920
rect 68352 18880 68392 18920
rect 68434 18880 68474 18920
rect 68516 18880 68556 18920
rect 68598 18880 68638 18920
rect 68680 18880 68720 18920
rect 72352 18880 72392 18920
rect 72434 18880 72474 18920
rect 72516 18880 72556 18920
rect 72598 18880 72638 18920
rect 72680 18880 72720 18920
rect 76352 18880 76392 18920
rect 76434 18880 76474 18920
rect 76516 18880 76556 18920
rect 76598 18880 76638 18920
rect 76680 18880 76720 18920
rect 80352 18880 80392 18920
rect 80434 18880 80474 18920
rect 80516 18880 80556 18920
rect 80598 18880 80638 18920
rect 80680 18880 80720 18920
rect 84352 18880 84392 18920
rect 84434 18880 84474 18920
rect 84516 18880 84556 18920
rect 84598 18880 84638 18920
rect 84680 18880 84720 18920
rect 88352 18880 88392 18920
rect 88434 18880 88474 18920
rect 88516 18880 88556 18920
rect 88598 18880 88638 18920
rect 88680 18880 88720 18920
rect 92352 18880 92392 18920
rect 92434 18880 92474 18920
rect 92516 18880 92556 18920
rect 92598 18880 92638 18920
rect 92680 18880 92720 18920
rect 96352 18880 96392 18920
rect 96434 18880 96474 18920
rect 96516 18880 96556 18920
rect 96598 18880 96638 18920
rect 96680 18880 96720 18920
rect 74956 18712 74996 18752
rect 72940 18544 72980 18584
rect 74284 18544 74324 18584
rect 76492 18544 76532 18584
rect 77452 18544 77492 18584
rect 78124 18544 78164 18584
rect 85036 18544 85076 18584
rect 86284 18544 86324 18584
rect 89452 18555 89492 18595
rect 92908 18544 92948 18584
rect 95116 18544 95156 18584
rect 95980 18544 96020 18584
rect 96940 18544 96980 18584
rect 97612 18544 97652 18584
rect 74572 18460 74612 18500
rect 75148 18460 75188 18500
rect 75820 18460 75860 18500
rect 78412 18460 78452 18500
rect 78988 18460 79028 18500
rect 79372 18460 79412 18500
rect 79852 18460 79892 18500
rect 81004 18460 81044 18500
rect 81388 18460 81428 18500
rect 81772 18460 81812 18500
rect 82252 18460 82292 18500
rect 83020 18460 83060 18500
rect 83404 18460 83444 18500
rect 83788 18460 83828 18500
rect 84268 18460 84308 18500
rect 84652 18460 84692 18500
rect 85516 18460 85556 18500
rect 85900 18460 85940 18500
rect 86572 18460 86612 18500
rect 87052 18460 87092 18500
rect 87724 18460 87764 18500
rect 88204 18460 88244 18500
rect 88588 18460 88628 18500
rect 88972 18460 89012 18500
rect 89740 18460 89780 18500
rect 90124 18460 90164 18500
rect 90604 18460 90644 18500
rect 91276 18460 91316 18500
rect 91852 18460 91892 18500
rect 92236 18460 92276 18500
rect 92620 18460 92660 18500
rect 93100 18460 93140 18500
rect 93868 18460 93908 18500
rect 94252 18460 94292 18500
rect 94924 18460 94964 18500
rect 95500 18460 95540 18500
rect 96268 18460 96308 18500
rect 97132 18460 97172 18500
rect 652 18376 692 18416
rect 78796 18376 78836 18416
rect 73036 18292 73076 18332
rect 74188 18292 74228 18332
rect 74764 18292 74804 18332
rect 74956 18292 74996 18332
rect 76012 18292 76052 18332
rect 76588 18292 76628 18332
rect 77548 18292 77588 18332
rect 78220 18292 78260 18332
rect 78604 18292 78644 18332
rect 79564 18292 79604 18332
rect 80044 18292 80084 18332
rect 81196 18292 81236 18332
rect 81580 18292 81620 18332
rect 81964 18292 82004 18332
rect 82444 18292 82484 18332
rect 83212 18292 83252 18332
rect 83596 18292 83636 18332
rect 83980 18292 84020 18332
rect 84460 18292 84500 18332
rect 84844 18292 84884 18332
rect 85132 18292 85172 18332
rect 85708 18292 85748 18332
rect 86092 18292 86132 18332
rect 86380 18292 86420 18332
rect 86764 18292 86804 18332
rect 87244 18292 87284 18332
rect 87916 18292 87956 18332
rect 88396 18292 88436 18332
rect 88780 18292 88820 18332
rect 89164 18292 89204 18332
rect 89548 18292 89588 18332
rect 89932 18292 89972 18332
rect 90316 18292 90356 18332
rect 90796 18292 90836 18332
rect 91468 18292 91508 18332
rect 91660 18292 91700 18332
rect 92044 18292 92084 18332
rect 92428 18292 92468 18332
rect 92812 18292 92852 18332
rect 93292 18292 93332 18332
rect 94060 18292 94100 18332
rect 94444 18292 94484 18332
rect 94732 18292 94772 18332
rect 95212 18292 95252 18332
rect 95692 18292 95732 18332
rect 95884 18292 95924 18332
rect 96460 18292 96500 18332
rect 96844 18292 96884 18332
rect 97324 18292 97364 18332
rect 97516 18292 97556 18332
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 7112 18124 7152 18164
rect 7194 18124 7234 18164
rect 7276 18124 7316 18164
rect 7358 18124 7398 18164
rect 7440 18124 7480 18164
rect 11112 18124 11152 18164
rect 11194 18124 11234 18164
rect 11276 18124 11316 18164
rect 11358 18124 11398 18164
rect 11440 18124 11480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 19112 18124 19152 18164
rect 19194 18124 19234 18164
rect 19276 18124 19316 18164
rect 19358 18124 19398 18164
rect 19440 18124 19480 18164
rect 23112 18124 23152 18164
rect 23194 18124 23234 18164
rect 23276 18124 23316 18164
rect 23358 18124 23398 18164
rect 23440 18124 23480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 31112 18124 31152 18164
rect 31194 18124 31234 18164
rect 31276 18124 31316 18164
rect 31358 18124 31398 18164
rect 31440 18124 31480 18164
rect 35112 18124 35152 18164
rect 35194 18124 35234 18164
rect 35276 18124 35316 18164
rect 35358 18124 35398 18164
rect 35440 18124 35480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 43112 18124 43152 18164
rect 43194 18124 43234 18164
rect 43276 18124 43316 18164
rect 43358 18124 43398 18164
rect 43440 18124 43480 18164
rect 47112 18124 47152 18164
rect 47194 18124 47234 18164
rect 47276 18124 47316 18164
rect 47358 18124 47398 18164
rect 47440 18124 47480 18164
rect 51112 18124 51152 18164
rect 51194 18124 51234 18164
rect 51276 18124 51316 18164
rect 51358 18124 51398 18164
rect 51440 18124 51480 18164
rect 55112 18124 55152 18164
rect 55194 18124 55234 18164
rect 55276 18124 55316 18164
rect 55358 18124 55398 18164
rect 55440 18124 55480 18164
rect 59112 18124 59152 18164
rect 59194 18124 59234 18164
rect 59276 18124 59316 18164
rect 59358 18124 59398 18164
rect 59440 18124 59480 18164
rect 63112 18124 63152 18164
rect 63194 18124 63234 18164
rect 63276 18124 63316 18164
rect 63358 18124 63398 18164
rect 63440 18124 63480 18164
rect 67112 18124 67152 18164
rect 67194 18124 67234 18164
rect 67276 18124 67316 18164
rect 67358 18124 67398 18164
rect 67440 18124 67480 18164
rect 71112 18124 71152 18164
rect 71194 18124 71234 18164
rect 71276 18124 71316 18164
rect 71358 18124 71398 18164
rect 71440 18124 71480 18164
rect 75112 18124 75152 18164
rect 75194 18124 75234 18164
rect 75276 18124 75316 18164
rect 75358 18124 75398 18164
rect 75440 18124 75480 18164
rect 79112 18124 79152 18164
rect 79194 18124 79234 18164
rect 79276 18124 79316 18164
rect 79358 18124 79398 18164
rect 79440 18124 79480 18164
rect 83112 18124 83152 18164
rect 83194 18124 83234 18164
rect 83276 18124 83316 18164
rect 83358 18124 83398 18164
rect 83440 18124 83480 18164
rect 87112 18124 87152 18164
rect 87194 18124 87234 18164
rect 87276 18124 87316 18164
rect 87358 18124 87398 18164
rect 87440 18124 87480 18164
rect 91112 18124 91152 18164
rect 91194 18124 91234 18164
rect 91276 18124 91316 18164
rect 91358 18124 91398 18164
rect 91440 18124 91480 18164
rect 95112 18124 95152 18164
rect 95194 18124 95234 18164
rect 95276 18124 95316 18164
rect 95358 18124 95398 18164
rect 95440 18124 95480 18164
rect 99112 18124 99152 18164
rect 99194 18124 99234 18164
rect 99276 18124 99316 18164
rect 99358 18124 99398 18164
rect 99440 18124 99480 18164
rect 652 17872 692 17912
rect 98284 17872 98324 17912
rect 73708 17788 73748 17828
rect 74092 17788 74132 17828
rect 74476 17788 74516 17828
rect 75340 17788 75380 17828
rect 76204 17788 76244 17828
rect 76588 17788 76628 17828
rect 76972 17788 77012 17828
rect 77356 17788 77396 17828
rect 78220 17788 78260 17828
rect 78700 17788 78740 17828
rect 80140 17788 80180 17828
rect 80524 17788 80564 17828
rect 82636 17788 82676 17828
rect 84940 17788 84980 17828
rect 86188 17788 86228 17828
rect 89452 17788 89492 17828
rect 93772 17788 93812 17828
rect 95020 17788 95060 17828
rect 95884 17788 95924 17828
rect 96652 17788 96692 17828
rect 97036 17788 97076 17828
rect 97900 17788 97940 17828
rect 98476 17788 98516 17828
rect 75052 17704 75092 17744
rect 75820 17704 75860 17744
rect 77740 17704 77780 17744
rect 79180 17704 79220 17744
rect 79468 17704 79508 17744
rect 79852 17704 79892 17744
rect 81004 17704 81044 17744
rect 81292 17704 81332 17744
rect 81484 17704 81524 17744
rect 81964 17704 82004 17744
rect 82252 17704 82292 17744
rect 83020 17704 83060 17744
rect 83404 17704 83444 17744
rect 83788 17704 83828 17744
rect 84172 17704 84212 17744
rect 84748 17704 84788 17744
rect 85420 17704 85460 17744
rect 85804 17704 85844 17744
rect 86572 17704 86612 17744
rect 87052 17704 87092 17744
rect 87436 17704 87476 17744
rect 88204 17704 88244 17744
rect 88588 17704 88628 17744
rect 89068 17704 89108 17744
rect 89932 17704 89972 17744
rect 90220 17704 90260 17744
rect 90604 17704 90644 17744
rect 90988 17704 91028 17744
rect 91372 17704 91412 17744
rect 91852 17704 91892 17744
rect 92236 17704 92276 17744
rect 92812 17704 92852 17744
rect 93188 17709 93228 17749
rect 94060 17704 94100 17744
rect 94252 17704 94292 17744
rect 94732 17704 94772 17744
rect 95404 17704 95444 17744
rect 96364 17704 96404 17744
rect 97420 17704 97460 17744
rect 98668 17704 98708 17744
rect 81868 17620 81908 17660
rect 84652 17620 84692 17660
rect 92908 17620 92948 17660
rect 98764 17620 98804 17660
rect 73900 17536 73940 17576
rect 74284 17536 74324 17576
rect 74668 17536 74708 17576
rect 75148 17536 75188 17576
rect 75532 17536 75572 17576
rect 75724 17536 75764 17576
rect 76396 17536 76436 17576
rect 76780 17536 76820 17576
rect 77164 17536 77204 17576
rect 77548 17536 77588 17576
rect 77836 17536 77876 17576
rect 78412 17536 78452 17576
rect 78892 17536 78932 17576
rect 79084 17536 79124 17576
rect 79564 17536 79604 17576
rect 79948 17536 79988 17576
rect 80332 17536 80372 17576
rect 80716 17536 80756 17576
rect 80908 17536 80948 17576
rect 81196 17536 81236 17576
rect 81580 17536 81620 17576
rect 82348 17536 82388 17576
rect 82828 17536 82868 17576
rect 83116 17536 83156 17576
rect 83500 17536 83540 17576
rect 83884 17536 83924 17576
rect 84268 17536 84308 17576
rect 85132 17536 85172 17576
rect 85516 17536 85556 17576
rect 85900 17536 85940 17576
rect 86380 17536 86420 17576
rect 86668 17536 86708 17576
rect 87148 17536 87188 17576
rect 87532 17536 87572 17576
rect 88300 17536 88340 17576
rect 88684 17536 88724 17576
rect 89164 17536 89204 17576
rect 89644 17536 89684 17576
rect 89836 17536 89876 17576
rect 90316 17536 90356 17576
rect 90700 17536 90740 17576
rect 91084 17536 91124 17576
rect 91468 17536 91508 17576
rect 91948 17536 91988 17576
rect 92332 17536 92372 17576
rect 93100 17536 93140 17576
rect 93580 17536 93620 17576
rect 93964 17536 94004 17576
rect 94348 17536 94388 17576
rect 94828 17536 94868 17576
rect 95212 17536 95252 17576
rect 95500 17536 95540 17576
rect 96076 17536 96116 17576
rect 96268 17536 96308 17576
rect 96844 17536 96884 17576
rect 97228 17536 97268 17576
rect 97516 17536 97556 17576
rect 97708 17536 97748 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 8352 17368 8392 17408
rect 8434 17368 8474 17408
rect 8516 17368 8556 17408
rect 8598 17368 8638 17408
rect 8680 17368 8720 17408
rect 12352 17368 12392 17408
rect 12434 17368 12474 17408
rect 12516 17368 12556 17408
rect 12598 17368 12638 17408
rect 12680 17368 12720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 20352 17368 20392 17408
rect 20434 17368 20474 17408
rect 20516 17368 20556 17408
rect 20598 17368 20638 17408
rect 20680 17368 20720 17408
rect 24352 17368 24392 17408
rect 24434 17368 24474 17408
rect 24516 17368 24556 17408
rect 24598 17368 24638 17408
rect 24680 17368 24720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 32352 17368 32392 17408
rect 32434 17368 32474 17408
rect 32516 17368 32556 17408
rect 32598 17368 32638 17408
rect 32680 17368 32720 17408
rect 36352 17368 36392 17408
rect 36434 17368 36474 17408
rect 36516 17368 36556 17408
rect 36598 17368 36638 17408
rect 36680 17368 36720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 44352 17368 44392 17408
rect 44434 17368 44474 17408
rect 44516 17368 44556 17408
rect 44598 17368 44638 17408
rect 44680 17368 44720 17408
rect 48352 17368 48392 17408
rect 48434 17368 48474 17408
rect 48516 17368 48556 17408
rect 48598 17368 48638 17408
rect 48680 17368 48720 17408
rect 52352 17368 52392 17408
rect 52434 17368 52474 17408
rect 52516 17368 52556 17408
rect 52598 17368 52638 17408
rect 52680 17368 52720 17408
rect 56352 17368 56392 17408
rect 56434 17368 56474 17408
rect 56516 17368 56556 17408
rect 56598 17368 56638 17408
rect 56680 17368 56720 17408
rect 60352 17368 60392 17408
rect 60434 17368 60474 17408
rect 60516 17368 60556 17408
rect 60598 17368 60638 17408
rect 60680 17368 60720 17408
rect 64352 17368 64392 17408
rect 64434 17368 64474 17408
rect 64516 17368 64556 17408
rect 64598 17368 64638 17408
rect 64680 17368 64720 17408
rect 68352 17368 68392 17408
rect 68434 17368 68474 17408
rect 68516 17368 68556 17408
rect 68598 17368 68638 17408
rect 68680 17368 68720 17408
rect 72352 17368 72392 17408
rect 72434 17368 72474 17408
rect 72516 17368 72556 17408
rect 72598 17368 72638 17408
rect 72680 17368 72720 17408
rect 76352 17368 76392 17408
rect 76434 17368 76474 17408
rect 76516 17368 76556 17408
rect 76598 17368 76638 17408
rect 76680 17368 76720 17408
rect 80352 17368 80392 17408
rect 80434 17368 80474 17408
rect 80516 17368 80556 17408
rect 80598 17368 80638 17408
rect 80680 17368 80720 17408
rect 84352 17368 84392 17408
rect 84434 17368 84474 17408
rect 84516 17368 84556 17408
rect 84598 17368 84638 17408
rect 84680 17368 84720 17408
rect 88352 17368 88392 17408
rect 88434 17368 88474 17408
rect 88516 17368 88556 17408
rect 88598 17368 88638 17408
rect 88680 17368 88720 17408
rect 92352 17368 92392 17408
rect 92434 17368 92474 17408
rect 92516 17368 92556 17408
rect 92598 17368 92638 17408
rect 92680 17368 92720 17408
rect 96352 17368 96392 17408
rect 96434 17368 96474 17408
rect 96516 17368 96556 17408
rect 96598 17368 96638 17408
rect 96680 17368 96720 17408
rect 652 16864 692 16904
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 7112 16612 7152 16652
rect 7194 16612 7234 16652
rect 7276 16612 7316 16652
rect 7358 16612 7398 16652
rect 7440 16612 7480 16652
rect 11112 16612 11152 16652
rect 11194 16612 11234 16652
rect 11276 16612 11316 16652
rect 11358 16612 11398 16652
rect 11440 16612 11480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 19112 16612 19152 16652
rect 19194 16612 19234 16652
rect 19276 16612 19316 16652
rect 19358 16612 19398 16652
rect 19440 16612 19480 16652
rect 23112 16612 23152 16652
rect 23194 16612 23234 16652
rect 23276 16612 23316 16652
rect 23358 16612 23398 16652
rect 23440 16612 23480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 31112 16612 31152 16652
rect 31194 16612 31234 16652
rect 31276 16612 31316 16652
rect 31358 16612 31398 16652
rect 31440 16612 31480 16652
rect 35112 16612 35152 16652
rect 35194 16612 35234 16652
rect 35276 16612 35316 16652
rect 35358 16612 35398 16652
rect 35440 16612 35480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 43112 16612 43152 16652
rect 43194 16612 43234 16652
rect 43276 16612 43316 16652
rect 43358 16612 43398 16652
rect 43440 16612 43480 16652
rect 47112 16612 47152 16652
rect 47194 16612 47234 16652
rect 47276 16612 47316 16652
rect 47358 16612 47398 16652
rect 47440 16612 47480 16652
rect 51112 16612 51152 16652
rect 51194 16612 51234 16652
rect 51276 16612 51316 16652
rect 51358 16612 51398 16652
rect 51440 16612 51480 16652
rect 55112 16612 55152 16652
rect 55194 16612 55234 16652
rect 55276 16612 55316 16652
rect 55358 16612 55398 16652
rect 55440 16612 55480 16652
rect 59112 16612 59152 16652
rect 59194 16612 59234 16652
rect 59276 16612 59316 16652
rect 59358 16612 59398 16652
rect 59440 16612 59480 16652
rect 63112 16612 63152 16652
rect 63194 16612 63234 16652
rect 63276 16612 63316 16652
rect 63358 16612 63398 16652
rect 63440 16612 63480 16652
rect 67112 16612 67152 16652
rect 67194 16612 67234 16652
rect 67276 16612 67316 16652
rect 67358 16612 67398 16652
rect 67440 16612 67480 16652
rect 652 16360 692 16400
rect 69100 16276 69140 16316
rect 69292 16024 69332 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 8352 15856 8392 15896
rect 8434 15856 8474 15896
rect 8516 15856 8556 15896
rect 8598 15856 8638 15896
rect 8680 15856 8720 15896
rect 12352 15856 12392 15896
rect 12434 15856 12474 15896
rect 12516 15856 12556 15896
rect 12598 15856 12638 15896
rect 12680 15856 12720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 20352 15856 20392 15896
rect 20434 15856 20474 15896
rect 20516 15856 20556 15896
rect 20598 15856 20638 15896
rect 20680 15856 20720 15896
rect 24352 15856 24392 15896
rect 24434 15856 24474 15896
rect 24516 15856 24556 15896
rect 24598 15856 24638 15896
rect 24680 15856 24720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 32352 15856 32392 15896
rect 32434 15856 32474 15896
rect 32516 15856 32556 15896
rect 32598 15856 32638 15896
rect 32680 15856 32720 15896
rect 36352 15856 36392 15896
rect 36434 15856 36474 15896
rect 36516 15856 36556 15896
rect 36598 15856 36638 15896
rect 36680 15856 36720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 44352 15856 44392 15896
rect 44434 15856 44474 15896
rect 44516 15856 44556 15896
rect 44598 15856 44638 15896
rect 44680 15856 44720 15896
rect 48352 15856 48392 15896
rect 48434 15856 48474 15896
rect 48516 15856 48556 15896
rect 48598 15856 48638 15896
rect 48680 15856 48720 15896
rect 52352 15856 52392 15896
rect 52434 15856 52474 15896
rect 52516 15856 52556 15896
rect 52598 15856 52638 15896
rect 52680 15856 52720 15896
rect 56352 15856 56392 15896
rect 56434 15856 56474 15896
rect 56516 15856 56556 15896
rect 56598 15856 56638 15896
rect 56680 15856 56720 15896
rect 60352 15856 60392 15896
rect 60434 15856 60474 15896
rect 60516 15856 60556 15896
rect 60598 15856 60638 15896
rect 60680 15856 60720 15896
rect 64352 15856 64392 15896
rect 64434 15856 64474 15896
rect 64516 15856 64556 15896
rect 64598 15856 64638 15896
rect 64680 15856 64720 15896
rect 68352 15856 68392 15896
rect 68434 15856 68474 15896
rect 68516 15856 68556 15896
rect 68598 15856 68638 15896
rect 68680 15856 68720 15896
rect 67372 15688 67412 15728
rect 68236 15520 68276 15560
rect 68428 15520 68468 15560
rect 844 15436 884 15476
rect 1996 15436 2036 15476
rect 67180 15436 67220 15476
rect 67756 15436 67796 15476
rect 67564 15352 67604 15392
rect 652 15268 692 15308
rect 1804 15268 1844 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 7112 15100 7152 15140
rect 7194 15100 7234 15140
rect 7276 15100 7316 15140
rect 7358 15100 7398 15140
rect 7440 15100 7480 15140
rect 11112 15100 11152 15140
rect 11194 15100 11234 15140
rect 11276 15100 11316 15140
rect 11358 15100 11398 15140
rect 11440 15100 11480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 19112 15100 19152 15140
rect 19194 15100 19234 15140
rect 19276 15100 19316 15140
rect 19358 15100 19398 15140
rect 19440 15100 19480 15140
rect 23112 15100 23152 15140
rect 23194 15100 23234 15140
rect 23276 15100 23316 15140
rect 23358 15100 23398 15140
rect 23440 15100 23480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 31112 15100 31152 15140
rect 31194 15100 31234 15140
rect 31276 15100 31316 15140
rect 31358 15100 31398 15140
rect 31440 15100 31480 15140
rect 35112 15100 35152 15140
rect 35194 15100 35234 15140
rect 35276 15100 35316 15140
rect 35358 15100 35398 15140
rect 35440 15100 35480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 43112 15100 43152 15140
rect 43194 15100 43234 15140
rect 43276 15100 43316 15140
rect 43358 15100 43398 15140
rect 43440 15100 43480 15140
rect 47112 15100 47152 15140
rect 47194 15100 47234 15140
rect 47276 15100 47316 15140
rect 47358 15100 47398 15140
rect 47440 15100 47480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 55112 15100 55152 15140
rect 55194 15100 55234 15140
rect 55276 15100 55316 15140
rect 55358 15100 55398 15140
rect 55440 15100 55480 15140
rect 59112 15100 59152 15140
rect 59194 15100 59234 15140
rect 59276 15100 59316 15140
rect 59358 15100 59398 15140
rect 59440 15100 59480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 67112 15100 67152 15140
rect 67194 15100 67234 15140
rect 67276 15100 67316 15140
rect 67358 15100 67398 15140
rect 67440 15100 67480 15140
rect 1708 14932 1748 14972
rect 68716 14932 68756 14972
rect 69100 14932 69140 14972
rect 69484 14932 69524 14972
rect 69868 14932 69908 14972
rect 844 14764 884 14804
rect 1900 14764 1940 14804
rect 68044 14764 68084 14804
rect 69676 14764 69716 14804
rect 68140 14680 68180 14720
rect 68620 14680 68660 14720
rect 69004 14680 69044 14720
rect 69388 14680 69428 14720
rect 652 14512 692 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 8352 14344 8392 14384
rect 8434 14344 8474 14384
rect 8516 14344 8556 14384
rect 8598 14344 8638 14384
rect 8680 14344 8720 14384
rect 12352 14344 12392 14384
rect 12434 14344 12474 14384
rect 12516 14344 12556 14384
rect 12598 14344 12638 14384
rect 12680 14344 12720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 20352 14344 20392 14384
rect 20434 14344 20474 14384
rect 20516 14344 20556 14384
rect 20598 14344 20638 14384
rect 20680 14344 20720 14384
rect 24352 14344 24392 14384
rect 24434 14344 24474 14384
rect 24516 14344 24556 14384
rect 24598 14344 24638 14384
rect 24680 14344 24720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 32352 14344 32392 14384
rect 32434 14344 32474 14384
rect 32516 14344 32556 14384
rect 32598 14344 32638 14384
rect 32680 14344 32720 14384
rect 36352 14344 36392 14384
rect 36434 14344 36474 14384
rect 36516 14344 36556 14384
rect 36598 14344 36638 14384
rect 36680 14344 36720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 44352 14344 44392 14384
rect 44434 14344 44474 14384
rect 44516 14344 44556 14384
rect 44598 14344 44638 14384
rect 44680 14344 44720 14384
rect 48352 14344 48392 14384
rect 48434 14344 48474 14384
rect 48516 14344 48556 14384
rect 48598 14344 48638 14384
rect 48680 14344 48720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 56352 14344 56392 14384
rect 56434 14344 56474 14384
rect 56516 14344 56556 14384
rect 56598 14344 56638 14384
rect 56680 14344 56720 14384
rect 60352 14344 60392 14384
rect 60434 14344 60474 14384
rect 60516 14344 60556 14384
rect 60598 14344 60638 14384
rect 60680 14344 60720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 68352 14344 68392 14384
rect 68434 14344 68474 14384
rect 68516 14344 68556 14384
rect 68598 14344 68638 14384
rect 68680 14344 68720 14384
rect 1324 14176 1364 14216
rect 69388 14176 69428 14216
rect 69868 14176 69908 14216
rect 69772 14008 69812 14048
rect 1516 13924 1556 13964
rect 69196 13924 69236 13964
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 7112 13588 7152 13628
rect 7194 13588 7234 13628
rect 7276 13588 7316 13628
rect 7358 13588 7398 13628
rect 7440 13588 7480 13628
rect 11112 13588 11152 13628
rect 11194 13588 11234 13628
rect 11276 13588 11316 13628
rect 11358 13588 11398 13628
rect 11440 13588 11480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 19112 13588 19152 13628
rect 19194 13588 19234 13628
rect 19276 13588 19316 13628
rect 19358 13588 19398 13628
rect 19440 13588 19480 13628
rect 23112 13588 23152 13628
rect 23194 13588 23234 13628
rect 23276 13588 23316 13628
rect 23358 13588 23398 13628
rect 23440 13588 23480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 31112 13588 31152 13628
rect 31194 13588 31234 13628
rect 31276 13588 31316 13628
rect 31358 13588 31398 13628
rect 31440 13588 31480 13628
rect 35112 13588 35152 13628
rect 35194 13588 35234 13628
rect 35276 13588 35316 13628
rect 35358 13588 35398 13628
rect 35440 13588 35480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 43112 13588 43152 13628
rect 43194 13588 43234 13628
rect 43276 13588 43316 13628
rect 43358 13588 43398 13628
rect 43440 13588 43480 13628
rect 47112 13588 47152 13628
rect 47194 13588 47234 13628
rect 47276 13588 47316 13628
rect 47358 13588 47398 13628
rect 47440 13588 47480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 55112 13588 55152 13628
rect 55194 13588 55234 13628
rect 55276 13588 55316 13628
rect 55358 13588 55398 13628
rect 55440 13588 55480 13628
rect 59112 13588 59152 13628
rect 59194 13588 59234 13628
rect 59276 13588 59316 13628
rect 59358 13588 59398 13628
rect 59440 13588 59480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 67112 13588 67152 13628
rect 67194 13588 67234 13628
rect 67276 13588 67316 13628
rect 67358 13588 67398 13628
rect 67440 13588 67480 13628
rect 1708 13336 1748 13376
rect 844 13252 884 13292
rect 1900 13252 1940 13292
rect 652 13000 692 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 8352 12832 8392 12872
rect 8434 12832 8474 12872
rect 8516 12832 8556 12872
rect 8598 12832 8638 12872
rect 8680 12832 8720 12872
rect 12352 12832 12392 12872
rect 12434 12832 12474 12872
rect 12516 12832 12556 12872
rect 12598 12832 12638 12872
rect 12680 12832 12720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 20352 12832 20392 12872
rect 20434 12832 20474 12872
rect 20516 12832 20556 12872
rect 20598 12832 20638 12872
rect 20680 12832 20720 12872
rect 24352 12832 24392 12872
rect 24434 12832 24474 12872
rect 24516 12832 24556 12872
rect 24598 12832 24638 12872
rect 24680 12832 24720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 32352 12832 32392 12872
rect 32434 12832 32474 12872
rect 32516 12832 32556 12872
rect 32598 12832 32638 12872
rect 32680 12832 32720 12872
rect 36352 12832 36392 12872
rect 36434 12832 36474 12872
rect 36516 12832 36556 12872
rect 36598 12832 36638 12872
rect 36680 12832 36720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 44352 12832 44392 12872
rect 44434 12832 44474 12872
rect 44516 12832 44556 12872
rect 44598 12832 44638 12872
rect 44680 12832 44720 12872
rect 48352 12832 48392 12872
rect 48434 12832 48474 12872
rect 48516 12832 48556 12872
rect 48598 12832 48638 12872
rect 48680 12832 48720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 56352 12832 56392 12872
rect 56434 12832 56474 12872
rect 56516 12832 56556 12872
rect 56598 12832 56638 12872
rect 56680 12832 56720 12872
rect 60352 12832 60392 12872
rect 60434 12832 60474 12872
rect 60516 12832 60556 12872
rect 60598 12832 60638 12872
rect 60680 12832 60720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 68352 12832 68392 12872
rect 68434 12832 68474 12872
rect 68516 12832 68556 12872
rect 68598 12832 68638 12872
rect 68680 12832 68720 12872
rect 844 12412 884 12452
rect 1804 12412 1844 12452
rect 652 12328 692 12368
rect 1612 12244 1652 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 7112 12076 7152 12116
rect 7194 12076 7234 12116
rect 7276 12076 7316 12116
rect 7358 12076 7398 12116
rect 7440 12076 7480 12116
rect 11112 12076 11152 12116
rect 11194 12076 11234 12116
rect 11276 12076 11316 12116
rect 11358 12076 11398 12116
rect 11440 12076 11480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 19112 12076 19152 12116
rect 19194 12076 19234 12116
rect 19276 12076 19316 12116
rect 19358 12076 19398 12116
rect 19440 12076 19480 12116
rect 23112 12076 23152 12116
rect 23194 12076 23234 12116
rect 23276 12076 23316 12116
rect 23358 12076 23398 12116
rect 23440 12076 23480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 31112 12076 31152 12116
rect 31194 12076 31234 12116
rect 31276 12076 31316 12116
rect 31358 12076 31398 12116
rect 31440 12076 31480 12116
rect 35112 12076 35152 12116
rect 35194 12076 35234 12116
rect 35276 12076 35316 12116
rect 35358 12076 35398 12116
rect 35440 12076 35480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 43112 12076 43152 12116
rect 43194 12076 43234 12116
rect 43276 12076 43316 12116
rect 43358 12076 43398 12116
rect 43440 12076 43480 12116
rect 47112 12076 47152 12116
rect 47194 12076 47234 12116
rect 47276 12076 47316 12116
rect 47358 12076 47398 12116
rect 47440 12076 47480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 55112 12076 55152 12116
rect 55194 12076 55234 12116
rect 55276 12076 55316 12116
rect 55358 12076 55398 12116
rect 55440 12076 55480 12116
rect 59112 12076 59152 12116
rect 59194 12076 59234 12116
rect 59276 12076 59316 12116
rect 59358 12076 59398 12116
rect 59440 12076 59480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 67112 12076 67152 12116
rect 67194 12076 67234 12116
rect 67276 12076 67316 12116
rect 67358 12076 67398 12116
rect 67440 12076 67480 12116
rect 1996 11908 2036 11948
rect 844 11740 884 11780
rect 2188 11740 2228 11780
rect 652 11488 692 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 8352 11320 8392 11360
rect 8434 11320 8474 11360
rect 8516 11320 8556 11360
rect 8598 11320 8638 11360
rect 8680 11320 8720 11360
rect 12352 11320 12392 11360
rect 12434 11320 12474 11360
rect 12516 11320 12556 11360
rect 12598 11320 12638 11360
rect 12680 11320 12720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 20352 11320 20392 11360
rect 20434 11320 20474 11360
rect 20516 11320 20556 11360
rect 20598 11320 20638 11360
rect 20680 11320 20720 11360
rect 24352 11320 24392 11360
rect 24434 11320 24474 11360
rect 24516 11320 24556 11360
rect 24598 11320 24638 11360
rect 24680 11320 24720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 32352 11320 32392 11360
rect 32434 11320 32474 11360
rect 32516 11320 32556 11360
rect 32598 11320 32638 11360
rect 32680 11320 32720 11360
rect 36352 11320 36392 11360
rect 36434 11320 36474 11360
rect 36516 11320 36556 11360
rect 36598 11320 36638 11360
rect 36680 11320 36720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 44352 11320 44392 11360
rect 44434 11320 44474 11360
rect 44516 11320 44556 11360
rect 44598 11320 44638 11360
rect 44680 11320 44720 11360
rect 48352 11320 48392 11360
rect 48434 11320 48474 11360
rect 48516 11320 48556 11360
rect 48598 11320 48638 11360
rect 48680 11320 48720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 56352 11320 56392 11360
rect 56434 11320 56474 11360
rect 56516 11320 56556 11360
rect 56598 11320 56638 11360
rect 56680 11320 56720 11360
rect 60352 11320 60392 11360
rect 60434 11320 60474 11360
rect 60516 11320 60556 11360
rect 60598 11320 60638 11360
rect 60680 11320 60720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 68352 11320 68392 11360
rect 68434 11320 68474 11360
rect 68516 11320 68556 11360
rect 68598 11320 68638 11360
rect 68680 11320 68720 11360
rect 69772 10984 69812 11024
rect 844 10900 884 10940
rect 1612 10900 1652 10940
rect 69292 10900 69332 10940
rect 1420 10816 1460 10856
rect 652 10732 692 10772
rect 69484 10732 69524 10772
rect 69868 10732 69908 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 7112 10564 7152 10604
rect 7194 10564 7234 10604
rect 7276 10564 7316 10604
rect 7358 10564 7398 10604
rect 7440 10564 7480 10604
rect 11112 10564 11152 10604
rect 11194 10564 11234 10604
rect 11276 10564 11316 10604
rect 11358 10564 11398 10604
rect 11440 10564 11480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 19112 10564 19152 10604
rect 19194 10564 19234 10604
rect 19276 10564 19316 10604
rect 19358 10564 19398 10604
rect 19440 10564 19480 10604
rect 23112 10564 23152 10604
rect 23194 10564 23234 10604
rect 23276 10564 23316 10604
rect 23358 10564 23398 10604
rect 23440 10564 23480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 31112 10564 31152 10604
rect 31194 10564 31234 10604
rect 31276 10564 31316 10604
rect 31358 10564 31398 10604
rect 31440 10564 31480 10604
rect 35112 10564 35152 10604
rect 35194 10564 35234 10604
rect 35276 10564 35316 10604
rect 35358 10564 35398 10604
rect 35440 10564 35480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 43112 10564 43152 10604
rect 43194 10564 43234 10604
rect 43276 10564 43316 10604
rect 43358 10564 43398 10604
rect 43440 10564 43480 10604
rect 47112 10564 47152 10604
rect 47194 10564 47234 10604
rect 47276 10564 47316 10604
rect 47358 10564 47398 10604
rect 47440 10564 47480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 55112 10564 55152 10604
rect 55194 10564 55234 10604
rect 55276 10564 55316 10604
rect 55358 10564 55398 10604
rect 55440 10564 55480 10604
rect 59112 10564 59152 10604
rect 59194 10564 59234 10604
rect 59276 10564 59316 10604
rect 59358 10564 59398 10604
rect 59440 10564 59480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 67112 10564 67152 10604
rect 67194 10564 67234 10604
rect 67276 10564 67316 10604
rect 67358 10564 67398 10604
rect 67440 10564 67480 10604
rect 1324 10312 1364 10352
rect 67660 10312 67700 10352
rect 69196 10312 69236 10352
rect 844 10228 884 10268
rect 1516 10228 1556 10268
rect 67468 10228 67508 10268
rect 69004 10228 69044 10268
rect 68332 10144 68372 10184
rect 68524 10144 68564 10184
rect 68716 10144 68756 10184
rect 69388 10144 69428 10184
rect 69676 10144 69716 10184
rect 68236 10060 68276 10100
rect 69484 10060 69524 10100
rect 69772 10060 69812 10100
rect 652 9976 692 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 8352 9808 8392 9848
rect 8434 9808 8474 9848
rect 8516 9808 8556 9848
rect 8598 9808 8638 9848
rect 8680 9808 8720 9848
rect 12352 9808 12392 9848
rect 12434 9808 12474 9848
rect 12516 9808 12556 9848
rect 12598 9808 12638 9848
rect 12680 9808 12720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 20352 9808 20392 9848
rect 20434 9808 20474 9848
rect 20516 9808 20556 9848
rect 20598 9808 20638 9848
rect 20680 9808 20720 9848
rect 24352 9808 24392 9848
rect 24434 9808 24474 9848
rect 24516 9808 24556 9848
rect 24598 9808 24638 9848
rect 24680 9808 24720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 32352 9808 32392 9848
rect 32434 9808 32474 9848
rect 32516 9808 32556 9848
rect 32598 9808 32638 9848
rect 32680 9808 32720 9848
rect 36352 9808 36392 9848
rect 36434 9808 36474 9848
rect 36516 9808 36556 9848
rect 36598 9808 36638 9848
rect 36680 9808 36720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 44352 9808 44392 9848
rect 44434 9808 44474 9848
rect 44516 9808 44556 9848
rect 44598 9808 44638 9848
rect 44680 9808 44720 9848
rect 48352 9808 48392 9848
rect 48434 9808 48474 9848
rect 48516 9808 48556 9848
rect 48598 9808 48638 9848
rect 48680 9808 48720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 56352 9808 56392 9848
rect 56434 9808 56474 9848
rect 56516 9808 56556 9848
rect 56598 9808 56638 9848
rect 56680 9808 56720 9848
rect 60352 9808 60392 9848
rect 60434 9808 60474 9848
rect 60516 9808 60556 9848
rect 60598 9808 60638 9848
rect 60680 9808 60720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 68352 9808 68392 9848
rect 68434 9808 68474 9848
rect 68516 9808 68556 9848
rect 68598 9808 68638 9848
rect 68680 9808 68720 9848
rect 69580 9640 69620 9680
rect 69868 9640 69908 9680
rect 69772 9472 69812 9512
rect 844 9388 884 9428
rect 1516 9388 1556 9428
rect 69004 9388 69044 9428
rect 69388 9388 69428 9428
rect 1324 9304 1364 9344
rect 69196 9304 69236 9344
rect 652 9220 692 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 7112 9052 7152 9092
rect 7194 9052 7234 9092
rect 7276 9052 7316 9092
rect 7358 9052 7398 9092
rect 7440 9052 7480 9092
rect 11112 9052 11152 9092
rect 11194 9052 11234 9092
rect 11276 9052 11316 9092
rect 11358 9052 11398 9092
rect 11440 9052 11480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 19112 9052 19152 9092
rect 19194 9052 19234 9092
rect 19276 9052 19316 9092
rect 19358 9052 19398 9092
rect 19440 9052 19480 9092
rect 23112 9052 23152 9092
rect 23194 9052 23234 9092
rect 23276 9052 23316 9092
rect 23358 9052 23398 9092
rect 23440 9052 23480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 31112 9052 31152 9092
rect 31194 9052 31234 9092
rect 31276 9052 31316 9092
rect 31358 9052 31398 9092
rect 31440 9052 31480 9092
rect 35112 9052 35152 9092
rect 35194 9052 35234 9092
rect 35276 9052 35316 9092
rect 35358 9052 35398 9092
rect 35440 9052 35480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 43112 9052 43152 9092
rect 43194 9052 43234 9092
rect 43276 9052 43316 9092
rect 43358 9052 43398 9092
rect 43440 9052 43480 9092
rect 47112 9052 47152 9092
rect 47194 9052 47234 9092
rect 47276 9052 47316 9092
rect 47358 9052 47398 9092
rect 47440 9052 47480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 55112 9052 55152 9092
rect 55194 9052 55234 9092
rect 55276 9052 55316 9092
rect 55358 9052 55398 9092
rect 55440 9052 55480 9092
rect 59112 9052 59152 9092
rect 59194 9052 59234 9092
rect 59276 9052 59316 9092
rect 59358 9052 59398 9092
rect 59440 9052 59480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 67112 9052 67152 9092
rect 67194 9052 67234 9092
rect 67276 9052 67316 9092
rect 67358 9052 67398 9092
rect 67440 9052 67480 9092
rect 1420 8800 1460 8840
rect 844 8716 884 8756
rect 1612 8716 1652 8756
rect 1996 8716 2036 8756
rect 652 8464 692 8504
rect 1804 8464 1844 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 8352 8296 8392 8336
rect 8434 8296 8474 8336
rect 8516 8296 8556 8336
rect 8598 8296 8638 8336
rect 8680 8296 8720 8336
rect 12352 8296 12392 8336
rect 12434 8296 12474 8336
rect 12516 8296 12556 8336
rect 12598 8296 12638 8336
rect 12680 8296 12720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 20352 8296 20392 8336
rect 20434 8296 20474 8336
rect 20516 8296 20556 8336
rect 20598 8296 20638 8336
rect 20680 8296 20720 8336
rect 24352 8296 24392 8336
rect 24434 8296 24474 8336
rect 24516 8296 24556 8336
rect 24598 8296 24638 8336
rect 24680 8296 24720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 32352 8296 32392 8336
rect 32434 8296 32474 8336
rect 32516 8296 32556 8336
rect 32598 8296 32638 8336
rect 32680 8296 32720 8336
rect 36352 8296 36392 8336
rect 36434 8296 36474 8336
rect 36516 8296 36556 8336
rect 36598 8296 36638 8336
rect 36680 8296 36720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 44352 8296 44392 8336
rect 44434 8296 44474 8336
rect 44516 8296 44556 8336
rect 44598 8296 44638 8336
rect 44680 8296 44720 8336
rect 48352 8296 48392 8336
rect 48434 8296 48474 8336
rect 48516 8296 48556 8336
rect 48598 8296 48638 8336
rect 48680 8296 48720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 56352 8296 56392 8336
rect 56434 8296 56474 8336
rect 56516 8296 56556 8336
rect 56598 8296 56638 8336
rect 56680 8296 56720 8336
rect 60352 8296 60392 8336
rect 60434 8296 60474 8336
rect 60516 8296 60556 8336
rect 60598 8296 60638 8336
rect 60680 8296 60720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 68352 8296 68392 8336
rect 68434 8296 68474 8336
rect 68516 8296 68556 8336
rect 68598 8296 68638 8336
rect 68680 8296 68720 8336
rect 844 7876 884 7916
rect 1708 7876 1748 7916
rect 1516 7792 1556 7832
rect 652 7708 692 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 7112 7540 7152 7580
rect 7194 7540 7234 7580
rect 7276 7540 7316 7580
rect 7358 7540 7398 7580
rect 7440 7540 7480 7580
rect 11112 7540 11152 7580
rect 11194 7540 11234 7580
rect 11276 7540 11316 7580
rect 11358 7540 11398 7580
rect 11440 7540 11480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 19112 7540 19152 7580
rect 19194 7540 19234 7580
rect 19276 7540 19316 7580
rect 19358 7540 19398 7580
rect 19440 7540 19480 7580
rect 23112 7540 23152 7580
rect 23194 7540 23234 7580
rect 23276 7540 23316 7580
rect 23358 7540 23398 7580
rect 23440 7540 23480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 31112 7540 31152 7580
rect 31194 7540 31234 7580
rect 31276 7540 31316 7580
rect 31358 7540 31398 7580
rect 31440 7540 31480 7580
rect 35112 7540 35152 7580
rect 35194 7540 35234 7580
rect 35276 7540 35316 7580
rect 35358 7540 35398 7580
rect 35440 7540 35480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 43112 7540 43152 7580
rect 43194 7540 43234 7580
rect 43276 7540 43316 7580
rect 43358 7540 43398 7580
rect 43440 7540 43480 7580
rect 47112 7540 47152 7580
rect 47194 7540 47234 7580
rect 47276 7540 47316 7580
rect 47358 7540 47398 7580
rect 47440 7540 47480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 55112 7540 55152 7580
rect 55194 7540 55234 7580
rect 55276 7540 55316 7580
rect 55358 7540 55398 7580
rect 55440 7540 55480 7580
rect 59112 7540 59152 7580
rect 59194 7540 59234 7580
rect 59276 7540 59316 7580
rect 59358 7540 59398 7580
rect 59440 7540 59480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 67112 7540 67152 7580
rect 67194 7540 67234 7580
rect 67276 7540 67316 7580
rect 67358 7540 67398 7580
rect 67440 7540 67480 7580
rect 71112 7540 71152 7580
rect 71194 7540 71234 7580
rect 71276 7540 71316 7580
rect 71358 7540 71398 7580
rect 71440 7540 71480 7580
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 79112 7540 79152 7580
rect 79194 7540 79234 7580
rect 79276 7540 79316 7580
rect 79358 7540 79398 7580
rect 79440 7540 79480 7580
rect 83112 7540 83152 7580
rect 83194 7540 83234 7580
rect 83276 7540 83316 7580
rect 83358 7540 83398 7580
rect 83440 7540 83480 7580
rect 87112 7540 87152 7580
rect 87194 7540 87234 7580
rect 87276 7540 87316 7580
rect 87358 7540 87398 7580
rect 87440 7540 87480 7580
rect 91112 7540 91152 7580
rect 91194 7540 91234 7580
rect 91276 7540 91316 7580
rect 91358 7540 91398 7580
rect 91440 7540 91480 7580
rect 95112 7540 95152 7580
rect 95194 7540 95234 7580
rect 95276 7540 95316 7580
rect 95358 7540 95398 7580
rect 95440 7540 95480 7580
rect 99112 7540 99152 7580
rect 99194 7540 99234 7580
rect 99276 7540 99316 7580
rect 99358 7540 99398 7580
rect 99440 7540 99480 7580
rect 73420 7372 73460 7412
rect 73804 7372 73844 7412
rect 75244 7372 75284 7412
rect 75916 7372 75956 7412
rect 76300 7372 76340 7412
rect 77068 7372 77108 7412
rect 78028 7372 78068 7412
rect 78316 7372 78356 7412
rect 78796 7372 78836 7412
rect 79180 7372 79220 7412
rect 79468 7372 79508 7412
rect 79852 7372 79892 7412
rect 81484 7372 81524 7412
rect 81676 7372 81716 7412
rect 82348 7372 82388 7412
rect 83404 7372 83444 7412
rect 83884 7372 83924 7412
rect 84652 7372 84692 7412
rect 85036 7372 85076 7412
rect 85708 7372 85748 7412
rect 87148 7372 87188 7412
rect 87724 7372 87764 7412
rect 88780 7372 88820 7412
rect 88972 7372 89012 7412
rect 89644 7372 89684 7412
rect 90412 7372 90452 7412
rect 90604 7372 90644 7412
rect 91852 7372 91892 7412
rect 92908 7372 92948 7412
rect 93292 7372 93332 7412
rect 94732 7372 94772 7412
rect 95116 7372 95156 7412
rect 95884 7372 95924 7412
rect 96844 7372 96884 7412
rect 97132 7372 97172 7412
rect 97420 7372 97460 7412
rect 97996 7372 98036 7412
rect 98476 7372 98516 7412
rect 74476 7288 74516 7328
rect 80044 7288 80084 7328
rect 80716 7288 80756 7328
rect 86284 7288 86324 7328
rect 86476 7288 86516 7328
rect 91180 7288 91220 7328
rect 92332 7288 92372 7328
rect 92524 7288 92564 7328
rect 93964 7288 94004 7328
rect 96652 7288 96692 7328
rect 844 7204 884 7244
rect 73612 7204 73652 7244
rect 74284 7204 74324 7244
rect 74668 7204 74708 7244
rect 75052 7204 75092 7244
rect 75436 7204 75476 7244
rect 75724 7204 75764 7244
rect 76108 7204 76148 7244
rect 76876 7204 76916 7244
rect 77452 7204 77492 7244
rect 77836 7204 77876 7244
rect 79660 7204 79700 7244
rect 80236 7204 80276 7244
rect 80524 7204 80564 7244
rect 81100 7204 81140 7244
rect 81292 7204 81332 7244
rect 82828 7204 82868 7244
rect 83020 7204 83060 7244
rect 84268 7204 84308 7244
rect 84844 7204 84884 7244
rect 85228 7204 85268 7244
rect 86092 7204 86132 7244
rect 86668 7204 86708 7244
rect 88012 7204 88052 7244
rect 88588 7204 88628 7244
rect 89452 7204 89492 7244
rect 90028 7204 90068 7244
rect 90988 7204 91028 7244
rect 91372 7204 91412 7244
rect 92140 7204 92180 7244
rect 92716 7204 92756 7244
rect 93100 7204 93140 7244
rect 94156 7204 94196 7244
rect 94348 7204 94388 7244
rect 94924 7204 94964 7244
rect 95308 7204 95348 7244
rect 95692 7204 95732 7244
rect 96268 7204 96308 7244
rect 96460 7204 96500 7244
rect 97612 7204 97652 7244
rect 98188 7204 98228 7244
rect 98668 7204 98708 7244
rect 73324 7120 73364 7160
rect 76684 7120 76724 7160
rect 78124 7120 78164 7160
rect 78412 7120 78452 7160
rect 78700 7109 78740 7149
rect 79084 7120 79124 7160
rect 79372 7120 79412 7160
rect 81772 7120 81812 7160
rect 81964 7109 82004 7149
rect 82060 7120 82100 7160
rect 82252 7120 82292 7160
rect 83116 7120 83156 7160
rect 83308 7120 83348 7160
rect 83788 7120 83828 7160
rect 84556 7120 84596 7160
rect 85612 7120 85652 7160
rect 86860 7120 86900 7160
rect 87244 7120 87284 7160
rect 87436 7120 87476 7160
rect 87532 7120 87572 7160
rect 87820 7120 87860 7160
rect 89068 7120 89108 7160
rect 90316 7120 90356 7160
rect 90713 7120 90753 7160
rect 91756 7120 91796 7160
rect 93388 7120 93428 7160
rect 93676 7120 93716 7160
rect 96940 7120 96980 7160
rect 97228 7120 97268 7160
rect 76588 7036 76628 7076
rect 652 6952 692 6992
rect 74092 6952 74132 6992
rect 74860 6952 74900 6992
rect 77260 6952 77300 6992
rect 77644 6952 77684 6992
rect 80908 6952 80948 6992
rect 82636 6952 82676 6992
rect 84076 6952 84116 6992
rect 85420 6952 85460 6992
rect 86956 6952 86996 6992
rect 88204 6952 88244 6992
rect 89836 6952 89876 6992
rect 91564 6952 91604 6992
rect 93772 6952 93812 6992
rect 94540 6952 94580 6992
rect 96076 6952 96116 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 8352 6784 8392 6824
rect 8434 6784 8474 6824
rect 8516 6784 8556 6824
rect 8598 6784 8638 6824
rect 8680 6784 8720 6824
rect 12352 6784 12392 6824
rect 12434 6784 12474 6824
rect 12516 6784 12556 6824
rect 12598 6784 12638 6824
rect 12680 6784 12720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 20352 6784 20392 6824
rect 20434 6784 20474 6824
rect 20516 6784 20556 6824
rect 20598 6784 20638 6824
rect 20680 6784 20720 6824
rect 24352 6784 24392 6824
rect 24434 6784 24474 6824
rect 24516 6784 24556 6824
rect 24598 6784 24638 6824
rect 24680 6784 24720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 32352 6784 32392 6824
rect 32434 6784 32474 6824
rect 32516 6784 32556 6824
rect 32598 6784 32638 6824
rect 32680 6784 32720 6824
rect 36352 6784 36392 6824
rect 36434 6784 36474 6824
rect 36516 6784 36556 6824
rect 36598 6784 36638 6824
rect 36680 6784 36720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 44352 6784 44392 6824
rect 44434 6784 44474 6824
rect 44516 6784 44556 6824
rect 44598 6784 44638 6824
rect 44680 6784 44720 6824
rect 48352 6784 48392 6824
rect 48434 6784 48474 6824
rect 48516 6784 48556 6824
rect 48598 6784 48638 6824
rect 48680 6784 48720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 56352 6784 56392 6824
rect 56434 6784 56474 6824
rect 56516 6784 56556 6824
rect 56598 6784 56638 6824
rect 56680 6784 56720 6824
rect 60352 6784 60392 6824
rect 60434 6784 60474 6824
rect 60516 6784 60556 6824
rect 60598 6784 60638 6824
rect 60680 6784 60720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 68352 6784 68392 6824
rect 68434 6784 68474 6824
rect 68516 6784 68556 6824
rect 68598 6784 68638 6824
rect 68680 6784 68720 6824
rect 72352 6784 72392 6824
rect 72434 6784 72474 6824
rect 72516 6784 72556 6824
rect 72598 6784 72638 6824
rect 72680 6784 72720 6824
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 80352 6784 80392 6824
rect 80434 6784 80474 6824
rect 80516 6784 80556 6824
rect 80598 6784 80638 6824
rect 80680 6784 80720 6824
rect 84352 6784 84392 6824
rect 84434 6784 84474 6824
rect 84516 6784 84556 6824
rect 84598 6784 84638 6824
rect 84680 6784 84720 6824
rect 88352 6784 88392 6824
rect 88434 6784 88474 6824
rect 88516 6784 88556 6824
rect 88598 6784 88638 6824
rect 88680 6784 88720 6824
rect 92352 6784 92392 6824
rect 92434 6784 92474 6824
rect 92516 6784 92556 6824
rect 92598 6784 92638 6824
rect 92680 6784 92720 6824
rect 96352 6784 96392 6824
rect 96434 6784 96474 6824
rect 96516 6784 96556 6824
rect 96598 6784 96638 6824
rect 96680 6784 96720 6824
rect 1324 6616 1364 6656
rect 74188 6616 74228 6656
rect 75244 6616 75284 6656
rect 75532 6616 75572 6656
rect 75820 6616 75860 6656
rect 76396 6616 76436 6656
rect 76780 6616 76820 6656
rect 77164 6616 77204 6656
rect 77932 6616 77972 6656
rect 78316 6616 78356 6656
rect 79084 6616 79124 6656
rect 80044 6616 80084 6656
rect 80620 6616 80660 6656
rect 81100 6616 81140 6656
rect 81484 6616 81524 6656
rect 81868 6616 81908 6656
rect 82252 6616 82292 6656
rect 82924 6616 82964 6656
rect 83404 6616 83444 6656
rect 83884 6616 83924 6656
rect 84364 6616 84404 6656
rect 84748 6616 84788 6656
rect 84940 6616 84980 6656
rect 85420 6616 85460 6656
rect 85804 6616 85844 6656
rect 86284 6616 86324 6656
rect 87052 6616 87092 6656
rect 87532 6616 87572 6656
rect 87916 6616 87956 6656
rect 88300 6616 88340 6656
rect 88492 6616 88532 6656
rect 89260 6616 89300 6656
rect 90604 6616 90644 6656
rect 91084 6616 91124 6656
rect 91276 6616 91316 6656
rect 91852 6616 91892 6656
rect 92332 6616 92372 6656
rect 92620 6616 92660 6656
rect 93196 6616 93236 6656
rect 93580 6616 93620 6656
rect 94060 6616 94100 6656
rect 94252 6616 94292 6656
rect 94828 6616 94868 6656
rect 95308 6616 95348 6656
rect 95596 6616 95636 6656
rect 96556 6616 96596 6656
rect 97132 6616 97172 6656
rect 97420 6616 97460 6656
rect 97708 6616 97748 6656
rect 98092 6616 98132 6656
rect 74092 6448 74132 6488
rect 75145 6435 75185 6475
rect 75436 6448 75476 6488
rect 75724 6448 75764 6488
rect 76300 6448 76340 6488
rect 76684 6448 76724 6488
rect 79948 6448 79988 6488
rect 81388 6448 81428 6488
rect 85036 6448 85076 6488
rect 88588 6448 88628 6488
rect 88780 6448 88820 6488
rect 88876 6448 88916 6488
rect 89164 6448 89204 6488
rect 91372 6448 91412 6488
rect 92524 6448 92564 6488
rect 94732 6448 94772 6488
rect 95692 6448 95732 6488
rect 95884 6448 95924 6488
rect 97324 6448 97364 6488
rect 97804 6448 97844 6488
rect 97996 6448 98036 6488
rect 1516 6364 1556 6404
rect 74380 6364 74420 6404
rect 74764 6364 74804 6404
rect 76972 6364 77012 6404
rect 77740 6364 77780 6404
rect 78124 6364 78164 6404
rect 78892 6364 78932 6404
rect 79564 6364 79604 6404
rect 80428 6364 80468 6404
rect 80908 6364 80948 6404
rect 81676 6364 81716 6404
rect 82060 6364 82100 6404
rect 82732 6364 82772 6404
rect 83212 6364 83252 6404
rect 83692 6364 83732 6404
rect 84172 6364 84212 6404
rect 84556 6364 84596 6404
rect 85228 6364 85268 6404
rect 85612 6364 85652 6404
rect 86092 6364 86132 6404
rect 86860 6364 86900 6404
rect 87340 6364 87380 6404
rect 87724 6364 87764 6404
rect 88108 6364 88148 6404
rect 89644 6364 89684 6404
rect 90412 6364 90452 6404
rect 90892 6364 90932 6404
rect 91660 6364 91700 6404
rect 92140 6364 92180 6404
rect 93004 6364 93044 6404
rect 93388 6364 93428 6404
rect 93868 6364 93908 6404
rect 94444 6364 94484 6404
rect 95116 6364 95156 6404
rect 96364 6364 96404 6404
rect 96940 6364 96980 6404
rect 74956 6280 74996 6320
rect 79372 6280 79412 6320
rect 89452 6280 89492 6320
rect 74572 6196 74612 6236
rect 95980 6196 96020 6236
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 7112 6028 7152 6068
rect 7194 6028 7234 6068
rect 7276 6028 7316 6068
rect 7358 6028 7398 6068
rect 7440 6028 7480 6068
rect 11112 6028 11152 6068
rect 11194 6028 11234 6068
rect 11276 6028 11316 6068
rect 11358 6028 11398 6068
rect 11440 6028 11480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 19112 6028 19152 6068
rect 19194 6028 19234 6068
rect 19276 6028 19316 6068
rect 19358 6028 19398 6068
rect 19440 6028 19480 6068
rect 23112 6028 23152 6068
rect 23194 6028 23234 6068
rect 23276 6028 23316 6068
rect 23358 6028 23398 6068
rect 23440 6028 23480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 31112 6028 31152 6068
rect 31194 6028 31234 6068
rect 31276 6028 31316 6068
rect 31358 6028 31398 6068
rect 31440 6028 31480 6068
rect 35112 6028 35152 6068
rect 35194 6028 35234 6068
rect 35276 6028 35316 6068
rect 35358 6028 35398 6068
rect 35440 6028 35480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 43112 6028 43152 6068
rect 43194 6028 43234 6068
rect 43276 6028 43316 6068
rect 43358 6028 43398 6068
rect 43440 6028 43480 6068
rect 47112 6028 47152 6068
rect 47194 6028 47234 6068
rect 47276 6028 47316 6068
rect 47358 6028 47398 6068
rect 47440 6028 47480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 55112 6028 55152 6068
rect 55194 6028 55234 6068
rect 55276 6028 55316 6068
rect 55358 6028 55398 6068
rect 55440 6028 55480 6068
rect 59112 6028 59152 6068
rect 59194 6028 59234 6068
rect 59276 6028 59316 6068
rect 59358 6028 59398 6068
rect 59440 6028 59480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 67112 6028 67152 6068
rect 67194 6028 67234 6068
rect 67276 6028 67316 6068
rect 67358 6028 67398 6068
rect 67440 6028 67480 6068
rect 71112 6028 71152 6068
rect 71194 6028 71234 6068
rect 71276 6028 71316 6068
rect 71358 6028 71398 6068
rect 71440 6028 71480 6068
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 79112 6028 79152 6068
rect 79194 6028 79234 6068
rect 79276 6028 79316 6068
rect 79358 6028 79398 6068
rect 79440 6028 79480 6068
rect 83112 6028 83152 6068
rect 83194 6028 83234 6068
rect 83276 6028 83316 6068
rect 83358 6028 83398 6068
rect 83440 6028 83480 6068
rect 87112 6028 87152 6068
rect 87194 6028 87234 6068
rect 87276 6028 87316 6068
rect 87358 6028 87398 6068
rect 87440 6028 87480 6068
rect 91112 6028 91152 6068
rect 91194 6028 91234 6068
rect 91276 6028 91316 6068
rect 91358 6028 91398 6068
rect 91440 6028 91480 6068
rect 95112 6028 95152 6068
rect 95194 6028 95234 6068
rect 95276 6028 95316 6068
rect 95358 6028 95398 6068
rect 95440 6028 95480 6068
rect 99112 6028 99152 6068
rect 99194 6028 99234 6068
rect 99276 6028 99316 6068
rect 99358 6028 99398 6068
rect 99440 6028 99480 6068
rect 75340 5860 75380 5900
rect 76684 5860 76724 5900
rect 78316 5860 78356 5900
rect 78796 5860 78836 5900
rect 80140 5860 80180 5900
rect 80332 5860 80372 5900
rect 81196 5860 81236 5900
rect 82636 5860 82676 5900
rect 83596 5860 83636 5900
rect 85516 5860 85556 5900
rect 86764 5860 86804 5900
rect 87628 5860 87668 5900
rect 89068 5860 89108 5900
rect 89644 5860 89684 5900
rect 90220 5860 90260 5900
rect 91660 5860 91700 5900
rect 92812 5860 92852 5900
rect 93196 5860 93236 5900
rect 93580 5860 93620 5900
rect 93964 5860 94004 5900
rect 95692 5860 95732 5900
rect 95980 5860 96020 5900
rect 98764 5860 98804 5900
rect 1804 5776 1844 5816
rect 844 5692 884 5732
rect 1612 5692 1652 5732
rect 1996 5692 2036 5732
rect 75148 5692 75188 5732
rect 76492 5692 76532 5732
rect 78604 5692 78644 5732
rect 79948 5692 79988 5732
rect 82444 5692 82484 5732
rect 86572 5692 86612 5732
rect 88876 5692 88916 5732
rect 90412 5692 90452 5732
rect 95500 5692 95540 5732
rect 78220 5608 78260 5648
rect 80428 5608 80468 5648
rect 81100 5608 81140 5648
rect 83500 5608 83540 5648
rect 85420 5608 85460 5648
rect 87532 5608 87572 5648
rect 89548 5608 89588 5648
rect 91564 5608 91604 5648
rect 92908 5608 92948 5648
rect 93292 5608 93332 5648
rect 93676 5608 93716 5648
rect 93868 5608 93908 5648
rect 95884 5608 95924 5648
rect 98380 5608 98420 5648
rect 98668 5608 98708 5648
rect 652 5440 692 5480
rect 1420 5440 1460 5480
rect 98284 5440 98324 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 8352 5272 8392 5312
rect 8434 5272 8474 5312
rect 8516 5272 8556 5312
rect 8598 5272 8638 5312
rect 8680 5272 8720 5312
rect 12352 5272 12392 5312
rect 12434 5272 12474 5312
rect 12516 5272 12556 5312
rect 12598 5272 12638 5312
rect 12680 5272 12720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 20352 5272 20392 5312
rect 20434 5272 20474 5312
rect 20516 5272 20556 5312
rect 20598 5272 20638 5312
rect 20680 5272 20720 5312
rect 24352 5272 24392 5312
rect 24434 5272 24474 5312
rect 24516 5272 24556 5312
rect 24598 5272 24638 5312
rect 24680 5272 24720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 32352 5272 32392 5312
rect 32434 5272 32474 5312
rect 32516 5272 32556 5312
rect 32598 5272 32638 5312
rect 32680 5272 32720 5312
rect 36352 5272 36392 5312
rect 36434 5272 36474 5312
rect 36516 5272 36556 5312
rect 36598 5272 36638 5312
rect 36680 5272 36720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 44352 5272 44392 5312
rect 44434 5272 44474 5312
rect 44516 5272 44556 5312
rect 44598 5272 44638 5312
rect 44680 5272 44720 5312
rect 48352 5272 48392 5312
rect 48434 5272 48474 5312
rect 48516 5272 48556 5312
rect 48598 5272 48638 5312
rect 48680 5272 48720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 56352 5272 56392 5312
rect 56434 5272 56474 5312
rect 56516 5272 56556 5312
rect 56598 5272 56638 5312
rect 56680 5272 56720 5312
rect 60352 5272 60392 5312
rect 60434 5272 60474 5312
rect 60516 5272 60556 5312
rect 60598 5272 60638 5312
rect 60680 5272 60720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 68352 5272 68392 5312
rect 68434 5272 68474 5312
rect 68516 5272 68556 5312
rect 68598 5272 68638 5312
rect 68680 5272 68720 5312
rect 72352 5272 72392 5312
rect 72434 5272 72474 5312
rect 72516 5272 72556 5312
rect 72598 5272 72638 5312
rect 72680 5272 72720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 80352 5272 80392 5312
rect 80434 5272 80474 5312
rect 80516 5272 80556 5312
rect 80598 5272 80638 5312
rect 80680 5272 80720 5312
rect 84352 5272 84392 5312
rect 84434 5272 84474 5312
rect 84516 5272 84556 5312
rect 84598 5272 84638 5312
rect 84680 5272 84720 5312
rect 88352 5272 88392 5312
rect 88434 5272 88474 5312
rect 88516 5272 88556 5312
rect 88598 5272 88638 5312
rect 88680 5272 88720 5312
rect 92352 5272 92392 5312
rect 92434 5272 92474 5312
rect 92516 5272 92556 5312
rect 92598 5272 92638 5312
rect 92680 5272 92720 5312
rect 96352 5272 96392 5312
rect 96434 5272 96474 5312
rect 96516 5272 96556 5312
rect 96598 5272 96638 5312
rect 96680 5272 96720 5312
rect 844 4852 884 4892
rect 1420 4852 1460 4892
rect 1804 4852 1844 4892
rect 2188 4852 2228 4892
rect 96940 4852 96980 4892
rect 652 4768 692 4808
rect 97132 4768 97172 4808
rect 1228 4684 1268 4724
rect 1612 4684 1652 4724
rect 1996 4684 2036 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 7112 4516 7152 4556
rect 7194 4516 7234 4556
rect 7276 4516 7316 4556
rect 7358 4516 7398 4556
rect 7440 4516 7480 4556
rect 11112 4516 11152 4556
rect 11194 4516 11234 4556
rect 11276 4516 11316 4556
rect 11358 4516 11398 4556
rect 11440 4516 11480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 19112 4516 19152 4556
rect 19194 4516 19234 4556
rect 19276 4516 19316 4556
rect 19358 4516 19398 4556
rect 19440 4516 19480 4556
rect 23112 4516 23152 4556
rect 23194 4516 23234 4556
rect 23276 4516 23316 4556
rect 23358 4516 23398 4556
rect 23440 4516 23480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 31112 4516 31152 4556
rect 31194 4516 31234 4556
rect 31276 4516 31316 4556
rect 31358 4516 31398 4556
rect 31440 4516 31480 4556
rect 35112 4516 35152 4556
rect 35194 4516 35234 4556
rect 35276 4516 35316 4556
rect 35358 4516 35398 4556
rect 35440 4516 35480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 43112 4516 43152 4556
rect 43194 4516 43234 4556
rect 43276 4516 43316 4556
rect 43358 4516 43398 4556
rect 43440 4516 43480 4556
rect 47112 4516 47152 4556
rect 47194 4516 47234 4556
rect 47276 4516 47316 4556
rect 47358 4516 47398 4556
rect 47440 4516 47480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 55112 4516 55152 4556
rect 55194 4516 55234 4556
rect 55276 4516 55316 4556
rect 55358 4516 55398 4556
rect 55440 4516 55480 4556
rect 59112 4516 59152 4556
rect 59194 4516 59234 4556
rect 59276 4516 59316 4556
rect 59358 4516 59398 4556
rect 59440 4516 59480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 67112 4516 67152 4556
rect 67194 4516 67234 4556
rect 67276 4516 67316 4556
rect 67358 4516 67398 4556
rect 67440 4516 67480 4556
rect 71112 4516 71152 4556
rect 71194 4516 71234 4556
rect 71276 4516 71316 4556
rect 71358 4516 71398 4556
rect 71440 4516 71480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 79112 4516 79152 4556
rect 79194 4516 79234 4556
rect 79276 4516 79316 4556
rect 79358 4516 79398 4556
rect 79440 4516 79480 4556
rect 83112 4516 83152 4556
rect 83194 4516 83234 4556
rect 83276 4516 83316 4556
rect 83358 4516 83398 4556
rect 83440 4516 83480 4556
rect 87112 4516 87152 4556
rect 87194 4516 87234 4556
rect 87276 4516 87316 4556
rect 87358 4516 87398 4556
rect 87440 4516 87480 4556
rect 91112 4516 91152 4556
rect 91194 4516 91234 4556
rect 91276 4516 91316 4556
rect 91358 4516 91398 4556
rect 91440 4516 91480 4556
rect 95112 4516 95152 4556
rect 95194 4516 95234 4556
rect 95276 4516 95316 4556
rect 95358 4516 95398 4556
rect 95440 4516 95480 4556
rect 99112 4516 99152 4556
rect 99194 4516 99234 4556
rect 99276 4516 99316 4556
rect 99358 4516 99398 4556
rect 99440 4516 99480 4556
rect 844 4180 884 4220
rect 652 3928 692 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 8352 3760 8392 3800
rect 8434 3760 8474 3800
rect 8516 3760 8556 3800
rect 8598 3760 8638 3800
rect 8680 3760 8720 3800
rect 12352 3760 12392 3800
rect 12434 3760 12474 3800
rect 12516 3760 12556 3800
rect 12598 3760 12638 3800
rect 12680 3760 12720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 20352 3760 20392 3800
rect 20434 3760 20474 3800
rect 20516 3760 20556 3800
rect 20598 3760 20638 3800
rect 20680 3760 20720 3800
rect 24352 3760 24392 3800
rect 24434 3760 24474 3800
rect 24516 3760 24556 3800
rect 24598 3760 24638 3800
rect 24680 3760 24720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 32352 3760 32392 3800
rect 32434 3760 32474 3800
rect 32516 3760 32556 3800
rect 32598 3760 32638 3800
rect 32680 3760 32720 3800
rect 36352 3760 36392 3800
rect 36434 3760 36474 3800
rect 36516 3760 36556 3800
rect 36598 3760 36638 3800
rect 36680 3760 36720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 44352 3760 44392 3800
rect 44434 3760 44474 3800
rect 44516 3760 44556 3800
rect 44598 3760 44638 3800
rect 44680 3760 44720 3800
rect 48352 3760 48392 3800
rect 48434 3760 48474 3800
rect 48516 3760 48556 3800
rect 48598 3760 48638 3800
rect 48680 3760 48720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 56352 3760 56392 3800
rect 56434 3760 56474 3800
rect 56516 3760 56556 3800
rect 56598 3760 56638 3800
rect 56680 3760 56720 3800
rect 60352 3760 60392 3800
rect 60434 3760 60474 3800
rect 60516 3760 60556 3800
rect 60598 3760 60638 3800
rect 60680 3760 60720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 68352 3760 68392 3800
rect 68434 3760 68474 3800
rect 68516 3760 68556 3800
rect 68598 3760 68638 3800
rect 68680 3760 68720 3800
rect 72352 3760 72392 3800
rect 72434 3760 72474 3800
rect 72516 3760 72556 3800
rect 72598 3760 72638 3800
rect 72680 3760 72720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 80352 3760 80392 3800
rect 80434 3760 80474 3800
rect 80516 3760 80556 3800
rect 80598 3760 80638 3800
rect 80680 3760 80720 3800
rect 84352 3760 84392 3800
rect 84434 3760 84474 3800
rect 84516 3760 84556 3800
rect 84598 3760 84638 3800
rect 84680 3760 84720 3800
rect 88352 3760 88392 3800
rect 88434 3760 88474 3800
rect 88516 3760 88556 3800
rect 88598 3760 88638 3800
rect 88680 3760 88720 3800
rect 92352 3760 92392 3800
rect 92434 3760 92474 3800
rect 92516 3760 92556 3800
rect 92598 3760 92638 3800
rect 92680 3760 92720 3800
rect 96352 3760 96392 3800
rect 96434 3760 96474 3800
rect 96516 3760 96556 3800
rect 96598 3760 96638 3800
rect 96680 3760 96720 3800
rect 844 3340 884 3380
rect 652 3172 692 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 7112 3004 7152 3044
rect 7194 3004 7234 3044
rect 7276 3004 7316 3044
rect 7358 3004 7398 3044
rect 7440 3004 7480 3044
rect 11112 3004 11152 3044
rect 11194 3004 11234 3044
rect 11276 3004 11316 3044
rect 11358 3004 11398 3044
rect 11440 3004 11480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 19112 3004 19152 3044
rect 19194 3004 19234 3044
rect 19276 3004 19316 3044
rect 19358 3004 19398 3044
rect 19440 3004 19480 3044
rect 23112 3004 23152 3044
rect 23194 3004 23234 3044
rect 23276 3004 23316 3044
rect 23358 3004 23398 3044
rect 23440 3004 23480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 31112 3004 31152 3044
rect 31194 3004 31234 3044
rect 31276 3004 31316 3044
rect 31358 3004 31398 3044
rect 31440 3004 31480 3044
rect 35112 3004 35152 3044
rect 35194 3004 35234 3044
rect 35276 3004 35316 3044
rect 35358 3004 35398 3044
rect 35440 3004 35480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 43112 3004 43152 3044
rect 43194 3004 43234 3044
rect 43276 3004 43316 3044
rect 43358 3004 43398 3044
rect 43440 3004 43480 3044
rect 47112 3004 47152 3044
rect 47194 3004 47234 3044
rect 47276 3004 47316 3044
rect 47358 3004 47398 3044
rect 47440 3004 47480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 55112 3004 55152 3044
rect 55194 3004 55234 3044
rect 55276 3004 55316 3044
rect 55358 3004 55398 3044
rect 55440 3004 55480 3044
rect 59112 3004 59152 3044
rect 59194 3004 59234 3044
rect 59276 3004 59316 3044
rect 59358 3004 59398 3044
rect 59440 3004 59480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 67112 3004 67152 3044
rect 67194 3004 67234 3044
rect 67276 3004 67316 3044
rect 67358 3004 67398 3044
rect 67440 3004 67480 3044
rect 71112 3004 71152 3044
rect 71194 3004 71234 3044
rect 71276 3004 71316 3044
rect 71358 3004 71398 3044
rect 71440 3004 71480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 79112 3004 79152 3044
rect 79194 3004 79234 3044
rect 79276 3004 79316 3044
rect 79358 3004 79398 3044
rect 79440 3004 79480 3044
rect 83112 3004 83152 3044
rect 83194 3004 83234 3044
rect 83276 3004 83316 3044
rect 83358 3004 83398 3044
rect 83440 3004 83480 3044
rect 87112 3004 87152 3044
rect 87194 3004 87234 3044
rect 87276 3004 87316 3044
rect 87358 3004 87398 3044
rect 87440 3004 87480 3044
rect 91112 3004 91152 3044
rect 91194 3004 91234 3044
rect 91276 3004 91316 3044
rect 91358 3004 91398 3044
rect 91440 3004 91480 3044
rect 95112 3004 95152 3044
rect 95194 3004 95234 3044
rect 95276 3004 95316 3044
rect 95358 3004 95398 3044
rect 95440 3004 95480 3044
rect 99112 3004 99152 3044
rect 99194 3004 99234 3044
rect 99276 3004 99316 3044
rect 99358 3004 99398 3044
rect 99440 3004 99480 3044
rect 844 2668 884 2708
rect 652 2416 692 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 8352 2248 8392 2288
rect 8434 2248 8474 2288
rect 8516 2248 8556 2288
rect 8598 2248 8638 2288
rect 8680 2248 8720 2288
rect 12352 2248 12392 2288
rect 12434 2248 12474 2288
rect 12516 2248 12556 2288
rect 12598 2248 12638 2288
rect 12680 2248 12720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 20352 2248 20392 2288
rect 20434 2248 20474 2288
rect 20516 2248 20556 2288
rect 20598 2248 20638 2288
rect 20680 2248 20720 2288
rect 24352 2248 24392 2288
rect 24434 2248 24474 2288
rect 24516 2248 24556 2288
rect 24598 2248 24638 2288
rect 24680 2248 24720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 32352 2248 32392 2288
rect 32434 2248 32474 2288
rect 32516 2248 32556 2288
rect 32598 2248 32638 2288
rect 32680 2248 32720 2288
rect 36352 2248 36392 2288
rect 36434 2248 36474 2288
rect 36516 2248 36556 2288
rect 36598 2248 36638 2288
rect 36680 2248 36720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 44352 2248 44392 2288
rect 44434 2248 44474 2288
rect 44516 2248 44556 2288
rect 44598 2248 44638 2288
rect 44680 2248 44720 2288
rect 48352 2248 48392 2288
rect 48434 2248 48474 2288
rect 48516 2248 48556 2288
rect 48598 2248 48638 2288
rect 48680 2248 48720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 56352 2248 56392 2288
rect 56434 2248 56474 2288
rect 56516 2248 56556 2288
rect 56598 2248 56638 2288
rect 56680 2248 56720 2288
rect 60352 2248 60392 2288
rect 60434 2248 60474 2288
rect 60516 2248 60556 2288
rect 60598 2248 60638 2288
rect 60680 2248 60720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 68352 2248 68392 2288
rect 68434 2248 68474 2288
rect 68516 2248 68556 2288
rect 68598 2248 68638 2288
rect 68680 2248 68720 2288
rect 72352 2248 72392 2288
rect 72434 2248 72474 2288
rect 72516 2248 72556 2288
rect 72598 2248 72638 2288
rect 72680 2248 72720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 80352 2248 80392 2288
rect 80434 2248 80474 2288
rect 80516 2248 80556 2288
rect 80598 2248 80638 2288
rect 80680 2248 80720 2288
rect 84352 2248 84392 2288
rect 84434 2248 84474 2288
rect 84516 2248 84556 2288
rect 84598 2248 84638 2288
rect 84680 2248 84720 2288
rect 88352 2248 88392 2288
rect 88434 2248 88474 2288
rect 88516 2248 88556 2288
rect 88598 2248 88638 2288
rect 88680 2248 88720 2288
rect 92352 2248 92392 2288
rect 92434 2248 92474 2288
rect 92516 2248 92556 2288
rect 92598 2248 92638 2288
rect 92680 2248 92720 2288
rect 96352 2248 96392 2288
rect 96434 2248 96474 2288
rect 96516 2248 96556 2288
rect 96598 2248 96638 2288
rect 96680 2248 96720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 7112 1492 7152 1532
rect 7194 1492 7234 1532
rect 7276 1492 7316 1532
rect 7358 1492 7398 1532
rect 7440 1492 7480 1532
rect 11112 1492 11152 1532
rect 11194 1492 11234 1532
rect 11276 1492 11316 1532
rect 11358 1492 11398 1532
rect 11440 1492 11480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 19112 1492 19152 1532
rect 19194 1492 19234 1532
rect 19276 1492 19316 1532
rect 19358 1492 19398 1532
rect 19440 1492 19480 1532
rect 23112 1492 23152 1532
rect 23194 1492 23234 1532
rect 23276 1492 23316 1532
rect 23358 1492 23398 1532
rect 23440 1492 23480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 31112 1492 31152 1532
rect 31194 1492 31234 1532
rect 31276 1492 31316 1532
rect 31358 1492 31398 1532
rect 31440 1492 31480 1532
rect 35112 1492 35152 1532
rect 35194 1492 35234 1532
rect 35276 1492 35316 1532
rect 35358 1492 35398 1532
rect 35440 1492 35480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 43112 1492 43152 1532
rect 43194 1492 43234 1532
rect 43276 1492 43316 1532
rect 43358 1492 43398 1532
rect 43440 1492 43480 1532
rect 47112 1492 47152 1532
rect 47194 1492 47234 1532
rect 47276 1492 47316 1532
rect 47358 1492 47398 1532
rect 47440 1492 47480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 55112 1492 55152 1532
rect 55194 1492 55234 1532
rect 55276 1492 55316 1532
rect 55358 1492 55398 1532
rect 55440 1492 55480 1532
rect 59112 1492 59152 1532
rect 59194 1492 59234 1532
rect 59276 1492 59316 1532
rect 59358 1492 59398 1532
rect 59440 1492 59480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 67112 1492 67152 1532
rect 67194 1492 67234 1532
rect 67276 1492 67316 1532
rect 67358 1492 67398 1532
rect 67440 1492 67480 1532
rect 71112 1492 71152 1532
rect 71194 1492 71234 1532
rect 71276 1492 71316 1532
rect 71358 1492 71398 1532
rect 71440 1492 71480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 79112 1492 79152 1532
rect 79194 1492 79234 1532
rect 79276 1492 79316 1532
rect 79358 1492 79398 1532
rect 79440 1492 79480 1532
rect 83112 1492 83152 1532
rect 83194 1492 83234 1532
rect 83276 1492 83316 1532
rect 83358 1492 83398 1532
rect 83440 1492 83480 1532
rect 87112 1492 87152 1532
rect 87194 1492 87234 1532
rect 87276 1492 87316 1532
rect 87358 1492 87398 1532
rect 87440 1492 87480 1532
rect 91112 1492 91152 1532
rect 91194 1492 91234 1532
rect 91276 1492 91316 1532
rect 91358 1492 91398 1532
rect 91440 1492 91480 1532
rect 95112 1492 95152 1532
rect 95194 1492 95234 1532
rect 95276 1492 95316 1532
rect 95358 1492 95398 1532
rect 95440 1492 95480 1532
rect 99112 1492 99152 1532
rect 99194 1492 99234 1532
rect 99276 1492 99316 1532
rect 99358 1492 99398 1532
rect 99440 1492 99480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 8352 736 8392 776
rect 8434 736 8474 776
rect 8516 736 8556 776
rect 8598 736 8638 776
rect 8680 736 8720 776
rect 12352 736 12392 776
rect 12434 736 12474 776
rect 12516 736 12556 776
rect 12598 736 12638 776
rect 12680 736 12720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 20352 736 20392 776
rect 20434 736 20474 776
rect 20516 736 20556 776
rect 20598 736 20638 776
rect 20680 736 20720 776
rect 24352 736 24392 776
rect 24434 736 24474 776
rect 24516 736 24556 776
rect 24598 736 24638 776
rect 24680 736 24720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 32352 736 32392 776
rect 32434 736 32474 776
rect 32516 736 32556 776
rect 32598 736 32638 776
rect 32680 736 32720 776
rect 36352 736 36392 776
rect 36434 736 36474 776
rect 36516 736 36556 776
rect 36598 736 36638 776
rect 36680 736 36720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 44352 736 44392 776
rect 44434 736 44474 776
rect 44516 736 44556 776
rect 44598 736 44638 776
rect 44680 736 44720 776
rect 48352 736 48392 776
rect 48434 736 48474 776
rect 48516 736 48556 776
rect 48598 736 48638 776
rect 48680 736 48720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 56352 736 56392 776
rect 56434 736 56474 776
rect 56516 736 56556 776
rect 56598 736 56638 776
rect 56680 736 56720 776
rect 60352 736 60392 776
rect 60434 736 60474 776
rect 60516 736 60556 776
rect 60598 736 60638 776
rect 60680 736 60720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 68352 736 68392 776
rect 68434 736 68474 776
rect 68516 736 68556 776
rect 68598 736 68638 776
rect 68680 736 68720 776
rect 72352 736 72392 776
rect 72434 736 72474 776
rect 72516 736 72556 776
rect 72598 736 72638 776
rect 72680 736 72720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
rect 80352 736 80392 776
rect 80434 736 80474 776
rect 80516 736 80556 776
rect 80598 736 80638 776
rect 80680 736 80720 776
rect 84352 736 84392 776
rect 84434 736 84474 776
rect 84516 736 84556 776
rect 84598 736 84638 776
rect 84680 736 84720 776
rect 88352 736 88392 776
rect 88434 736 88474 776
rect 88516 736 88556 776
rect 88598 736 88638 776
rect 88680 736 88720 776
rect 92352 736 92392 776
rect 92434 736 92474 776
rect 92516 736 92556 776
rect 92598 736 92638 776
rect 92680 736 92720 776
rect 96352 736 96392 776
rect 96434 736 96474 776
rect 96516 736 96556 776
rect 96598 736 96638 776
rect 96680 736 96720 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 8352 38576 8720 38585
rect 8392 38536 8434 38576
rect 8474 38536 8516 38576
rect 8556 38536 8598 38576
rect 8638 38536 8680 38576
rect 8352 38527 8720 38536
rect 12352 38576 12720 38585
rect 12392 38536 12434 38576
rect 12474 38536 12516 38576
rect 12556 38536 12598 38576
rect 12638 38536 12680 38576
rect 12352 38527 12720 38536
rect 16352 38576 16720 38585
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16352 38527 16720 38536
rect 20352 38576 20720 38585
rect 20392 38536 20434 38576
rect 20474 38536 20516 38576
rect 20556 38536 20598 38576
rect 20638 38536 20680 38576
rect 20352 38527 20720 38536
rect 24352 38576 24720 38585
rect 24392 38536 24434 38576
rect 24474 38536 24516 38576
rect 24556 38536 24598 38576
rect 24638 38536 24680 38576
rect 24352 38527 24720 38536
rect 28352 38576 28720 38585
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28352 38527 28720 38536
rect 32352 38576 32720 38585
rect 32392 38536 32434 38576
rect 32474 38536 32516 38576
rect 32556 38536 32598 38576
rect 32638 38536 32680 38576
rect 32352 38527 32720 38536
rect 36352 38576 36720 38585
rect 36392 38536 36434 38576
rect 36474 38536 36516 38576
rect 36556 38536 36598 38576
rect 36638 38536 36680 38576
rect 36352 38527 36720 38536
rect 40352 38576 40720 38585
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40352 38527 40720 38536
rect 44352 38576 44720 38585
rect 44392 38536 44434 38576
rect 44474 38536 44516 38576
rect 44556 38536 44598 38576
rect 44638 38536 44680 38576
rect 44352 38527 44720 38536
rect 48352 38576 48720 38585
rect 48392 38536 48434 38576
rect 48474 38536 48516 38576
rect 48556 38536 48598 38576
rect 48638 38536 48680 38576
rect 48352 38527 48720 38536
rect 52352 38576 52720 38585
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52352 38527 52720 38536
rect 56352 38576 56720 38585
rect 56392 38536 56434 38576
rect 56474 38536 56516 38576
rect 56556 38536 56598 38576
rect 56638 38536 56680 38576
rect 56352 38527 56720 38536
rect 60352 38576 60720 38585
rect 60392 38536 60434 38576
rect 60474 38536 60516 38576
rect 60556 38536 60598 38576
rect 60638 38536 60680 38576
rect 60352 38527 60720 38536
rect 64352 38576 64720 38585
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64352 38527 64720 38536
rect 68352 38576 68720 38585
rect 68392 38536 68434 38576
rect 68474 38536 68516 38576
rect 68556 38536 68598 38576
rect 68638 38536 68680 38576
rect 68352 38527 68720 38536
rect 72352 38576 72720 38585
rect 72392 38536 72434 38576
rect 72474 38536 72516 38576
rect 72556 38536 72598 38576
rect 72638 38536 72680 38576
rect 72352 38527 72720 38536
rect 76352 38576 76720 38585
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76352 38527 76720 38536
rect 80352 38576 80720 38585
rect 80392 38536 80434 38576
rect 80474 38536 80516 38576
rect 80556 38536 80598 38576
rect 80638 38536 80680 38576
rect 80352 38527 80720 38536
rect 84352 38576 84720 38585
rect 84392 38536 84434 38576
rect 84474 38536 84516 38576
rect 84556 38536 84598 38576
rect 84638 38536 84680 38576
rect 84352 38527 84720 38536
rect 88352 38576 88720 38585
rect 88392 38536 88434 38576
rect 88474 38536 88516 38576
rect 88556 38536 88598 38576
rect 88638 38536 88680 38576
rect 88352 38527 88720 38536
rect 92352 38576 92720 38585
rect 92392 38536 92434 38576
rect 92474 38536 92516 38576
rect 92556 38536 92598 38576
rect 92638 38536 92680 38576
rect 92352 38527 92720 38536
rect 96352 38576 96720 38585
rect 96392 38536 96434 38576
rect 96474 38536 96516 38576
rect 96556 38536 96598 38576
rect 96638 38536 96680 38576
rect 96352 38527 96720 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 7112 37820 7480 37829
rect 7152 37780 7194 37820
rect 7234 37780 7276 37820
rect 7316 37780 7358 37820
rect 7398 37780 7440 37820
rect 7112 37771 7480 37780
rect 11112 37820 11480 37829
rect 11152 37780 11194 37820
rect 11234 37780 11276 37820
rect 11316 37780 11358 37820
rect 11398 37780 11440 37820
rect 11112 37771 11480 37780
rect 15112 37820 15480 37829
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15112 37771 15480 37780
rect 19112 37820 19480 37829
rect 19152 37780 19194 37820
rect 19234 37780 19276 37820
rect 19316 37780 19358 37820
rect 19398 37780 19440 37820
rect 19112 37771 19480 37780
rect 23112 37820 23480 37829
rect 23152 37780 23194 37820
rect 23234 37780 23276 37820
rect 23316 37780 23358 37820
rect 23398 37780 23440 37820
rect 23112 37771 23480 37780
rect 27112 37820 27480 37829
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27112 37771 27480 37780
rect 31112 37820 31480 37829
rect 31152 37780 31194 37820
rect 31234 37780 31276 37820
rect 31316 37780 31358 37820
rect 31398 37780 31440 37820
rect 31112 37771 31480 37780
rect 35112 37820 35480 37829
rect 35152 37780 35194 37820
rect 35234 37780 35276 37820
rect 35316 37780 35358 37820
rect 35398 37780 35440 37820
rect 35112 37771 35480 37780
rect 39112 37820 39480 37829
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39112 37771 39480 37780
rect 43112 37820 43480 37829
rect 43152 37780 43194 37820
rect 43234 37780 43276 37820
rect 43316 37780 43358 37820
rect 43398 37780 43440 37820
rect 43112 37771 43480 37780
rect 47112 37820 47480 37829
rect 47152 37780 47194 37820
rect 47234 37780 47276 37820
rect 47316 37780 47358 37820
rect 47398 37780 47440 37820
rect 47112 37771 47480 37780
rect 51112 37820 51480 37829
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51112 37771 51480 37780
rect 55112 37820 55480 37829
rect 55152 37780 55194 37820
rect 55234 37780 55276 37820
rect 55316 37780 55358 37820
rect 55398 37780 55440 37820
rect 55112 37771 55480 37780
rect 59112 37820 59480 37829
rect 59152 37780 59194 37820
rect 59234 37780 59276 37820
rect 59316 37780 59358 37820
rect 59398 37780 59440 37820
rect 59112 37771 59480 37780
rect 63112 37820 63480 37829
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63112 37771 63480 37780
rect 67112 37820 67480 37829
rect 67152 37780 67194 37820
rect 67234 37780 67276 37820
rect 67316 37780 67358 37820
rect 67398 37780 67440 37820
rect 67112 37771 67480 37780
rect 71112 37820 71480 37829
rect 71152 37780 71194 37820
rect 71234 37780 71276 37820
rect 71316 37780 71358 37820
rect 71398 37780 71440 37820
rect 71112 37771 71480 37780
rect 75112 37820 75480 37829
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75112 37771 75480 37780
rect 79112 37820 79480 37829
rect 79152 37780 79194 37820
rect 79234 37780 79276 37820
rect 79316 37780 79358 37820
rect 79398 37780 79440 37820
rect 79112 37771 79480 37780
rect 83112 37820 83480 37829
rect 83152 37780 83194 37820
rect 83234 37780 83276 37820
rect 83316 37780 83358 37820
rect 83398 37780 83440 37820
rect 83112 37771 83480 37780
rect 87112 37820 87480 37829
rect 87152 37780 87194 37820
rect 87234 37780 87276 37820
rect 87316 37780 87358 37820
rect 87398 37780 87440 37820
rect 87112 37771 87480 37780
rect 91112 37820 91480 37829
rect 91152 37780 91194 37820
rect 91234 37780 91276 37820
rect 91316 37780 91358 37820
rect 91398 37780 91440 37820
rect 91112 37771 91480 37780
rect 95112 37820 95480 37829
rect 95152 37780 95194 37820
rect 95234 37780 95276 37820
rect 95316 37780 95358 37820
rect 95398 37780 95440 37820
rect 95112 37771 95480 37780
rect 99112 37820 99480 37829
rect 99152 37780 99194 37820
rect 99234 37780 99276 37820
rect 99316 37780 99358 37820
rect 99398 37780 99440 37820
rect 99112 37771 99480 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 8352 37064 8720 37073
rect 8392 37024 8434 37064
rect 8474 37024 8516 37064
rect 8556 37024 8598 37064
rect 8638 37024 8680 37064
rect 8352 37015 8720 37024
rect 12352 37064 12720 37073
rect 12392 37024 12434 37064
rect 12474 37024 12516 37064
rect 12556 37024 12598 37064
rect 12638 37024 12680 37064
rect 12352 37015 12720 37024
rect 16352 37064 16720 37073
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16352 37015 16720 37024
rect 20352 37064 20720 37073
rect 20392 37024 20434 37064
rect 20474 37024 20516 37064
rect 20556 37024 20598 37064
rect 20638 37024 20680 37064
rect 20352 37015 20720 37024
rect 24352 37064 24720 37073
rect 24392 37024 24434 37064
rect 24474 37024 24516 37064
rect 24556 37024 24598 37064
rect 24638 37024 24680 37064
rect 24352 37015 24720 37024
rect 28352 37064 28720 37073
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28352 37015 28720 37024
rect 32352 37064 32720 37073
rect 32392 37024 32434 37064
rect 32474 37024 32516 37064
rect 32556 37024 32598 37064
rect 32638 37024 32680 37064
rect 32352 37015 32720 37024
rect 36352 37064 36720 37073
rect 36392 37024 36434 37064
rect 36474 37024 36516 37064
rect 36556 37024 36598 37064
rect 36638 37024 36680 37064
rect 36352 37015 36720 37024
rect 40352 37064 40720 37073
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40352 37015 40720 37024
rect 44352 37064 44720 37073
rect 44392 37024 44434 37064
rect 44474 37024 44516 37064
rect 44556 37024 44598 37064
rect 44638 37024 44680 37064
rect 44352 37015 44720 37024
rect 48352 37064 48720 37073
rect 48392 37024 48434 37064
rect 48474 37024 48516 37064
rect 48556 37024 48598 37064
rect 48638 37024 48680 37064
rect 48352 37015 48720 37024
rect 52352 37064 52720 37073
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52352 37015 52720 37024
rect 56352 37064 56720 37073
rect 56392 37024 56434 37064
rect 56474 37024 56516 37064
rect 56556 37024 56598 37064
rect 56638 37024 56680 37064
rect 56352 37015 56720 37024
rect 60352 37064 60720 37073
rect 60392 37024 60434 37064
rect 60474 37024 60516 37064
rect 60556 37024 60598 37064
rect 60638 37024 60680 37064
rect 60352 37015 60720 37024
rect 64352 37064 64720 37073
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64352 37015 64720 37024
rect 68352 37064 68720 37073
rect 68392 37024 68434 37064
rect 68474 37024 68516 37064
rect 68556 37024 68598 37064
rect 68638 37024 68680 37064
rect 68352 37015 68720 37024
rect 72352 37064 72720 37073
rect 72392 37024 72434 37064
rect 72474 37024 72516 37064
rect 72556 37024 72598 37064
rect 72638 37024 72680 37064
rect 72352 37015 72720 37024
rect 76352 37064 76720 37073
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76352 37015 76720 37024
rect 80352 37064 80720 37073
rect 80392 37024 80434 37064
rect 80474 37024 80516 37064
rect 80556 37024 80598 37064
rect 80638 37024 80680 37064
rect 80352 37015 80720 37024
rect 84352 37064 84720 37073
rect 84392 37024 84434 37064
rect 84474 37024 84516 37064
rect 84556 37024 84598 37064
rect 84638 37024 84680 37064
rect 84352 37015 84720 37024
rect 88352 37064 88720 37073
rect 88392 37024 88434 37064
rect 88474 37024 88516 37064
rect 88556 37024 88598 37064
rect 88638 37024 88680 37064
rect 88352 37015 88720 37024
rect 92352 37064 92720 37073
rect 92392 37024 92434 37064
rect 92474 37024 92516 37064
rect 92556 37024 92598 37064
rect 92638 37024 92680 37064
rect 92352 37015 92720 37024
rect 96352 37064 96720 37073
rect 96392 37024 96434 37064
rect 96474 37024 96516 37064
rect 96556 37024 96598 37064
rect 96638 37024 96680 37064
rect 96352 37015 96720 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 7112 36308 7480 36317
rect 7152 36268 7194 36308
rect 7234 36268 7276 36308
rect 7316 36268 7358 36308
rect 7398 36268 7440 36308
rect 7112 36259 7480 36268
rect 11112 36308 11480 36317
rect 11152 36268 11194 36308
rect 11234 36268 11276 36308
rect 11316 36268 11358 36308
rect 11398 36268 11440 36308
rect 11112 36259 11480 36268
rect 15112 36308 15480 36317
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15112 36259 15480 36268
rect 19112 36308 19480 36317
rect 19152 36268 19194 36308
rect 19234 36268 19276 36308
rect 19316 36268 19358 36308
rect 19398 36268 19440 36308
rect 19112 36259 19480 36268
rect 23112 36308 23480 36317
rect 23152 36268 23194 36308
rect 23234 36268 23276 36308
rect 23316 36268 23358 36308
rect 23398 36268 23440 36308
rect 23112 36259 23480 36268
rect 27112 36308 27480 36317
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27112 36259 27480 36268
rect 31112 36308 31480 36317
rect 31152 36268 31194 36308
rect 31234 36268 31276 36308
rect 31316 36268 31358 36308
rect 31398 36268 31440 36308
rect 31112 36259 31480 36268
rect 35112 36308 35480 36317
rect 35152 36268 35194 36308
rect 35234 36268 35276 36308
rect 35316 36268 35358 36308
rect 35398 36268 35440 36308
rect 35112 36259 35480 36268
rect 39112 36308 39480 36317
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39112 36259 39480 36268
rect 43112 36308 43480 36317
rect 43152 36268 43194 36308
rect 43234 36268 43276 36308
rect 43316 36268 43358 36308
rect 43398 36268 43440 36308
rect 43112 36259 43480 36268
rect 47112 36308 47480 36317
rect 47152 36268 47194 36308
rect 47234 36268 47276 36308
rect 47316 36268 47358 36308
rect 47398 36268 47440 36308
rect 47112 36259 47480 36268
rect 51112 36308 51480 36317
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51112 36259 51480 36268
rect 55112 36308 55480 36317
rect 55152 36268 55194 36308
rect 55234 36268 55276 36308
rect 55316 36268 55358 36308
rect 55398 36268 55440 36308
rect 55112 36259 55480 36268
rect 59112 36308 59480 36317
rect 59152 36268 59194 36308
rect 59234 36268 59276 36308
rect 59316 36268 59358 36308
rect 59398 36268 59440 36308
rect 59112 36259 59480 36268
rect 63112 36308 63480 36317
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63112 36259 63480 36268
rect 67112 36308 67480 36317
rect 67152 36268 67194 36308
rect 67234 36268 67276 36308
rect 67316 36268 67358 36308
rect 67398 36268 67440 36308
rect 67112 36259 67480 36268
rect 71112 36308 71480 36317
rect 71152 36268 71194 36308
rect 71234 36268 71276 36308
rect 71316 36268 71358 36308
rect 71398 36268 71440 36308
rect 71112 36259 71480 36268
rect 75112 36308 75480 36317
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75112 36259 75480 36268
rect 79112 36308 79480 36317
rect 79152 36268 79194 36308
rect 79234 36268 79276 36308
rect 79316 36268 79358 36308
rect 79398 36268 79440 36308
rect 79112 36259 79480 36268
rect 83112 36308 83480 36317
rect 83152 36268 83194 36308
rect 83234 36268 83276 36308
rect 83316 36268 83358 36308
rect 83398 36268 83440 36308
rect 83112 36259 83480 36268
rect 87112 36308 87480 36317
rect 87152 36268 87194 36308
rect 87234 36268 87276 36308
rect 87316 36268 87358 36308
rect 87398 36268 87440 36308
rect 87112 36259 87480 36268
rect 91112 36308 91480 36317
rect 91152 36268 91194 36308
rect 91234 36268 91276 36308
rect 91316 36268 91358 36308
rect 91398 36268 91440 36308
rect 91112 36259 91480 36268
rect 95112 36308 95480 36317
rect 95152 36268 95194 36308
rect 95234 36268 95276 36308
rect 95316 36268 95358 36308
rect 95398 36268 95440 36308
rect 95112 36259 95480 36268
rect 99112 36308 99480 36317
rect 99152 36268 99194 36308
rect 99234 36268 99276 36308
rect 99316 36268 99358 36308
rect 99398 36268 99440 36308
rect 99112 36259 99480 36268
rect 74860 35972 74900 35981
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 8352 35552 8720 35561
rect 8392 35512 8434 35552
rect 8474 35512 8516 35552
rect 8556 35512 8598 35552
rect 8638 35512 8680 35552
rect 8352 35503 8720 35512
rect 12352 35552 12720 35561
rect 12392 35512 12434 35552
rect 12474 35512 12516 35552
rect 12556 35512 12598 35552
rect 12638 35512 12680 35552
rect 12352 35503 12720 35512
rect 16352 35552 16720 35561
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16352 35503 16720 35512
rect 20352 35552 20720 35561
rect 20392 35512 20434 35552
rect 20474 35512 20516 35552
rect 20556 35512 20598 35552
rect 20638 35512 20680 35552
rect 20352 35503 20720 35512
rect 24352 35552 24720 35561
rect 24392 35512 24434 35552
rect 24474 35512 24516 35552
rect 24556 35512 24598 35552
rect 24638 35512 24680 35552
rect 24352 35503 24720 35512
rect 28352 35552 28720 35561
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28352 35503 28720 35512
rect 32352 35552 32720 35561
rect 32392 35512 32434 35552
rect 32474 35512 32516 35552
rect 32556 35512 32598 35552
rect 32638 35512 32680 35552
rect 32352 35503 32720 35512
rect 36352 35552 36720 35561
rect 36392 35512 36434 35552
rect 36474 35512 36516 35552
rect 36556 35512 36598 35552
rect 36638 35512 36680 35552
rect 36352 35503 36720 35512
rect 40352 35552 40720 35561
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40352 35503 40720 35512
rect 44352 35552 44720 35561
rect 44392 35512 44434 35552
rect 44474 35512 44516 35552
rect 44556 35512 44598 35552
rect 44638 35512 44680 35552
rect 44352 35503 44720 35512
rect 48352 35552 48720 35561
rect 48392 35512 48434 35552
rect 48474 35512 48516 35552
rect 48556 35512 48598 35552
rect 48638 35512 48680 35552
rect 48352 35503 48720 35512
rect 52352 35552 52720 35561
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52352 35503 52720 35512
rect 56352 35552 56720 35561
rect 56392 35512 56434 35552
rect 56474 35512 56516 35552
rect 56556 35512 56598 35552
rect 56638 35512 56680 35552
rect 56352 35503 56720 35512
rect 60352 35552 60720 35561
rect 60392 35512 60434 35552
rect 60474 35512 60516 35552
rect 60556 35512 60598 35552
rect 60638 35512 60680 35552
rect 60352 35503 60720 35512
rect 64352 35552 64720 35561
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64352 35503 64720 35512
rect 68352 35552 68720 35561
rect 68392 35512 68434 35552
rect 68474 35512 68516 35552
rect 68556 35512 68598 35552
rect 68638 35512 68680 35552
rect 68352 35503 68720 35512
rect 72352 35552 72720 35561
rect 72392 35512 72434 35552
rect 72474 35512 72516 35552
rect 72556 35512 72598 35552
rect 72638 35512 72680 35552
rect 72352 35503 72720 35512
rect 73708 35132 73748 35143
rect 74860 35141 74900 35932
rect 76588 35972 76628 35981
rect 77452 35972 77492 35981
rect 78604 35972 78644 35981
rect 79372 35972 79412 35981
rect 76628 35932 76820 35972
rect 76588 35923 76628 35932
rect 76780 35888 76820 35932
rect 77492 35932 77588 35972
rect 77452 35923 77492 35932
rect 76780 35848 76916 35888
rect 75052 35720 75092 35729
rect 74956 35680 75052 35720
rect 73708 35057 73748 35092
rect 73899 35132 73941 35141
rect 73899 35092 73900 35132
rect 73940 35092 73941 35132
rect 73899 35083 73941 35092
rect 74091 35132 74133 35141
rect 74091 35092 74092 35132
rect 74132 35092 74133 35132
rect 74091 35083 74133 35092
rect 74668 35132 74708 35141
rect 74859 35132 74901 35141
rect 74708 35092 74804 35132
rect 74668 35083 74708 35092
rect 73707 35048 73749 35057
rect 73707 35008 73708 35048
rect 73748 35008 73749 35048
rect 73707 34999 73749 35008
rect 73900 34964 73940 35083
rect 74092 34998 74132 35083
rect 74475 35048 74517 35057
rect 74475 35008 74476 35048
rect 74516 35008 74517 35048
rect 74475 34999 74517 35008
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 7112 34796 7480 34805
rect 7152 34756 7194 34796
rect 7234 34756 7276 34796
rect 7316 34756 7358 34796
rect 7398 34756 7440 34796
rect 7112 34747 7480 34756
rect 11112 34796 11480 34805
rect 11152 34756 11194 34796
rect 11234 34756 11276 34796
rect 11316 34756 11358 34796
rect 11398 34756 11440 34796
rect 11112 34747 11480 34756
rect 15112 34796 15480 34805
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15112 34747 15480 34756
rect 19112 34796 19480 34805
rect 19152 34756 19194 34796
rect 19234 34756 19276 34796
rect 19316 34756 19358 34796
rect 19398 34756 19440 34796
rect 19112 34747 19480 34756
rect 23112 34796 23480 34805
rect 23152 34756 23194 34796
rect 23234 34756 23276 34796
rect 23316 34756 23358 34796
rect 23398 34756 23440 34796
rect 23112 34747 23480 34756
rect 27112 34796 27480 34805
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27112 34747 27480 34756
rect 31112 34796 31480 34805
rect 31152 34756 31194 34796
rect 31234 34756 31276 34796
rect 31316 34756 31358 34796
rect 31398 34756 31440 34796
rect 31112 34747 31480 34756
rect 35112 34796 35480 34805
rect 35152 34756 35194 34796
rect 35234 34756 35276 34796
rect 35316 34756 35358 34796
rect 35398 34756 35440 34796
rect 35112 34747 35480 34756
rect 39112 34796 39480 34805
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39112 34747 39480 34756
rect 43112 34796 43480 34805
rect 43152 34756 43194 34796
rect 43234 34756 43276 34796
rect 43316 34756 43358 34796
rect 43398 34756 43440 34796
rect 43112 34747 43480 34756
rect 47112 34796 47480 34805
rect 47152 34756 47194 34796
rect 47234 34756 47276 34796
rect 47316 34756 47358 34796
rect 47398 34756 47440 34796
rect 47112 34747 47480 34756
rect 51112 34796 51480 34805
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51112 34747 51480 34756
rect 55112 34796 55480 34805
rect 55152 34756 55194 34796
rect 55234 34756 55276 34796
rect 55316 34756 55358 34796
rect 55398 34756 55440 34796
rect 55112 34747 55480 34756
rect 59112 34796 59480 34805
rect 59152 34756 59194 34796
rect 59234 34756 59276 34796
rect 59316 34756 59358 34796
rect 59398 34756 59440 34796
rect 59112 34747 59480 34756
rect 63112 34796 63480 34805
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63112 34747 63480 34756
rect 67112 34796 67480 34805
rect 67152 34756 67194 34796
rect 67234 34756 67276 34796
rect 67316 34756 67358 34796
rect 67398 34756 67440 34796
rect 67112 34747 67480 34756
rect 71112 34796 71480 34805
rect 71152 34756 71194 34796
rect 71234 34756 71276 34796
rect 71316 34756 71358 34796
rect 71398 34756 71440 34796
rect 71112 34747 71480 34756
rect 69771 34460 69813 34469
rect 69771 34420 69772 34460
rect 69812 34420 69813 34460
rect 69771 34411 69813 34420
rect 73419 34460 73461 34469
rect 73419 34420 73420 34460
rect 73460 34420 73461 34460
rect 73419 34411 73461 34420
rect 73900 34460 73940 34924
rect 73900 34411 73940 34420
rect 74284 34964 74324 34973
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 8352 34040 8720 34049
rect 8392 34000 8434 34040
rect 8474 34000 8516 34040
rect 8556 34000 8598 34040
rect 8638 34000 8680 34040
rect 8352 33991 8720 34000
rect 12352 34040 12720 34049
rect 12392 34000 12434 34040
rect 12474 34000 12516 34040
rect 12556 34000 12598 34040
rect 12638 34000 12680 34040
rect 12352 33991 12720 34000
rect 16352 34040 16720 34049
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16352 33991 16720 34000
rect 20352 34040 20720 34049
rect 20392 34000 20434 34040
rect 20474 34000 20516 34040
rect 20556 34000 20598 34040
rect 20638 34000 20680 34040
rect 20352 33991 20720 34000
rect 24352 34040 24720 34049
rect 24392 34000 24434 34040
rect 24474 34000 24516 34040
rect 24556 34000 24598 34040
rect 24638 34000 24680 34040
rect 24352 33991 24720 34000
rect 28352 34040 28720 34049
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28352 33991 28720 34000
rect 32352 34040 32720 34049
rect 32392 34000 32434 34040
rect 32474 34000 32516 34040
rect 32556 34000 32598 34040
rect 32638 34000 32680 34040
rect 32352 33991 32720 34000
rect 36352 34040 36720 34049
rect 36392 34000 36434 34040
rect 36474 34000 36516 34040
rect 36556 34000 36598 34040
rect 36638 34000 36680 34040
rect 36352 33991 36720 34000
rect 40352 34040 40720 34049
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40352 33991 40720 34000
rect 44352 34040 44720 34049
rect 44392 34000 44434 34040
rect 44474 34000 44516 34040
rect 44556 34000 44598 34040
rect 44638 34000 44680 34040
rect 44352 33991 44720 34000
rect 48352 34040 48720 34049
rect 48392 34000 48434 34040
rect 48474 34000 48516 34040
rect 48556 34000 48598 34040
rect 48638 34000 48680 34040
rect 48352 33991 48720 34000
rect 52352 34040 52720 34049
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52352 33991 52720 34000
rect 56352 34040 56720 34049
rect 56392 34000 56434 34040
rect 56474 34000 56516 34040
rect 56556 34000 56598 34040
rect 56638 34000 56680 34040
rect 56352 33991 56720 34000
rect 60352 34040 60720 34049
rect 60392 34000 60434 34040
rect 60474 34000 60516 34040
rect 60556 34000 60598 34040
rect 60638 34000 60680 34040
rect 60352 33991 60720 34000
rect 64352 34040 64720 34049
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64352 33991 64720 34000
rect 68352 34040 68720 34049
rect 68392 34000 68434 34040
rect 68474 34000 68516 34040
rect 68556 34000 68598 34040
rect 68638 34000 68680 34040
rect 68352 33991 68720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 7112 33284 7480 33293
rect 7152 33244 7194 33284
rect 7234 33244 7276 33284
rect 7316 33244 7358 33284
rect 7398 33244 7440 33284
rect 7112 33235 7480 33244
rect 11112 33284 11480 33293
rect 11152 33244 11194 33284
rect 11234 33244 11276 33284
rect 11316 33244 11358 33284
rect 11398 33244 11440 33284
rect 11112 33235 11480 33244
rect 15112 33284 15480 33293
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15112 33235 15480 33244
rect 19112 33284 19480 33293
rect 19152 33244 19194 33284
rect 19234 33244 19276 33284
rect 19316 33244 19358 33284
rect 19398 33244 19440 33284
rect 19112 33235 19480 33244
rect 23112 33284 23480 33293
rect 23152 33244 23194 33284
rect 23234 33244 23276 33284
rect 23316 33244 23358 33284
rect 23398 33244 23440 33284
rect 23112 33235 23480 33244
rect 27112 33284 27480 33293
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27112 33235 27480 33244
rect 31112 33284 31480 33293
rect 31152 33244 31194 33284
rect 31234 33244 31276 33284
rect 31316 33244 31358 33284
rect 31398 33244 31440 33284
rect 31112 33235 31480 33244
rect 35112 33284 35480 33293
rect 35152 33244 35194 33284
rect 35234 33244 35276 33284
rect 35316 33244 35358 33284
rect 35398 33244 35440 33284
rect 35112 33235 35480 33244
rect 39112 33284 39480 33293
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39112 33235 39480 33244
rect 43112 33284 43480 33293
rect 43152 33244 43194 33284
rect 43234 33244 43276 33284
rect 43316 33244 43358 33284
rect 43398 33244 43440 33284
rect 43112 33235 43480 33244
rect 47112 33284 47480 33293
rect 47152 33244 47194 33284
rect 47234 33244 47276 33284
rect 47316 33244 47358 33284
rect 47398 33244 47440 33284
rect 47112 33235 47480 33244
rect 51112 33284 51480 33293
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51112 33235 51480 33244
rect 55112 33284 55480 33293
rect 55152 33244 55194 33284
rect 55234 33244 55276 33284
rect 55316 33244 55358 33284
rect 55398 33244 55440 33284
rect 55112 33235 55480 33244
rect 59112 33284 59480 33293
rect 59152 33244 59194 33284
rect 59234 33244 59276 33284
rect 59316 33244 59358 33284
rect 59398 33244 59440 33284
rect 59112 33235 59480 33244
rect 63112 33284 63480 33293
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63112 33235 63480 33244
rect 67112 33284 67480 33293
rect 67152 33244 67194 33284
rect 67234 33244 67276 33284
rect 67316 33244 67358 33284
rect 67398 33244 67440 33284
rect 67112 33235 67480 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 8352 32528 8720 32537
rect 8392 32488 8434 32528
rect 8474 32488 8516 32528
rect 8556 32488 8598 32528
rect 8638 32488 8680 32528
rect 8352 32479 8720 32488
rect 12352 32528 12720 32537
rect 12392 32488 12434 32528
rect 12474 32488 12516 32528
rect 12556 32488 12598 32528
rect 12638 32488 12680 32528
rect 12352 32479 12720 32488
rect 16352 32528 16720 32537
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16352 32479 16720 32488
rect 20352 32528 20720 32537
rect 20392 32488 20434 32528
rect 20474 32488 20516 32528
rect 20556 32488 20598 32528
rect 20638 32488 20680 32528
rect 20352 32479 20720 32488
rect 24352 32528 24720 32537
rect 24392 32488 24434 32528
rect 24474 32488 24516 32528
rect 24556 32488 24598 32528
rect 24638 32488 24680 32528
rect 24352 32479 24720 32488
rect 28352 32528 28720 32537
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28352 32479 28720 32488
rect 32352 32528 32720 32537
rect 32392 32488 32434 32528
rect 32474 32488 32516 32528
rect 32556 32488 32598 32528
rect 32638 32488 32680 32528
rect 32352 32479 32720 32488
rect 36352 32528 36720 32537
rect 36392 32488 36434 32528
rect 36474 32488 36516 32528
rect 36556 32488 36598 32528
rect 36638 32488 36680 32528
rect 36352 32479 36720 32488
rect 40352 32528 40720 32537
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40352 32479 40720 32488
rect 44352 32528 44720 32537
rect 44392 32488 44434 32528
rect 44474 32488 44516 32528
rect 44556 32488 44598 32528
rect 44638 32488 44680 32528
rect 44352 32479 44720 32488
rect 48352 32528 48720 32537
rect 48392 32488 48434 32528
rect 48474 32488 48516 32528
rect 48556 32488 48598 32528
rect 48638 32488 48680 32528
rect 48352 32479 48720 32488
rect 52352 32528 52720 32537
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52352 32479 52720 32488
rect 56352 32528 56720 32537
rect 56392 32488 56434 32528
rect 56474 32488 56516 32528
rect 56556 32488 56598 32528
rect 56638 32488 56680 32528
rect 56352 32479 56720 32488
rect 60352 32528 60720 32537
rect 60392 32488 60434 32528
rect 60474 32488 60516 32528
rect 60556 32488 60598 32528
rect 60638 32488 60680 32528
rect 60352 32479 60720 32488
rect 64352 32528 64720 32537
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64352 32479 64720 32488
rect 68352 32528 68720 32537
rect 68392 32488 68434 32528
rect 68474 32488 68516 32528
rect 68556 32488 68598 32528
rect 68638 32488 68680 32528
rect 68352 32479 68720 32488
rect 69772 32192 69812 34411
rect 73420 34326 73460 34411
rect 73612 34208 73652 34217
rect 74092 34208 74132 34217
rect 73652 34168 74036 34208
rect 73612 34159 73652 34168
rect 72352 34040 72720 34049
rect 72392 34000 72434 34040
rect 72474 34000 72516 34040
rect 72556 34000 72598 34040
rect 72638 34000 72680 34040
rect 72352 33991 72720 34000
rect 71787 32780 71829 32789
rect 71787 32740 71788 32780
rect 71828 32740 71829 32780
rect 71787 32731 71829 32740
rect 67563 32108 67605 32117
rect 67563 32068 67564 32108
rect 67604 32068 67605 32108
rect 67563 32059 67605 32068
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 7112 31772 7480 31781
rect 7152 31732 7194 31772
rect 7234 31732 7276 31772
rect 7316 31732 7358 31772
rect 7398 31732 7440 31772
rect 7112 31723 7480 31732
rect 11112 31772 11480 31781
rect 11152 31732 11194 31772
rect 11234 31732 11276 31772
rect 11316 31732 11358 31772
rect 11398 31732 11440 31772
rect 11112 31723 11480 31732
rect 15112 31772 15480 31781
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15112 31723 15480 31732
rect 19112 31772 19480 31781
rect 19152 31732 19194 31772
rect 19234 31732 19276 31772
rect 19316 31732 19358 31772
rect 19398 31732 19440 31772
rect 19112 31723 19480 31732
rect 23112 31772 23480 31781
rect 23152 31732 23194 31772
rect 23234 31732 23276 31772
rect 23316 31732 23358 31772
rect 23398 31732 23440 31772
rect 23112 31723 23480 31732
rect 27112 31772 27480 31781
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27112 31723 27480 31732
rect 31112 31772 31480 31781
rect 31152 31732 31194 31772
rect 31234 31732 31276 31772
rect 31316 31732 31358 31772
rect 31398 31732 31440 31772
rect 31112 31723 31480 31732
rect 35112 31772 35480 31781
rect 35152 31732 35194 31772
rect 35234 31732 35276 31772
rect 35316 31732 35358 31772
rect 35398 31732 35440 31772
rect 35112 31723 35480 31732
rect 39112 31772 39480 31781
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39112 31723 39480 31732
rect 43112 31772 43480 31781
rect 43152 31732 43194 31772
rect 43234 31732 43276 31772
rect 43316 31732 43358 31772
rect 43398 31732 43440 31772
rect 43112 31723 43480 31732
rect 47112 31772 47480 31781
rect 47152 31732 47194 31772
rect 47234 31732 47276 31772
rect 47316 31732 47358 31772
rect 47398 31732 47440 31772
rect 47112 31723 47480 31732
rect 51112 31772 51480 31781
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51112 31723 51480 31732
rect 55112 31772 55480 31781
rect 55152 31732 55194 31772
rect 55234 31732 55276 31772
rect 55316 31732 55358 31772
rect 55398 31732 55440 31772
rect 55112 31723 55480 31732
rect 59112 31772 59480 31781
rect 59152 31732 59194 31772
rect 59234 31732 59276 31772
rect 59316 31732 59358 31772
rect 59398 31732 59440 31772
rect 59112 31723 59480 31732
rect 63112 31772 63480 31781
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63112 31723 63480 31732
rect 67112 31772 67480 31781
rect 67152 31732 67194 31772
rect 67234 31732 67276 31772
rect 67316 31732 67358 31772
rect 67398 31732 67440 31772
rect 67112 31723 67480 31732
rect 67564 31613 67604 32059
rect 68907 31856 68949 31865
rect 68907 31816 68908 31856
rect 68948 31816 68949 31856
rect 68907 31807 68949 31816
rect 67179 31604 67221 31613
rect 67179 31564 67180 31604
rect 67220 31564 67221 31604
rect 67179 31555 67221 31564
rect 67563 31604 67605 31613
rect 67563 31564 67564 31604
rect 67604 31564 67605 31604
rect 67563 31555 67605 31564
rect 68811 31604 68853 31613
rect 68811 31564 68812 31604
rect 68852 31564 68853 31604
rect 68811 31555 68853 31564
rect 67180 31520 67220 31555
rect 67180 31469 67220 31480
rect 67659 31520 67701 31529
rect 67659 31480 67660 31520
rect 67700 31480 67701 31520
rect 67659 31471 67701 31480
rect 67276 31352 67316 31363
rect 67276 31277 67316 31312
rect 67564 31352 67604 31363
rect 67564 31277 67604 31312
rect 67275 31268 67317 31277
rect 67275 31228 67276 31268
rect 67316 31228 67317 31268
rect 67275 31219 67317 31228
rect 67563 31268 67605 31277
rect 67563 31228 67564 31268
rect 67604 31228 67605 31268
rect 67563 31219 67605 31228
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 8352 31016 8720 31025
rect 8392 30976 8434 31016
rect 8474 30976 8516 31016
rect 8556 30976 8598 31016
rect 8638 30976 8680 31016
rect 8352 30967 8720 30976
rect 12352 31016 12720 31025
rect 12392 30976 12434 31016
rect 12474 30976 12516 31016
rect 12556 30976 12598 31016
rect 12638 30976 12680 31016
rect 12352 30967 12720 30976
rect 16352 31016 16720 31025
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16352 30967 16720 30976
rect 20352 31016 20720 31025
rect 20392 30976 20434 31016
rect 20474 30976 20516 31016
rect 20556 30976 20598 31016
rect 20638 30976 20680 31016
rect 20352 30967 20720 30976
rect 24352 31016 24720 31025
rect 24392 30976 24434 31016
rect 24474 30976 24516 31016
rect 24556 30976 24598 31016
rect 24638 30976 24680 31016
rect 24352 30967 24720 30976
rect 28352 31016 28720 31025
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28352 30967 28720 30976
rect 32352 31016 32720 31025
rect 32392 30976 32434 31016
rect 32474 30976 32516 31016
rect 32556 30976 32598 31016
rect 32638 30976 32680 31016
rect 32352 30967 32720 30976
rect 36352 31016 36720 31025
rect 36392 30976 36434 31016
rect 36474 30976 36516 31016
rect 36556 30976 36598 31016
rect 36638 30976 36680 31016
rect 36352 30967 36720 30976
rect 40352 31016 40720 31025
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40352 30967 40720 30976
rect 44352 31016 44720 31025
rect 44392 30976 44434 31016
rect 44474 30976 44516 31016
rect 44556 30976 44598 31016
rect 44638 30976 44680 31016
rect 44352 30967 44720 30976
rect 48352 31016 48720 31025
rect 48392 30976 48434 31016
rect 48474 30976 48516 31016
rect 48556 30976 48598 31016
rect 48638 30976 48680 31016
rect 48352 30967 48720 30976
rect 52352 31016 52720 31025
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52352 30967 52720 30976
rect 56352 31016 56720 31025
rect 56392 30976 56434 31016
rect 56474 30976 56516 31016
rect 56556 30976 56598 31016
rect 56638 30976 56680 31016
rect 56352 30967 56720 30976
rect 60352 31016 60720 31025
rect 60392 30976 60434 31016
rect 60474 30976 60516 31016
rect 60556 30976 60598 31016
rect 60638 30976 60680 31016
rect 60352 30967 60720 30976
rect 64352 31016 64720 31025
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64352 30967 64720 30976
rect 67276 30596 67316 31219
rect 67564 30848 67604 30857
rect 67660 30848 67700 31471
rect 68812 31470 68852 31555
rect 68620 31436 68660 31445
rect 67604 30808 67700 30848
rect 67756 31352 67796 31361
rect 67564 30799 67604 30808
rect 67756 30689 67796 31312
rect 68620 31277 68660 31396
rect 68619 31268 68661 31277
rect 68619 31228 68620 31268
rect 68660 31228 68661 31268
rect 68619 31219 68661 31228
rect 68352 31016 68720 31025
rect 68392 30976 68434 31016
rect 68474 30976 68516 31016
rect 68556 30976 68598 31016
rect 68638 30976 68680 31016
rect 68352 30967 68720 30976
rect 68620 30848 68660 30857
rect 68908 30848 68948 31807
rect 69483 31772 69525 31781
rect 69483 31732 69484 31772
rect 69524 31732 69525 31772
rect 69483 31723 69525 31732
rect 69195 31520 69237 31529
rect 69195 31480 69196 31520
rect 69236 31480 69237 31520
rect 69195 31471 69237 31480
rect 68660 30808 68948 30848
rect 69004 31436 69044 31445
rect 68620 30799 68660 30808
rect 68523 30764 68565 30773
rect 68523 30724 68524 30764
rect 68564 30724 68565 30764
rect 68523 30715 68565 30724
rect 67755 30680 67797 30689
rect 67755 30640 67756 30680
rect 67796 30640 67797 30680
rect 67755 30631 67797 30640
rect 68043 30680 68085 30689
rect 68043 30640 68044 30680
rect 68084 30640 68085 30680
rect 68043 30631 68085 30640
rect 68524 30680 68564 30715
rect 69004 30689 69044 31396
rect 69196 31386 69236 31471
rect 69388 31436 69428 31445
rect 69291 31268 69333 31277
rect 69291 31228 69292 31268
rect 69332 31228 69333 31268
rect 69291 31219 69333 31228
rect 69099 30848 69141 30857
rect 69099 30808 69100 30848
rect 69140 30808 69141 30848
rect 69099 30799 69141 30808
rect 69100 30714 69140 30799
rect 69292 30773 69332 31219
rect 69388 31193 69428 31396
rect 69387 31184 69429 31193
rect 69387 31144 69388 31184
rect 69428 31144 69429 31184
rect 69387 31135 69429 31144
rect 69388 30848 69428 30857
rect 69484 30848 69524 31723
rect 69579 31520 69621 31529
rect 69579 31480 69580 31520
rect 69620 31480 69621 31520
rect 69579 31471 69621 31480
rect 69580 31386 69620 31471
rect 69675 31352 69717 31361
rect 69675 31312 69676 31352
rect 69716 31312 69717 31352
rect 69675 31303 69717 31312
rect 69772 31352 69812 32152
rect 69867 31940 69909 31949
rect 69867 31900 69868 31940
rect 69908 31900 69909 31940
rect 69867 31891 69909 31900
rect 69868 31806 69908 31891
rect 69867 31604 69909 31613
rect 69867 31564 69868 31604
rect 69908 31564 69909 31604
rect 69867 31555 69909 31564
rect 69868 31470 69908 31555
rect 69579 31184 69621 31193
rect 69579 31144 69580 31184
rect 69620 31144 69621 31184
rect 69579 31135 69621 31144
rect 69428 30808 69524 30848
rect 69388 30799 69428 30808
rect 69291 30764 69333 30773
rect 69291 30724 69292 30764
rect 69332 30724 69333 30764
rect 69291 30715 69333 30724
rect 67372 30596 67412 30605
rect 67276 30556 67372 30596
rect 67372 30547 67412 30556
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 7112 30260 7480 30269
rect 7152 30220 7194 30260
rect 7234 30220 7276 30260
rect 7316 30220 7358 30260
rect 7398 30220 7440 30260
rect 7112 30211 7480 30220
rect 11112 30260 11480 30269
rect 11152 30220 11194 30260
rect 11234 30220 11276 30260
rect 11316 30220 11358 30260
rect 11398 30220 11440 30260
rect 11112 30211 11480 30220
rect 15112 30260 15480 30269
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15112 30211 15480 30220
rect 19112 30260 19480 30269
rect 19152 30220 19194 30260
rect 19234 30220 19276 30260
rect 19316 30220 19358 30260
rect 19398 30220 19440 30260
rect 19112 30211 19480 30220
rect 23112 30260 23480 30269
rect 23152 30220 23194 30260
rect 23234 30220 23276 30260
rect 23316 30220 23358 30260
rect 23398 30220 23440 30260
rect 23112 30211 23480 30220
rect 27112 30260 27480 30269
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27112 30211 27480 30220
rect 31112 30260 31480 30269
rect 31152 30220 31194 30260
rect 31234 30220 31276 30260
rect 31316 30220 31358 30260
rect 31398 30220 31440 30260
rect 31112 30211 31480 30220
rect 35112 30260 35480 30269
rect 35152 30220 35194 30260
rect 35234 30220 35276 30260
rect 35316 30220 35358 30260
rect 35398 30220 35440 30260
rect 35112 30211 35480 30220
rect 39112 30260 39480 30269
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39112 30211 39480 30220
rect 43112 30260 43480 30269
rect 43152 30220 43194 30260
rect 43234 30220 43276 30260
rect 43316 30220 43358 30260
rect 43398 30220 43440 30260
rect 43112 30211 43480 30220
rect 47112 30260 47480 30269
rect 47152 30220 47194 30260
rect 47234 30220 47276 30260
rect 47316 30220 47358 30260
rect 47398 30220 47440 30260
rect 47112 30211 47480 30220
rect 51112 30260 51480 30269
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51112 30211 51480 30220
rect 55112 30260 55480 30269
rect 55152 30220 55194 30260
rect 55234 30220 55276 30260
rect 55316 30220 55358 30260
rect 55398 30220 55440 30260
rect 55112 30211 55480 30220
rect 59112 30260 59480 30269
rect 59152 30220 59194 30260
rect 59234 30220 59276 30260
rect 59316 30220 59358 30260
rect 59398 30220 59440 30260
rect 59112 30211 59480 30220
rect 63112 30260 63480 30269
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63112 30211 63480 30220
rect 67112 30260 67480 30269
rect 67152 30220 67194 30260
rect 67234 30220 67276 30260
rect 67316 30220 67358 30260
rect 67398 30220 67440 30260
rect 67112 30211 67480 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 8352 29504 8720 29513
rect 8392 29464 8434 29504
rect 8474 29464 8516 29504
rect 8556 29464 8598 29504
rect 8638 29464 8680 29504
rect 8352 29455 8720 29464
rect 12352 29504 12720 29513
rect 12392 29464 12434 29504
rect 12474 29464 12516 29504
rect 12556 29464 12598 29504
rect 12638 29464 12680 29504
rect 12352 29455 12720 29464
rect 16352 29504 16720 29513
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16352 29455 16720 29464
rect 20352 29504 20720 29513
rect 20392 29464 20434 29504
rect 20474 29464 20516 29504
rect 20556 29464 20598 29504
rect 20638 29464 20680 29504
rect 20352 29455 20720 29464
rect 24352 29504 24720 29513
rect 24392 29464 24434 29504
rect 24474 29464 24516 29504
rect 24556 29464 24598 29504
rect 24638 29464 24680 29504
rect 24352 29455 24720 29464
rect 28352 29504 28720 29513
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28352 29455 28720 29464
rect 32352 29504 32720 29513
rect 32392 29464 32434 29504
rect 32474 29464 32516 29504
rect 32556 29464 32598 29504
rect 32638 29464 32680 29504
rect 32352 29455 32720 29464
rect 36352 29504 36720 29513
rect 36392 29464 36434 29504
rect 36474 29464 36516 29504
rect 36556 29464 36598 29504
rect 36638 29464 36680 29504
rect 36352 29455 36720 29464
rect 40352 29504 40720 29513
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40352 29455 40720 29464
rect 44352 29504 44720 29513
rect 44392 29464 44434 29504
rect 44474 29464 44516 29504
rect 44556 29464 44598 29504
rect 44638 29464 44680 29504
rect 44352 29455 44720 29464
rect 48352 29504 48720 29513
rect 48392 29464 48434 29504
rect 48474 29464 48516 29504
rect 48556 29464 48598 29504
rect 48638 29464 48680 29504
rect 48352 29455 48720 29464
rect 52352 29504 52720 29513
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52352 29455 52720 29464
rect 56352 29504 56720 29513
rect 56392 29464 56434 29504
rect 56474 29464 56516 29504
rect 56556 29464 56598 29504
rect 56638 29464 56680 29504
rect 56352 29455 56720 29464
rect 60352 29504 60720 29513
rect 60392 29464 60434 29504
rect 60474 29464 60516 29504
rect 60556 29464 60598 29504
rect 60638 29464 60680 29504
rect 60352 29455 60720 29464
rect 64352 29504 64720 29513
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64352 29455 64720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 7112 28748 7480 28757
rect 7152 28708 7194 28748
rect 7234 28708 7276 28748
rect 7316 28708 7358 28748
rect 7398 28708 7440 28748
rect 7112 28699 7480 28708
rect 11112 28748 11480 28757
rect 11152 28708 11194 28748
rect 11234 28708 11276 28748
rect 11316 28708 11358 28748
rect 11398 28708 11440 28748
rect 11112 28699 11480 28708
rect 15112 28748 15480 28757
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15112 28699 15480 28708
rect 19112 28748 19480 28757
rect 19152 28708 19194 28748
rect 19234 28708 19276 28748
rect 19316 28708 19358 28748
rect 19398 28708 19440 28748
rect 19112 28699 19480 28708
rect 23112 28748 23480 28757
rect 23152 28708 23194 28748
rect 23234 28708 23276 28748
rect 23316 28708 23358 28748
rect 23398 28708 23440 28748
rect 23112 28699 23480 28708
rect 27112 28748 27480 28757
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27112 28699 27480 28708
rect 31112 28748 31480 28757
rect 31152 28708 31194 28748
rect 31234 28708 31276 28748
rect 31316 28708 31358 28748
rect 31398 28708 31440 28748
rect 31112 28699 31480 28708
rect 35112 28748 35480 28757
rect 35152 28708 35194 28748
rect 35234 28708 35276 28748
rect 35316 28708 35358 28748
rect 35398 28708 35440 28748
rect 35112 28699 35480 28708
rect 39112 28748 39480 28757
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39112 28699 39480 28708
rect 43112 28748 43480 28757
rect 43152 28708 43194 28748
rect 43234 28708 43276 28748
rect 43316 28708 43358 28748
rect 43398 28708 43440 28748
rect 43112 28699 43480 28708
rect 47112 28748 47480 28757
rect 47152 28708 47194 28748
rect 47234 28708 47276 28748
rect 47316 28708 47358 28748
rect 47398 28708 47440 28748
rect 47112 28699 47480 28708
rect 51112 28748 51480 28757
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51112 28699 51480 28708
rect 55112 28748 55480 28757
rect 55152 28708 55194 28748
rect 55234 28708 55276 28748
rect 55316 28708 55358 28748
rect 55398 28708 55440 28748
rect 55112 28699 55480 28708
rect 59112 28748 59480 28757
rect 59152 28708 59194 28748
rect 59234 28708 59276 28748
rect 59316 28708 59358 28748
rect 59398 28708 59440 28748
rect 59112 28699 59480 28708
rect 63112 28748 63480 28757
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63112 28699 63480 28708
rect 67112 28748 67480 28757
rect 67152 28708 67194 28748
rect 67234 28708 67276 28748
rect 67316 28708 67358 28748
rect 67398 28708 67440 28748
rect 67112 28699 67480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 8352 27992 8720 28001
rect 8392 27952 8434 27992
rect 8474 27952 8516 27992
rect 8556 27952 8598 27992
rect 8638 27952 8680 27992
rect 8352 27943 8720 27952
rect 12352 27992 12720 28001
rect 12392 27952 12434 27992
rect 12474 27952 12516 27992
rect 12556 27952 12598 27992
rect 12638 27952 12680 27992
rect 12352 27943 12720 27952
rect 16352 27992 16720 28001
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16352 27943 16720 27952
rect 20352 27992 20720 28001
rect 20392 27952 20434 27992
rect 20474 27952 20516 27992
rect 20556 27952 20598 27992
rect 20638 27952 20680 27992
rect 20352 27943 20720 27952
rect 24352 27992 24720 28001
rect 24392 27952 24434 27992
rect 24474 27952 24516 27992
rect 24556 27952 24598 27992
rect 24638 27952 24680 27992
rect 24352 27943 24720 27952
rect 28352 27992 28720 28001
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28352 27943 28720 27952
rect 32352 27992 32720 28001
rect 32392 27952 32434 27992
rect 32474 27952 32516 27992
rect 32556 27952 32598 27992
rect 32638 27952 32680 27992
rect 32352 27943 32720 27952
rect 36352 27992 36720 28001
rect 36392 27952 36434 27992
rect 36474 27952 36516 27992
rect 36556 27952 36598 27992
rect 36638 27952 36680 27992
rect 36352 27943 36720 27952
rect 40352 27992 40720 28001
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40352 27943 40720 27952
rect 44352 27992 44720 28001
rect 44392 27952 44434 27992
rect 44474 27952 44516 27992
rect 44556 27952 44598 27992
rect 44638 27952 44680 27992
rect 44352 27943 44720 27952
rect 48352 27992 48720 28001
rect 48392 27952 48434 27992
rect 48474 27952 48516 27992
rect 48556 27952 48598 27992
rect 48638 27952 48680 27992
rect 48352 27943 48720 27952
rect 52352 27992 52720 28001
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52352 27943 52720 27952
rect 56352 27992 56720 28001
rect 56392 27952 56434 27992
rect 56474 27952 56516 27992
rect 56556 27952 56598 27992
rect 56638 27952 56680 27992
rect 56352 27943 56720 27952
rect 60352 27992 60720 28001
rect 60392 27952 60434 27992
rect 60474 27952 60516 27992
rect 60556 27952 60598 27992
rect 60638 27952 60680 27992
rect 60352 27943 60720 27952
rect 64352 27992 64720 28001
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64352 27943 64720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 7112 27236 7480 27245
rect 7152 27196 7194 27236
rect 7234 27196 7276 27236
rect 7316 27196 7358 27236
rect 7398 27196 7440 27236
rect 7112 27187 7480 27196
rect 11112 27236 11480 27245
rect 11152 27196 11194 27236
rect 11234 27196 11276 27236
rect 11316 27196 11358 27236
rect 11398 27196 11440 27236
rect 11112 27187 11480 27196
rect 15112 27236 15480 27245
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15112 27187 15480 27196
rect 19112 27236 19480 27245
rect 19152 27196 19194 27236
rect 19234 27196 19276 27236
rect 19316 27196 19358 27236
rect 19398 27196 19440 27236
rect 19112 27187 19480 27196
rect 23112 27236 23480 27245
rect 23152 27196 23194 27236
rect 23234 27196 23276 27236
rect 23316 27196 23358 27236
rect 23398 27196 23440 27236
rect 23112 27187 23480 27196
rect 27112 27236 27480 27245
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27112 27187 27480 27196
rect 31112 27236 31480 27245
rect 31152 27196 31194 27236
rect 31234 27196 31276 27236
rect 31316 27196 31358 27236
rect 31398 27196 31440 27236
rect 31112 27187 31480 27196
rect 35112 27236 35480 27245
rect 35152 27196 35194 27236
rect 35234 27196 35276 27236
rect 35316 27196 35358 27236
rect 35398 27196 35440 27236
rect 35112 27187 35480 27196
rect 39112 27236 39480 27245
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39112 27187 39480 27196
rect 43112 27236 43480 27245
rect 43152 27196 43194 27236
rect 43234 27196 43276 27236
rect 43316 27196 43358 27236
rect 43398 27196 43440 27236
rect 43112 27187 43480 27196
rect 47112 27236 47480 27245
rect 47152 27196 47194 27236
rect 47234 27196 47276 27236
rect 47316 27196 47358 27236
rect 47398 27196 47440 27236
rect 47112 27187 47480 27196
rect 51112 27236 51480 27245
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51112 27187 51480 27196
rect 55112 27236 55480 27245
rect 55152 27196 55194 27236
rect 55234 27196 55276 27236
rect 55316 27196 55358 27236
rect 55398 27196 55440 27236
rect 55112 27187 55480 27196
rect 59112 27236 59480 27245
rect 59152 27196 59194 27236
rect 59234 27196 59276 27236
rect 59316 27196 59358 27236
rect 59398 27196 59440 27236
rect 59112 27187 59480 27196
rect 63112 27236 63480 27245
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63112 27187 63480 27196
rect 67112 27236 67480 27245
rect 67152 27196 67194 27236
rect 67234 27196 67276 27236
rect 67316 27196 67358 27236
rect 67398 27196 67440 27236
rect 67112 27187 67480 27196
rect 68044 26984 68084 30631
rect 68524 30629 68564 30640
rect 69003 30680 69045 30689
rect 69003 30640 69004 30680
rect 69044 30640 69045 30680
rect 69003 30631 69045 30640
rect 69292 30680 69332 30715
rect 69004 30546 69044 30631
rect 69292 30630 69332 30640
rect 69580 30680 69620 31135
rect 69676 30848 69716 31303
rect 69772 31277 69812 31312
rect 69771 31268 69813 31277
rect 69771 31228 69772 31268
rect 69812 31228 69813 31268
rect 69771 31219 69813 31228
rect 69772 31188 69812 31219
rect 69676 30799 69716 30808
rect 68352 29504 68720 29513
rect 68392 29464 68434 29504
rect 68474 29464 68516 29504
rect 68556 29464 68598 29504
rect 68638 29464 68680 29504
rect 68352 29455 68720 29464
rect 68352 27992 68720 28001
rect 68392 27952 68434 27992
rect 68474 27952 68516 27992
rect 68556 27952 68598 27992
rect 68638 27952 68680 27992
rect 68352 27943 68720 27952
rect 68812 27572 68852 27581
rect 68140 26984 68180 26993
rect 67948 26944 68140 26984
rect 67948 26900 67988 26944
rect 68140 26935 68180 26944
rect 68332 26900 68372 26909
rect 67948 26851 67988 26860
rect 68236 26860 68332 26900
rect 67756 26648 67796 26657
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 8352 26480 8720 26489
rect 8392 26440 8434 26480
rect 8474 26440 8516 26480
rect 8556 26440 8598 26480
rect 8638 26440 8680 26480
rect 8352 26431 8720 26440
rect 12352 26480 12720 26489
rect 12392 26440 12434 26480
rect 12474 26440 12516 26480
rect 12556 26440 12598 26480
rect 12638 26440 12680 26480
rect 12352 26431 12720 26440
rect 16352 26480 16720 26489
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16352 26431 16720 26440
rect 20352 26480 20720 26489
rect 20392 26440 20434 26480
rect 20474 26440 20516 26480
rect 20556 26440 20598 26480
rect 20638 26440 20680 26480
rect 20352 26431 20720 26440
rect 24352 26480 24720 26489
rect 24392 26440 24434 26480
rect 24474 26440 24516 26480
rect 24556 26440 24598 26480
rect 24638 26440 24680 26480
rect 24352 26431 24720 26440
rect 28352 26480 28720 26489
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28352 26431 28720 26440
rect 32352 26480 32720 26489
rect 32392 26440 32434 26480
rect 32474 26440 32516 26480
rect 32556 26440 32598 26480
rect 32638 26440 32680 26480
rect 32352 26431 32720 26440
rect 36352 26480 36720 26489
rect 36392 26440 36434 26480
rect 36474 26440 36516 26480
rect 36556 26440 36598 26480
rect 36638 26440 36680 26480
rect 36352 26431 36720 26440
rect 40352 26480 40720 26489
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40352 26431 40720 26440
rect 44352 26480 44720 26489
rect 44392 26440 44434 26480
rect 44474 26440 44516 26480
rect 44556 26440 44598 26480
rect 44638 26440 44680 26480
rect 44352 26431 44720 26440
rect 48352 26480 48720 26489
rect 48392 26440 48434 26480
rect 48474 26440 48516 26480
rect 48556 26440 48598 26480
rect 48638 26440 48680 26480
rect 48352 26431 48720 26440
rect 52352 26480 52720 26489
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52352 26431 52720 26440
rect 56352 26480 56720 26489
rect 56392 26440 56434 26480
rect 56474 26440 56516 26480
rect 56556 26440 56598 26480
rect 56638 26440 56680 26480
rect 56352 26431 56720 26440
rect 60352 26480 60720 26489
rect 60392 26440 60434 26480
rect 60474 26440 60516 26480
rect 60556 26440 60598 26480
rect 60638 26440 60680 26480
rect 60352 26431 60720 26440
rect 64352 26480 64720 26489
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64352 26431 64720 26440
rect 67564 26144 67604 26153
rect 67564 26060 67604 26104
rect 67756 26060 67796 26608
rect 67564 26020 67756 26060
rect 67468 25892 67508 25901
rect 67508 25852 67604 25892
rect 67468 25843 67508 25852
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 7112 25724 7480 25733
rect 7152 25684 7194 25724
rect 7234 25684 7276 25724
rect 7316 25684 7358 25724
rect 7398 25684 7440 25724
rect 7112 25675 7480 25684
rect 11112 25724 11480 25733
rect 11152 25684 11194 25724
rect 11234 25684 11276 25724
rect 11316 25684 11358 25724
rect 11398 25684 11440 25724
rect 11112 25675 11480 25684
rect 15112 25724 15480 25733
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15112 25675 15480 25684
rect 19112 25724 19480 25733
rect 19152 25684 19194 25724
rect 19234 25684 19276 25724
rect 19316 25684 19358 25724
rect 19398 25684 19440 25724
rect 19112 25675 19480 25684
rect 23112 25724 23480 25733
rect 23152 25684 23194 25724
rect 23234 25684 23276 25724
rect 23316 25684 23358 25724
rect 23398 25684 23440 25724
rect 23112 25675 23480 25684
rect 27112 25724 27480 25733
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27112 25675 27480 25684
rect 31112 25724 31480 25733
rect 31152 25684 31194 25724
rect 31234 25684 31276 25724
rect 31316 25684 31358 25724
rect 31398 25684 31440 25724
rect 31112 25675 31480 25684
rect 35112 25724 35480 25733
rect 35152 25684 35194 25724
rect 35234 25684 35276 25724
rect 35316 25684 35358 25724
rect 35398 25684 35440 25724
rect 35112 25675 35480 25684
rect 39112 25724 39480 25733
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39112 25675 39480 25684
rect 43112 25724 43480 25733
rect 43152 25684 43194 25724
rect 43234 25684 43276 25724
rect 43316 25684 43358 25724
rect 43398 25684 43440 25724
rect 43112 25675 43480 25684
rect 47112 25724 47480 25733
rect 47152 25684 47194 25724
rect 47234 25684 47276 25724
rect 47316 25684 47358 25724
rect 47398 25684 47440 25724
rect 47112 25675 47480 25684
rect 51112 25724 51480 25733
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51112 25675 51480 25684
rect 55112 25724 55480 25733
rect 55152 25684 55194 25724
rect 55234 25684 55276 25724
rect 55316 25684 55358 25724
rect 55398 25684 55440 25724
rect 55112 25675 55480 25684
rect 59112 25724 59480 25733
rect 59152 25684 59194 25724
rect 59234 25684 59276 25724
rect 59316 25684 59358 25724
rect 59398 25684 59440 25724
rect 59112 25675 59480 25684
rect 63112 25724 63480 25733
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63112 25675 63480 25684
rect 67112 25724 67480 25733
rect 67152 25684 67194 25724
rect 67234 25684 67276 25724
rect 67316 25684 67358 25724
rect 67398 25684 67440 25724
rect 67112 25675 67480 25684
rect 652 25304 692 25313
rect 652 24977 692 25264
rect 843 25304 885 25313
rect 843 25264 844 25304
rect 884 25264 885 25304
rect 843 25255 885 25264
rect 844 25170 884 25255
rect 651 24968 693 24977
rect 651 24928 652 24968
rect 692 24928 693 24968
rect 651 24919 693 24928
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 8352 24968 8720 24977
rect 8392 24928 8434 24968
rect 8474 24928 8516 24968
rect 8556 24928 8598 24968
rect 8638 24928 8680 24968
rect 8352 24919 8720 24928
rect 12352 24968 12720 24977
rect 12392 24928 12434 24968
rect 12474 24928 12516 24968
rect 12556 24928 12598 24968
rect 12638 24928 12680 24968
rect 12352 24919 12720 24928
rect 16352 24968 16720 24977
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16352 24919 16720 24928
rect 20352 24968 20720 24977
rect 20392 24928 20434 24968
rect 20474 24928 20516 24968
rect 20556 24928 20598 24968
rect 20638 24928 20680 24968
rect 20352 24919 20720 24928
rect 24352 24968 24720 24977
rect 24392 24928 24434 24968
rect 24474 24928 24516 24968
rect 24556 24928 24598 24968
rect 24638 24928 24680 24968
rect 24352 24919 24720 24928
rect 28352 24968 28720 24977
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28352 24919 28720 24928
rect 32352 24968 32720 24977
rect 32392 24928 32434 24968
rect 32474 24928 32516 24968
rect 32556 24928 32598 24968
rect 32638 24928 32680 24968
rect 32352 24919 32720 24928
rect 36352 24968 36720 24977
rect 36392 24928 36434 24968
rect 36474 24928 36516 24968
rect 36556 24928 36598 24968
rect 36638 24928 36680 24968
rect 36352 24919 36720 24928
rect 40352 24968 40720 24977
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40352 24919 40720 24928
rect 44352 24968 44720 24977
rect 44392 24928 44434 24968
rect 44474 24928 44516 24968
rect 44556 24928 44598 24968
rect 44638 24928 44680 24968
rect 44352 24919 44720 24928
rect 48352 24968 48720 24977
rect 48392 24928 48434 24968
rect 48474 24928 48516 24968
rect 48556 24928 48598 24968
rect 48638 24928 48680 24968
rect 48352 24919 48720 24928
rect 52352 24968 52720 24977
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52352 24919 52720 24928
rect 56352 24968 56720 24977
rect 56392 24928 56434 24968
rect 56474 24928 56516 24968
rect 56556 24928 56598 24968
rect 56638 24928 56680 24968
rect 56352 24919 56720 24928
rect 60352 24968 60720 24977
rect 60392 24928 60434 24968
rect 60474 24928 60516 24968
rect 60556 24928 60598 24968
rect 60638 24928 60680 24968
rect 60352 24919 60720 24928
rect 64352 24968 64720 24977
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64352 24919 64720 24928
rect 67564 24893 67604 25852
rect 67756 25313 67796 26020
rect 67948 25892 67988 25901
rect 67948 25649 67988 25852
rect 67947 25640 67989 25649
rect 67947 25600 67948 25640
rect 67988 25600 67989 25640
rect 67947 25591 67989 25600
rect 67755 25304 67797 25313
rect 67755 25264 67756 25304
rect 67796 25264 67797 25304
rect 67755 25255 67797 25264
rect 67563 24884 67605 24893
rect 67563 24844 67564 24884
rect 67604 24844 67605 24884
rect 67563 24835 67605 24844
rect 652 24632 692 24641
rect 652 24137 692 24592
rect 844 24632 884 24641
rect 651 24128 693 24137
rect 651 24088 652 24128
rect 692 24088 693 24128
rect 651 24079 693 24088
rect 844 23960 884 24592
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 7112 24212 7480 24221
rect 7152 24172 7194 24212
rect 7234 24172 7276 24212
rect 7316 24172 7358 24212
rect 7398 24172 7440 24212
rect 7112 24163 7480 24172
rect 11112 24212 11480 24221
rect 11152 24172 11194 24212
rect 11234 24172 11276 24212
rect 11316 24172 11358 24212
rect 11398 24172 11440 24212
rect 11112 24163 11480 24172
rect 15112 24212 15480 24221
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15112 24163 15480 24172
rect 19112 24212 19480 24221
rect 19152 24172 19194 24212
rect 19234 24172 19276 24212
rect 19316 24172 19358 24212
rect 19398 24172 19440 24212
rect 19112 24163 19480 24172
rect 23112 24212 23480 24221
rect 23152 24172 23194 24212
rect 23234 24172 23276 24212
rect 23316 24172 23358 24212
rect 23398 24172 23440 24212
rect 23112 24163 23480 24172
rect 27112 24212 27480 24221
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27112 24163 27480 24172
rect 31112 24212 31480 24221
rect 31152 24172 31194 24212
rect 31234 24172 31276 24212
rect 31316 24172 31358 24212
rect 31398 24172 31440 24212
rect 31112 24163 31480 24172
rect 35112 24212 35480 24221
rect 35152 24172 35194 24212
rect 35234 24172 35276 24212
rect 35316 24172 35358 24212
rect 35398 24172 35440 24212
rect 35112 24163 35480 24172
rect 39112 24212 39480 24221
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39112 24163 39480 24172
rect 43112 24212 43480 24221
rect 43152 24172 43194 24212
rect 43234 24172 43276 24212
rect 43316 24172 43358 24212
rect 43398 24172 43440 24212
rect 43112 24163 43480 24172
rect 47112 24212 47480 24221
rect 47152 24172 47194 24212
rect 47234 24172 47276 24212
rect 47316 24172 47358 24212
rect 47398 24172 47440 24212
rect 47112 24163 47480 24172
rect 51112 24212 51480 24221
rect 51152 24172 51194 24212
rect 51234 24172 51276 24212
rect 51316 24172 51358 24212
rect 51398 24172 51440 24212
rect 51112 24163 51480 24172
rect 55112 24212 55480 24221
rect 55152 24172 55194 24212
rect 55234 24172 55276 24212
rect 55316 24172 55358 24212
rect 55398 24172 55440 24212
rect 55112 24163 55480 24172
rect 59112 24212 59480 24221
rect 59152 24172 59194 24212
rect 59234 24172 59276 24212
rect 59316 24172 59358 24212
rect 59398 24172 59440 24212
rect 59112 24163 59480 24172
rect 63112 24212 63480 24221
rect 63152 24172 63194 24212
rect 63234 24172 63276 24212
rect 63316 24172 63358 24212
rect 63398 24172 63440 24212
rect 63112 24163 63480 24172
rect 67112 24212 67480 24221
rect 67152 24172 67194 24212
rect 67234 24172 67276 24212
rect 67316 24172 67358 24212
rect 67398 24172 67440 24212
rect 67112 24163 67480 24172
rect 844 23920 980 23960
rect 652 23792 692 23801
rect 652 23297 692 23752
rect 843 23792 885 23801
rect 843 23752 844 23792
rect 884 23752 885 23792
rect 843 23743 885 23752
rect 844 23658 884 23743
rect 651 23288 693 23297
rect 651 23248 652 23288
rect 692 23248 693 23288
rect 651 23239 693 23248
rect 652 23120 692 23129
rect 556 23080 652 23120
rect 556 22457 596 23080
rect 652 23071 692 23080
rect 843 23120 885 23129
rect 843 23080 844 23120
rect 884 23080 885 23120
rect 843 23071 885 23080
rect 844 22986 884 23071
rect 555 22448 597 22457
rect 555 22408 556 22448
rect 596 22408 597 22448
rect 555 22399 597 22408
rect 652 22448 692 22457
rect 652 21617 692 22408
rect 940 22037 980 23920
rect 2091 23792 2133 23801
rect 2091 23752 2092 23792
rect 2132 23752 2133 23792
rect 2091 23743 2133 23752
rect 2092 23297 2132 23743
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 8352 23456 8720 23465
rect 8392 23416 8434 23456
rect 8474 23416 8516 23456
rect 8556 23416 8598 23456
rect 8638 23416 8680 23456
rect 8352 23407 8720 23416
rect 12352 23456 12720 23465
rect 12392 23416 12434 23456
rect 12474 23416 12516 23456
rect 12556 23416 12598 23456
rect 12638 23416 12680 23456
rect 12352 23407 12720 23416
rect 16352 23456 16720 23465
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16352 23407 16720 23416
rect 20352 23456 20720 23465
rect 20392 23416 20434 23456
rect 20474 23416 20516 23456
rect 20556 23416 20598 23456
rect 20638 23416 20680 23456
rect 20352 23407 20720 23416
rect 24352 23456 24720 23465
rect 24392 23416 24434 23456
rect 24474 23416 24516 23456
rect 24556 23416 24598 23456
rect 24638 23416 24680 23456
rect 24352 23407 24720 23416
rect 28352 23456 28720 23465
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28352 23407 28720 23416
rect 32352 23456 32720 23465
rect 32392 23416 32434 23456
rect 32474 23416 32516 23456
rect 32556 23416 32598 23456
rect 32638 23416 32680 23456
rect 32352 23407 32720 23416
rect 36352 23456 36720 23465
rect 36392 23416 36434 23456
rect 36474 23416 36516 23456
rect 36556 23416 36598 23456
rect 36638 23416 36680 23456
rect 36352 23407 36720 23416
rect 40352 23456 40720 23465
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40352 23407 40720 23416
rect 44352 23456 44720 23465
rect 44392 23416 44434 23456
rect 44474 23416 44516 23456
rect 44556 23416 44598 23456
rect 44638 23416 44680 23456
rect 44352 23407 44720 23416
rect 48352 23456 48720 23465
rect 48392 23416 48434 23456
rect 48474 23416 48516 23456
rect 48556 23416 48598 23456
rect 48638 23416 48680 23456
rect 48352 23407 48720 23416
rect 52352 23456 52720 23465
rect 52392 23416 52434 23456
rect 52474 23416 52516 23456
rect 52556 23416 52598 23456
rect 52638 23416 52680 23456
rect 52352 23407 52720 23416
rect 56352 23456 56720 23465
rect 56392 23416 56434 23456
rect 56474 23416 56516 23456
rect 56556 23416 56598 23456
rect 56638 23416 56680 23456
rect 56352 23407 56720 23416
rect 60352 23456 60720 23465
rect 60392 23416 60434 23456
rect 60474 23416 60516 23456
rect 60556 23416 60598 23456
rect 60638 23416 60680 23456
rect 60352 23407 60720 23416
rect 64352 23456 64720 23465
rect 64392 23416 64434 23456
rect 64474 23416 64516 23456
rect 64556 23416 64598 23456
rect 64638 23416 64680 23456
rect 64352 23407 64720 23416
rect 68236 23297 68276 26860
rect 68332 26851 68372 26860
rect 68352 26480 68720 26489
rect 68392 26440 68434 26480
rect 68474 26440 68516 26480
rect 68556 26440 68598 26480
rect 68638 26440 68680 26480
rect 68352 26431 68720 26440
rect 68812 26153 68852 27532
rect 69004 27404 69044 27413
rect 68619 26144 68661 26153
rect 68619 26104 68620 26144
rect 68660 26104 68661 26144
rect 68619 26095 68661 26104
rect 68811 26144 68853 26153
rect 68811 26104 68812 26144
rect 68852 26104 68853 26144
rect 68811 26095 68853 26104
rect 68331 26060 68373 26069
rect 68331 26020 68332 26060
rect 68372 26020 68373 26060
rect 68331 26011 68373 26020
rect 68332 25397 68372 26011
rect 68620 26010 68660 26095
rect 68811 25976 68853 25985
rect 68811 25936 68812 25976
rect 68852 25936 68853 25976
rect 68811 25927 68853 25936
rect 68524 25892 68564 25901
rect 68524 25649 68564 25852
rect 68523 25640 68565 25649
rect 68523 25600 68524 25640
rect 68564 25600 68565 25640
rect 68523 25591 68565 25600
rect 68812 25556 68852 25927
rect 68812 25507 68852 25516
rect 68908 25892 68948 25901
rect 68331 25388 68373 25397
rect 68331 25348 68332 25388
rect 68372 25348 68373 25388
rect 68331 25339 68373 25348
rect 68620 25388 68660 25399
rect 68620 25313 68660 25348
rect 68619 25304 68661 25313
rect 68619 25264 68620 25304
rect 68660 25264 68661 25304
rect 68619 25255 68661 25264
rect 68908 25145 68948 25852
rect 69004 25733 69044 27364
rect 69484 26900 69524 26909
rect 69100 26144 69140 26155
rect 69484 26153 69524 26860
rect 69100 26069 69140 26104
rect 69291 26144 69333 26153
rect 69291 26104 69292 26144
rect 69332 26104 69333 26144
rect 69291 26095 69333 26104
rect 69483 26144 69525 26153
rect 69483 26104 69484 26144
rect 69524 26104 69525 26144
rect 69483 26095 69525 26104
rect 69099 26060 69141 26069
rect 69099 26020 69100 26060
rect 69140 26020 69141 26060
rect 69099 26011 69141 26020
rect 69196 25892 69236 25903
rect 69196 25817 69236 25852
rect 69195 25808 69237 25817
rect 69195 25768 69196 25808
rect 69236 25768 69237 25808
rect 69195 25759 69237 25768
rect 69003 25724 69045 25733
rect 69003 25684 69004 25724
rect 69044 25684 69045 25724
rect 69003 25675 69045 25684
rect 69292 25304 69332 26095
rect 69580 26069 69620 30640
rect 69676 26648 69716 26657
rect 69387 26060 69429 26069
rect 69387 26020 69388 26060
rect 69428 26020 69429 26060
rect 69387 26011 69429 26020
rect 69579 26060 69621 26069
rect 69579 26020 69580 26060
rect 69620 26020 69621 26060
rect 69579 26011 69621 26020
rect 69388 25926 69428 26011
rect 69579 25892 69621 25901
rect 69579 25852 69580 25892
rect 69620 25852 69621 25892
rect 69579 25843 69621 25852
rect 69580 25758 69620 25843
rect 69676 25556 69716 26608
rect 69771 26144 69813 26153
rect 69771 26104 69772 26144
rect 69812 26104 69813 26144
rect 69771 26095 69813 26104
rect 69772 26010 69812 26095
rect 69868 25892 69908 25901
rect 69908 25852 70004 25892
rect 69868 25843 69908 25852
rect 69867 25556 69909 25565
rect 69676 25516 69812 25556
rect 69676 25388 69716 25397
rect 68907 25136 68949 25145
rect 68907 25096 68908 25136
rect 68948 25096 68949 25136
rect 68907 25087 68949 25096
rect 69292 25061 69332 25264
rect 69483 25304 69525 25313
rect 69483 25264 69484 25304
rect 69524 25264 69525 25304
rect 69483 25255 69525 25264
rect 69484 25170 69524 25255
rect 69676 25061 69716 25348
rect 69772 25229 69812 25516
rect 69867 25516 69868 25556
rect 69908 25516 69909 25556
rect 69867 25507 69909 25516
rect 69868 25422 69908 25507
rect 69964 25481 70004 25852
rect 69963 25472 70005 25481
rect 69963 25432 69964 25472
rect 70004 25432 70005 25472
rect 69963 25423 70005 25432
rect 69771 25220 69813 25229
rect 69771 25180 69772 25220
rect 69812 25180 69813 25220
rect 69771 25171 69813 25180
rect 69291 25052 69333 25061
rect 69291 25012 69292 25052
rect 69332 25012 69333 25052
rect 69291 25003 69333 25012
rect 69675 25052 69717 25061
rect 69675 25012 69676 25052
rect 69716 25012 69717 25052
rect 69675 25003 69717 25012
rect 68352 24968 68720 24977
rect 68392 24928 68434 24968
rect 68474 24928 68516 24968
rect 68556 24928 68598 24968
rect 68638 24928 68680 24968
rect 68352 24919 68720 24928
rect 68352 23456 68720 23465
rect 68392 23416 68434 23456
rect 68474 23416 68516 23456
rect 68556 23416 68598 23456
rect 68638 23416 68680 23456
rect 68352 23407 68720 23416
rect 71788 23381 71828 32731
rect 73899 32108 73941 32117
rect 73899 32068 73900 32108
rect 73940 32068 73941 32108
rect 73899 32059 73941 32068
rect 73611 32024 73653 32033
rect 73611 31984 73612 32024
rect 73652 31984 73653 32024
rect 73611 31975 73653 31984
rect 73227 31772 73269 31781
rect 73132 31732 73228 31772
rect 73268 31732 73269 31772
rect 73132 31688 73172 31732
rect 73227 31723 73269 31732
rect 72268 31648 72596 31688
rect 72268 31520 72308 31648
rect 71884 31480 72308 31520
rect 72414 31520 72456 31529
rect 72414 31480 72415 31520
rect 72455 31480 72456 31520
rect 72556 31520 72596 31648
rect 73105 31648 73172 31688
rect 73612 31688 73652 31975
rect 73900 31688 73940 32059
rect 73996 31688 74036 34168
rect 74132 34168 74228 34208
rect 74092 34159 74132 34168
rect 74188 32780 74228 34168
rect 74284 32957 74324 34924
rect 74476 34914 74516 34999
rect 74667 34628 74709 34637
rect 74667 34588 74668 34628
rect 74708 34588 74709 34628
rect 74667 34579 74709 34588
rect 74668 34460 74708 34579
rect 74475 34292 74517 34301
rect 74475 34252 74476 34292
rect 74516 34252 74517 34292
rect 74475 34243 74517 34252
rect 74476 34208 74516 34243
rect 74476 34157 74516 34168
rect 74283 32948 74325 32957
rect 74283 32908 74284 32948
rect 74324 32908 74325 32948
rect 74283 32899 74325 32908
rect 74668 32789 74708 34420
rect 74764 34292 74804 35092
rect 74859 35092 74860 35132
rect 74900 35092 74901 35132
rect 74859 35083 74901 35092
rect 74860 34553 74900 35083
rect 74859 34544 74901 34553
rect 74859 34504 74860 34544
rect 74900 34504 74901 34544
rect 74859 34495 74901 34504
rect 74857 34365 74897 34384
rect 74956 34376 74996 35680
rect 75052 35671 75092 35680
rect 76779 35720 76821 35729
rect 76779 35680 76780 35720
rect 76820 35680 76821 35720
rect 76779 35671 76821 35680
rect 76780 35586 76820 35671
rect 76352 35552 76720 35561
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76352 35503 76720 35512
rect 76876 35468 76916 35848
rect 76780 35428 76916 35468
rect 76108 35216 76148 35227
rect 76108 35141 76148 35176
rect 76203 35216 76245 35225
rect 76203 35176 76204 35216
rect 76244 35176 76245 35216
rect 76203 35167 76245 35176
rect 76683 35216 76725 35225
rect 76780 35216 76820 35428
rect 77548 35225 77588 35932
rect 78508 35932 78604 35972
rect 78644 35932 79372 35972
rect 77644 35720 77684 35729
rect 76683 35176 76684 35216
rect 76724 35176 76820 35216
rect 77259 35216 77301 35225
rect 77259 35176 77260 35216
rect 77300 35176 77301 35216
rect 76683 35167 76725 35176
rect 77259 35167 77301 35176
rect 77547 35216 77589 35225
rect 77547 35176 77548 35216
rect 77588 35176 77589 35216
rect 77547 35167 77589 35176
rect 75627 35132 75669 35141
rect 75627 35092 75628 35132
rect 75668 35092 75669 35132
rect 75627 35083 75669 35092
rect 76107 35132 76149 35141
rect 76107 35092 76108 35132
rect 76148 35092 76149 35132
rect 76107 35083 76149 35092
rect 75628 34998 75668 35083
rect 75820 34964 75860 34973
rect 76012 34964 76052 34973
rect 75724 34924 75820 34964
rect 75112 34796 75480 34805
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75112 34747 75480 34756
rect 75148 34469 75188 34554
rect 75147 34460 75189 34469
rect 75147 34420 75148 34460
rect 75188 34420 75189 34460
rect 75147 34411 75189 34420
rect 75627 34376 75669 34385
rect 74956 34336 75092 34376
rect 74857 34301 74897 34325
rect 74857 34292 74901 34301
rect 74764 34252 74860 34292
rect 74900 34252 74901 34292
rect 75052 34292 75092 34336
rect 75627 34336 75628 34376
rect 75668 34336 75669 34376
rect 75627 34327 75669 34336
rect 75052 34252 75188 34292
rect 74859 34243 74901 34252
rect 74956 34208 74996 34217
rect 74996 34168 75092 34208
rect 74956 34159 74996 34168
rect 74763 32948 74805 32957
rect 74763 32908 74764 32948
rect 74804 32908 74805 32948
rect 74763 32899 74805 32908
rect 74667 32780 74709 32789
rect 74188 32740 74420 32780
rect 74283 31856 74325 31865
rect 74283 31816 74284 31856
rect 74324 31816 74325 31856
rect 74283 31807 74325 31816
rect 73612 31648 73655 31688
rect 73900 31648 73945 31688
rect 73996 31648 74055 31688
rect 72556 31480 72745 31520
rect 71884 30857 71924 31480
rect 72414 31471 72456 31480
rect 72304 31352 72346 31361
rect 72304 31312 72305 31352
rect 72345 31312 72346 31352
rect 72304 31303 72346 31312
rect 72305 31248 72345 31303
rect 72415 31248 72455 31471
rect 72705 31248 72745 31480
rect 72814 31436 72856 31445
rect 72814 31396 72815 31436
rect 72855 31396 72856 31436
rect 72814 31387 72856 31396
rect 72815 31248 72855 31387
rect 73105 31248 73145 31648
rect 73214 31604 73256 31613
rect 73214 31564 73215 31604
rect 73255 31564 73256 31604
rect 73214 31555 73256 31564
rect 73215 31248 73255 31555
rect 73504 31520 73546 31529
rect 73504 31480 73505 31520
rect 73545 31480 73546 31520
rect 73504 31471 73546 31480
rect 73505 31248 73545 31471
rect 73615 31248 73655 31648
rect 73905 31248 73945 31648
rect 74015 31248 74055 31648
rect 74284 31604 74324 31807
rect 74380 31688 74420 32740
rect 74667 32740 74668 32780
rect 74708 32740 74709 32780
rect 74667 32731 74709 32740
rect 74667 31940 74709 31949
rect 74667 31900 74668 31940
rect 74708 31900 74709 31940
rect 74667 31891 74709 31900
rect 74380 31648 74455 31688
rect 74284 31564 74345 31604
rect 74305 31248 74345 31564
rect 74415 31248 74455 31648
rect 74668 31436 74708 31891
rect 74764 31520 74804 32899
rect 75052 31688 75092 34168
rect 75148 31772 75188 34252
rect 75628 34242 75668 34327
rect 75340 34208 75380 34217
rect 75340 32789 75380 34168
rect 75532 34208 75572 34217
rect 75339 32780 75381 32789
rect 75339 32740 75340 32780
rect 75380 32740 75381 32780
rect 75339 32731 75381 32740
rect 75148 31732 75255 31772
rect 75052 31648 75145 31688
rect 74764 31480 74855 31520
rect 74668 31396 74745 31436
rect 74705 31248 74745 31396
rect 74815 31248 74855 31480
rect 75105 31248 75145 31648
rect 75215 31248 75255 31732
rect 75532 31688 75572 34168
rect 75627 32780 75669 32789
rect 75627 32740 75628 32780
rect 75668 32740 75669 32780
rect 75627 32731 75669 32740
rect 75628 31688 75668 32731
rect 75505 31648 75572 31688
rect 75615 31648 75668 31688
rect 75505 31248 75545 31648
rect 75615 31248 75655 31648
rect 75724 31361 75764 34924
rect 75820 34915 75860 34924
rect 75916 34924 76012 34964
rect 75916 34544 75956 34924
rect 76012 34915 76052 34924
rect 75820 34504 75956 34544
rect 75820 31688 75860 34504
rect 76204 34460 76244 35167
rect 76587 35132 76629 35141
rect 76587 35092 76588 35132
rect 76628 35092 76629 35132
rect 76587 35083 76629 35092
rect 75916 34376 75956 34387
rect 76204 34385 76244 34420
rect 75916 34301 75956 34336
rect 76203 34376 76245 34385
rect 76203 34336 76204 34376
rect 76244 34336 76245 34376
rect 76588 34376 76628 35083
rect 76684 35082 76724 35167
rect 77067 35132 77109 35141
rect 77067 35092 77068 35132
rect 77108 35092 77109 35132
rect 77067 35083 77109 35092
rect 77068 34998 77108 35083
rect 77260 35048 77300 35167
rect 77548 35082 77588 35167
rect 77260 34999 77300 35008
rect 76780 34964 76820 34973
rect 77452 34964 77492 34973
rect 76780 34460 76820 34924
rect 77356 34924 77452 34964
rect 76972 34460 77012 34471
rect 76780 34420 76916 34460
rect 76684 34376 76724 34385
rect 76588 34336 76684 34376
rect 76203 34327 76245 34336
rect 76684 34327 76724 34336
rect 75915 34292 75957 34301
rect 76204 34296 76244 34327
rect 75915 34252 75916 34292
rect 75956 34252 75957 34292
rect 75915 34243 75957 34252
rect 76780 34217 76820 34302
rect 76012 34208 76052 34217
rect 76396 34208 76436 34217
rect 76052 34168 76148 34208
rect 76012 34159 76052 34168
rect 75820 31648 75945 31688
rect 75723 31352 75765 31361
rect 75723 31312 75724 31352
rect 75764 31312 75765 31352
rect 75723 31303 75765 31312
rect 75905 31248 75945 31648
rect 76108 31604 76148 34168
rect 76204 34168 76396 34208
rect 76204 31688 76244 34168
rect 76396 34159 76436 34168
rect 76779 34208 76821 34217
rect 76779 34168 76780 34208
rect 76820 34168 76821 34208
rect 76779 34159 76821 34168
rect 76352 34040 76720 34049
rect 76876 34040 76916 34420
rect 76972 34385 77012 34420
rect 76971 34376 77013 34385
rect 77356 34376 77396 34924
rect 77452 34915 77492 34924
rect 77644 34544 77684 35680
rect 77835 35216 77877 35225
rect 77835 35176 77836 35216
rect 77876 35176 77877 35216
rect 77835 35167 77877 35176
rect 78508 35216 78548 35932
rect 78604 35923 78644 35932
rect 78508 35167 78548 35176
rect 78796 35720 78836 35729
rect 76971 34336 76972 34376
rect 77012 34336 77013 34376
rect 76971 34327 77013 34336
rect 77068 34336 77396 34376
rect 77452 34504 77684 34544
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76352 33991 76720 34000
rect 76780 34000 76916 34040
rect 76683 33872 76725 33881
rect 76683 33832 76684 33872
rect 76724 33832 76725 33872
rect 76683 33823 76725 33832
rect 76684 32537 76724 33823
rect 76683 32528 76725 32537
rect 76683 32488 76684 32528
rect 76724 32488 76725 32528
rect 76683 32479 76725 32488
rect 76780 31688 76820 34000
rect 76204 31648 76455 31688
rect 76108 31564 76345 31604
rect 76014 31352 76056 31361
rect 76014 31312 76015 31352
rect 76055 31312 76056 31352
rect 76014 31303 76056 31312
rect 76015 31248 76055 31303
rect 76305 31248 76345 31564
rect 76415 31248 76455 31648
rect 76705 31648 76820 31688
rect 76705 31248 76745 31648
rect 76814 31520 76856 31529
rect 76814 31480 76815 31520
rect 76855 31480 76856 31520
rect 76814 31471 76856 31480
rect 76815 31248 76855 31471
rect 77068 31352 77108 34336
rect 77164 34208 77204 34217
rect 77204 34168 77300 34208
rect 77164 34159 77204 34168
rect 77260 31352 77300 34168
rect 77355 32528 77397 32537
rect 77355 32488 77356 32528
rect 77396 32488 77397 32528
rect 77355 32479 77397 32488
rect 77356 31604 77396 32479
rect 77452 31688 77492 34504
rect 77836 34460 77876 35167
rect 78604 34964 78644 34973
rect 78508 34924 78604 34964
rect 77548 34376 77588 34387
rect 77836 34385 77876 34420
rect 78220 34460 78260 34471
rect 78220 34385 78260 34420
rect 77548 34301 77588 34336
rect 77835 34376 77877 34385
rect 77835 34336 77836 34376
rect 77876 34336 77877 34376
rect 77835 34327 77877 34336
rect 78219 34376 78261 34385
rect 78219 34336 78220 34376
rect 78260 34336 78261 34376
rect 78219 34327 78261 34336
rect 77547 34292 77589 34301
rect 77547 34252 77548 34292
rect 77588 34252 77589 34292
rect 77547 34243 77589 34252
rect 77644 34208 77684 34217
rect 78028 34208 78068 34217
rect 77684 34168 77876 34208
rect 77644 34159 77684 34168
rect 77836 31688 77876 34168
rect 78028 31688 78068 34168
rect 78315 34208 78357 34217
rect 78315 34168 78316 34208
rect 78356 34168 78357 34208
rect 78315 34159 78357 34168
rect 78412 34208 78452 34217
rect 78316 31688 78356 34159
rect 77452 31648 77655 31688
rect 77836 31648 77945 31688
rect 77356 31564 77545 31604
rect 77068 31312 77145 31352
rect 77105 31248 77145 31312
rect 77215 31312 77300 31352
rect 77215 31248 77255 31312
rect 77505 31248 77545 31564
rect 77615 31248 77655 31648
rect 77905 31248 77945 31648
rect 78015 31648 78068 31688
rect 78305 31648 78356 31688
rect 78412 31688 78452 34168
rect 78508 31688 78548 34924
rect 78604 34915 78644 34924
rect 78699 34376 78741 34385
rect 78699 34336 78700 34376
rect 78740 34336 78741 34376
rect 78699 34327 78741 34336
rect 78700 34242 78740 34327
rect 78603 34208 78645 34217
rect 78603 34168 78604 34208
rect 78644 34168 78645 34208
rect 78603 34159 78645 34168
rect 78604 34074 78644 34159
rect 78796 31688 78836 35680
rect 78892 34376 78932 35932
rect 79180 35720 79220 35729
rect 79084 35680 79180 35720
rect 78988 35141 79028 35226
rect 78987 35132 79029 35141
rect 78987 35092 78988 35132
rect 79028 35092 79029 35132
rect 78987 35083 79029 35092
rect 79084 34964 79124 35680
rect 79180 35671 79220 35680
rect 79180 35384 79220 35393
rect 79276 35384 79316 35932
rect 79372 35923 79412 35932
rect 81388 35972 81428 35981
rect 80236 35888 80276 35897
rect 79220 35344 79316 35384
rect 79180 35335 79220 35344
rect 79276 35132 79316 35344
rect 80140 35848 80236 35888
rect 79756 35216 79796 35225
rect 79372 35132 79412 35141
rect 79276 35092 79372 35132
rect 79372 35083 79412 35092
rect 78988 34924 79124 34964
rect 79564 34964 79604 34973
rect 79604 34924 79700 34964
rect 78988 34376 79028 34924
rect 79564 34915 79604 34924
rect 79112 34796 79480 34805
rect 79152 34756 79194 34796
rect 79234 34756 79276 34796
rect 79316 34756 79358 34796
rect 79398 34756 79440 34796
rect 79112 34747 79480 34756
rect 79372 34376 79412 34385
rect 78988 34336 79220 34376
rect 78892 34327 78932 34336
rect 78988 34208 79028 34217
rect 79028 34168 79124 34208
rect 78988 34159 79028 34168
rect 79084 31688 79124 34168
rect 79180 31772 79220 34336
rect 79275 34292 79317 34301
rect 79372 34292 79412 34336
rect 79275 34252 79276 34292
rect 79316 34252 79412 34292
rect 79275 34243 79317 34252
rect 79468 34208 79508 34217
rect 79180 31732 79255 31772
rect 78412 31648 78455 31688
rect 78508 31648 78745 31688
rect 78796 31648 78855 31688
rect 79084 31648 79145 31688
rect 78015 31248 78055 31648
rect 78305 31248 78345 31648
rect 78415 31248 78455 31648
rect 78705 31248 78745 31648
rect 78815 31248 78855 31648
rect 79105 31248 79145 31648
rect 79215 31248 79255 31732
rect 79468 31688 79508 34168
rect 79660 31688 79700 34924
rect 79756 34460 79796 35176
rect 80140 35132 80180 35848
rect 80236 35839 80276 35848
rect 80332 35720 80372 35729
rect 80140 35057 80180 35092
rect 80236 35680 80332 35720
rect 80139 35048 80181 35057
rect 80044 35008 80140 35048
rect 80180 35008 80181 35048
rect 79756 34385 79796 34420
rect 79852 34964 79892 34973
rect 79755 34376 79797 34385
rect 79755 34336 79756 34376
rect 79796 34336 79797 34376
rect 79755 34327 79797 34336
rect 79756 34296 79796 34327
rect 79468 31648 79545 31688
rect 79505 31248 79545 31648
rect 79615 31648 79700 31688
rect 79615 31248 79655 31648
rect 79852 31352 79892 34924
rect 80044 34376 80084 35008
rect 80139 34999 80181 35008
rect 80236 34721 80276 35680
rect 80332 35671 80372 35680
rect 80352 35552 80720 35561
rect 80392 35512 80434 35552
rect 80474 35512 80516 35552
rect 80556 35512 80598 35552
rect 80638 35512 80680 35552
rect 80352 35503 80720 35512
rect 80620 35216 80660 35225
rect 80620 35057 80660 35176
rect 80908 35132 80948 35143
rect 80908 35057 80948 35092
rect 81388 35057 81428 35932
rect 85036 35972 85076 35981
rect 85420 35972 85460 35981
rect 85076 35932 85420 35972
rect 81580 35720 81620 35729
rect 81620 35680 81716 35720
rect 81580 35671 81620 35680
rect 81580 35216 81620 35227
rect 81580 35141 81620 35176
rect 81579 35132 81621 35141
rect 81579 35092 81580 35132
rect 81620 35092 81621 35132
rect 81579 35083 81621 35092
rect 80427 35048 80469 35057
rect 80427 35008 80428 35048
rect 80468 35008 80469 35048
rect 80427 34999 80469 35008
rect 80619 35048 80661 35057
rect 80619 35008 80620 35048
rect 80660 35008 80661 35048
rect 80619 34999 80661 35008
rect 80907 35048 80949 35057
rect 80907 35008 80908 35048
rect 80948 35008 80949 35048
rect 80907 34999 80949 35008
rect 81387 35048 81429 35057
rect 81387 35008 81388 35048
rect 81428 35008 81429 35048
rect 81387 34999 81429 35008
rect 80332 34964 80372 34973
rect 80235 34712 80277 34721
rect 80235 34672 80236 34712
rect 80276 34672 80277 34712
rect 80235 34663 80277 34672
rect 80127 34376 80167 34382
rect 80044 34373 80167 34376
rect 80044 34336 80127 34373
rect 80127 34324 80167 34333
rect 80236 34292 80276 34301
rect 80276 34252 80284 34292
rect 80236 34243 80284 34252
rect 79948 34208 79988 34217
rect 79988 34168 80084 34208
rect 79948 34159 79988 34168
rect 80044 31352 80084 34168
rect 80244 34124 80284 34243
rect 80332 34217 80372 34924
rect 80428 34460 80468 34999
rect 80716 34964 80756 34973
rect 80716 34721 80756 34924
rect 81100 34964 81140 34973
rect 80715 34712 80757 34721
rect 80715 34672 80716 34712
rect 80756 34672 80757 34712
rect 80715 34663 80757 34672
rect 80620 34544 80660 34553
rect 80660 34504 80948 34544
rect 80620 34495 80660 34504
rect 80331 34208 80373 34217
rect 80331 34168 80332 34208
rect 80372 34168 80373 34208
rect 80428 34208 80468 34420
rect 80812 34208 80852 34217
rect 80428 34168 80812 34208
rect 80331 34159 80373 34168
rect 80812 34159 80852 34168
rect 80236 34084 80284 34124
rect 80236 32789 80276 34084
rect 80352 34040 80720 34049
rect 80392 34000 80434 34040
rect 80474 34000 80516 34040
rect 80556 34000 80598 34040
rect 80638 34000 80680 34040
rect 80352 33991 80720 34000
rect 80427 33872 80469 33881
rect 80427 33832 80428 33872
rect 80468 33832 80469 33872
rect 80427 33823 80469 33832
rect 80331 33788 80373 33797
rect 80331 33748 80332 33788
rect 80372 33748 80373 33788
rect 80331 33739 80373 33748
rect 80235 32780 80277 32789
rect 80235 32740 80236 32780
rect 80276 32740 80277 32780
rect 80235 32731 80277 32740
rect 80332 31688 80372 33739
rect 80428 31688 80468 33823
rect 80715 32780 80757 32789
rect 80715 32740 80716 32780
rect 80756 32740 80757 32780
rect 80715 32731 80757 32740
rect 80716 31688 80756 32731
rect 80908 31688 80948 34504
rect 81004 34469 81044 34554
rect 81003 34460 81045 34469
rect 81003 34420 81004 34460
rect 81044 34420 81045 34460
rect 81003 34411 81045 34420
rect 81003 34292 81045 34301
rect 81003 34252 81004 34292
rect 81044 34252 81045 34292
rect 81003 34243 81045 34252
rect 79852 31312 79945 31352
rect 79905 31248 79945 31312
rect 80015 31312 80084 31352
rect 80305 31648 80372 31688
rect 80415 31648 80468 31688
rect 80705 31648 80756 31688
rect 80815 31648 80948 31688
rect 80015 31248 80055 31312
rect 80305 31248 80345 31648
rect 80415 31248 80455 31648
rect 80705 31248 80745 31648
rect 80815 31248 80855 31648
rect 81004 31604 81044 34243
rect 81100 31688 81140 34924
rect 81484 34964 81524 34973
rect 81524 34924 81620 34964
rect 81484 34915 81524 34924
rect 81195 34460 81237 34469
rect 81195 34420 81196 34460
rect 81236 34420 81237 34460
rect 81195 34411 81237 34420
rect 81483 34460 81525 34469
rect 81483 34420 81484 34460
rect 81524 34420 81525 34460
rect 81483 34411 81525 34420
rect 81196 34376 81236 34411
rect 81196 34325 81236 34336
rect 81484 34326 81524 34411
rect 81292 34208 81332 34217
rect 81292 32789 81332 34168
rect 81291 32780 81333 32789
rect 81291 32740 81292 32780
rect 81332 32740 81333 32780
rect 81291 32731 81333 32740
rect 81580 31688 81620 34924
rect 81676 34544 81716 35680
rect 84352 35552 84720 35561
rect 84392 35512 84434 35552
rect 84474 35512 84516 35552
rect 84556 35512 84598 35552
rect 84638 35512 84680 35552
rect 84352 35503 84720 35512
rect 82348 35216 82388 35225
rect 82348 35141 82388 35176
rect 83883 35216 83925 35225
rect 83883 35176 83884 35216
rect 83924 35176 83925 35216
rect 83883 35167 83925 35176
rect 84267 35216 84309 35225
rect 84267 35176 84268 35216
rect 84308 35176 84309 35216
rect 84267 35167 84309 35176
rect 84651 35216 84693 35225
rect 84651 35176 84652 35216
rect 84692 35176 84693 35216
rect 84651 35167 84693 35176
rect 85036 35216 85076 35932
rect 85420 35923 85460 35932
rect 92236 35972 92276 35981
rect 86572 35888 86612 35897
rect 85227 35720 85269 35729
rect 85227 35680 85228 35720
rect 85268 35680 85269 35720
rect 85227 35671 85269 35680
rect 85612 35720 85652 35729
rect 85228 35586 85268 35671
rect 81771 35132 81813 35141
rect 81771 35092 81772 35132
rect 81812 35092 81813 35132
rect 81771 35083 81813 35092
rect 82347 35132 82389 35141
rect 82347 35092 82348 35132
rect 82388 35092 82389 35132
rect 82347 35083 82389 35092
rect 82635 35132 82677 35141
rect 82635 35092 82636 35132
rect 82676 35092 82677 35132
rect 82635 35083 82677 35092
rect 83307 35132 83349 35141
rect 83307 35092 83308 35132
rect 83348 35092 83349 35132
rect 83307 35083 83349 35092
rect 83499 35132 83541 35141
rect 83499 35092 83500 35132
rect 83540 35092 83541 35132
rect 83499 35083 83541 35092
rect 83884 35132 83924 35167
rect 81772 34998 81812 35083
rect 81964 34964 82004 34973
rect 81868 34544 81908 34555
rect 81676 34504 81812 34544
rect 81675 34376 81717 34385
rect 81675 34336 81676 34376
rect 81716 34336 81717 34376
rect 81675 34327 81717 34336
rect 81676 34208 81716 34327
rect 81676 34159 81716 34168
rect 81100 31648 81255 31688
rect 81004 31564 81145 31604
rect 81105 31248 81145 31564
rect 81215 31248 81255 31648
rect 81505 31648 81620 31688
rect 81505 31248 81545 31648
rect 81772 31604 81812 34504
rect 81868 34469 81908 34504
rect 81867 34460 81909 34469
rect 81867 34420 81868 34460
rect 81908 34420 81909 34460
rect 81867 34411 81909 34420
rect 81964 32864 82004 34924
rect 82252 34553 82292 34566
rect 82251 34544 82293 34553
rect 82348 34544 82388 35083
rect 82636 34998 82676 35083
rect 83308 34998 83348 35083
rect 83500 34998 83540 35083
rect 82444 34964 82484 34973
rect 82828 34964 82868 34973
rect 83116 34964 83156 34973
rect 82484 34924 82580 34964
rect 82444 34915 82484 34924
rect 82156 34504 82252 34544
rect 82292 34504 82388 34544
rect 82060 34460 82100 34469
rect 82060 34133 82100 34420
rect 82156 34385 82196 34504
rect 82251 34495 82293 34504
rect 82252 34471 82292 34495
rect 82252 34422 82292 34431
rect 82155 34376 82197 34385
rect 82155 34336 82156 34376
rect 82196 34336 82197 34376
rect 82155 34327 82197 34336
rect 82444 34208 82484 34217
rect 82059 34124 82101 34133
rect 82059 34084 82060 34124
rect 82100 34084 82101 34124
rect 82059 34075 82101 34084
rect 81964 32824 82100 32864
rect 81867 32780 81909 32789
rect 81867 32740 81868 32780
rect 81908 32740 81920 32780
rect 81867 32731 81920 32740
rect 81880 32696 81920 32731
rect 81880 32656 82004 32696
rect 81964 31688 82004 32656
rect 81615 31564 81812 31604
rect 81905 31648 82004 31688
rect 81615 31248 81655 31564
rect 81905 31248 81945 31648
rect 82060 31604 82100 32824
rect 82444 31688 82484 34168
rect 82415 31648 82484 31688
rect 82015 31564 82100 31604
rect 82304 31604 82346 31613
rect 82304 31564 82305 31604
rect 82345 31564 82346 31604
rect 82015 31248 82055 31564
rect 82304 31555 82346 31564
rect 82305 31248 82345 31555
rect 82415 31248 82455 31648
rect 82540 31604 82580 34924
rect 82635 34544 82677 34553
rect 82635 34504 82636 34544
rect 82676 34504 82677 34544
rect 82635 34495 82677 34504
rect 82636 34376 82676 34495
rect 82636 34327 82676 34336
rect 82732 34208 82772 34217
rect 82732 31781 82772 34168
rect 82731 31772 82773 31781
rect 82731 31732 82732 31772
rect 82772 31732 82773 31772
rect 82731 31723 82773 31732
rect 82828 31688 82868 34924
rect 83020 34924 83116 34964
rect 83020 34040 83060 34924
rect 83116 34915 83156 34924
rect 83692 34964 83732 34973
rect 83112 34796 83480 34805
rect 83152 34756 83194 34796
rect 83234 34756 83276 34796
rect 83316 34756 83358 34796
rect 83398 34756 83440 34796
rect 83112 34747 83480 34756
rect 83307 34628 83349 34637
rect 83307 34588 83308 34628
rect 83348 34588 83349 34628
rect 83307 34579 83349 34588
rect 83595 34628 83637 34637
rect 83595 34588 83596 34628
rect 83636 34588 83637 34628
rect 83595 34579 83637 34588
rect 83308 34494 83348 34579
rect 83115 34460 83157 34469
rect 83115 34420 83116 34460
rect 83156 34420 83157 34460
rect 83115 34411 83157 34420
rect 83116 34326 83156 34411
rect 83596 34376 83636 34579
rect 83596 34327 83636 34336
rect 83500 34208 83540 34217
rect 83500 34049 83540 34168
rect 83499 34040 83541 34049
rect 83020 34000 83252 34040
rect 83115 33872 83157 33881
rect 83115 33832 83116 33872
rect 83156 33832 83157 33872
rect 83115 33823 83157 33832
rect 83116 31688 83156 33823
rect 82815 31648 82868 31688
rect 83105 31648 83156 31688
rect 83212 31688 83252 34000
rect 83499 34000 83500 34040
rect 83540 34000 83541 34040
rect 83499 33991 83541 34000
rect 83212 31648 83255 31688
rect 82540 31564 82745 31604
rect 82705 31248 82745 31564
rect 82815 31248 82855 31648
rect 83105 31248 83145 31648
rect 83215 31248 83255 31648
rect 83504 31604 83546 31613
rect 83504 31564 83505 31604
rect 83545 31564 83546 31604
rect 83504 31555 83546 31564
rect 83505 31248 83545 31555
rect 83692 31352 83732 34924
rect 83884 34637 83924 35092
rect 84268 35132 84308 35167
rect 84268 35081 84308 35092
rect 84652 35082 84692 35167
rect 84076 34964 84116 34973
rect 83980 34924 84076 34964
rect 83883 34628 83925 34637
rect 83883 34588 83884 34628
rect 83924 34588 83925 34628
rect 83883 34579 83925 34588
rect 83884 34376 83924 34579
rect 83884 34327 83924 34336
rect 83788 34208 83828 34217
rect 83788 31613 83828 34168
rect 83883 34208 83925 34217
rect 83883 34168 83884 34208
rect 83924 34168 83925 34208
rect 83883 34159 83925 34168
rect 83787 31604 83829 31613
rect 83787 31564 83788 31604
rect 83828 31564 83829 31604
rect 83884 31604 83924 34159
rect 83980 31688 84020 34924
rect 84076 34915 84116 34924
rect 84460 34964 84500 34973
rect 84171 34628 84213 34637
rect 84171 34588 84172 34628
rect 84212 34588 84213 34628
rect 84171 34579 84213 34588
rect 84172 34376 84212 34579
rect 84460 34544 84500 34924
rect 84748 34964 84788 34973
rect 84652 34553 84692 34584
rect 84172 34327 84212 34336
rect 84268 34504 84500 34544
rect 84651 34544 84693 34553
rect 84651 34504 84652 34544
rect 84692 34504 84693 34544
rect 84075 34208 84117 34217
rect 84075 34168 84076 34208
rect 84116 34168 84117 34208
rect 84075 34159 84117 34168
rect 84076 34074 84116 34159
rect 84171 34124 84213 34133
rect 84171 34084 84172 34124
rect 84212 34084 84213 34124
rect 84171 34075 84213 34084
rect 84172 31688 84212 34075
rect 84268 33872 84308 34504
rect 84651 34495 84693 34504
rect 84652 34460 84692 34495
rect 84460 34376 84500 34385
rect 84652 34376 84692 34420
rect 84748 34385 84788 34924
rect 85036 34637 85076 35176
rect 85132 34964 85172 34973
rect 85035 34628 85077 34637
rect 85035 34588 85036 34628
rect 85076 34588 85077 34628
rect 85035 34579 85077 34588
rect 85035 34460 85077 34469
rect 85035 34420 85036 34460
rect 85076 34420 85077 34460
rect 85035 34411 85077 34420
rect 84500 34336 84692 34376
rect 84747 34376 84789 34385
rect 84747 34336 84748 34376
rect 84788 34336 84789 34376
rect 84460 34327 84500 34336
rect 84747 34327 84789 34336
rect 85036 34326 85076 34411
rect 84364 34217 84404 34302
rect 84363 34208 84405 34217
rect 84363 34168 84364 34208
rect 84404 34168 84405 34208
rect 84363 34159 84405 34168
rect 84844 34208 84884 34217
rect 84352 34040 84720 34049
rect 84392 34000 84434 34040
rect 84474 34000 84516 34040
rect 84556 34000 84598 34040
rect 84638 34000 84680 34040
rect 84352 33991 84720 34000
rect 84268 33832 84500 33872
rect 84460 31688 84500 33832
rect 84844 31688 84884 34168
rect 84939 34208 84981 34217
rect 84939 34168 84940 34208
rect 84980 34168 84981 34208
rect 84939 34159 84981 34168
rect 83980 31648 84055 31688
rect 84172 31648 84345 31688
rect 83884 31564 83945 31604
rect 83787 31555 83829 31564
rect 83615 31312 83732 31352
rect 83615 31248 83655 31312
rect 83905 31248 83945 31564
rect 84015 31248 84055 31648
rect 84305 31248 84345 31648
rect 84415 31648 84500 31688
rect 84815 31648 84884 31688
rect 84415 31248 84455 31648
rect 84704 31604 84746 31613
rect 84704 31564 84705 31604
rect 84745 31564 84746 31604
rect 84704 31555 84746 31564
rect 84705 31248 84745 31555
rect 84815 31248 84855 31648
rect 84940 31613 84980 34159
rect 85132 31688 85172 34924
rect 85227 34544 85269 34553
rect 85227 34504 85228 34544
rect 85268 34504 85269 34544
rect 85227 34495 85269 34504
rect 85419 34544 85461 34553
rect 85419 34504 85420 34544
rect 85460 34504 85461 34544
rect 85419 34495 85461 34504
rect 85228 34410 85268 34495
rect 85420 34376 85460 34495
rect 85420 34327 85460 34336
rect 85516 34208 85556 34217
rect 85516 31688 85556 34168
rect 85105 31648 85172 31688
rect 85505 31648 85556 31688
rect 85612 31688 85652 35680
rect 85804 35216 85844 35225
rect 85804 34553 85844 35176
rect 86572 35141 86612 35848
rect 87820 35888 87860 35897
rect 89836 35888 89876 35897
rect 90220 35888 90260 35897
rect 87860 35848 88148 35888
rect 87820 35839 87860 35848
rect 86668 35720 86708 35729
rect 87916 35720 87956 35729
rect 86708 35680 86804 35720
rect 86668 35671 86708 35680
rect 86091 35132 86133 35141
rect 86091 35092 86092 35132
rect 86132 35092 86133 35132
rect 86091 35083 86133 35092
rect 86379 35132 86421 35141
rect 86379 35092 86380 35132
rect 86420 35092 86421 35132
rect 86379 35083 86421 35092
rect 86571 35132 86613 35141
rect 86571 35092 86572 35132
rect 86612 35092 86613 35132
rect 86571 35083 86613 35092
rect 86668 35132 86708 35141
rect 86092 34998 86132 35083
rect 85900 34964 85940 34973
rect 85803 34544 85845 34553
rect 85803 34504 85804 34544
rect 85844 34504 85845 34544
rect 85803 34495 85845 34504
rect 85804 34460 85844 34495
rect 85804 34409 85844 34420
rect 85900 31688 85940 34924
rect 86284 34964 86324 34973
rect 85996 34208 86036 34217
rect 85996 31688 86036 34168
rect 86187 34208 86229 34217
rect 86187 34168 86188 34208
rect 86228 34168 86229 34208
rect 86187 34159 86229 34168
rect 85612 31648 85655 31688
rect 85900 31648 85945 31688
rect 85996 31648 86055 31688
rect 84939 31604 84981 31613
rect 84939 31564 84940 31604
rect 84980 31564 84981 31604
rect 84939 31555 84981 31564
rect 85105 31248 85145 31648
rect 85214 31520 85256 31529
rect 85214 31480 85215 31520
rect 85255 31480 85256 31520
rect 85214 31471 85256 31480
rect 85215 31248 85255 31471
rect 85505 31248 85545 31648
rect 85615 31248 85655 31648
rect 85905 31248 85945 31648
rect 86015 31248 86055 31648
rect 86188 31604 86228 34159
rect 86284 31688 86324 34924
rect 86380 34628 86420 35083
rect 86475 35048 86517 35057
rect 86475 35008 86476 35048
rect 86516 35008 86517 35048
rect 86475 34999 86517 35008
rect 86380 34579 86420 34588
rect 86476 34460 86516 34999
rect 86668 34973 86708 35092
rect 86667 34964 86709 34973
rect 86667 34924 86668 34964
rect 86708 34924 86709 34964
rect 86667 34915 86709 34924
rect 86572 34460 86612 34469
rect 86476 34420 86572 34460
rect 86572 34411 86612 34420
rect 86764 34376 86804 35680
rect 87956 35680 88052 35720
rect 87916 35671 87956 35680
rect 87627 35216 87669 35225
rect 87724 35216 87764 35225
rect 87627 35176 87628 35216
rect 87668 35176 87724 35216
rect 87627 35167 87669 35176
rect 87724 35167 87764 35176
rect 87051 35132 87093 35141
rect 86956 35092 87052 35132
rect 87092 35092 87093 35132
rect 86860 34964 86900 34973
rect 86860 34637 86900 34924
rect 86859 34628 86901 34637
rect 86859 34588 86860 34628
rect 86900 34588 86901 34628
rect 86859 34579 86901 34588
rect 86956 34460 86996 35092
rect 87051 35083 87093 35092
rect 87435 35132 87477 35141
rect 87435 35092 87436 35132
rect 87476 35092 87477 35132
rect 87435 35083 87477 35092
rect 87916 35132 87956 35143
rect 87052 34998 87092 35083
rect 87244 34973 87284 35058
rect 87436 34998 87476 35083
rect 87916 35057 87956 35092
rect 87915 35048 87957 35057
rect 87915 35008 87916 35048
rect 87956 35008 87957 35048
rect 87915 34999 87957 35008
rect 87243 34964 87285 34973
rect 87243 34924 87244 34964
rect 87284 34924 87285 34964
rect 87243 34915 87285 34924
rect 87628 34964 87668 34973
rect 87112 34796 87480 34805
rect 87152 34756 87194 34796
rect 87234 34756 87276 34796
rect 87316 34756 87358 34796
rect 87398 34756 87440 34796
rect 87112 34747 87480 34756
rect 86668 34336 86804 34376
rect 86860 34420 87092 34460
rect 86860 34376 86900 34420
rect 86668 31688 86708 34336
rect 86860 34327 86900 34336
rect 87052 34376 87092 34420
rect 87340 34376 87380 34385
rect 87092 34336 87340 34376
rect 87052 34327 87092 34336
rect 87340 34327 87380 34336
rect 86763 34208 86805 34217
rect 86763 34168 86764 34208
rect 86804 34168 86805 34208
rect 86763 34159 86805 34168
rect 87148 34208 87188 34217
rect 86764 34074 86804 34159
rect 87148 31772 87188 34168
rect 87052 31732 87188 31772
rect 87436 34208 87476 34217
rect 86284 31648 86455 31688
rect 86668 31648 86745 31688
rect 86188 31564 86345 31604
rect 86305 31248 86345 31564
rect 86415 31248 86455 31648
rect 86705 31248 86745 31648
rect 86814 31520 86856 31529
rect 86814 31480 86815 31520
rect 86855 31480 86856 31520
rect 87052 31520 87092 31732
rect 87214 31604 87256 31613
rect 87214 31564 87215 31604
rect 87255 31564 87256 31604
rect 87214 31555 87256 31564
rect 87052 31480 87145 31520
rect 86814 31471 86856 31480
rect 86815 31248 86855 31471
rect 87105 31248 87145 31480
rect 87215 31248 87255 31555
rect 87436 31352 87476 34168
rect 87628 34049 87668 34924
rect 87723 34964 87765 34973
rect 87723 34924 87724 34964
rect 87764 34924 87765 34964
rect 87723 34915 87765 34924
rect 87627 34040 87669 34049
rect 87627 34000 87628 34040
rect 87668 34000 87669 34040
rect 87627 33991 87669 34000
rect 87724 31688 87764 34915
rect 87819 34460 87861 34469
rect 87819 34420 87820 34460
rect 87860 34420 87861 34460
rect 87819 34411 87861 34420
rect 87820 34326 87860 34411
rect 88012 34376 88052 35680
rect 88108 35384 88148 35848
rect 89876 35848 90220 35888
rect 88352 35552 88720 35561
rect 88392 35512 88434 35552
rect 88474 35512 88516 35552
rect 88556 35512 88598 35552
rect 88638 35512 88680 35552
rect 88352 35503 88720 35512
rect 88108 35225 88148 35344
rect 88107 35216 88149 35225
rect 88107 35176 88108 35216
rect 88148 35176 88149 35216
rect 88107 35167 88149 35176
rect 88491 35216 88533 35225
rect 88491 35176 88492 35216
rect 88532 35176 88533 35216
rect 88491 35167 88533 35176
rect 88108 34469 88148 35167
rect 88492 35132 88532 35167
rect 88492 35081 88532 35092
rect 88683 35132 88725 35141
rect 88683 35092 88684 35132
rect 88724 35092 88725 35132
rect 88683 35083 88725 35092
rect 89068 35132 89108 35141
rect 88684 34998 88724 35083
rect 88299 34964 88341 34973
rect 88299 34924 88300 34964
rect 88340 34924 88341 34964
rect 88299 34915 88341 34924
rect 88876 34964 88916 34973
rect 88300 34830 88340 34915
rect 88107 34460 88149 34469
rect 88107 34420 88108 34460
rect 88148 34420 88149 34460
rect 88107 34411 88149 34420
rect 88299 34460 88341 34469
rect 88299 34420 88300 34460
rect 88340 34420 88341 34460
rect 88299 34411 88341 34420
rect 88683 34460 88725 34469
rect 88683 34420 88684 34460
rect 88724 34420 88725 34460
rect 88683 34411 88725 34420
rect 87916 34336 88052 34376
rect 87916 31688 87956 34336
rect 88300 34326 88340 34411
rect 88684 34376 88724 34411
rect 88684 34325 88724 34336
rect 87615 31648 87764 31688
rect 87905 31648 87956 31688
rect 88012 34208 88052 34217
rect 88492 34208 88532 34217
rect 88012 31688 88052 34168
rect 88204 34168 88492 34208
rect 88012 31648 88055 31688
rect 87436 31312 87545 31352
rect 87505 31248 87545 31312
rect 87615 31248 87655 31648
rect 87905 31248 87945 31648
rect 88015 31248 88055 31648
rect 88204 31613 88244 34168
rect 88492 34159 88532 34168
rect 88780 34208 88820 34217
rect 88352 34040 88720 34049
rect 88392 34000 88434 34040
rect 88474 34000 88516 34040
rect 88556 34000 88598 34040
rect 88638 34000 88680 34040
rect 88352 33991 88720 34000
rect 88299 33872 88341 33881
rect 88299 33832 88300 33872
rect 88340 33832 88341 33872
rect 88299 33823 88341 33832
rect 88203 31604 88245 31613
rect 88203 31564 88204 31604
rect 88244 31564 88245 31604
rect 88300 31604 88340 33823
rect 88780 32528 88820 34168
rect 88684 32488 88820 32528
rect 88414 31604 88456 31613
rect 88300 31564 88345 31604
rect 88203 31555 88245 31564
rect 88305 31248 88345 31564
rect 88414 31564 88415 31604
rect 88455 31564 88456 31604
rect 88414 31555 88456 31564
rect 88415 31248 88455 31555
rect 88684 31352 88724 32488
rect 88876 31352 88916 34924
rect 89068 34544 89108 35092
rect 89452 35132 89492 35141
rect 89355 35048 89397 35057
rect 89355 35008 89356 35048
rect 89396 35008 89397 35048
rect 89355 34999 89397 35008
rect 89260 34964 89300 34973
rect 89164 34544 89204 34553
rect 89068 34504 89164 34544
rect 89164 34385 89204 34504
rect 89163 34376 89205 34385
rect 89163 34336 89164 34376
rect 89204 34336 89205 34376
rect 89163 34327 89205 34336
rect 89067 34208 89109 34217
rect 89067 34168 89068 34208
rect 89108 34168 89109 34208
rect 89067 34159 89109 34168
rect 89068 31688 89108 34159
rect 89068 31648 89145 31688
rect 88684 31312 88745 31352
rect 88705 31248 88745 31312
rect 88815 31312 88916 31352
rect 88815 31248 88855 31312
rect 89105 31248 89145 31648
rect 89260 31352 89300 34924
rect 89356 34460 89396 34999
rect 89356 34301 89396 34420
rect 89452 34385 89492 35092
rect 89836 35132 89876 35848
rect 90220 35839 90260 35848
rect 89932 35720 89972 35729
rect 90316 35720 90356 35729
rect 89932 35309 89972 35680
rect 90124 35680 90316 35720
rect 89931 35300 89973 35309
rect 89931 35260 89932 35300
rect 89972 35260 89973 35300
rect 89931 35251 89973 35260
rect 89931 35132 89973 35141
rect 89876 35092 89932 35132
rect 89972 35092 89973 35132
rect 89836 35083 89876 35092
rect 89931 35083 89973 35092
rect 89644 34964 89684 34973
rect 89684 34924 89780 34964
rect 89644 34915 89684 34924
rect 89451 34376 89493 34385
rect 89451 34336 89452 34376
rect 89492 34336 89493 34376
rect 89451 34327 89493 34336
rect 89643 34376 89685 34385
rect 89643 34336 89644 34376
rect 89684 34336 89685 34376
rect 89643 34327 89685 34336
rect 89355 34292 89397 34301
rect 89355 34252 89356 34292
rect 89396 34252 89397 34292
rect 89355 34243 89397 34252
rect 89644 34242 89684 34327
rect 89547 34208 89589 34217
rect 89547 34168 89548 34208
rect 89588 34168 89589 34208
rect 89547 34159 89589 34168
rect 89548 34074 89588 34159
rect 89740 31688 89780 34924
rect 89932 34385 89972 35083
rect 90028 34964 90068 34973
rect 89931 34377 89973 34385
rect 89931 34336 89932 34377
rect 89972 34336 89973 34377
rect 89931 34327 89973 34336
rect 89836 34208 89876 34217
rect 89836 31772 89876 34168
rect 89615 31648 89780 31688
rect 89823 31732 89876 31772
rect 89504 31436 89546 31445
rect 89504 31396 89505 31436
rect 89545 31396 89546 31436
rect 89504 31387 89546 31396
rect 89215 31312 89300 31352
rect 89215 31248 89255 31312
rect 89505 31248 89545 31387
rect 89615 31248 89655 31648
rect 89823 31604 89863 31732
rect 90028 31688 90068 34924
rect 89740 31564 89863 31604
rect 90015 31648 90068 31688
rect 90124 31688 90164 35680
rect 90316 35671 90356 35680
rect 90220 35141 90260 35226
rect 90682 35141 90722 35253
rect 91084 35141 91124 35226
rect 91468 35216 91508 35227
rect 91468 35141 91508 35176
rect 91756 35141 91796 35226
rect 92236 35216 92276 35932
rect 93964 35888 94004 35897
rect 94924 35888 94964 35897
rect 94004 35848 94924 35888
rect 92428 35729 92468 35814
rect 92427 35720 92469 35729
rect 92427 35680 92428 35720
rect 92468 35680 92469 35720
rect 92427 35671 92469 35680
rect 93868 35720 93908 35729
rect 92352 35552 92720 35561
rect 92392 35512 92434 35552
rect 92474 35512 92516 35552
rect 92556 35512 92598 35552
rect 92638 35512 92680 35552
rect 92352 35503 92720 35512
rect 92236 35141 92276 35176
rect 93100 35216 93140 35225
rect 93100 35141 93140 35176
rect 90219 35132 90261 35141
rect 90219 35092 90220 35132
rect 90260 35092 90261 35132
rect 90219 35083 90261 35092
rect 90681 35132 90723 35141
rect 90681 35089 90682 35132
rect 90722 35089 90723 35132
rect 90681 35083 90723 35089
rect 91083 35132 91125 35141
rect 91083 35092 91084 35132
rect 91124 35092 91125 35132
rect 91083 35083 91125 35092
rect 91467 35132 91509 35141
rect 91467 35092 91468 35132
rect 91508 35092 91509 35132
rect 91467 35083 91509 35092
rect 91755 35132 91797 35141
rect 91755 35092 91756 35132
rect 91796 35092 91797 35132
rect 91755 35083 91797 35092
rect 92235 35132 92277 35141
rect 92235 35092 92236 35132
rect 92276 35092 92277 35132
rect 92235 35083 92277 35092
rect 92427 35132 92469 35141
rect 92427 35092 92428 35132
rect 92468 35092 92469 35132
rect 92427 35083 92469 35092
rect 92619 35132 92661 35141
rect 92619 35092 92620 35132
rect 92660 35092 92661 35132
rect 92619 35083 92661 35092
rect 93099 35132 93141 35141
rect 93388 35132 93428 35141
rect 93099 35092 93100 35132
rect 93140 35092 93388 35132
rect 93099 35083 93141 35092
rect 93388 35083 93428 35092
rect 90412 34964 90452 34973
rect 90219 34880 90261 34889
rect 90219 34840 90220 34880
rect 90260 34840 90261 34880
rect 90219 34831 90261 34840
rect 90220 34553 90260 34831
rect 90219 34544 90261 34553
rect 90219 34504 90220 34544
rect 90260 34504 90261 34544
rect 90219 34495 90261 34504
rect 90220 34376 90260 34495
rect 90220 34327 90260 34336
rect 90315 34208 90357 34217
rect 90315 34168 90316 34208
rect 90356 34168 90357 34208
rect 90315 34159 90357 34168
rect 90316 34074 90356 34159
rect 90412 31688 90452 34924
rect 90682 34796 90722 35083
rect 90604 34756 90722 34796
rect 90892 34964 90932 34973
rect 91276 34964 91316 34973
rect 90604 34469 90644 34756
rect 90508 34460 90548 34469
rect 90603 34460 90645 34469
rect 90548 34420 90604 34460
rect 90644 34420 90645 34460
rect 90508 34411 90548 34420
rect 90603 34411 90645 34420
rect 90603 34208 90645 34217
rect 90603 34168 90604 34208
rect 90644 34168 90645 34208
rect 90603 34159 90645 34168
rect 90700 34208 90740 34217
rect 90740 34168 90836 34208
rect 90604 31688 90644 34159
rect 90700 34140 90740 34168
rect 90796 31688 90836 34168
rect 90892 32780 90932 34924
rect 90988 34924 91276 34964
rect 90988 34628 91028 34924
rect 91276 34915 91316 34924
rect 91564 34964 91604 34973
rect 91948 34964 91988 34973
rect 92332 34964 92372 34973
rect 91604 34924 91892 34964
rect 91564 34915 91604 34924
rect 91112 34796 91480 34805
rect 91152 34756 91194 34796
rect 91234 34756 91276 34796
rect 91316 34756 91358 34796
rect 91398 34756 91440 34796
rect 91112 34747 91480 34756
rect 90988 34588 91124 34628
rect 90988 34460 91028 34469
rect 90988 34301 91028 34420
rect 90987 34292 91029 34301
rect 90987 34252 90988 34292
rect 91028 34252 91029 34292
rect 90987 34243 91029 34252
rect 90892 32740 91028 32780
rect 90124 31648 90345 31688
rect 90412 31648 90455 31688
rect 90604 31648 90745 31688
rect 90796 31648 90855 31688
rect 89740 31445 89780 31564
rect 89904 31520 89946 31529
rect 89904 31480 89905 31520
rect 89945 31480 89946 31520
rect 89904 31471 89946 31480
rect 89739 31436 89781 31445
rect 89739 31396 89740 31436
rect 89780 31396 89781 31436
rect 89739 31387 89781 31396
rect 89905 31248 89945 31471
rect 90015 31248 90055 31648
rect 90305 31248 90345 31648
rect 90415 31248 90455 31648
rect 90705 31248 90745 31648
rect 90815 31248 90855 31648
rect 90988 31445 91028 32740
rect 91084 31688 91124 34588
rect 91180 34544 91220 34555
rect 91180 34469 91220 34504
rect 91179 34460 91221 34469
rect 91179 34420 91180 34460
rect 91220 34420 91221 34460
rect 91179 34411 91221 34420
rect 91467 34460 91509 34469
rect 91467 34420 91468 34460
rect 91508 34420 91509 34460
rect 91467 34411 91509 34420
rect 91755 34460 91797 34469
rect 91755 34420 91756 34460
rect 91796 34420 91797 34460
rect 91755 34411 91797 34420
rect 91468 34376 91508 34411
rect 91468 34325 91508 34336
rect 91756 34376 91796 34411
rect 91756 34325 91796 34336
rect 91372 34208 91412 34217
rect 91084 31648 91255 31688
rect 91104 31520 91146 31529
rect 91104 31480 91105 31520
rect 91145 31480 91146 31520
rect 91104 31471 91146 31480
rect 90987 31436 91029 31445
rect 90987 31396 90988 31436
rect 91028 31396 91029 31436
rect 90987 31387 91029 31396
rect 91105 31248 91145 31471
rect 91215 31248 91255 31648
rect 91372 31529 91412 34168
rect 91660 34208 91700 34217
rect 91660 32780 91700 34168
rect 91564 32740 91700 32780
rect 91564 31688 91604 32740
rect 91505 31648 91604 31688
rect 91852 31688 91892 34924
rect 91988 34924 92180 34964
rect 91948 34915 91988 34924
rect 92043 34376 92085 34385
rect 92043 34336 92044 34376
rect 92084 34336 92085 34376
rect 92043 34327 92085 34336
rect 92044 34242 92084 34327
rect 91947 34208 91989 34217
rect 91947 34168 91948 34208
rect 91988 34168 91989 34208
rect 91947 34159 91989 34168
rect 91948 34074 91988 34159
rect 92140 32780 92180 34924
rect 92236 34460 92276 34471
rect 92236 34385 92276 34420
rect 92235 34376 92277 34385
rect 92235 34336 92236 34376
rect 92276 34336 92277 34376
rect 92235 34327 92277 34336
rect 92332 34208 92372 34924
rect 92428 34628 92468 35083
rect 92620 34998 92660 35083
rect 92812 34964 92852 34973
rect 92852 34924 92948 34964
rect 92812 34915 92852 34924
rect 92428 34579 92468 34588
rect 92619 34544 92661 34553
rect 92619 34504 92620 34544
rect 92660 34504 92661 34544
rect 92619 34495 92661 34504
rect 92620 34376 92660 34495
rect 92812 34385 92852 34470
rect 92620 34327 92660 34336
rect 92811 34376 92853 34385
rect 92811 34336 92812 34376
rect 92852 34336 92853 34376
rect 92811 34327 92853 34336
rect 92044 32740 92180 32780
rect 92236 34168 92372 34208
rect 92811 34208 92853 34217
rect 92811 34168 92812 34208
rect 92852 34168 92853 34208
rect 92044 31688 92084 32740
rect 91852 31648 91945 31688
rect 91371 31520 91413 31529
rect 91371 31480 91372 31520
rect 91412 31480 91413 31520
rect 91371 31471 91413 31480
rect 91505 31248 91545 31648
rect 91614 31436 91656 31445
rect 91614 31396 91615 31436
rect 91655 31396 91656 31436
rect 91614 31387 91656 31396
rect 91615 31248 91655 31387
rect 91905 31248 91945 31648
rect 92015 31648 92084 31688
rect 92236 31688 92276 34168
rect 92811 34159 92853 34168
rect 92352 34040 92720 34049
rect 92392 34000 92434 34040
rect 92474 34000 92516 34040
rect 92556 34000 92598 34040
rect 92638 34000 92680 34040
rect 92352 33991 92720 34000
rect 92812 32780 92852 34159
rect 92716 32740 92852 32780
rect 92716 31688 92756 32740
rect 92908 31688 92948 34924
rect 93100 34469 93140 35083
rect 93196 34964 93236 34973
rect 93580 34964 93620 34973
rect 93236 34924 93428 34964
rect 93196 34915 93236 34924
rect 93099 34460 93141 34469
rect 93099 34420 93100 34460
rect 93140 34420 93141 34460
rect 93099 34411 93141 34420
rect 93099 34208 93141 34217
rect 93292 34208 93332 34217
rect 93099 34168 93100 34208
rect 93140 34168 93141 34208
rect 93099 34159 93141 34168
rect 93196 34168 93292 34208
rect 92236 31648 92345 31688
rect 92015 31248 92055 31648
rect 92305 31248 92345 31648
rect 92705 31648 92756 31688
rect 92815 31648 92948 31688
rect 93100 31688 93140 34159
rect 93196 31688 93236 34168
rect 93292 34159 93332 34168
rect 93388 31688 93428 34924
rect 93620 34924 93716 34964
rect 93580 34915 93620 34924
rect 93580 34469 93620 34500
rect 93579 34460 93621 34469
rect 93579 34420 93580 34460
rect 93620 34420 93621 34460
rect 93579 34411 93621 34420
rect 93580 34376 93620 34411
rect 93580 34301 93620 34336
rect 93579 34292 93621 34301
rect 93579 34252 93580 34292
rect 93620 34252 93621 34292
rect 93579 34243 93621 34252
rect 93483 34208 93525 34217
rect 93483 34168 93484 34208
rect 93524 34168 93525 34208
rect 93483 34159 93525 34168
rect 93484 34074 93524 34159
rect 93676 31688 93716 34924
rect 93868 34628 93908 35680
rect 93964 35384 94004 35848
rect 93964 35335 94004 35344
rect 94156 35132 94196 35141
rect 94540 35132 94580 35848
rect 94828 35216 94868 35848
rect 94924 35839 94964 35848
rect 94828 35167 94868 35176
rect 95020 35720 95060 35729
rect 94196 35092 94292 35132
rect 94156 35083 94196 35092
rect 93964 34964 94004 34973
rect 94004 34924 94100 34964
rect 93964 34915 94004 34924
rect 93868 34588 94004 34628
rect 93867 34460 93909 34469
rect 93867 34420 93868 34460
rect 93908 34420 93909 34460
rect 93867 34411 93909 34420
rect 93868 34326 93908 34411
rect 93964 31772 94004 34588
rect 94060 34469 94100 34924
rect 94059 34460 94101 34469
rect 94059 34420 94060 34460
rect 94100 34420 94101 34460
rect 94059 34411 94101 34420
rect 94252 34385 94292 35092
rect 94540 35083 94580 35092
rect 94348 34964 94388 34973
rect 94732 34964 94772 34973
rect 94388 34924 94484 34964
rect 94348 34915 94388 34924
rect 94251 34376 94293 34385
rect 94251 34336 94252 34376
rect 94292 34336 94293 34376
rect 94251 34327 94293 34336
rect 94252 34242 94292 34327
rect 93100 31648 93145 31688
rect 93196 31648 93255 31688
rect 93388 31648 93545 31688
rect 92414 31520 92456 31529
rect 92414 31480 92415 31520
rect 92455 31480 92456 31520
rect 92414 31471 92456 31480
rect 92415 31248 92455 31471
rect 92705 31248 92745 31648
rect 92815 31248 92855 31648
rect 93105 31248 93145 31648
rect 93215 31248 93255 31648
rect 93505 31248 93545 31648
rect 93615 31648 93716 31688
rect 93905 31732 94004 31772
rect 94060 34208 94100 34217
rect 93615 31248 93655 31648
rect 93905 31248 93945 31732
rect 94060 31688 94100 34168
rect 94348 34208 94388 34217
rect 94348 31688 94388 34168
rect 94015 31648 94100 31688
rect 94305 31648 94388 31688
rect 94015 31248 94055 31648
rect 94305 31248 94345 31648
rect 94444 31604 94484 34924
rect 94635 34460 94677 34469
rect 94635 34420 94636 34460
rect 94676 34420 94677 34460
rect 94635 34411 94677 34420
rect 94636 34326 94676 34411
rect 94732 31688 94772 34924
rect 95020 34628 95060 35680
rect 96352 35552 96720 35561
rect 96392 35512 96434 35552
rect 96474 35512 96516 35552
rect 96556 35512 96598 35552
rect 96638 35512 96680 35552
rect 96352 35503 96720 35512
rect 95212 35216 95252 35227
rect 95212 35141 95252 35176
rect 95211 35132 95253 35141
rect 95211 35092 95212 35132
rect 95252 35092 95253 35132
rect 95211 35083 95253 35092
rect 95403 35132 95445 35141
rect 95403 35092 95404 35132
rect 95444 35092 95445 35132
rect 95403 35083 95445 35092
rect 95788 35132 95828 35160
rect 96172 35141 96212 35226
rect 97036 35216 97076 35225
rect 95883 35132 95925 35141
rect 95828 35092 95884 35132
rect 95924 35092 95925 35132
rect 95788 35083 95828 35092
rect 95883 35083 95925 35092
rect 96171 35132 96213 35141
rect 96556 35132 96596 35141
rect 96171 35092 96172 35132
rect 96212 35092 96213 35132
rect 96171 35083 96213 35092
rect 96460 35092 96556 35132
rect 95116 34973 95156 35058
rect 95404 34998 95444 35083
rect 95115 34964 95157 34973
rect 95115 34924 95116 34964
rect 95156 34924 95157 34964
rect 95115 34915 95157 34924
rect 95596 34964 95636 34973
rect 95787 34964 95829 34973
rect 95636 34924 95732 34964
rect 95596 34915 95636 34924
rect 95112 34796 95480 34805
rect 95152 34756 95194 34796
rect 95234 34756 95276 34796
rect 95316 34756 95358 34796
rect 95398 34756 95440 34796
rect 95112 34747 95480 34756
rect 95020 34588 95156 34628
rect 95020 34460 95060 34469
rect 95020 34301 95060 34420
rect 95019 34292 95061 34301
rect 95019 34252 95020 34292
rect 95060 34252 95061 34292
rect 95019 34243 95061 34252
rect 94828 34208 94868 34217
rect 94828 31688 94868 34168
rect 95116 31688 95156 34588
rect 95595 34376 95637 34385
rect 95595 34336 95596 34376
rect 95636 34336 95637 34376
rect 95595 34327 95637 34336
rect 95596 34242 95636 34327
rect 94415 31564 94484 31604
rect 94705 31648 94772 31688
rect 94815 31648 94868 31688
rect 95105 31648 95156 31688
rect 95212 34208 95252 34217
rect 95212 31688 95252 34168
rect 95500 34208 95540 34217
rect 95500 31688 95540 34168
rect 95212 31648 95255 31688
rect 95500 31648 95545 31688
rect 94415 31248 94455 31564
rect 94705 31248 94745 31648
rect 94815 31248 94855 31648
rect 95105 31248 95145 31648
rect 95215 31248 95255 31648
rect 95505 31248 95545 31648
rect 95692 31604 95732 34924
rect 95787 34924 95788 34964
rect 95828 34924 95829 34964
rect 95787 34915 95829 34924
rect 95615 31564 95732 31604
rect 95788 31604 95828 34915
rect 95884 34628 95924 35083
rect 95884 34579 95924 34588
rect 95980 34964 96020 34973
rect 95980 31688 96020 34924
rect 96171 34964 96213 34973
rect 96171 34924 96172 34964
rect 96212 34924 96213 34964
rect 96171 34915 96213 34924
rect 96364 34964 96404 34973
rect 96075 34460 96117 34469
rect 96075 34420 96076 34460
rect 96116 34420 96117 34460
rect 96075 34411 96117 34420
rect 96076 34326 96116 34411
rect 96172 31688 96212 34915
rect 96268 34460 96308 34471
rect 96268 34385 96308 34420
rect 96267 34376 96309 34385
rect 96267 34336 96268 34376
rect 96308 34336 96309 34376
rect 96267 34327 96309 34336
rect 96364 34208 96404 34924
rect 96460 34544 96500 35092
rect 96556 35083 96596 35092
rect 96748 34964 96788 34973
rect 96460 34469 96500 34504
rect 96652 34924 96748 34964
rect 96459 34460 96501 34469
rect 96459 34420 96460 34460
rect 96500 34420 96501 34460
rect 96459 34411 96501 34420
rect 96652 34217 96692 34924
rect 96748 34915 96788 34924
rect 96939 34964 96981 34973
rect 96939 34924 96940 34964
rect 96980 34924 96981 34964
rect 96939 34915 96981 34924
rect 96940 34830 96980 34915
rect 96844 34553 96884 34638
rect 96843 34544 96885 34553
rect 96843 34504 96844 34544
rect 96884 34504 96885 34544
rect 96843 34495 96885 34504
rect 97036 34460 97076 35176
rect 97803 35132 97845 35141
rect 97803 35092 97804 35132
rect 97844 35092 97845 35132
rect 97803 35083 97845 35092
rect 97131 34544 97173 34553
rect 97131 34504 97132 34544
rect 97172 34504 97173 34544
rect 97131 34495 97173 34504
rect 97036 34385 97076 34420
rect 96747 34376 96789 34385
rect 96747 34336 96748 34376
rect 96788 34336 96789 34376
rect 96747 34327 96789 34336
rect 97035 34376 97077 34385
rect 97035 34336 97036 34376
rect 97076 34336 97077 34376
rect 97035 34327 97077 34336
rect 96748 34242 96788 34327
rect 96268 34168 96404 34208
rect 96651 34208 96693 34217
rect 96651 34168 96652 34208
rect 96692 34168 96693 34208
rect 96268 31772 96308 34168
rect 96651 34159 96693 34168
rect 96939 34124 96981 34133
rect 96939 34084 96940 34124
rect 96980 34084 96981 34124
rect 96939 34075 96981 34084
rect 96352 34040 96720 34049
rect 96392 34000 96434 34040
rect 96474 34000 96516 34040
rect 96556 34000 96598 34040
rect 96638 34000 96680 34040
rect 96352 33991 96720 34000
rect 96843 34040 96885 34049
rect 96843 34000 96844 34040
rect 96884 34000 96885 34040
rect 96843 33991 96885 34000
rect 96844 31772 96884 33991
rect 96268 31732 96455 31772
rect 95980 31648 96055 31688
rect 96172 31648 96345 31688
rect 95788 31564 95945 31604
rect 95615 31248 95655 31564
rect 95905 31248 95945 31564
rect 96015 31248 96055 31648
rect 96305 31248 96345 31648
rect 96415 31248 96455 31732
rect 96705 31732 96884 31772
rect 96705 31248 96745 31732
rect 96940 31688 96980 34075
rect 97132 31688 97172 34495
rect 97804 34469 97844 35083
rect 97996 34964 98036 34973
rect 98036 34924 98132 34964
rect 97996 34915 98036 34924
rect 97515 34460 97557 34469
rect 97515 34420 97516 34460
rect 97556 34420 97557 34460
rect 97515 34411 97557 34420
rect 97803 34460 97845 34469
rect 97803 34420 97804 34460
rect 97844 34420 97845 34460
rect 97803 34411 97845 34420
rect 97516 34326 97556 34411
rect 97900 34385 97940 34470
rect 97899 34376 97941 34385
rect 97899 34336 97900 34376
rect 97940 34336 97941 34376
rect 97899 34327 97941 34336
rect 97228 34208 97268 34217
rect 97228 31688 97268 34168
rect 96815 31648 96980 31688
rect 97105 31648 97172 31688
rect 97215 31648 97268 31688
rect 97708 34208 97748 34217
rect 96815 31248 96855 31648
rect 97105 31248 97145 31648
rect 97215 31248 97255 31648
rect 97504 31604 97546 31613
rect 97708 31604 97748 34168
rect 97899 34208 97941 34217
rect 97899 34168 97900 34208
rect 97940 34168 97941 34208
rect 97899 34159 97941 34168
rect 97996 34208 98036 34217
rect 97900 31688 97940 34159
rect 97996 34049 98036 34168
rect 97995 34040 98037 34049
rect 97995 34000 97996 34040
rect 98036 34000 98037 34040
rect 97995 33991 98037 34000
rect 97900 31648 97945 31688
rect 97504 31564 97505 31604
rect 97545 31564 97546 31604
rect 97504 31555 97546 31564
rect 97615 31564 97748 31604
rect 97505 31248 97545 31555
rect 97615 31248 97655 31564
rect 97905 31248 97945 31648
rect 98092 31604 98132 34924
rect 99112 34796 99480 34805
rect 99152 34756 99194 34796
rect 99234 34756 99276 34796
rect 99316 34756 99358 34796
rect 99398 34756 99440 34796
rect 99112 34747 99480 34756
rect 98668 34504 98996 34544
rect 98668 34460 98708 34504
rect 98668 34411 98708 34420
rect 98283 34376 98325 34385
rect 98283 34336 98284 34376
rect 98324 34336 98325 34376
rect 98283 34327 98325 34336
rect 98859 34376 98901 34385
rect 98859 34336 98860 34376
rect 98900 34336 98901 34376
rect 98956 34376 98996 34504
rect 99148 34376 99188 34385
rect 98956 34336 99148 34376
rect 98859 34327 98901 34336
rect 98284 34242 98324 34327
rect 98860 34242 98900 34327
rect 98188 34208 98228 34217
rect 98188 31613 98228 34168
rect 98476 34208 98516 34217
rect 98476 31688 98516 34168
rect 98955 34208 98997 34217
rect 98955 34168 98956 34208
rect 98996 34168 98997 34208
rect 98955 34159 98997 34168
rect 98956 34074 98996 34159
rect 98415 31648 98516 31688
rect 98015 31564 98132 31604
rect 98187 31604 98229 31613
rect 98187 31564 98188 31604
rect 98228 31564 98229 31604
rect 98015 31248 98055 31564
rect 98187 31555 98229 31564
rect 98304 31604 98346 31613
rect 98304 31564 98305 31604
rect 98345 31564 98346 31604
rect 98304 31555 98346 31564
rect 98305 31248 98345 31555
rect 98415 31248 98455 31648
rect 71883 30848 71925 30857
rect 71883 30808 71884 30848
rect 71924 30808 71925 30848
rect 71883 30799 71925 30808
rect 72305 25901 72345 26040
rect 72304 25892 72346 25901
rect 72304 25852 72305 25892
rect 72345 25852 72346 25892
rect 72304 25843 72346 25852
rect 72415 25817 72455 26040
rect 72705 25817 72745 26040
rect 72414 25808 72456 25817
rect 72414 25768 72415 25808
rect 72455 25768 72456 25808
rect 72414 25759 72456 25768
rect 72704 25808 72746 25817
rect 72704 25768 72705 25808
rect 72745 25768 72746 25808
rect 72704 25759 72746 25768
rect 72815 25733 72855 26040
rect 72815 25724 72885 25733
rect 72815 25684 72844 25724
rect 72884 25684 72885 25724
rect 73105 25724 73145 26040
rect 73215 25808 73255 26040
rect 73215 25768 73364 25808
rect 73105 25684 73268 25724
rect 72843 25675 72885 25684
rect 73228 25565 73268 25684
rect 73227 25556 73269 25565
rect 73227 25516 73228 25556
rect 73268 25516 73269 25556
rect 73227 25507 73269 25516
rect 73035 25304 73077 25313
rect 73035 25264 73036 25304
rect 73076 25264 73077 25304
rect 73035 25255 73077 25264
rect 72352 23456 72720 23465
rect 72392 23416 72434 23456
rect 72474 23416 72516 23456
rect 72556 23416 72598 23456
rect 72638 23416 72680 23456
rect 72352 23407 72720 23416
rect 71787 23372 71829 23381
rect 71787 23332 71788 23372
rect 71828 23332 71829 23372
rect 71787 23323 71829 23332
rect 2091 23288 2133 23297
rect 2091 23248 2092 23288
rect 2132 23248 2133 23288
rect 2091 23239 2133 23248
rect 68235 23288 68277 23297
rect 68235 23248 68236 23288
rect 68276 23248 68277 23288
rect 68235 23239 68277 23248
rect 1995 23120 2037 23129
rect 1995 23080 1996 23120
rect 2036 23080 2037 23120
rect 1995 23071 2037 23080
rect 939 22028 981 22037
rect 939 21988 940 22028
rect 980 21988 981 22028
rect 939 21979 981 21988
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 652 20936 692 20945
rect 652 20777 692 20896
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 652 19794 692 19879
rect 652 19424 692 19433
rect 652 19097 692 19384
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 652 18416 692 18425
rect 652 18257 692 18376
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17912 692 17921
rect 652 17417 692 17872
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 652 16904 692 16913
rect 652 16577 692 16864
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 652 16400 692 16409
rect 652 15737 692 16360
rect 651 15728 693 15737
rect 651 15688 652 15728
rect 692 15688 693 15728
rect 651 15679 693 15688
rect 1996 15485 2036 23071
rect 844 15476 884 15485
rect 652 15308 692 15317
rect 652 14897 692 15268
rect 844 14981 884 15436
rect 1995 15476 2037 15485
rect 1995 15436 1996 15476
rect 2036 15436 2037 15476
rect 1995 15427 2037 15436
rect 1996 15342 2036 15427
rect 1804 15308 1844 15317
rect 843 14972 885 14981
rect 843 14932 844 14972
rect 884 14932 885 14972
rect 843 14923 885 14932
rect 1707 14972 1749 14981
rect 1707 14932 1708 14972
rect 1748 14932 1749 14972
rect 1707 14923 1749 14932
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 1708 14838 1748 14923
rect 844 14804 884 14813
rect 652 14552 692 14561
rect 652 14057 692 14512
rect 844 14225 884 14764
rect 1804 14804 1844 15268
rect 1900 14804 1940 14813
rect 1804 14764 1900 14804
rect 843 14216 885 14225
rect 843 14176 844 14216
rect 884 14176 885 14216
rect 843 14167 885 14176
rect 1323 14216 1365 14225
rect 1323 14176 1324 14216
rect 1364 14176 1365 14216
rect 1323 14167 1365 14176
rect 1324 14082 1364 14167
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 1516 13964 1556 13973
rect 1804 13964 1844 14764
rect 1900 14755 1940 14764
rect 1556 13924 1844 13964
rect 1516 13915 1556 13924
rect 843 13376 885 13385
rect 843 13336 844 13376
rect 884 13336 885 13376
rect 843 13327 885 13336
rect 1707 13376 1749 13385
rect 1707 13336 1708 13376
rect 1748 13336 1749 13376
rect 1707 13327 1749 13336
rect 844 13292 884 13327
rect 844 13241 884 13252
rect 1708 13242 1748 13327
rect 1804 13292 1844 13924
rect 1900 13292 1940 13301
rect 1804 13252 1900 13292
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 844 12452 884 12461
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 652 12234 692 12319
rect 844 11957 884 12412
rect 1804 12452 1844 13252
rect 1900 13243 1940 13252
rect 1612 12284 1652 12293
rect 843 11948 885 11957
rect 843 11908 844 11948
rect 884 11908 885 11948
rect 843 11899 885 11908
rect 1612 11789 1652 12244
rect 843 11780 885 11789
rect 843 11740 844 11780
rect 884 11740 885 11780
rect 843 11731 885 11740
rect 1611 11780 1653 11789
rect 1611 11740 1612 11780
rect 1652 11740 1653 11780
rect 1611 11731 1653 11740
rect 844 11646 884 11731
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 844 10940 884 10951
rect 1804 10949 1844 12412
rect 1995 11948 2037 11957
rect 1995 11908 1996 11948
rect 2036 11908 2037 11948
rect 1995 11899 2037 11908
rect 1996 11814 2036 11899
rect 1611 10940 1653 10949
rect 844 10865 884 10900
rect 1516 10900 1612 10940
rect 1652 10900 1653 10940
rect 843 10856 885 10865
rect 843 10816 844 10856
rect 884 10816 885 10856
rect 843 10807 885 10816
rect 1419 10856 1461 10865
rect 1419 10816 1420 10856
rect 1460 10816 1461 10856
rect 1419 10807 1461 10816
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 652 10638 692 10723
rect 1420 10722 1460 10807
rect 843 10352 885 10361
rect 843 10312 844 10352
rect 884 10312 885 10352
rect 843 10303 885 10312
rect 1323 10352 1365 10361
rect 1323 10312 1324 10352
rect 1364 10312 1365 10352
rect 1323 10303 1365 10312
rect 844 10268 884 10303
rect 844 10217 884 10228
rect 1324 10218 1364 10303
rect 1516 10268 1556 10900
rect 1611 10891 1653 10900
rect 1803 10940 1845 10949
rect 1803 10900 1804 10940
rect 1844 10900 1845 10940
rect 1803 10891 1845 10900
rect 1612 10806 1652 10891
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 844 9428 884 9439
rect 844 9353 884 9388
rect 1516 9428 1556 10228
rect 1516 9379 1556 9388
rect 843 9344 885 9353
rect 843 9304 844 9344
rect 884 9304 885 9344
rect 843 9295 885 9304
rect 1323 9344 1365 9353
rect 1323 9304 1324 9344
rect 1364 9304 1365 9344
rect 1323 9295 1365 9304
rect 652 9260 692 9269
rect 652 9017 692 9220
rect 1324 9210 1364 9295
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 843 8840 885 8849
rect 843 8800 844 8840
rect 884 8800 885 8840
rect 843 8791 885 8800
rect 1419 8840 1461 8849
rect 1419 8800 1420 8840
rect 1460 8800 1461 8840
rect 1419 8791 1461 8800
rect 844 8756 884 8791
rect 844 8705 884 8716
rect 1420 8706 1460 8791
rect 1612 8756 1652 8765
rect 1996 8756 2036 8765
rect 2092 8756 2132 23239
rect 73036 23120 73076 25255
rect 73324 25229 73364 25768
rect 73505 25724 73545 26040
rect 73505 25684 73556 25724
rect 73516 25229 73556 25684
rect 73615 25640 73655 26040
rect 73905 25892 73945 26040
rect 73612 25600 73655 25640
rect 73804 25852 73945 25892
rect 73323 25220 73365 25229
rect 73323 25180 73324 25220
rect 73364 25180 73365 25220
rect 73323 25171 73365 25180
rect 73515 25220 73557 25229
rect 73515 25180 73516 25220
rect 73556 25180 73557 25220
rect 73515 25171 73557 25180
rect 73323 25052 73365 25061
rect 73323 25012 73324 25052
rect 73364 25012 73365 25052
rect 73323 25003 73365 25012
rect 73131 24128 73173 24137
rect 73131 24088 73132 24128
rect 73172 24088 73173 24128
rect 73131 24079 73173 24088
rect 73132 23288 73172 24079
rect 73132 23239 73172 23248
rect 73036 23071 73076 23080
rect 73324 23120 73364 25003
rect 73420 23288 73460 23297
rect 73612 23288 73652 25600
rect 73804 25397 73844 25852
rect 74015 25808 74055 26040
rect 74305 25901 74345 26040
rect 74304 25892 74346 25901
rect 74304 25852 74305 25892
rect 74345 25852 74346 25892
rect 74304 25843 74346 25852
rect 73996 25768 74055 25808
rect 73899 25724 73941 25733
rect 73899 25684 73900 25724
rect 73940 25684 73941 25724
rect 73899 25675 73941 25684
rect 73803 25388 73845 25397
rect 73803 25348 73804 25388
rect 73844 25348 73845 25388
rect 73803 25339 73845 25348
rect 73460 23248 73652 23288
rect 73420 23239 73460 23248
rect 73364 23080 73844 23120
rect 73324 23071 73364 23080
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 7112 22700 7480 22709
rect 7152 22660 7194 22700
rect 7234 22660 7276 22700
rect 7316 22660 7358 22700
rect 7398 22660 7440 22700
rect 7112 22651 7480 22660
rect 11112 22700 11480 22709
rect 11152 22660 11194 22700
rect 11234 22660 11276 22700
rect 11316 22660 11358 22700
rect 11398 22660 11440 22700
rect 11112 22651 11480 22660
rect 15112 22700 15480 22709
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15112 22651 15480 22660
rect 19112 22700 19480 22709
rect 19152 22660 19194 22700
rect 19234 22660 19276 22700
rect 19316 22660 19358 22700
rect 19398 22660 19440 22700
rect 19112 22651 19480 22660
rect 23112 22700 23480 22709
rect 23152 22660 23194 22700
rect 23234 22660 23276 22700
rect 23316 22660 23358 22700
rect 23398 22660 23440 22700
rect 23112 22651 23480 22660
rect 27112 22700 27480 22709
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27112 22651 27480 22660
rect 31112 22700 31480 22709
rect 31152 22660 31194 22700
rect 31234 22660 31276 22700
rect 31316 22660 31358 22700
rect 31398 22660 31440 22700
rect 31112 22651 31480 22660
rect 35112 22700 35480 22709
rect 35152 22660 35194 22700
rect 35234 22660 35276 22700
rect 35316 22660 35358 22700
rect 35398 22660 35440 22700
rect 35112 22651 35480 22660
rect 39112 22700 39480 22709
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39112 22651 39480 22660
rect 43112 22700 43480 22709
rect 43152 22660 43194 22700
rect 43234 22660 43276 22700
rect 43316 22660 43358 22700
rect 43398 22660 43440 22700
rect 43112 22651 43480 22660
rect 47112 22700 47480 22709
rect 47152 22660 47194 22700
rect 47234 22660 47276 22700
rect 47316 22660 47358 22700
rect 47398 22660 47440 22700
rect 47112 22651 47480 22660
rect 51112 22700 51480 22709
rect 51152 22660 51194 22700
rect 51234 22660 51276 22700
rect 51316 22660 51358 22700
rect 51398 22660 51440 22700
rect 51112 22651 51480 22660
rect 55112 22700 55480 22709
rect 55152 22660 55194 22700
rect 55234 22660 55276 22700
rect 55316 22660 55358 22700
rect 55398 22660 55440 22700
rect 55112 22651 55480 22660
rect 59112 22700 59480 22709
rect 59152 22660 59194 22700
rect 59234 22660 59276 22700
rect 59316 22660 59358 22700
rect 59398 22660 59440 22700
rect 59112 22651 59480 22660
rect 63112 22700 63480 22709
rect 63152 22660 63194 22700
rect 63234 22660 63276 22700
rect 63316 22660 63358 22700
rect 63398 22660 63440 22700
rect 63112 22651 63480 22660
rect 67112 22700 67480 22709
rect 67152 22660 67194 22700
rect 67234 22660 67276 22700
rect 67316 22660 67358 22700
rect 67398 22660 67440 22700
rect 67112 22651 67480 22660
rect 71112 22700 71480 22709
rect 71152 22660 71194 22700
rect 71234 22660 71276 22700
rect 71316 22660 71358 22700
rect 71398 22660 71440 22700
rect 71112 22651 71480 22660
rect 73804 22280 73844 23080
rect 73900 22532 73940 25675
rect 73996 25481 74036 25768
rect 74415 25733 74455 26040
rect 74414 25724 74456 25733
rect 74414 25684 74415 25724
rect 74455 25684 74456 25724
rect 74414 25675 74456 25684
rect 74705 25640 74745 26040
rect 74668 25600 74745 25640
rect 74815 25640 74855 26040
rect 75105 25640 75145 26040
rect 74815 25600 74900 25640
rect 73995 25472 74037 25481
rect 73995 25432 73996 25472
rect 74036 25432 74037 25472
rect 73995 25423 74037 25432
rect 74091 25220 74133 25229
rect 74091 25180 74092 25220
rect 74132 25180 74133 25220
rect 74091 25171 74133 25180
rect 74092 23288 74132 25171
rect 74092 23239 74132 23248
rect 74188 23120 74228 23129
rect 74188 23036 74228 23080
rect 74380 23036 74420 23045
rect 74188 22996 74380 23036
rect 73900 22483 73940 22492
rect 74380 22289 74420 22996
rect 74571 22868 74613 22877
rect 74571 22828 74572 22868
rect 74612 22828 74613 22868
rect 74571 22819 74613 22828
rect 74572 22734 74612 22819
rect 74572 22532 74612 22541
rect 74668 22532 74708 25600
rect 74860 24137 74900 25600
rect 74956 25600 75145 25640
rect 75215 25640 75255 26040
rect 75505 25640 75545 26040
rect 75615 25640 75655 26040
rect 75819 25724 75861 25733
rect 75819 25684 75820 25724
rect 75860 25684 75861 25724
rect 75819 25675 75861 25684
rect 75215 25600 75284 25640
rect 75505 25600 75572 25640
rect 75615 25600 75668 25640
rect 74859 24128 74901 24137
rect 74859 24088 74860 24128
rect 74900 24088 74901 24128
rect 74859 24079 74901 24088
rect 74956 23288 74996 25600
rect 75244 24893 75284 25600
rect 75243 24884 75285 24893
rect 75243 24844 75244 24884
rect 75284 24844 75285 24884
rect 75243 24835 75285 24844
rect 74956 23239 74996 23248
rect 75532 23288 75572 25600
rect 75628 25229 75668 25600
rect 75627 25220 75669 25229
rect 75627 25180 75628 25220
rect 75668 25180 75669 25220
rect 75627 25171 75669 25180
rect 75627 23372 75669 23381
rect 75627 23332 75628 23372
rect 75668 23332 75669 23372
rect 75627 23323 75669 23332
rect 75532 23239 75572 23248
rect 74763 23036 74805 23045
rect 74763 22996 74764 23036
rect 74804 22996 74805 23036
rect 74763 22987 74805 22996
rect 75147 23036 75189 23045
rect 75147 22996 75148 23036
rect 75188 22996 75189 23036
rect 75147 22987 75189 22996
rect 75340 23036 75380 23045
rect 74612 22492 74708 22532
rect 74572 22483 74612 22492
rect 74764 22364 74804 22987
rect 75148 22952 75188 22987
rect 75148 22901 75188 22912
rect 75340 22877 75380 22996
rect 75628 22961 75668 23323
rect 75723 23036 75765 23045
rect 75723 22996 75724 23036
rect 75764 22996 75765 23036
rect 75723 22987 75765 22996
rect 75627 22952 75669 22961
rect 75627 22912 75628 22952
rect 75668 22912 75669 22952
rect 75627 22903 75669 22912
rect 75339 22868 75381 22877
rect 75339 22828 75340 22868
rect 75380 22828 75381 22868
rect 75339 22819 75381 22828
rect 75112 22700 75480 22709
rect 75152 22660 75194 22700
rect 75234 22660 75276 22700
rect 75316 22660 75358 22700
rect 75398 22660 75440 22700
rect 75112 22651 75480 22660
rect 75243 22532 75285 22541
rect 75243 22492 75244 22532
rect 75284 22492 75285 22532
rect 75243 22483 75285 22492
rect 75435 22532 75477 22541
rect 75435 22492 75436 22532
rect 75476 22492 75477 22532
rect 75435 22483 75477 22492
rect 74764 22315 74804 22324
rect 75052 22448 75092 22457
rect 75052 22289 75092 22408
rect 75244 22364 75284 22483
rect 75436 22398 75476 22483
rect 75244 22315 75284 22324
rect 75628 22364 75668 22903
rect 75628 22315 75668 22324
rect 73804 22231 73844 22240
rect 74379 22280 74421 22289
rect 74379 22240 74380 22280
rect 74420 22240 74421 22280
rect 74379 22231 74421 22240
rect 75051 22280 75093 22289
rect 75051 22240 75052 22280
rect 75092 22240 75093 22280
rect 75051 22231 75093 22240
rect 75724 22121 75764 22987
rect 75820 22532 75860 25675
rect 75905 25640 75945 26040
rect 76015 25640 76055 26040
rect 76305 25640 76345 26040
rect 76415 25733 76455 26040
rect 76587 25808 76629 25817
rect 76587 25768 76588 25808
rect 76628 25768 76629 25808
rect 76587 25759 76629 25768
rect 76414 25724 76456 25733
rect 76414 25684 76415 25724
rect 76455 25684 76456 25724
rect 76414 25675 76456 25684
rect 75905 25600 75956 25640
rect 75916 23288 75956 25600
rect 75916 23239 75956 23248
rect 76012 25600 76055 25640
rect 76204 25600 76345 25640
rect 75916 22532 75956 22541
rect 75820 22492 75916 22532
rect 75916 22483 75956 22492
rect 75819 22280 75861 22289
rect 75819 22240 75820 22280
rect 75860 22240 75861 22280
rect 75819 22231 75861 22240
rect 75820 22146 75860 22231
rect 75723 22112 75765 22121
rect 75723 22072 75724 22112
rect 75764 22072 75765 22112
rect 75723 22063 75765 22072
rect 9387 22028 9429 22037
rect 9387 21988 9388 22028
rect 9428 21988 9429 22028
rect 9387 21979 9429 21988
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 8352 21944 8720 21953
rect 8392 21904 8434 21944
rect 8474 21904 8516 21944
rect 8556 21904 8598 21944
rect 8638 21904 8680 21944
rect 8352 21895 8720 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 7112 21188 7480 21197
rect 7152 21148 7194 21188
rect 7234 21148 7276 21188
rect 7316 21148 7358 21188
rect 7398 21148 7440 21188
rect 7112 21139 7480 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 8352 20432 8720 20441
rect 8392 20392 8434 20432
rect 8474 20392 8516 20432
rect 8556 20392 8598 20432
rect 8638 20392 8680 20432
rect 8352 20383 8720 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 7112 19676 7480 19685
rect 7152 19636 7194 19676
rect 7234 19636 7276 19676
rect 7316 19636 7358 19676
rect 7398 19636 7440 19676
rect 7112 19627 7480 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 8352 18920 8720 18929
rect 8392 18880 8434 18920
rect 8474 18880 8516 18920
rect 8556 18880 8598 18920
rect 8638 18880 8680 18920
rect 8352 18871 8720 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 7112 18164 7480 18173
rect 7152 18124 7194 18164
rect 7234 18124 7276 18164
rect 7316 18124 7358 18164
rect 7398 18124 7440 18164
rect 7112 18115 7480 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 8352 17408 8720 17417
rect 8392 17368 8434 17408
rect 8474 17368 8516 17408
rect 8556 17368 8598 17408
rect 8638 17368 8680 17408
rect 8352 17359 8720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 7112 16652 7480 16661
rect 7152 16612 7194 16652
rect 7234 16612 7276 16652
rect 7316 16612 7358 16652
rect 7398 16612 7440 16652
rect 7112 16603 7480 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 8352 15896 8720 15905
rect 8392 15856 8434 15896
rect 8474 15856 8516 15896
rect 8556 15856 8598 15896
rect 8638 15856 8680 15896
rect 8352 15847 8720 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 7112 15140 7480 15149
rect 7152 15100 7194 15140
rect 7234 15100 7276 15140
rect 7316 15100 7358 15140
rect 7398 15100 7440 15140
rect 7112 15091 7480 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 8352 14384 8720 14393
rect 8392 14344 8434 14384
rect 8474 14344 8516 14384
rect 8556 14344 8598 14384
rect 8638 14344 8680 14384
rect 8352 14335 8720 14344
rect 9388 13973 9428 21979
rect 12352 21944 12720 21953
rect 12392 21904 12434 21944
rect 12474 21904 12516 21944
rect 12556 21904 12598 21944
rect 12638 21904 12680 21944
rect 12352 21895 12720 21904
rect 16352 21944 16720 21953
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16352 21895 16720 21904
rect 20352 21944 20720 21953
rect 20392 21904 20434 21944
rect 20474 21904 20516 21944
rect 20556 21904 20598 21944
rect 20638 21904 20680 21944
rect 20352 21895 20720 21904
rect 24352 21944 24720 21953
rect 24392 21904 24434 21944
rect 24474 21904 24516 21944
rect 24556 21904 24598 21944
rect 24638 21904 24680 21944
rect 24352 21895 24720 21904
rect 28352 21944 28720 21953
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28352 21895 28720 21904
rect 32352 21944 32720 21953
rect 32392 21904 32434 21944
rect 32474 21904 32516 21944
rect 32556 21904 32598 21944
rect 32638 21904 32680 21944
rect 32352 21895 32720 21904
rect 36352 21944 36720 21953
rect 36392 21904 36434 21944
rect 36474 21904 36516 21944
rect 36556 21904 36598 21944
rect 36638 21904 36680 21944
rect 36352 21895 36720 21904
rect 40352 21944 40720 21953
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40352 21895 40720 21904
rect 44352 21944 44720 21953
rect 44392 21904 44434 21944
rect 44474 21904 44516 21944
rect 44556 21904 44598 21944
rect 44638 21904 44680 21944
rect 44352 21895 44720 21904
rect 48352 21944 48720 21953
rect 48392 21904 48434 21944
rect 48474 21904 48516 21944
rect 48556 21904 48598 21944
rect 48638 21904 48680 21944
rect 48352 21895 48720 21904
rect 52352 21944 52720 21953
rect 52392 21904 52434 21944
rect 52474 21904 52516 21944
rect 52556 21904 52598 21944
rect 52638 21904 52680 21944
rect 52352 21895 52720 21904
rect 56352 21944 56720 21953
rect 56392 21904 56434 21944
rect 56474 21904 56516 21944
rect 56556 21904 56598 21944
rect 56638 21904 56680 21944
rect 56352 21895 56720 21904
rect 60352 21944 60720 21953
rect 60392 21904 60434 21944
rect 60474 21904 60516 21944
rect 60556 21904 60598 21944
rect 60638 21904 60680 21944
rect 60352 21895 60720 21904
rect 64352 21944 64720 21953
rect 64392 21904 64434 21944
rect 64474 21904 64516 21944
rect 64556 21904 64598 21944
rect 64638 21904 64680 21944
rect 64352 21895 64720 21904
rect 68352 21944 68720 21953
rect 68392 21904 68434 21944
rect 68474 21904 68516 21944
rect 68556 21904 68598 21944
rect 68638 21904 68680 21944
rect 68352 21895 68720 21904
rect 72352 21944 72720 21953
rect 72392 21904 72434 21944
rect 72474 21904 72516 21944
rect 72556 21904 72598 21944
rect 72638 21904 72680 21944
rect 72352 21895 72720 21904
rect 75724 21608 75764 22063
rect 75820 21776 75860 21785
rect 76012 21776 76052 25600
rect 76108 23036 76148 23045
rect 76108 22877 76148 22996
rect 76107 22868 76149 22877
rect 76107 22828 76108 22868
rect 76148 22828 76149 22868
rect 76107 22819 76149 22828
rect 76204 22532 76244 25600
rect 76588 23633 76628 25759
rect 76705 25640 76745 26040
rect 76815 25817 76855 26040
rect 76814 25808 76856 25817
rect 76814 25768 76815 25808
rect 76855 25768 76856 25808
rect 76814 25759 76856 25768
rect 77105 25640 77145 26040
rect 76705 25600 76820 25640
rect 76587 23624 76629 23633
rect 76587 23584 76588 23624
rect 76628 23584 76629 23624
rect 76587 23575 76629 23584
rect 76352 23456 76720 23465
rect 76392 23416 76434 23456
rect 76474 23416 76516 23456
rect 76556 23416 76598 23456
rect 76638 23416 76680 23456
rect 76352 23407 76720 23416
rect 76299 23288 76341 23297
rect 76299 23248 76300 23288
rect 76340 23248 76341 23288
rect 76299 23239 76341 23248
rect 76683 23288 76725 23297
rect 76683 23248 76684 23288
rect 76724 23248 76725 23288
rect 76683 23239 76725 23248
rect 76300 23036 76340 23239
rect 76300 22987 76340 22996
rect 76491 22952 76533 22961
rect 76491 22912 76492 22952
rect 76532 22912 76533 22952
rect 76491 22903 76533 22912
rect 76492 22818 76532 22903
rect 76300 22532 76340 22541
rect 76204 22492 76300 22532
rect 76300 22483 76340 22492
rect 76684 22532 76724 23239
rect 76684 22483 76724 22492
rect 76108 22364 76148 22373
rect 76108 22121 76148 22324
rect 76588 22280 76628 22289
rect 76588 22121 76628 22240
rect 76107 22112 76149 22121
rect 76107 22072 76108 22112
rect 76148 22072 76149 22112
rect 76107 22063 76149 22072
rect 76587 22112 76629 22121
rect 76587 22072 76588 22112
rect 76628 22072 76629 22112
rect 76587 22063 76629 22072
rect 76352 21944 76720 21953
rect 76392 21904 76434 21944
rect 76474 21904 76516 21944
rect 76556 21904 76598 21944
rect 76638 21904 76680 21944
rect 76352 21895 76720 21904
rect 75860 21736 76052 21776
rect 76587 21776 76629 21785
rect 76587 21736 76588 21776
rect 76628 21736 76629 21776
rect 75820 21727 75860 21736
rect 76587 21727 76629 21736
rect 76780 21776 76820 25600
rect 77068 25600 77145 25640
rect 77068 23288 77108 25600
rect 77215 25556 77255 26040
rect 77505 25640 77545 26040
rect 77068 23239 77108 23248
rect 77164 25516 77255 25556
rect 77452 25600 77545 25640
rect 76875 23036 76917 23045
rect 76875 22996 76876 23036
rect 76916 22996 76917 23036
rect 76875 22987 76917 22996
rect 76876 22902 76916 22987
rect 77164 22532 77204 25516
rect 77452 23288 77492 25600
rect 77615 25556 77655 26040
rect 77905 25640 77945 26040
rect 78015 25640 78055 26040
rect 78305 25640 78345 26040
rect 78415 25640 78455 26040
rect 78705 25808 78745 26040
rect 77905 25600 77972 25640
rect 78015 25600 78068 25640
rect 78305 25600 78356 25640
rect 77452 23239 77492 23248
rect 77548 25516 77655 25556
rect 77260 23036 77300 23045
rect 77260 22709 77300 22996
rect 77259 22700 77301 22709
rect 77259 22660 77260 22700
rect 77300 22660 77301 22700
rect 77259 22651 77301 22660
rect 77260 22532 77300 22541
rect 77164 22492 77260 22532
rect 77260 22483 77300 22492
rect 77163 22280 77205 22289
rect 77163 22240 77164 22280
rect 77204 22240 77205 22280
rect 77163 22231 77205 22240
rect 77164 22146 77204 22231
rect 77548 21776 77588 25516
rect 77836 23036 77876 23045
rect 77836 22877 77876 22996
rect 77644 22868 77684 22877
rect 77835 22868 77877 22877
rect 77684 22828 77780 22868
rect 77644 22819 77684 22828
rect 77740 22709 77780 22828
rect 77835 22828 77836 22868
rect 77876 22828 77877 22868
rect 77835 22819 77877 22828
rect 77739 22700 77781 22709
rect 77739 22660 77740 22700
rect 77780 22660 77781 22700
rect 77739 22651 77781 22660
rect 77740 22373 77780 22651
rect 77932 22532 77972 25600
rect 78028 23288 78068 25600
rect 78028 23239 78068 23248
rect 78124 23120 78164 23129
rect 78124 22709 78164 23080
rect 78123 22700 78165 22709
rect 78123 22660 78124 22700
rect 78164 22660 78165 22700
rect 78123 22651 78165 22660
rect 77932 22483 77972 22492
rect 78124 22373 78164 22651
rect 78316 22532 78356 25600
rect 78412 25600 78455 25640
rect 78604 25768 78745 25808
rect 78412 23297 78452 25600
rect 78411 23288 78453 23297
rect 78411 23248 78412 23288
rect 78452 23248 78453 23288
rect 78411 23239 78453 23248
rect 78604 23288 78644 25768
rect 78815 25724 78855 26040
rect 78604 23239 78644 23248
rect 78700 25684 78855 25724
rect 78411 23036 78453 23045
rect 78411 22996 78412 23036
rect 78452 22996 78453 23036
rect 78411 22987 78453 22996
rect 78412 22902 78452 22987
rect 78316 22483 78356 22492
rect 77739 22364 77781 22373
rect 77739 22324 77740 22364
rect 77780 22324 77781 22364
rect 77739 22315 77781 22324
rect 78123 22364 78165 22373
rect 78123 22324 78124 22364
rect 78164 22324 78165 22364
rect 78123 22315 78165 22324
rect 77644 21776 77684 21785
rect 77548 21736 77644 21776
rect 76780 21727 76820 21736
rect 77644 21727 77684 21736
rect 75724 21559 75764 21568
rect 76588 21524 76628 21727
rect 77548 21608 77588 21619
rect 77548 21533 77588 21568
rect 77740 21533 77780 22315
rect 78124 22230 78164 22315
rect 78700 22112 78740 25684
rect 79105 25640 79145 26040
rect 78892 25600 79145 25640
rect 79215 25640 79255 26040
rect 79505 25640 79545 26040
rect 79615 25724 79655 26040
rect 79905 25808 79945 26040
rect 80015 25892 80055 26040
rect 80015 25852 80084 25892
rect 79905 25768 79988 25808
rect 79615 25684 79892 25724
rect 79215 25600 79316 25640
rect 79505 25600 79700 25640
rect 78796 23036 78836 23045
rect 78796 22877 78836 22996
rect 78795 22868 78837 22877
rect 78795 22828 78796 22868
rect 78836 22828 78837 22868
rect 78795 22819 78837 22828
rect 78796 22289 78836 22374
rect 78892 22364 78932 25600
rect 79276 24464 79316 25600
rect 79276 24424 79508 24464
rect 79179 23288 79221 23297
rect 79179 23248 79180 23288
rect 79220 23248 79221 23288
rect 79179 23239 79221 23248
rect 79468 23288 79508 24424
rect 79468 23239 79508 23248
rect 79180 23154 79220 23239
rect 79276 23120 79316 23129
rect 78987 23036 79029 23045
rect 78987 22996 78988 23036
rect 79028 22996 79029 23036
rect 78987 22987 79029 22996
rect 78988 22952 79028 22987
rect 78988 22901 79028 22912
rect 79276 22877 79316 23080
rect 79564 23120 79604 23131
rect 79564 23045 79604 23080
rect 79563 23036 79605 23045
rect 79563 22996 79564 23036
rect 79604 22996 79605 23036
rect 79563 22987 79605 22996
rect 79275 22868 79317 22877
rect 79275 22828 79276 22868
rect 79316 22828 79317 22868
rect 79275 22819 79317 22828
rect 79112 22700 79480 22709
rect 79152 22660 79194 22700
rect 79234 22660 79276 22700
rect 79316 22660 79358 22700
rect 79398 22660 79440 22700
rect 79112 22651 79480 22660
rect 79564 22364 79604 22987
rect 78892 22324 79124 22364
rect 78795 22280 78837 22289
rect 78795 22240 78796 22280
rect 78836 22240 78837 22280
rect 78795 22231 78837 22240
rect 78892 22112 78932 22121
rect 78700 22072 78892 22112
rect 78892 22063 78932 22072
rect 79084 21776 79124 22324
rect 79564 22315 79604 22324
rect 79084 21727 79124 21736
rect 79468 21776 79508 21785
rect 79660 21776 79700 25600
rect 79852 23288 79892 25684
rect 79852 23239 79892 23248
rect 79756 23120 79796 23131
rect 79756 23045 79796 23080
rect 79755 23036 79797 23045
rect 79755 22996 79756 23036
rect 79796 22996 79797 23036
rect 79755 22987 79797 22996
rect 79756 22532 79796 22541
rect 79948 22532 79988 25768
rect 80044 24473 80084 25852
rect 80305 25640 80345 26040
rect 80140 25600 80345 25640
rect 80415 25640 80455 26040
rect 80705 25640 80745 26040
rect 80815 25640 80855 26040
rect 81105 25640 81145 26040
rect 80415 25600 80468 25640
rect 80705 25600 80756 25640
rect 80043 24464 80085 24473
rect 80043 24424 80044 24464
rect 80084 24424 80085 24464
rect 80043 24415 80085 24424
rect 79796 22492 79988 22532
rect 80044 23120 80084 23129
rect 79756 22483 79796 22492
rect 79947 22364 79989 22373
rect 80044 22364 80084 23080
rect 80140 22532 80180 25600
rect 80428 24389 80468 25600
rect 80427 24380 80469 24389
rect 80427 24340 80428 24380
rect 80468 24340 80469 24380
rect 80427 24331 80469 24340
rect 80716 23633 80756 25600
rect 80812 25600 80855 25640
rect 81100 25600 81145 25640
rect 81215 25640 81255 26040
rect 81505 25640 81545 26040
rect 81215 25600 81332 25640
rect 80715 23624 80757 23633
rect 80715 23584 80716 23624
rect 80756 23584 80757 23624
rect 80715 23575 80757 23584
rect 80352 23456 80720 23465
rect 80392 23416 80434 23456
rect 80474 23416 80516 23456
rect 80556 23416 80598 23456
rect 80638 23416 80680 23456
rect 80352 23407 80720 23416
rect 80619 23288 80661 23297
rect 80619 23248 80620 23288
rect 80660 23248 80661 23288
rect 80619 23239 80661 23248
rect 80235 23120 80277 23129
rect 80235 23080 80236 23120
rect 80276 23080 80277 23120
rect 80235 23071 80277 23080
rect 80236 22986 80276 23071
rect 80524 22868 80564 22877
rect 80140 22483 80180 22492
rect 80428 22828 80524 22868
rect 80428 22373 80468 22828
rect 80524 22819 80564 22828
rect 80620 22532 80660 23239
rect 80715 23204 80757 23213
rect 80715 23164 80716 23204
rect 80756 23164 80757 23204
rect 80715 23155 80757 23164
rect 80716 23036 80756 23155
rect 80716 22541 80756 22996
rect 80620 22483 80660 22492
rect 80715 22532 80757 22541
rect 80715 22492 80716 22532
rect 80756 22492 80757 22532
rect 80715 22483 80757 22492
rect 80812 22532 80852 25600
rect 80907 24464 80949 24473
rect 80907 24424 80908 24464
rect 80948 24424 80949 24464
rect 80907 24415 80949 24424
rect 80908 23288 80948 24415
rect 80908 23239 80948 23248
rect 81003 23120 81045 23129
rect 81003 23080 81004 23120
rect 81044 23080 81045 23120
rect 81003 23071 81045 23080
rect 80812 22483 80852 22492
rect 79947 22324 79948 22364
rect 79988 22324 80084 22364
rect 80427 22364 80469 22373
rect 80427 22324 80428 22364
rect 80468 22324 80469 22364
rect 79947 22315 79989 22324
rect 80427 22315 80469 22324
rect 79948 22230 79988 22315
rect 80428 22230 80468 22315
rect 80908 22280 80948 22289
rect 81004 22280 81044 23071
rect 80948 22240 81044 22280
rect 80908 22231 80948 22240
rect 80352 21944 80720 21953
rect 80392 21904 80434 21944
rect 80474 21904 80516 21944
rect 80556 21904 80598 21944
rect 80638 21904 80680 21944
rect 80352 21895 80720 21904
rect 79508 21736 79700 21776
rect 81004 21776 81044 21785
rect 81100 21776 81140 25600
rect 81195 24380 81237 24389
rect 81195 24340 81196 24380
rect 81236 24340 81237 24380
rect 81195 24331 81237 24340
rect 81196 23288 81236 24331
rect 81292 23288 81332 25600
rect 81484 25600 81545 25640
rect 81615 25640 81655 26040
rect 81615 25600 81812 25640
rect 81484 23540 81524 25600
rect 81484 23500 81716 23540
rect 81484 23288 81524 23297
rect 81292 23248 81484 23288
rect 81196 23239 81236 23248
rect 81484 23239 81524 23248
rect 81291 23120 81333 23129
rect 81291 23080 81292 23120
rect 81332 23080 81333 23120
rect 81291 23071 81333 23080
rect 81579 23120 81621 23129
rect 81579 23080 81580 23120
rect 81620 23080 81621 23120
rect 81579 23071 81621 23080
rect 81292 22364 81332 23071
rect 81580 22986 81620 23071
rect 81484 22532 81524 22541
rect 81676 22532 81716 23500
rect 81772 23288 81812 25600
rect 81905 25556 81945 26040
rect 82015 25640 82055 26040
rect 82305 25640 82345 26040
rect 82415 25724 82455 26040
rect 82415 25684 82580 25724
rect 82015 25600 82100 25640
rect 82305 25600 82388 25640
rect 81905 25516 82004 25556
rect 81772 23239 81812 23248
rect 81867 23120 81909 23129
rect 81867 23080 81868 23120
rect 81908 23080 81909 23120
rect 81867 23071 81909 23080
rect 81868 22986 81908 23071
rect 81524 22492 81716 22532
rect 81868 22532 81908 22560
rect 81964 22532 82004 25516
rect 82060 23288 82100 25600
rect 82060 23239 82100 23248
rect 82155 23120 82197 23129
rect 82155 23080 82156 23120
rect 82196 23080 82197 23120
rect 82155 23071 82197 23080
rect 82156 22986 82196 23071
rect 81908 22492 82004 22532
rect 81484 22483 81524 22492
rect 81868 22483 81908 22492
rect 81292 22315 81332 22324
rect 81675 22364 81717 22373
rect 81675 22324 81676 22364
rect 81716 22324 81717 22364
rect 81675 22315 81717 22324
rect 81676 22230 81716 22315
rect 81044 21736 81140 21776
rect 82348 21776 82388 25600
rect 82443 23120 82485 23129
rect 82443 23080 82444 23120
rect 82484 23080 82485 23120
rect 82443 23071 82485 23080
rect 82444 23036 82484 23071
rect 82444 22985 82484 22996
rect 79468 21727 79508 21736
rect 81004 21727 81044 21736
rect 82348 21727 82388 21736
rect 82540 21776 82580 25684
rect 82705 25640 82745 26040
rect 82636 25600 82745 25640
rect 82815 25640 82855 26040
rect 83105 25640 83145 26040
rect 82815 25600 82964 25640
rect 82636 23288 82676 25600
rect 82636 23239 82676 23248
rect 82924 23288 82964 25600
rect 82924 23239 82964 23248
rect 83020 25600 83145 25640
rect 83215 25640 83255 26040
rect 83505 25640 83545 26040
rect 83215 25600 83348 25640
rect 82828 23120 82868 23129
rect 82636 23080 82828 23120
rect 82636 22373 82676 23080
rect 82828 23071 82868 23080
rect 82923 23120 82965 23129
rect 82923 23080 82924 23120
rect 82964 23080 82965 23120
rect 82923 23071 82965 23080
rect 82635 22364 82677 22373
rect 82635 22324 82636 22364
rect 82676 22324 82677 22364
rect 82924 22364 82964 23071
rect 83020 22532 83060 25600
rect 83211 23120 83253 23129
rect 83211 23080 83212 23120
rect 83252 23080 83253 23120
rect 83211 23071 83253 23080
rect 83212 22986 83252 23071
rect 83308 22877 83348 25600
rect 83500 25600 83545 25640
rect 83615 25640 83655 26040
rect 83905 25640 83945 26040
rect 83615 25600 83732 25640
rect 83500 23297 83540 25600
rect 83499 23288 83541 23297
rect 83499 23248 83500 23288
rect 83540 23248 83541 23288
rect 83499 23239 83541 23248
rect 83404 23120 83444 23129
rect 83404 22952 83444 23080
rect 83596 22952 83636 22961
rect 83404 22912 83596 22952
rect 83307 22868 83349 22877
rect 83307 22828 83308 22868
rect 83348 22828 83349 22868
rect 83307 22819 83349 22828
rect 83596 22709 83636 22912
rect 83112 22700 83480 22709
rect 83152 22660 83194 22700
rect 83234 22660 83276 22700
rect 83316 22660 83358 22700
rect 83398 22660 83440 22700
rect 83112 22651 83480 22660
rect 83595 22700 83637 22709
rect 83595 22660 83596 22700
rect 83636 22660 83637 22700
rect 83595 22651 83637 22660
rect 83020 22483 83060 22492
rect 83596 22532 83636 22541
rect 83692 22532 83732 25600
rect 83884 25600 83945 25640
rect 83787 23204 83829 23213
rect 83787 23164 83788 23204
rect 83828 23164 83829 23204
rect 83787 23155 83829 23164
rect 83788 23036 83828 23155
rect 83788 22987 83828 22996
rect 83787 22700 83829 22709
rect 83787 22660 83788 22700
rect 83828 22660 83829 22700
rect 83787 22651 83829 22660
rect 83636 22492 83732 22532
rect 83596 22483 83636 22492
rect 83788 22373 83828 22651
rect 83884 22532 83924 25600
rect 84015 25556 84055 26040
rect 84305 25640 84345 26040
rect 83980 25516 84055 25556
rect 84268 25600 84345 25640
rect 84415 25640 84455 26040
rect 84705 25733 84745 26040
rect 84704 25724 84746 25733
rect 84704 25684 84705 25724
rect 84745 25684 84746 25724
rect 84704 25675 84746 25684
rect 84815 25640 84855 26040
rect 84939 25724 84981 25733
rect 84939 25684 84940 25724
rect 84980 25684 84981 25724
rect 84939 25675 84981 25684
rect 84415 25600 84500 25640
rect 84815 25600 84884 25640
rect 83980 23045 84020 25516
rect 84268 23801 84308 25600
rect 84267 23792 84309 23801
rect 84267 23752 84268 23792
rect 84308 23752 84309 23792
rect 84267 23743 84309 23752
rect 84460 23624 84500 25600
rect 84268 23584 84500 23624
rect 84268 23288 84308 23584
rect 84352 23456 84720 23465
rect 84392 23416 84434 23456
rect 84474 23416 84516 23456
rect 84556 23416 84598 23456
rect 84638 23416 84680 23456
rect 84352 23407 84720 23416
rect 84460 23288 84500 23297
rect 84268 23248 84460 23288
rect 84460 23239 84500 23248
rect 84844 23288 84884 25600
rect 84844 23239 84884 23248
rect 84075 23120 84117 23129
rect 84363 23120 84405 23129
rect 84075 23080 84076 23120
rect 84116 23080 84212 23120
rect 84075 23071 84117 23080
rect 83979 23036 84021 23045
rect 83979 22996 83980 23036
rect 84020 22996 84021 23036
rect 83979 22987 84021 22996
rect 84076 22986 84116 23071
rect 83979 22868 84021 22877
rect 83979 22828 83980 22868
rect 84020 22828 84021 22868
rect 83979 22819 84021 22828
rect 83980 22734 84020 22819
rect 83980 22532 84020 22541
rect 83884 22492 83980 22532
rect 83980 22483 84020 22492
rect 83212 22364 83252 22373
rect 83595 22364 83637 22373
rect 82924 22324 83212 22364
rect 83252 22324 83540 22364
rect 82635 22315 82677 22324
rect 83212 22315 83252 22324
rect 82540 21727 82580 21736
rect 82636 21608 82676 22315
rect 83500 22280 83540 22324
rect 83595 22324 83596 22364
rect 83636 22324 83637 22364
rect 83595 22315 83637 22324
rect 83787 22364 83829 22373
rect 83787 22324 83788 22364
rect 83828 22324 83829 22364
rect 83787 22315 83829 22324
rect 83500 22231 83540 22240
rect 83596 21776 83636 22315
rect 83596 21727 83636 21736
rect 82636 21533 82676 21568
rect 83788 21533 83828 22315
rect 84172 22280 84212 23080
rect 84363 23080 84364 23120
rect 84404 23080 84405 23120
rect 84363 23071 84405 23080
rect 84747 23120 84789 23129
rect 84747 23080 84748 23120
rect 84788 23080 84789 23120
rect 84747 23071 84789 23080
rect 84267 23036 84309 23045
rect 84267 22996 84268 23036
rect 84308 22996 84309 23036
rect 84267 22987 84309 22996
rect 84268 22448 84308 22987
rect 84364 22986 84404 23071
rect 84748 22986 84788 23071
rect 84748 22532 84788 22541
rect 84940 22532 84980 25675
rect 85105 25640 85145 26040
rect 84788 22492 84980 22532
rect 85036 25600 85145 25640
rect 85215 25640 85255 26040
rect 85505 25724 85545 26040
rect 85420 25684 85545 25724
rect 85215 25600 85268 25640
rect 85036 22532 85076 25600
rect 85228 23288 85268 25600
rect 85420 23969 85460 25684
rect 85615 25640 85655 26040
rect 85516 25600 85655 25640
rect 85905 25640 85945 26040
rect 86015 25724 86055 26040
rect 86305 25724 86345 26040
rect 86015 25684 86228 25724
rect 85905 25600 86036 25640
rect 85419 23960 85461 23969
rect 85419 23920 85420 23960
rect 85460 23920 85461 23960
rect 85419 23911 85461 23920
rect 85228 23239 85268 23248
rect 85516 23288 85556 25600
rect 85516 23239 85556 23248
rect 85803 23204 85845 23213
rect 85803 23164 85804 23204
rect 85844 23164 85845 23204
rect 85803 23155 85845 23164
rect 85131 23120 85173 23129
rect 85131 23080 85132 23120
rect 85172 23080 85173 23120
rect 85131 23071 85173 23080
rect 85419 23120 85461 23129
rect 85419 23080 85420 23120
rect 85460 23080 85461 23120
rect 85419 23071 85461 23080
rect 85132 22986 85172 23071
rect 85420 22986 85460 23071
rect 85707 23036 85749 23045
rect 85707 22996 85708 23036
rect 85748 22996 85749 23036
rect 85707 22987 85749 22996
rect 85708 22902 85748 22987
rect 85132 22532 85172 22541
rect 85036 22492 85132 22532
rect 84748 22483 84788 22492
rect 85132 22483 85172 22492
rect 85419 22532 85461 22541
rect 85419 22492 85420 22532
rect 85460 22492 85461 22532
rect 85804 22532 85844 23155
rect 85900 22868 85940 22877
rect 85900 22709 85940 22828
rect 85899 22700 85941 22709
rect 85899 22660 85900 22700
rect 85940 22660 85941 22700
rect 85899 22651 85941 22660
rect 85996 22532 86036 25600
rect 86092 23036 86132 23045
rect 86092 22709 86132 22996
rect 86091 22700 86133 22709
rect 86091 22660 86092 22700
rect 86132 22660 86133 22700
rect 86091 22651 86133 22660
rect 85804 22492 85940 22532
rect 85419 22483 85461 22492
rect 84268 22408 84404 22448
rect 84268 22280 84308 22289
rect 84172 22240 84268 22280
rect 84268 22231 84308 22240
rect 84172 22112 84212 22121
rect 84364 22112 84404 22408
rect 85420 22398 85460 22483
rect 84555 22364 84597 22373
rect 84555 22324 84556 22364
rect 84596 22324 84597 22364
rect 84555 22315 84597 22324
rect 84939 22364 84981 22373
rect 84939 22324 84940 22364
rect 84980 22324 84981 22364
rect 84939 22315 84981 22324
rect 85611 22364 85653 22373
rect 85611 22324 85612 22364
rect 85652 22324 85653 22364
rect 85611 22315 85653 22324
rect 85803 22364 85845 22373
rect 85803 22324 85804 22364
rect 85844 22324 85845 22364
rect 85803 22315 85845 22324
rect 84556 22230 84596 22315
rect 84940 22230 84980 22315
rect 85612 22230 85652 22315
rect 85804 22230 85844 22315
rect 84212 22072 84404 22112
rect 84172 22063 84212 22072
rect 84352 21944 84720 21953
rect 84392 21904 84434 21944
rect 84474 21904 84516 21944
rect 84556 21904 84598 21944
rect 84638 21904 84680 21944
rect 84352 21895 84720 21904
rect 84363 21776 84405 21785
rect 84363 21736 84364 21776
rect 84404 21736 84405 21776
rect 84363 21727 84405 21736
rect 84364 21642 84404 21727
rect 85900 21608 85940 22492
rect 85996 22483 86036 22492
rect 86188 22364 86228 25684
rect 86284 25684 86345 25724
rect 86284 23288 86324 25684
rect 86415 25640 86455 26040
rect 86284 23239 86324 23248
rect 86380 25600 86455 25640
rect 86283 23036 86325 23045
rect 86283 22996 86284 23036
rect 86324 22996 86325 23036
rect 86283 22987 86325 22996
rect 85996 22324 86228 22364
rect 85996 21776 86036 22324
rect 86284 22289 86324 22987
rect 86380 22532 86420 25600
rect 86705 25556 86745 26040
rect 86815 25640 86855 26040
rect 87105 25640 87145 26040
rect 87215 25733 87255 26040
rect 87214 25724 87256 25733
rect 87214 25684 87215 25724
rect 87255 25684 87256 25724
rect 87214 25675 87256 25684
rect 87505 25640 87545 26040
rect 86815 25600 86900 25640
rect 87105 25600 87188 25640
rect 86705 25516 86804 25556
rect 86476 23120 86516 23129
rect 86476 22961 86516 23080
rect 86667 23120 86709 23129
rect 86667 23080 86668 23120
rect 86708 23080 86709 23120
rect 86667 23071 86709 23080
rect 86475 22952 86517 22961
rect 86475 22912 86476 22952
rect 86516 22912 86517 22952
rect 86475 22903 86517 22912
rect 86571 22700 86613 22709
rect 86571 22660 86572 22700
rect 86612 22660 86613 22700
rect 86571 22651 86613 22660
rect 86380 22492 86516 22532
rect 86379 22364 86421 22373
rect 86379 22324 86380 22364
rect 86420 22324 86421 22364
rect 86379 22315 86421 22324
rect 86283 22280 86325 22289
rect 86188 22240 86284 22280
rect 86324 22240 86325 22280
rect 86188 22112 86228 22240
rect 86283 22231 86325 22240
rect 86380 22230 86420 22315
rect 86188 22063 86228 22072
rect 85996 21727 86036 21736
rect 86380 21776 86420 21785
rect 86476 21776 86516 22492
rect 86572 22373 86612 22651
rect 86668 22457 86708 23071
rect 86764 22532 86804 25516
rect 86764 22483 86804 22492
rect 86667 22448 86709 22457
rect 86667 22408 86668 22448
rect 86708 22408 86709 22448
rect 86667 22399 86709 22408
rect 86571 22364 86613 22373
rect 86571 22324 86572 22364
rect 86612 22324 86613 22364
rect 86571 22315 86613 22324
rect 86420 21736 86516 21776
rect 86380 21727 86420 21736
rect 85900 21559 85940 21568
rect 86476 21608 86516 21617
rect 86572 21608 86612 22315
rect 86860 21776 86900 25600
rect 87148 23288 87188 25600
rect 87148 23239 87188 23248
rect 87436 25600 87545 25640
rect 87615 25640 87655 26040
rect 87723 25724 87765 25733
rect 87723 25684 87724 25724
rect 87764 25684 87765 25724
rect 87723 25675 87765 25684
rect 87615 25600 87668 25640
rect 86956 23036 86996 23045
rect 86956 22709 86996 22996
rect 87340 22877 87380 22962
rect 87339 22868 87381 22877
rect 87339 22828 87340 22868
rect 87380 22828 87381 22868
rect 87436 22868 87476 25600
rect 87532 23045 87572 23130
rect 87531 23036 87573 23045
rect 87531 22996 87532 23036
rect 87572 22996 87573 23036
rect 87531 22987 87573 22996
rect 87436 22828 87572 22868
rect 87339 22819 87381 22828
rect 86955 22700 86997 22709
rect 86955 22660 86956 22700
rect 86996 22660 86997 22700
rect 86955 22651 86997 22660
rect 87112 22700 87480 22709
rect 87152 22660 87194 22700
rect 87234 22660 87276 22700
rect 87316 22660 87358 22700
rect 87398 22660 87440 22700
rect 87112 22651 87480 22660
rect 87051 22532 87093 22541
rect 87051 22492 87052 22532
rect 87092 22492 87093 22532
rect 87051 22483 87093 22492
rect 87436 22532 87476 22541
rect 87532 22532 87572 22828
rect 87628 22541 87668 25600
rect 87724 23288 87764 25675
rect 87905 25640 87945 26040
rect 88015 25640 88055 26040
rect 88305 25808 88345 26040
rect 87905 25600 87956 25640
rect 87724 23239 87764 23248
rect 87820 23120 87860 23129
rect 87723 23036 87765 23045
rect 87723 22996 87724 23036
rect 87764 22996 87765 23036
rect 87723 22987 87765 22996
rect 87476 22492 87572 22532
rect 87627 22532 87669 22541
rect 87627 22492 87628 22532
rect 87668 22492 87669 22532
rect 87436 22483 87476 22492
rect 87627 22483 87669 22492
rect 87052 22398 87092 22483
rect 87244 22364 87284 22373
rect 86955 22280 86997 22289
rect 86955 22240 86956 22280
rect 86996 22240 86997 22280
rect 86955 22231 86997 22240
rect 86956 22146 86996 22231
rect 87244 22205 87284 22324
rect 87627 22364 87669 22373
rect 87627 22324 87628 22364
rect 87668 22324 87669 22364
rect 87627 22315 87669 22324
rect 87628 22230 87668 22315
rect 87724 22289 87764 22987
rect 87820 22877 87860 23080
rect 87819 22868 87861 22877
rect 87819 22828 87820 22868
rect 87860 22828 87861 22868
rect 87819 22819 87861 22828
rect 87820 22532 87860 22541
rect 87916 22532 87956 25600
rect 88012 25600 88055 25640
rect 88204 25768 88345 25808
rect 88012 23288 88052 25600
rect 88012 23239 88052 23248
rect 88108 23120 88148 23129
rect 88108 22877 88148 23080
rect 88107 22868 88149 22877
rect 88107 22828 88108 22868
rect 88148 22828 88149 22868
rect 88107 22819 88149 22828
rect 87860 22492 87956 22532
rect 88204 22532 88244 25768
rect 88415 25640 88455 26040
rect 88705 25640 88745 26040
rect 88396 25600 88455 25640
rect 88684 25600 88745 25640
rect 88815 25640 88855 26040
rect 89105 25640 89145 26040
rect 88815 25600 88916 25640
rect 88396 23633 88436 25600
rect 88395 23624 88437 23633
rect 88395 23584 88396 23624
rect 88436 23584 88437 23624
rect 88684 23624 88724 25600
rect 88684 23584 88820 23624
rect 88395 23575 88437 23584
rect 88352 23456 88720 23465
rect 88392 23416 88434 23456
rect 88474 23416 88516 23456
rect 88556 23416 88598 23456
rect 88638 23416 88680 23456
rect 88352 23407 88720 23416
rect 88395 23288 88437 23297
rect 88780 23288 88820 23584
rect 88395 23248 88396 23288
rect 88436 23248 88437 23288
rect 88395 23239 88437 23248
rect 88588 23248 88820 23288
rect 88876 23288 88916 25600
rect 88396 23154 88436 23239
rect 88492 23120 88532 23129
rect 88492 22877 88532 23080
rect 88491 22868 88533 22877
rect 88491 22828 88492 22868
rect 88532 22828 88533 22868
rect 88491 22819 88533 22828
rect 87820 22483 87860 22492
rect 88204 22483 88244 22492
rect 88588 22532 88628 23248
rect 88876 23239 88916 23248
rect 89068 25600 89145 25640
rect 88780 23120 88820 23129
rect 88780 22877 88820 23080
rect 88779 22868 88821 22877
rect 88779 22828 88780 22868
rect 88820 22828 88821 22868
rect 88779 22819 88821 22828
rect 88588 22483 88628 22492
rect 89068 22532 89108 25600
rect 89215 25556 89255 26040
rect 89505 25640 89545 26040
rect 89615 25724 89655 26040
rect 89615 25684 89684 25724
rect 89505 25600 89588 25640
rect 89068 22483 89108 22492
rect 89164 25516 89255 25556
rect 88012 22364 88052 22373
rect 87723 22280 87765 22289
rect 87723 22240 87724 22280
rect 87764 22240 87765 22280
rect 87723 22231 87765 22240
rect 88012 22205 88052 22324
rect 88395 22364 88437 22373
rect 88395 22324 88396 22364
rect 88436 22324 88437 22364
rect 88395 22315 88437 22324
rect 88875 22364 88917 22373
rect 88875 22324 88876 22364
rect 88916 22324 88917 22364
rect 88875 22315 88917 22324
rect 88396 22230 88436 22315
rect 88876 22230 88916 22315
rect 87243 22196 87285 22205
rect 87243 22156 87244 22196
rect 87284 22156 87285 22196
rect 87243 22147 87285 22156
rect 88011 22196 88053 22205
rect 88011 22156 88012 22196
rect 88052 22156 88053 22196
rect 88011 22147 88053 22156
rect 88352 21944 88720 21953
rect 88392 21904 88434 21944
rect 88474 21904 88516 21944
rect 88556 21904 88598 21944
rect 88638 21904 88680 21944
rect 88352 21895 88720 21904
rect 86860 21727 86900 21736
rect 89068 21776 89108 21785
rect 89164 21776 89204 25516
rect 89355 23288 89397 23297
rect 89355 23248 89356 23288
rect 89396 23248 89397 23288
rect 89355 23239 89397 23248
rect 89356 23154 89396 23239
rect 89451 23120 89493 23129
rect 89451 23080 89452 23120
rect 89492 23080 89493 23120
rect 89451 23071 89493 23080
rect 89452 22986 89492 23071
rect 89355 22532 89397 22541
rect 89355 22492 89356 22532
rect 89396 22492 89397 22532
rect 89355 22483 89397 22492
rect 89108 21736 89204 21776
rect 89068 21727 89108 21736
rect 86764 21608 86804 21617
rect 86516 21568 86764 21608
rect 86476 21559 86516 21568
rect 86764 21559 86804 21568
rect 89164 21608 89204 21617
rect 89356 21608 89396 22483
rect 89548 21776 89588 25600
rect 89644 23297 89684 25684
rect 89905 25640 89945 26040
rect 90015 25733 90055 26040
rect 90014 25724 90056 25733
rect 90014 25684 90015 25724
rect 90055 25684 90056 25724
rect 90014 25675 90056 25684
rect 90305 25640 90345 26040
rect 90415 25640 90455 26040
rect 90507 25724 90549 25733
rect 90507 25684 90508 25724
rect 90548 25684 90549 25724
rect 90507 25675 90549 25684
rect 89905 25600 89972 25640
rect 89643 23288 89685 23297
rect 89643 23248 89644 23288
rect 89684 23248 89685 23288
rect 89643 23239 89685 23248
rect 89644 23120 89684 23129
rect 89835 23120 89877 23129
rect 89684 23080 89780 23120
rect 89644 23071 89684 23080
rect 89740 22541 89780 23080
rect 89835 23080 89836 23120
rect 89876 23080 89877 23120
rect 89835 23071 89877 23080
rect 89836 22986 89876 23071
rect 89739 22532 89781 22541
rect 89739 22492 89740 22532
rect 89780 22492 89781 22532
rect 89739 22483 89781 22492
rect 89932 22532 89972 25600
rect 90220 25600 90345 25640
rect 90412 25600 90455 25640
rect 90124 22868 90164 22877
rect 90124 22541 90164 22828
rect 89932 22483 89972 22492
rect 90123 22532 90165 22541
rect 90123 22492 90124 22532
rect 90164 22492 90165 22532
rect 90123 22483 90165 22492
rect 90220 22532 90260 25600
rect 90412 23969 90452 25600
rect 90411 23960 90453 23969
rect 90411 23920 90412 23960
rect 90452 23920 90453 23960
rect 90411 23911 90453 23920
rect 90508 23288 90548 25675
rect 90705 25640 90745 26040
rect 90604 25600 90745 25640
rect 90815 25640 90855 26040
rect 91105 25640 91145 26040
rect 90815 25600 91028 25640
rect 90604 23288 90644 25600
rect 90988 23960 91028 25600
rect 91084 25600 91145 25640
rect 91215 25640 91255 26040
rect 91505 25640 91545 26040
rect 91615 25724 91655 26040
rect 91905 25901 91945 26040
rect 91904 25892 91946 25901
rect 91904 25852 91905 25892
rect 91945 25852 91946 25892
rect 92015 25892 92055 26040
rect 92139 25892 92181 25901
rect 92015 25852 92084 25892
rect 91904 25843 91946 25852
rect 91615 25684 91988 25724
rect 91215 25600 91316 25640
rect 91505 25600 91604 25640
rect 91084 24968 91124 25600
rect 91084 24928 91220 24968
rect 90988 23920 91124 23960
rect 90795 23876 90837 23885
rect 90795 23836 90796 23876
rect 90836 23836 90837 23876
rect 90795 23827 90837 23836
rect 90796 23288 90836 23827
rect 90604 23248 90740 23288
rect 90508 23239 90548 23248
rect 90507 23120 90549 23129
rect 90604 23120 90644 23148
rect 90507 23080 90508 23120
rect 90548 23080 90604 23120
rect 90507 23071 90549 23080
rect 90604 23071 90644 23080
rect 90315 23036 90357 23045
rect 90315 22996 90316 23036
rect 90356 22996 90357 23036
rect 90315 22987 90357 22996
rect 90316 22877 90356 22987
rect 90315 22868 90357 22877
rect 90315 22828 90316 22868
rect 90356 22828 90357 22868
rect 90315 22819 90357 22828
rect 90220 22483 90260 22492
rect 89740 22364 89780 22483
rect 89740 22315 89780 22324
rect 90412 22364 90452 22392
rect 90508 22373 90548 23071
rect 90603 22532 90645 22541
rect 90603 22492 90604 22532
rect 90644 22492 90645 22532
rect 90700 22532 90740 23248
rect 90796 23239 90836 23248
rect 91084 23288 91124 23920
rect 91180 23297 91220 24928
rect 91084 23239 91124 23248
rect 91179 23288 91221 23297
rect 91179 23248 91180 23288
rect 91220 23248 91221 23288
rect 91179 23239 91221 23248
rect 90892 23129 90932 23214
rect 90891 23120 90933 23129
rect 90891 23080 90892 23120
rect 90932 23080 90933 23120
rect 90891 23071 90933 23080
rect 91179 23120 91221 23129
rect 91179 23080 91180 23120
rect 91220 23080 91221 23120
rect 91179 23071 91221 23080
rect 91180 22986 91220 23071
rect 90891 22868 90933 22877
rect 91276 22868 91316 25600
rect 91371 25220 91413 25229
rect 91371 25180 91372 25220
rect 91412 25180 91413 25220
rect 91371 25171 91413 25180
rect 91372 23288 91412 25171
rect 91468 23288 91508 23297
rect 91372 23248 91468 23288
rect 91468 23239 91508 23248
rect 91372 23120 91412 23129
rect 91372 22877 91412 23080
rect 90891 22828 90892 22868
rect 90932 22828 90933 22868
rect 90891 22819 90933 22828
rect 90988 22828 91316 22868
rect 91371 22868 91413 22877
rect 91371 22828 91372 22868
rect 91412 22828 91413 22868
rect 90796 22532 90836 22541
rect 90700 22492 90796 22532
rect 90603 22483 90645 22492
rect 90796 22483 90836 22492
rect 90507 22364 90549 22373
rect 90452 22324 90508 22364
rect 90548 22324 90549 22364
rect 90412 22315 90452 22324
rect 90507 22315 90549 22324
rect 90604 22364 90644 22483
rect 90604 22315 90644 22324
rect 89548 21727 89588 21736
rect 89204 21568 89396 21608
rect 90892 21608 90932 22819
rect 90988 22532 91028 22828
rect 91371 22819 91413 22828
rect 91112 22700 91480 22709
rect 91152 22660 91194 22700
rect 91234 22660 91276 22700
rect 91316 22660 91358 22700
rect 91398 22660 91440 22700
rect 91112 22651 91480 22660
rect 91275 22532 91317 22541
rect 90988 22492 91220 22532
rect 90987 22364 91029 22373
rect 90987 22324 90988 22364
rect 91028 22324 91029 22364
rect 90987 22315 91029 22324
rect 90988 22280 91028 22315
rect 90988 22229 91028 22240
rect 91083 22280 91125 22289
rect 91083 22240 91084 22280
rect 91124 22240 91125 22280
rect 91083 22231 91125 22240
rect 91084 22146 91124 22231
rect 91180 21776 91220 22492
rect 91275 22492 91276 22532
rect 91316 22492 91317 22532
rect 91275 22483 91317 22492
rect 91468 22532 91508 22541
rect 91564 22532 91604 25600
rect 91755 23288 91797 23297
rect 91755 23248 91756 23288
rect 91796 23248 91797 23288
rect 91755 23239 91797 23248
rect 91659 23204 91701 23213
rect 91659 23164 91660 23204
rect 91700 23164 91701 23204
rect 91659 23155 91701 23164
rect 91660 23036 91700 23155
rect 91660 22987 91700 22996
rect 91508 22492 91604 22532
rect 91660 22532 91700 22541
rect 91756 22532 91796 23239
rect 91851 23036 91893 23045
rect 91851 22996 91852 23036
rect 91892 22996 91893 23036
rect 91851 22987 91893 22996
rect 91852 22952 91892 22987
rect 91852 22901 91892 22912
rect 91700 22492 91796 22532
rect 91468 22483 91508 22492
rect 91660 22483 91700 22492
rect 91276 22364 91316 22483
rect 91851 22448 91893 22457
rect 91851 22408 91852 22448
rect 91892 22408 91893 22448
rect 91851 22399 91893 22408
rect 91276 22315 91316 22324
rect 91852 22364 91892 22399
rect 91852 22313 91892 22324
rect 91948 22289 91988 25684
rect 92044 25229 92084 25852
rect 92139 25852 92140 25892
rect 92180 25852 92181 25892
rect 92139 25843 92181 25852
rect 92043 25220 92085 25229
rect 92043 25180 92044 25220
rect 92084 25180 92085 25220
rect 92043 25171 92085 25180
rect 92043 23036 92085 23045
rect 92043 22996 92044 23036
rect 92084 22996 92085 23036
rect 92043 22987 92085 22996
rect 92044 22902 92084 22987
rect 92044 22532 92084 22541
rect 92140 22532 92180 25843
rect 92305 25640 92345 26040
rect 92236 25600 92345 25640
rect 92415 25640 92455 26040
rect 92705 25640 92745 26040
rect 92815 25724 92855 26040
rect 92815 25684 93044 25724
rect 92415 25600 92468 25640
rect 92705 25600 92852 25640
rect 92236 23036 92276 25600
rect 92428 24053 92468 25600
rect 92427 24044 92469 24053
rect 92427 24004 92428 24044
rect 92468 24004 92469 24044
rect 92427 23995 92469 24004
rect 92352 23456 92720 23465
rect 92392 23416 92434 23456
rect 92474 23416 92516 23456
rect 92556 23416 92598 23456
rect 92638 23416 92680 23456
rect 92352 23407 92720 23416
rect 92428 23036 92468 23045
rect 92236 22996 92372 23036
rect 92236 22868 92276 22877
rect 92236 22625 92276 22828
rect 92235 22616 92277 22625
rect 92235 22576 92236 22616
rect 92276 22576 92277 22616
rect 92235 22567 92277 22576
rect 92084 22492 92180 22532
rect 92332 22532 92372 22996
rect 92468 22996 92564 23036
rect 92428 22987 92468 22996
rect 92524 22625 92564 22996
rect 92620 22868 92660 22877
rect 92620 22709 92660 22828
rect 92619 22700 92661 22709
rect 92619 22660 92620 22700
rect 92660 22660 92661 22700
rect 92619 22651 92661 22660
rect 92523 22616 92565 22625
rect 92523 22576 92524 22616
rect 92564 22576 92565 22616
rect 92523 22567 92565 22576
rect 92428 22532 92468 22541
rect 92332 22492 92428 22532
rect 92044 22483 92084 22492
rect 92428 22483 92468 22492
rect 92235 22364 92277 22373
rect 92235 22324 92236 22364
rect 92276 22324 92277 22364
rect 92524 22364 92564 22567
rect 92812 22532 92852 25600
rect 92908 23036 92948 23045
rect 92908 22709 92948 22996
rect 92907 22700 92949 22709
rect 92907 22660 92908 22700
rect 92948 22660 92949 22700
rect 92907 22651 92949 22660
rect 93004 22532 93044 25684
rect 93105 25640 93145 26040
rect 93100 25600 93145 25640
rect 93215 25640 93255 26040
rect 93505 25640 93545 26040
rect 93215 25600 93428 25640
rect 93100 23288 93140 25600
rect 93100 23239 93140 23248
rect 93292 23036 93332 23045
rect 93292 22709 93332 22996
rect 93099 22700 93141 22709
rect 93099 22660 93100 22700
rect 93140 22660 93141 22700
rect 93099 22651 93141 22660
rect 93291 22700 93333 22709
rect 93291 22660 93292 22700
rect 93332 22660 93333 22700
rect 93291 22651 93333 22660
rect 92812 22483 92852 22492
rect 92908 22492 93044 22532
rect 92620 22364 92660 22373
rect 92524 22324 92620 22364
rect 92235 22315 92277 22324
rect 91947 22280 91989 22289
rect 91947 22240 91948 22280
rect 91988 22240 91989 22280
rect 91947 22231 91989 22240
rect 92236 22230 92276 22315
rect 92620 22121 92660 22324
rect 92619 22112 92661 22121
rect 92619 22072 92620 22112
rect 92660 22072 92661 22112
rect 92619 22063 92661 22072
rect 92352 21944 92720 21953
rect 92392 21904 92434 21944
rect 92474 21904 92516 21944
rect 92556 21904 92598 21944
rect 92638 21904 92680 21944
rect 92352 21895 92720 21904
rect 91180 21727 91220 21736
rect 92812 21776 92852 21785
rect 92908 21776 92948 22492
rect 93004 22364 93044 22373
rect 93100 22364 93140 22651
rect 93044 22324 93140 22364
rect 93004 22315 93044 22324
rect 92852 21736 92948 21776
rect 93292 21776 93332 21785
rect 93388 21776 93428 25600
rect 93484 25600 93545 25640
rect 93615 25640 93655 26040
rect 93905 25640 93945 26040
rect 93615 25600 93716 25640
rect 93484 23288 93524 25600
rect 93579 23876 93621 23885
rect 93579 23836 93580 23876
rect 93620 23836 93621 23876
rect 93579 23827 93621 23836
rect 93484 23239 93524 23248
rect 93580 23120 93620 23827
rect 93676 23297 93716 25600
rect 93868 25600 93945 25640
rect 94015 25640 94055 26040
rect 94305 25640 94345 26040
rect 94415 25724 94455 26040
rect 94415 25684 94580 25724
rect 94015 25600 94196 25640
rect 94305 25600 94388 25640
rect 93675 23288 93717 23297
rect 93675 23248 93676 23288
rect 93716 23248 93717 23288
rect 93675 23239 93717 23248
rect 93676 23120 93716 23129
rect 93580 23080 93676 23120
rect 93676 23071 93716 23080
rect 93772 23120 93812 23129
rect 93483 23036 93525 23045
rect 93483 22996 93484 23036
rect 93524 22996 93525 23036
rect 93483 22987 93525 22996
rect 93484 22541 93524 22987
rect 93772 22709 93812 23080
rect 93771 22700 93813 22709
rect 93771 22660 93772 22700
rect 93812 22660 93813 22700
rect 93771 22651 93813 22660
rect 93483 22532 93525 22541
rect 93483 22492 93484 22532
rect 93524 22492 93525 22532
rect 93868 22532 93908 25600
rect 93963 23288 94005 23297
rect 93963 23248 93964 23288
rect 94004 23248 94005 23288
rect 93963 23239 94005 23248
rect 93964 23154 94004 23239
rect 94060 23120 94100 23129
rect 94060 22709 94100 23080
rect 94059 22700 94101 22709
rect 94059 22660 94060 22700
rect 94100 22660 94101 22700
rect 94059 22651 94101 22660
rect 93964 22532 94004 22541
rect 94156 22532 94196 25600
rect 93868 22492 93964 22532
rect 93483 22483 93525 22492
rect 93964 22483 94004 22492
rect 94060 22492 94196 22532
rect 94348 22532 94388 25600
rect 94444 23036 94484 23045
rect 94444 22709 94484 22996
rect 94443 22700 94485 22709
rect 94443 22660 94444 22700
rect 94484 22660 94485 22700
rect 94443 22651 94485 22660
rect 93484 22280 93524 22483
rect 93772 22373 93812 22458
rect 93771 22364 93813 22373
rect 93771 22324 93772 22364
rect 93812 22324 93813 22364
rect 93771 22315 93813 22324
rect 94060 22280 94100 22492
rect 94348 22483 94388 22492
rect 93484 22231 93524 22240
rect 93964 22240 94100 22280
rect 94156 22364 94196 22373
rect 94156 22280 94196 22324
rect 94444 22280 94484 22651
rect 94540 22532 94580 25684
rect 94705 25640 94745 26040
rect 94636 25600 94745 25640
rect 94815 25640 94855 26040
rect 95105 25817 95145 26040
rect 95104 25808 95146 25817
rect 95104 25768 95105 25808
rect 95145 25768 95146 25808
rect 95104 25759 95146 25768
rect 95215 25733 95255 26040
rect 95505 25808 95545 26040
rect 95615 25892 95655 26040
rect 95615 25852 95732 25892
rect 95505 25768 95636 25808
rect 95214 25724 95256 25733
rect 95214 25684 95215 25724
rect 95255 25684 95256 25724
rect 95214 25675 95256 25684
rect 94815 25600 94868 25640
rect 94636 23288 94676 25600
rect 94636 23239 94676 23248
rect 94828 23288 94868 25600
rect 95403 24716 95445 24725
rect 95403 24676 95404 24716
rect 95444 24676 95445 24716
rect 95403 24667 95445 24676
rect 94828 23239 94868 23248
rect 95404 23288 95444 24667
rect 95404 23239 95444 23248
rect 95308 23129 95348 23214
rect 94924 23120 94964 23129
rect 94828 23080 94924 23120
rect 94636 22532 94676 22541
rect 94540 22492 94636 22532
rect 94636 22483 94676 22492
rect 94828 22364 94868 23080
rect 94924 23071 94964 23080
rect 95307 23120 95349 23129
rect 95307 23080 95308 23120
rect 95348 23080 95349 23120
rect 95307 23071 95349 23080
rect 95112 22700 95480 22709
rect 95152 22660 95194 22700
rect 95234 22660 95276 22700
rect 95316 22660 95358 22700
rect 95398 22660 95440 22700
rect 95112 22651 95480 22660
rect 95403 22532 95445 22541
rect 95403 22492 95404 22532
rect 95444 22492 95445 22532
rect 95403 22483 95445 22492
rect 95500 22532 95540 22541
rect 95596 22532 95636 25768
rect 95692 24725 95732 25852
rect 95905 25640 95945 26040
rect 95884 25600 95945 25640
rect 96015 25640 96055 26040
rect 96305 25640 96345 26040
rect 96015 25600 96116 25640
rect 95691 24716 95733 24725
rect 95691 24676 95692 24716
rect 95732 24676 95733 24716
rect 95691 24667 95733 24676
rect 95884 23960 95924 25600
rect 95884 23920 96020 23960
rect 95691 23120 95733 23129
rect 95691 23080 95692 23120
rect 95732 23080 95733 23120
rect 95691 23071 95733 23080
rect 95884 23120 95924 23129
rect 95692 22961 95732 23071
rect 95691 22952 95733 22961
rect 95691 22912 95692 22952
rect 95732 22912 95828 22952
rect 95691 22903 95733 22912
rect 95540 22492 95636 22532
rect 95500 22483 95540 22492
rect 95115 22448 95157 22457
rect 95115 22408 95116 22448
rect 95156 22408 95157 22448
rect 95115 22399 95157 22408
rect 95307 22448 95349 22457
rect 95307 22408 95308 22448
rect 95348 22408 95349 22448
rect 95307 22399 95349 22408
rect 94923 22364 94965 22373
rect 94828 22324 94924 22364
rect 94964 22324 94965 22364
rect 94923 22315 94965 22324
rect 94540 22280 94580 22289
rect 94156 22240 94540 22280
rect 93580 22196 93620 22205
rect 93964 22196 94004 22240
rect 94540 22231 94580 22240
rect 94924 22230 94964 22315
rect 95116 22314 95156 22399
rect 95308 22364 95348 22399
rect 95308 22313 95348 22324
rect 93620 22156 94004 22196
rect 93580 22147 93620 22156
rect 93483 22112 93525 22121
rect 93483 22072 93484 22112
rect 93524 22072 93525 22112
rect 93483 22063 93525 22072
rect 93332 21736 93428 21776
rect 92812 21727 92852 21736
rect 93292 21727 93332 21736
rect 91084 21608 91124 21617
rect 90892 21568 91084 21608
rect 89164 21559 89204 21568
rect 76588 21475 76628 21484
rect 77547 21524 77589 21533
rect 77547 21484 77548 21524
rect 77588 21484 77589 21524
rect 77547 21475 77589 21484
rect 77739 21524 77781 21533
rect 77739 21484 77740 21524
rect 77780 21484 77781 21524
rect 77739 21475 77781 21484
rect 78891 21524 78933 21533
rect 78891 21484 78892 21524
rect 78932 21484 78933 21524
rect 78891 21475 78933 21484
rect 79275 21524 79317 21533
rect 79275 21484 79276 21524
rect 79316 21484 79317 21524
rect 79275 21475 79317 21484
rect 80811 21524 80853 21533
rect 80811 21484 80812 21524
rect 80852 21484 80853 21524
rect 80811 21475 80853 21484
rect 82155 21524 82197 21533
rect 82155 21484 82156 21524
rect 82196 21484 82197 21524
rect 82155 21475 82197 21484
rect 82635 21524 82677 21533
rect 82635 21484 82636 21524
rect 82676 21484 82677 21524
rect 82635 21475 82677 21484
rect 83403 21524 83445 21533
rect 83403 21484 83404 21524
rect 83444 21484 83445 21524
rect 83403 21475 83445 21484
rect 83787 21524 83829 21533
rect 83787 21484 83788 21524
rect 83828 21484 83829 21524
rect 83787 21475 83829 21484
rect 84171 21524 84213 21533
rect 84171 21484 84172 21524
rect 84212 21484 84213 21524
rect 84171 21475 84213 21484
rect 89356 21524 89396 21568
rect 91084 21559 91124 21568
rect 92715 21608 92757 21617
rect 92715 21568 92716 21608
rect 92756 21568 92757 21608
rect 92715 21559 92757 21568
rect 93387 21608 93429 21617
rect 93484 21608 93524 22063
rect 95211 21776 95253 21785
rect 95211 21736 95212 21776
rect 95252 21736 95253 21776
rect 95211 21727 95253 21736
rect 95212 21642 95252 21727
rect 93387 21568 93388 21608
rect 93428 21568 93524 21608
rect 95308 21608 95348 21617
rect 95404 21608 95444 22483
rect 95788 22457 95828 22912
rect 95884 22709 95924 23080
rect 95883 22700 95925 22709
rect 95883 22660 95884 22700
rect 95924 22660 95925 22700
rect 95883 22651 95925 22660
rect 95884 22532 95924 22541
rect 95980 22532 96020 23920
rect 96076 23297 96116 25600
rect 96172 25600 96345 25640
rect 96415 25640 96455 26040
rect 96415 25600 96596 25640
rect 96075 23288 96117 23297
rect 96075 23248 96076 23288
rect 96116 23248 96117 23288
rect 96075 23239 96117 23248
rect 96076 23036 96116 23045
rect 96076 22541 96116 22996
rect 95924 22492 96020 22532
rect 96075 22532 96117 22541
rect 96075 22492 96076 22532
rect 96116 22492 96117 22532
rect 96172 22532 96212 25600
rect 96556 23960 96596 25600
rect 96705 25556 96745 26040
rect 96815 25640 96855 26040
rect 97105 25640 97145 26040
rect 97215 25640 97255 26040
rect 97505 25640 97545 26040
rect 97615 25640 97655 26040
rect 97905 25640 97945 26040
rect 96815 25600 96980 25640
rect 97105 25600 97172 25640
rect 97215 25600 97364 25640
rect 97505 25600 97556 25640
rect 97615 25600 97748 25640
rect 96705 25516 96884 25556
rect 96844 24884 96884 25516
rect 96940 24968 96980 25600
rect 96940 24928 97076 24968
rect 96844 24844 96980 24884
rect 96556 23920 96884 23960
rect 96352 23456 96720 23465
rect 96392 23416 96434 23456
rect 96474 23416 96516 23456
rect 96556 23416 96598 23456
rect 96638 23416 96680 23456
rect 96352 23407 96720 23416
rect 96459 23288 96501 23297
rect 96459 23248 96460 23288
rect 96500 23248 96501 23288
rect 96459 23239 96501 23248
rect 96748 23288 96788 23297
rect 96844 23288 96884 23920
rect 96788 23248 96884 23288
rect 96748 23239 96788 23248
rect 96460 23154 96500 23239
rect 96556 23120 96596 23129
rect 96556 22961 96596 23080
rect 96844 23120 96884 23129
rect 96844 22961 96884 23080
rect 96555 22952 96597 22961
rect 96555 22912 96556 22952
rect 96596 22912 96597 22952
rect 96555 22903 96597 22912
rect 96843 22952 96885 22961
rect 96843 22912 96844 22952
rect 96884 22912 96885 22952
rect 96843 22903 96885 22912
rect 96268 22868 96308 22877
rect 96308 22828 96404 22868
rect 96268 22819 96308 22828
rect 96364 22709 96404 22828
rect 96363 22700 96405 22709
rect 96363 22660 96364 22700
rect 96404 22660 96405 22700
rect 96363 22651 96405 22660
rect 96268 22532 96308 22541
rect 96172 22492 96268 22532
rect 95884 22483 95924 22492
rect 96075 22483 96117 22492
rect 96268 22483 96308 22492
rect 95787 22448 95829 22457
rect 95787 22408 95788 22448
rect 95828 22408 95829 22448
rect 95787 22399 95829 22408
rect 96364 22373 96404 22651
rect 95691 22364 95733 22373
rect 95691 22324 95692 22364
rect 95732 22324 95733 22364
rect 95691 22315 95733 22324
rect 96075 22364 96117 22373
rect 96075 22324 96076 22364
rect 96116 22324 96117 22364
rect 96075 22315 96117 22324
rect 96363 22364 96405 22373
rect 96363 22324 96364 22364
rect 96404 22324 96405 22364
rect 96363 22315 96405 22324
rect 96556 22364 96596 22903
rect 96748 22532 96788 22541
rect 96940 22532 96980 24844
rect 97036 23288 97076 24928
rect 97132 23960 97172 25600
rect 97132 23920 97268 23960
rect 97036 23239 97076 23248
rect 97132 23120 97172 23129
rect 97132 22961 97172 23080
rect 97131 22952 97173 22961
rect 97131 22912 97132 22952
rect 97172 22912 97173 22952
rect 97131 22903 97173 22912
rect 96788 22492 96980 22532
rect 97036 22532 97076 22541
rect 97228 22532 97268 23920
rect 97324 23288 97364 25600
rect 97324 23239 97364 23248
rect 97420 23120 97460 23129
rect 97420 22961 97460 23080
rect 97419 22952 97461 22961
rect 97419 22912 97420 22952
rect 97460 22912 97461 22952
rect 97419 22903 97461 22912
rect 97076 22492 97268 22532
rect 97516 22532 97556 25600
rect 97708 23288 97748 25600
rect 97708 23239 97748 23248
rect 97900 25600 97945 25640
rect 98015 25640 98055 26040
rect 98305 25640 98345 26040
rect 98415 25724 98455 26040
rect 98415 25684 98900 25724
rect 98015 25600 98132 25640
rect 98305 25600 98516 25640
rect 97804 23129 97844 23214
rect 97803 23120 97845 23129
rect 97803 23080 97804 23120
rect 97844 23080 97845 23120
rect 97803 23071 97845 23080
rect 97803 22952 97845 22961
rect 97803 22912 97804 22952
rect 97844 22912 97845 22952
rect 97803 22903 97845 22912
rect 97612 22532 97652 22541
rect 97516 22492 97612 22532
rect 96748 22483 96788 22492
rect 97036 22483 97076 22492
rect 97612 22483 97652 22492
rect 96556 22315 96596 22324
rect 97227 22364 97269 22373
rect 97227 22324 97228 22364
rect 97268 22324 97269 22364
rect 97227 22315 97269 22324
rect 97804 22364 97844 22903
rect 97900 22532 97940 25600
rect 98092 23288 98132 25600
rect 98092 23239 98132 23248
rect 98476 23288 98516 25600
rect 98476 23239 98516 23248
rect 98860 23288 98900 25684
rect 99148 25481 99188 34336
rect 99244 34208 99284 34217
rect 99244 31613 99284 34168
rect 99243 31604 99285 31613
rect 99243 31564 99244 31604
rect 99284 31564 99285 31604
rect 99243 31555 99285 31564
rect 99147 25472 99189 25481
rect 99147 25432 99148 25472
rect 99188 25432 99189 25472
rect 99147 25423 99189 25432
rect 99148 23960 99188 25423
rect 98860 23239 98900 23248
rect 99052 23920 99188 23960
rect 98187 23120 98229 23129
rect 98956 23120 98996 23129
rect 99052 23120 99092 23920
rect 98187 23080 98188 23120
rect 98228 23080 98229 23120
rect 98187 23071 98229 23080
rect 98668 23080 98956 23120
rect 98996 23080 99092 23120
rect 97996 22532 98036 22541
rect 97900 22492 97996 22532
rect 97996 22483 98036 22492
rect 98188 22373 98228 23071
rect 98668 23036 98708 23080
rect 98956 23071 98996 23080
rect 98668 22987 98708 22996
rect 99112 22700 99480 22709
rect 99152 22660 99194 22700
rect 99234 22660 99276 22700
rect 99316 22660 99358 22700
rect 99398 22660 99440 22700
rect 99112 22651 99480 22660
rect 97804 22315 97844 22324
rect 98187 22364 98229 22373
rect 98187 22324 98188 22364
rect 98228 22324 98229 22364
rect 98187 22315 98229 22324
rect 95692 22230 95732 22315
rect 96076 22230 96116 22315
rect 97228 22230 97268 22315
rect 98188 22230 98228 22315
rect 96352 21944 96720 21953
rect 96392 21904 96434 21944
rect 96474 21904 96516 21944
rect 96556 21904 96598 21944
rect 96638 21904 96680 21944
rect 96352 21895 96720 21904
rect 95348 21568 95444 21608
rect 93387 21559 93429 21568
rect 95308 21559 95348 21568
rect 89356 21475 89396 21484
rect 78892 21390 78932 21475
rect 79276 21390 79316 21475
rect 80812 21390 80852 21475
rect 82156 21390 82196 21475
rect 82636 21444 82676 21475
rect 83404 21390 83444 21475
rect 84172 21390 84212 21475
rect 92716 21474 92756 21559
rect 93388 21474 93428 21559
rect 11112 21188 11480 21197
rect 11152 21148 11194 21188
rect 11234 21148 11276 21188
rect 11316 21148 11358 21188
rect 11398 21148 11440 21188
rect 11112 21139 11480 21148
rect 15112 21188 15480 21197
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15112 21139 15480 21148
rect 19112 21188 19480 21197
rect 19152 21148 19194 21188
rect 19234 21148 19276 21188
rect 19316 21148 19358 21188
rect 19398 21148 19440 21188
rect 19112 21139 19480 21148
rect 23112 21188 23480 21197
rect 23152 21148 23194 21188
rect 23234 21148 23276 21188
rect 23316 21148 23358 21188
rect 23398 21148 23440 21188
rect 23112 21139 23480 21148
rect 27112 21188 27480 21197
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27112 21139 27480 21148
rect 31112 21188 31480 21197
rect 31152 21148 31194 21188
rect 31234 21148 31276 21188
rect 31316 21148 31358 21188
rect 31398 21148 31440 21188
rect 31112 21139 31480 21148
rect 35112 21188 35480 21197
rect 35152 21148 35194 21188
rect 35234 21148 35276 21188
rect 35316 21148 35358 21188
rect 35398 21148 35440 21188
rect 35112 21139 35480 21148
rect 39112 21188 39480 21197
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39112 21139 39480 21148
rect 43112 21188 43480 21197
rect 43152 21148 43194 21188
rect 43234 21148 43276 21188
rect 43316 21148 43358 21188
rect 43398 21148 43440 21188
rect 43112 21139 43480 21148
rect 47112 21188 47480 21197
rect 47152 21148 47194 21188
rect 47234 21148 47276 21188
rect 47316 21148 47358 21188
rect 47398 21148 47440 21188
rect 47112 21139 47480 21148
rect 51112 21188 51480 21197
rect 51152 21148 51194 21188
rect 51234 21148 51276 21188
rect 51316 21148 51358 21188
rect 51398 21148 51440 21188
rect 51112 21139 51480 21148
rect 55112 21188 55480 21197
rect 55152 21148 55194 21188
rect 55234 21148 55276 21188
rect 55316 21148 55358 21188
rect 55398 21148 55440 21188
rect 55112 21139 55480 21148
rect 59112 21188 59480 21197
rect 59152 21148 59194 21188
rect 59234 21148 59276 21188
rect 59316 21148 59358 21188
rect 59398 21148 59440 21188
rect 59112 21139 59480 21148
rect 63112 21188 63480 21197
rect 63152 21148 63194 21188
rect 63234 21148 63276 21188
rect 63316 21148 63358 21188
rect 63398 21148 63440 21188
rect 63112 21139 63480 21148
rect 67112 21188 67480 21197
rect 67152 21148 67194 21188
rect 67234 21148 67276 21188
rect 67316 21148 67358 21188
rect 67398 21148 67440 21188
rect 67112 21139 67480 21148
rect 71112 21188 71480 21197
rect 71152 21148 71194 21188
rect 71234 21148 71276 21188
rect 71316 21148 71358 21188
rect 71398 21148 71440 21188
rect 71112 21139 71480 21148
rect 75112 21188 75480 21197
rect 75152 21148 75194 21188
rect 75234 21148 75276 21188
rect 75316 21148 75358 21188
rect 75398 21148 75440 21188
rect 75112 21139 75480 21148
rect 79112 21188 79480 21197
rect 79152 21148 79194 21188
rect 79234 21148 79276 21188
rect 79316 21148 79358 21188
rect 79398 21148 79440 21188
rect 79112 21139 79480 21148
rect 83112 21188 83480 21197
rect 83152 21148 83194 21188
rect 83234 21148 83276 21188
rect 83316 21148 83358 21188
rect 83398 21148 83440 21188
rect 83112 21139 83480 21148
rect 87112 21188 87480 21197
rect 87152 21148 87194 21188
rect 87234 21148 87276 21188
rect 87316 21148 87358 21188
rect 87398 21148 87440 21188
rect 87112 21139 87480 21148
rect 91112 21188 91480 21197
rect 91152 21148 91194 21188
rect 91234 21148 91276 21188
rect 91316 21148 91358 21188
rect 91398 21148 91440 21188
rect 91112 21139 91480 21148
rect 95112 21188 95480 21197
rect 95152 21148 95194 21188
rect 95234 21148 95276 21188
rect 95316 21148 95358 21188
rect 95398 21148 95440 21188
rect 95112 21139 95480 21148
rect 99112 21188 99480 21197
rect 99152 21148 99194 21188
rect 99234 21148 99276 21188
rect 99316 21148 99358 21188
rect 99398 21148 99440 21188
rect 99112 21139 99480 21148
rect 12352 20432 12720 20441
rect 12392 20392 12434 20432
rect 12474 20392 12516 20432
rect 12556 20392 12598 20432
rect 12638 20392 12680 20432
rect 12352 20383 12720 20392
rect 16352 20432 16720 20441
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16352 20383 16720 20392
rect 20352 20432 20720 20441
rect 20392 20392 20434 20432
rect 20474 20392 20516 20432
rect 20556 20392 20598 20432
rect 20638 20392 20680 20432
rect 20352 20383 20720 20392
rect 24352 20432 24720 20441
rect 24392 20392 24434 20432
rect 24474 20392 24516 20432
rect 24556 20392 24598 20432
rect 24638 20392 24680 20432
rect 24352 20383 24720 20392
rect 28352 20432 28720 20441
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28352 20383 28720 20392
rect 32352 20432 32720 20441
rect 32392 20392 32434 20432
rect 32474 20392 32516 20432
rect 32556 20392 32598 20432
rect 32638 20392 32680 20432
rect 32352 20383 32720 20392
rect 36352 20432 36720 20441
rect 36392 20392 36434 20432
rect 36474 20392 36516 20432
rect 36556 20392 36598 20432
rect 36638 20392 36680 20432
rect 36352 20383 36720 20392
rect 40352 20432 40720 20441
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40352 20383 40720 20392
rect 44352 20432 44720 20441
rect 44392 20392 44434 20432
rect 44474 20392 44516 20432
rect 44556 20392 44598 20432
rect 44638 20392 44680 20432
rect 44352 20383 44720 20392
rect 48352 20432 48720 20441
rect 48392 20392 48434 20432
rect 48474 20392 48516 20432
rect 48556 20392 48598 20432
rect 48638 20392 48680 20432
rect 48352 20383 48720 20392
rect 52352 20432 52720 20441
rect 52392 20392 52434 20432
rect 52474 20392 52516 20432
rect 52556 20392 52598 20432
rect 52638 20392 52680 20432
rect 52352 20383 52720 20392
rect 56352 20432 56720 20441
rect 56392 20392 56434 20432
rect 56474 20392 56516 20432
rect 56556 20392 56598 20432
rect 56638 20392 56680 20432
rect 56352 20383 56720 20392
rect 60352 20432 60720 20441
rect 60392 20392 60434 20432
rect 60474 20392 60516 20432
rect 60556 20392 60598 20432
rect 60638 20392 60680 20432
rect 60352 20383 60720 20392
rect 64352 20432 64720 20441
rect 64392 20392 64434 20432
rect 64474 20392 64516 20432
rect 64556 20392 64598 20432
rect 64638 20392 64680 20432
rect 64352 20383 64720 20392
rect 68352 20432 68720 20441
rect 68392 20392 68434 20432
rect 68474 20392 68516 20432
rect 68556 20392 68598 20432
rect 68638 20392 68680 20432
rect 68352 20383 68720 20392
rect 72352 20432 72720 20441
rect 72392 20392 72434 20432
rect 72474 20392 72516 20432
rect 72556 20392 72598 20432
rect 72638 20392 72680 20432
rect 72352 20383 72720 20392
rect 76352 20432 76720 20441
rect 76392 20392 76434 20432
rect 76474 20392 76516 20432
rect 76556 20392 76598 20432
rect 76638 20392 76680 20432
rect 76352 20383 76720 20392
rect 80352 20432 80720 20441
rect 80392 20392 80434 20432
rect 80474 20392 80516 20432
rect 80556 20392 80598 20432
rect 80638 20392 80680 20432
rect 80352 20383 80720 20392
rect 84352 20432 84720 20441
rect 84392 20392 84434 20432
rect 84474 20392 84516 20432
rect 84556 20392 84598 20432
rect 84638 20392 84680 20432
rect 84352 20383 84720 20392
rect 88352 20432 88720 20441
rect 88392 20392 88434 20432
rect 88474 20392 88516 20432
rect 88556 20392 88598 20432
rect 88638 20392 88680 20432
rect 88352 20383 88720 20392
rect 92352 20432 92720 20441
rect 92392 20392 92434 20432
rect 92474 20392 92516 20432
rect 92556 20392 92598 20432
rect 92638 20392 92680 20432
rect 92352 20383 92720 20392
rect 96352 20432 96720 20441
rect 96392 20392 96434 20432
rect 96474 20392 96516 20432
rect 96556 20392 96598 20432
rect 96638 20392 96680 20432
rect 96352 20383 96720 20392
rect 75532 20012 75572 20021
rect 11112 19676 11480 19685
rect 11152 19636 11194 19676
rect 11234 19636 11276 19676
rect 11316 19636 11358 19676
rect 11398 19636 11440 19676
rect 11112 19627 11480 19636
rect 15112 19676 15480 19685
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15112 19627 15480 19636
rect 19112 19676 19480 19685
rect 19152 19636 19194 19676
rect 19234 19636 19276 19676
rect 19316 19636 19358 19676
rect 19398 19636 19440 19676
rect 19112 19627 19480 19636
rect 23112 19676 23480 19685
rect 23152 19636 23194 19676
rect 23234 19636 23276 19676
rect 23316 19636 23358 19676
rect 23398 19636 23440 19676
rect 23112 19627 23480 19636
rect 27112 19676 27480 19685
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27112 19627 27480 19636
rect 31112 19676 31480 19685
rect 31152 19636 31194 19676
rect 31234 19636 31276 19676
rect 31316 19636 31358 19676
rect 31398 19636 31440 19676
rect 31112 19627 31480 19636
rect 35112 19676 35480 19685
rect 35152 19636 35194 19676
rect 35234 19636 35276 19676
rect 35316 19636 35358 19676
rect 35398 19636 35440 19676
rect 35112 19627 35480 19636
rect 39112 19676 39480 19685
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39112 19627 39480 19636
rect 43112 19676 43480 19685
rect 43152 19636 43194 19676
rect 43234 19636 43276 19676
rect 43316 19636 43358 19676
rect 43398 19636 43440 19676
rect 43112 19627 43480 19636
rect 47112 19676 47480 19685
rect 47152 19636 47194 19676
rect 47234 19636 47276 19676
rect 47316 19636 47358 19676
rect 47398 19636 47440 19676
rect 47112 19627 47480 19636
rect 51112 19676 51480 19685
rect 51152 19636 51194 19676
rect 51234 19636 51276 19676
rect 51316 19636 51358 19676
rect 51398 19636 51440 19676
rect 51112 19627 51480 19636
rect 55112 19676 55480 19685
rect 55152 19636 55194 19676
rect 55234 19636 55276 19676
rect 55316 19636 55358 19676
rect 55398 19636 55440 19676
rect 55112 19627 55480 19636
rect 59112 19676 59480 19685
rect 59152 19636 59194 19676
rect 59234 19636 59276 19676
rect 59316 19636 59358 19676
rect 59398 19636 59440 19676
rect 59112 19627 59480 19636
rect 63112 19676 63480 19685
rect 63152 19636 63194 19676
rect 63234 19636 63276 19676
rect 63316 19636 63358 19676
rect 63398 19636 63440 19676
rect 63112 19627 63480 19636
rect 67112 19676 67480 19685
rect 67152 19636 67194 19676
rect 67234 19636 67276 19676
rect 67316 19636 67358 19676
rect 67398 19636 67440 19676
rect 67112 19627 67480 19636
rect 71112 19676 71480 19685
rect 71152 19636 71194 19676
rect 71234 19636 71276 19676
rect 71316 19636 71358 19676
rect 71398 19636 71440 19676
rect 71112 19627 71480 19636
rect 75112 19676 75480 19685
rect 75152 19636 75194 19676
rect 75234 19636 75276 19676
rect 75316 19636 75358 19676
rect 75398 19636 75440 19676
rect 75112 19627 75480 19636
rect 74764 19340 74804 19349
rect 71787 19256 71829 19265
rect 71787 19216 71788 19256
rect 71828 19216 71829 19256
rect 74764 19256 74804 19300
rect 75244 19256 75284 19265
rect 74764 19216 75244 19256
rect 71787 19207 71829 19216
rect 12352 18920 12720 18929
rect 12392 18880 12434 18920
rect 12474 18880 12516 18920
rect 12556 18880 12598 18920
rect 12638 18880 12680 18920
rect 12352 18871 12720 18880
rect 16352 18920 16720 18929
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16352 18871 16720 18880
rect 20352 18920 20720 18929
rect 20392 18880 20434 18920
rect 20474 18880 20516 18920
rect 20556 18880 20598 18920
rect 20638 18880 20680 18920
rect 20352 18871 20720 18880
rect 24352 18920 24720 18929
rect 24392 18880 24434 18920
rect 24474 18880 24516 18920
rect 24556 18880 24598 18920
rect 24638 18880 24680 18920
rect 24352 18871 24720 18880
rect 28352 18920 28720 18929
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28352 18871 28720 18880
rect 32352 18920 32720 18929
rect 32392 18880 32434 18920
rect 32474 18880 32516 18920
rect 32556 18880 32598 18920
rect 32638 18880 32680 18920
rect 32352 18871 32720 18880
rect 36352 18920 36720 18929
rect 36392 18880 36434 18920
rect 36474 18880 36516 18920
rect 36556 18880 36598 18920
rect 36638 18880 36680 18920
rect 36352 18871 36720 18880
rect 40352 18920 40720 18929
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40352 18871 40720 18880
rect 44352 18920 44720 18929
rect 44392 18880 44434 18920
rect 44474 18880 44516 18920
rect 44556 18880 44598 18920
rect 44638 18880 44680 18920
rect 44352 18871 44720 18880
rect 48352 18920 48720 18929
rect 48392 18880 48434 18920
rect 48474 18880 48516 18920
rect 48556 18880 48598 18920
rect 48638 18880 48680 18920
rect 48352 18871 48720 18880
rect 52352 18920 52720 18929
rect 52392 18880 52434 18920
rect 52474 18880 52516 18920
rect 52556 18880 52598 18920
rect 52638 18880 52680 18920
rect 52352 18871 52720 18880
rect 56352 18920 56720 18929
rect 56392 18880 56434 18920
rect 56474 18880 56516 18920
rect 56556 18880 56598 18920
rect 56638 18880 56680 18920
rect 56352 18871 56720 18880
rect 60352 18920 60720 18929
rect 60392 18880 60434 18920
rect 60474 18880 60516 18920
rect 60556 18880 60598 18920
rect 60638 18880 60680 18920
rect 60352 18871 60720 18880
rect 64352 18920 64720 18929
rect 64392 18880 64434 18920
rect 64474 18880 64516 18920
rect 64556 18880 64598 18920
rect 64638 18880 64680 18920
rect 64352 18871 64720 18880
rect 68352 18920 68720 18929
rect 68392 18880 68434 18920
rect 68474 18880 68516 18920
rect 68556 18880 68598 18920
rect 68638 18880 68680 18920
rect 68352 18871 68720 18880
rect 68235 18584 68277 18593
rect 68235 18544 68236 18584
rect 68276 18544 68277 18584
rect 68235 18535 68277 18544
rect 11112 18164 11480 18173
rect 11152 18124 11194 18164
rect 11234 18124 11276 18164
rect 11316 18124 11358 18164
rect 11398 18124 11440 18164
rect 11112 18115 11480 18124
rect 15112 18164 15480 18173
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15112 18115 15480 18124
rect 19112 18164 19480 18173
rect 19152 18124 19194 18164
rect 19234 18124 19276 18164
rect 19316 18124 19358 18164
rect 19398 18124 19440 18164
rect 19112 18115 19480 18124
rect 23112 18164 23480 18173
rect 23152 18124 23194 18164
rect 23234 18124 23276 18164
rect 23316 18124 23358 18164
rect 23398 18124 23440 18164
rect 23112 18115 23480 18124
rect 27112 18164 27480 18173
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27112 18115 27480 18124
rect 31112 18164 31480 18173
rect 31152 18124 31194 18164
rect 31234 18124 31276 18164
rect 31316 18124 31358 18164
rect 31398 18124 31440 18164
rect 31112 18115 31480 18124
rect 35112 18164 35480 18173
rect 35152 18124 35194 18164
rect 35234 18124 35276 18164
rect 35316 18124 35358 18164
rect 35398 18124 35440 18164
rect 35112 18115 35480 18124
rect 39112 18164 39480 18173
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39112 18115 39480 18124
rect 43112 18164 43480 18173
rect 43152 18124 43194 18164
rect 43234 18124 43276 18164
rect 43316 18124 43358 18164
rect 43398 18124 43440 18164
rect 43112 18115 43480 18124
rect 47112 18164 47480 18173
rect 47152 18124 47194 18164
rect 47234 18124 47276 18164
rect 47316 18124 47358 18164
rect 47398 18124 47440 18164
rect 47112 18115 47480 18124
rect 51112 18164 51480 18173
rect 51152 18124 51194 18164
rect 51234 18124 51276 18164
rect 51316 18124 51358 18164
rect 51398 18124 51440 18164
rect 51112 18115 51480 18124
rect 55112 18164 55480 18173
rect 55152 18124 55194 18164
rect 55234 18124 55276 18164
rect 55316 18124 55358 18164
rect 55398 18124 55440 18164
rect 55112 18115 55480 18124
rect 59112 18164 59480 18173
rect 59152 18124 59194 18164
rect 59234 18124 59276 18164
rect 59316 18124 59358 18164
rect 59398 18124 59440 18164
rect 59112 18115 59480 18124
rect 63112 18164 63480 18173
rect 63152 18124 63194 18164
rect 63234 18124 63276 18164
rect 63316 18124 63358 18164
rect 63398 18124 63440 18164
rect 63112 18115 63480 18124
rect 67112 18164 67480 18173
rect 67152 18124 67194 18164
rect 67234 18124 67276 18164
rect 67316 18124 67358 18164
rect 67398 18124 67440 18164
rect 67112 18115 67480 18124
rect 12352 17408 12720 17417
rect 12392 17368 12434 17408
rect 12474 17368 12516 17408
rect 12556 17368 12598 17408
rect 12638 17368 12680 17408
rect 12352 17359 12720 17368
rect 16352 17408 16720 17417
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16352 17359 16720 17368
rect 20352 17408 20720 17417
rect 20392 17368 20434 17408
rect 20474 17368 20516 17408
rect 20556 17368 20598 17408
rect 20638 17368 20680 17408
rect 20352 17359 20720 17368
rect 24352 17408 24720 17417
rect 24392 17368 24434 17408
rect 24474 17368 24516 17408
rect 24556 17368 24598 17408
rect 24638 17368 24680 17408
rect 24352 17359 24720 17368
rect 28352 17408 28720 17417
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28352 17359 28720 17368
rect 32352 17408 32720 17417
rect 32392 17368 32434 17408
rect 32474 17368 32516 17408
rect 32556 17368 32598 17408
rect 32638 17368 32680 17408
rect 32352 17359 32720 17368
rect 36352 17408 36720 17417
rect 36392 17368 36434 17408
rect 36474 17368 36516 17408
rect 36556 17368 36598 17408
rect 36638 17368 36680 17408
rect 36352 17359 36720 17368
rect 40352 17408 40720 17417
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40352 17359 40720 17368
rect 44352 17408 44720 17417
rect 44392 17368 44434 17408
rect 44474 17368 44516 17408
rect 44556 17368 44598 17408
rect 44638 17368 44680 17408
rect 44352 17359 44720 17368
rect 48352 17408 48720 17417
rect 48392 17368 48434 17408
rect 48474 17368 48516 17408
rect 48556 17368 48598 17408
rect 48638 17368 48680 17408
rect 48352 17359 48720 17368
rect 52352 17408 52720 17417
rect 52392 17368 52434 17408
rect 52474 17368 52516 17408
rect 52556 17368 52598 17408
rect 52638 17368 52680 17408
rect 52352 17359 52720 17368
rect 56352 17408 56720 17417
rect 56392 17368 56434 17408
rect 56474 17368 56516 17408
rect 56556 17368 56598 17408
rect 56638 17368 56680 17408
rect 56352 17359 56720 17368
rect 60352 17408 60720 17417
rect 60392 17368 60434 17408
rect 60474 17368 60516 17408
rect 60556 17368 60598 17408
rect 60638 17368 60680 17408
rect 60352 17359 60720 17368
rect 64352 17408 64720 17417
rect 64392 17368 64434 17408
rect 64474 17368 64516 17408
rect 64556 17368 64598 17408
rect 64638 17368 64680 17408
rect 64352 17359 64720 17368
rect 11112 16652 11480 16661
rect 11152 16612 11194 16652
rect 11234 16612 11276 16652
rect 11316 16612 11358 16652
rect 11398 16612 11440 16652
rect 11112 16603 11480 16612
rect 15112 16652 15480 16661
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15112 16603 15480 16612
rect 19112 16652 19480 16661
rect 19152 16612 19194 16652
rect 19234 16612 19276 16652
rect 19316 16612 19358 16652
rect 19398 16612 19440 16652
rect 19112 16603 19480 16612
rect 23112 16652 23480 16661
rect 23152 16612 23194 16652
rect 23234 16612 23276 16652
rect 23316 16612 23358 16652
rect 23398 16612 23440 16652
rect 23112 16603 23480 16612
rect 27112 16652 27480 16661
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27112 16603 27480 16612
rect 31112 16652 31480 16661
rect 31152 16612 31194 16652
rect 31234 16612 31276 16652
rect 31316 16612 31358 16652
rect 31398 16612 31440 16652
rect 31112 16603 31480 16612
rect 35112 16652 35480 16661
rect 35152 16612 35194 16652
rect 35234 16612 35276 16652
rect 35316 16612 35358 16652
rect 35398 16612 35440 16652
rect 35112 16603 35480 16612
rect 39112 16652 39480 16661
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39112 16603 39480 16612
rect 43112 16652 43480 16661
rect 43152 16612 43194 16652
rect 43234 16612 43276 16652
rect 43316 16612 43358 16652
rect 43398 16612 43440 16652
rect 43112 16603 43480 16612
rect 47112 16652 47480 16661
rect 47152 16612 47194 16652
rect 47234 16612 47276 16652
rect 47316 16612 47358 16652
rect 47398 16612 47440 16652
rect 47112 16603 47480 16612
rect 51112 16652 51480 16661
rect 51152 16612 51194 16652
rect 51234 16612 51276 16652
rect 51316 16612 51358 16652
rect 51398 16612 51440 16652
rect 51112 16603 51480 16612
rect 55112 16652 55480 16661
rect 55152 16612 55194 16652
rect 55234 16612 55276 16652
rect 55316 16612 55358 16652
rect 55398 16612 55440 16652
rect 55112 16603 55480 16612
rect 59112 16652 59480 16661
rect 59152 16612 59194 16652
rect 59234 16612 59276 16652
rect 59316 16612 59358 16652
rect 59398 16612 59440 16652
rect 59112 16603 59480 16612
rect 63112 16652 63480 16661
rect 63152 16612 63194 16652
rect 63234 16612 63276 16652
rect 63316 16612 63358 16652
rect 63398 16612 63440 16652
rect 63112 16603 63480 16612
rect 67112 16652 67480 16661
rect 67152 16612 67194 16652
rect 67234 16612 67276 16652
rect 67316 16612 67358 16652
rect 67398 16612 67440 16652
rect 67112 16603 67480 16612
rect 67371 15980 67413 15989
rect 67371 15940 67372 15980
rect 67412 15940 67413 15980
rect 67371 15931 67413 15940
rect 12352 15896 12720 15905
rect 12392 15856 12434 15896
rect 12474 15856 12516 15896
rect 12556 15856 12598 15896
rect 12638 15856 12680 15896
rect 12352 15847 12720 15856
rect 16352 15896 16720 15905
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16352 15847 16720 15856
rect 20352 15896 20720 15905
rect 20392 15856 20434 15896
rect 20474 15856 20516 15896
rect 20556 15856 20598 15896
rect 20638 15856 20680 15896
rect 20352 15847 20720 15856
rect 24352 15896 24720 15905
rect 24392 15856 24434 15896
rect 24474 15856 24516 15896
rect 24556 15856 24598 15896
rect 24638 15856 24680 15896
rect 24352 15847 24720 15856
rect 28352 15896 28720 15905
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28352 15847 28720 15856
rect 32352 15896 32720 15905
rect 32392 15856 32434 15896
rect 32474 15856 32516 15896
rect 32556 15856 32598 15896
rect 32638 15856 32680 15896
rect 32352 15847 32720 15856
rect 36352 15896 36720 15905
rect 36392 15856 36434 15896
rect 36474 15856 36516 15896
rect 36556 15856 36598 15896
rect 36638 15856 36680 15896
rect 36352 15847 36720 15856
rect 40352 15896 40720 15905
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40352 15847 40720 15856
rect 44352 15896 44720 15905
rect 44392 15856 44434 15896
rect 44474 15856 44516 15896
rect 44556 15856 44598 15896
rect 44638 15856 44680 15896
rect 44352 15847 44720 15856
rect 48352 15896 48720 15905
rect 48392 15856 48434 15896
rect 48474 15856 48516 15896
rect 48556 15856 48598 15896
rect 48638 15856 48680 15896
rect 48352 15847 48720 15856
rect 52352 15896 52720 15905
rect 52392 15856 52434 15896
rect 52474 15856 52516 15896
rect 52556 15856 52598 15896
rect 52638 15856 52680 15896
rect 52352 15847 52720 15856
rect 56352 15896 56720 15905
rect 56392 15856 56434 15896
rect 56474 15856 56516 15896
rect 56556 15856 56598 15896
rect 56638 15856 56680 15896
rect 56352 15847 56720 15856
rect 60352 15896 60720 15905
rect 60392 15856 60434 15896
rect 60474 15856 60516 15896
rect 60556 15856 60598 15896
rect 60638 15856 60680 15896
rect 60352 15847 60720 15856
rect 64352 15896 64720 15905
rect 64392 15856 64434 15896
rect 64474 15856 64516 15896
rect 64556 15856 64598 15896
rect 64638 15856 64680 15896
rect 64352 15847 64720 15856
rect 67372 15728 67412 15931
rect 67372 15679 67412 15688
rect 67179 15560 67221 15569
rect 67179 15520 67180 15560
rect 67220 15520 67221 15560
rect 67179 15511 67221 15520
rect 67563 15560 67605 15569
rect 67563 15520 67564 15560
rect 67604 15520 67605 15560
rect 67563 15511 67605 15520
rect 68236 15560 68276 18535
rect 71112 18164 71480 18173
rect 71152 18124 71194 18164
rect 71234 18124 71276 18164
rect 71316 18124 71358 18164
rect 71398 18124 71440 18164
rect 71112 18115 71480 18124
rect 68352 17408 68720 17417
rect 68392 17368 68434 17408
rect 68474 17368 68516 17408
rect 68556 17368 68598 17408
rect 68638 17368 68680 17408
rect 68352 17359 68720 17368
rect 69100 16316 69140 16325
rect 68352 15896 68720 15905
rect 68392 15856 68434 15896
rect 68474 15856 68516 15896
rect 68556 15856 68598 15896
rect 68638 15856 68680 15896
rect 68352 15847 68720 15856
rect 68811 15896 68853 15905
rect 68811 15856 68812 15896
rect 68852 15856 68853 15896
rect 68811 15847 68853 15856
rect 67180 15476 67220 15511
rect 67180 15425 67220 15436
rect 67564 15392 67604 15511
rect 67755 15476 67797 15485
rect 67755 15436 67756 15476
rect 67796 15436 67797 15476
rect 67755 15427 67797 15436
rect 11112 15140 11480 15149
rect 11152 15100 11194 15140
rect 11234 15100 11276 15140
rect 11316 15100 11358 15140
rect 11398 15100 11440 15140
rect 11112 15091 11480 15100
rect 15112 15140 15480 15149
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15112 15091 15480 15100
rect 19112 15140 19480 15149
rect 19152 15100 19194 15140
rect 19234 15100 19276 15140
rect 19316 15100 19358 15140
rect 19398 15100 19440 15140
rect 19112 15091 19480 15100
rect 23112 15140 23480 15149
rect 23152 15100 23194 15140
rect 23234 15100 23276 15140
rect 23316 15100 23358 15140
rect 23398 15100 23440 15140
rect 23112 15091 23480 15100
rect 27112 15140 27480 15149
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27112 15091 27480 15100
rect 31112 15140 31480 15149
rect 31152 15100 31194 15140
rect 31234 15100 31276 15140
rect 31316 15100 31358 15140
rect 31398 15100 31440 15140
rect 31112 15091 31480 15100
rect 35112 15140 35480 15149
rect 35152 15100 35194 15140
rect 35234 15100 35276 15140
rect 35316 15100 35358 15140
rect 35398 15100 35440 15140
rect 35112 15091 35480 15100
rect 39112 15140 39480 15149
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39112 15091 39480 15100
rect 43112 15140 43480 15149
rect 43152 15100 43194 15140
rect 43234 15100 43276 15140
rect 43316 15100 43358 15140
rect 43398 15100 43440 15140
rect 43112 15091 43480 15100
rect 47112 15140 47480 15149
rect 47152 15100 47194 15140
rect 47234 15100 47276 15140
rect 47316 15100 47358 15140
rect 47398 15100 47440 15140
rect 47112 15091 47480 15100
rect 51112 15140 51480 15149
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51112 15091 51480 15100
rect 55112 15140 55480 15149
rect 55152 15100 55194 15140
rect 55234 15100 55276 15140
rect 55316 15100 55358 15140
rect 55398 15100 55440 15140
rect 55112 15091 55480 15100
rect 59112 15140 59480 15149
rect 59152 15100 59194 15140
rect 59234 15100 59276 15140
rect 59316 15100 59358 15140
rect 59398 15100 59440 15140
rect 59112 15091 59480 15100
rect 63112 15140 63480 15149
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63112 15091 63480 15100
rect 67112 15140 67480 15149
rect 67152 15100 67194 15140
rect 67234 15100 67276 15140
rect 67316 15100 67358 15140
rect 67398 15100 67440 15140
rect 67112 15091 67480 15100
rect 12352 14384 12720 14393
rect 12392 14344 12434 14384
rect 12474 14344 12516 14384
rect 12556 14344 12598 14384
rect 12638 14344 12680 14384
rect 12352 14335 12720 14344
rect 16352 14384 16720 14393
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16352 14335 16720 14344
rect 20352 14384 20720 14393
rect 20392 14344 20434 14384
rect 20474 14344 20516 14384
rect 20556 14344 20598 14384
rect 20638 14344 20680 14384
rect 20352 14335 20720 14344
rect 24352 14384 24720 14393
rect 24392 14344 24434 14384
rect 24474 14344 24516 14384
rect 24556 14344 24598 14384
rect 24638 14344 24680 14384
rect 24352 14335 24720 14344
rect 28352 14384 28720 14393
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28352 14335 28720 14344
rect 32352 14384 32720 14393
rect 32392 14344 32434 14384
rect 32474 14344 32516 14384
rect 32556 14344 32598 14384
rect 32638 14344 32680 14384
rect 32352 14335 32720 14344
rect 36352 14384 36720 14393
rect 36392 14344 36434 14384
rect 36474 14344 36516 14384
rect 36556 14344 36598 14384
rect 36638 14344 36680 14384
rect 36352 14335 36720 14344
rect 40352 14384 40720 14393
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40352 14335 40720 14344
rect 44352 14384 44720 14393
rect 44392 14344 44434 14384
rect 44474 14344 44516 14384
rect 44556 14344 44598 14384
rect 44638 14344 44680 14384
rect 44352 14335 44720 14344
rect 48352 14384 48720 14393
rect 48392 14344 48434 14384
rect 48474 14344 48516 14384
rect 48556 14344 48598 14384
rect 48638 14344 48680 14384
rect 48352 14335 48720 14344
rect 52352 14384 52720 14393
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52352 14335 52720 14344
rect 56352 14384 56720 14393
rect 56392 14344 56434 14384
rect 56474 14344 56516 14384
rect 56556 14344 56598 14384
rect 56638 14344 56680 14384
rect 56352 14335 56720 14344
rect 60352 14384 60720 14393
rect 60392 14344 60434 14384
rect 60474 14344 60516 14384
rect 60556 14344 60598 14384
rect 60638 14344 60680 14384
rect 60352 14335 60720 14344
rect 64352 14384 64720 14393
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64352 14335 64720 14344
rect 9387 13964 9429 13973
rect 9387 13924 9388 13964
rect 9428 13924 9429 13964
rect 9387 13915 9429 13924
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 7112 13628 7480 13637
rect 7152 13588 7194 13628
rect 7234 13588 7276 13628
rect 7316 13588 7358 13628
rect 7398 13588 7440 13628
rect 7112 13579 7480 13588
rect 11112 13628 11480 13637
rect 11152 13588 11194 13628
rect 11234 13588 11276 13628
rect 11316 13588 11358 13628
rect 11398 13588 11440 13628
rect 11112 13579 11480 13588
rect 15112 13628 15480 13637
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15112 13579 15480 13588
rect 19112 13628 19480 13637
rect 19152 13588 19194 13628
rect 19234 13588 19276 13628
rect 19316 13588 19358 13628
rect 19398 13588 19440 13628
rect 19112 13579 19480 13588
rect 23112 13628 23480 13637
rect 23152 13588 23194 13628
rect 23234 13588 23276 13628
rect 23316 13588 23358 13628
rect 23398 13588 23440 13628
rect 23112 13579 23480 13588
rect 27112 13628 27480 13637
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27112 13579 27480 13588
rect 31112 13628 31480 13637
rect 31152 13588 31194 13628
rect 31234 13588 31276 13628
rect 31316 13588 31358 13628
rect 31398 13588 31440 13628
rect 31112 13579 31480 13588
rect 35112 13628 35480 13637
rect 35152 13588 35194 13628
rect 35234 13588 35276 13628
rect 35316 13588 35358 13628
rect 35398 13588 35440 13628
rect 35112 13579 35480 13588
rect 39112 13628 39480 13637
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39112 13579 39480 13588
rect 43112 13628 43480 13637
rect 43152 13588 43194 13628
rect 43234 13588 43276 13628
rect 43316 13588 43358 13628
rect 43398 13588 43440 13628
rect 43112 13579 43480 13588
rect 47112 13628 47480 13637
rect 47152 13588 47194 13628
rect 47234 13588 47276 13628
rect 47316 13588 47358 13628
rect 47398 13588 47440 13628
rect 47112 13579 47480 13588
rect 51112 13628 51480 13637
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51112 13579 51480 13588
rect 55112 13628 55480 13637
rect 55152 13588 55194 13628
rect 55234 13588 55276 13628
rect 55316 13588 55358 13628
rect 55398 13588 55440 13628
rect 55112 13579 55480 13588
rect 59112 13628 59480 13637
rect 59152 13588 59194 13628
rect 59234 13588 59276 13628
rect 59316 13588 59358 13628
rect 59398 13588 59440 13628
rect 59112 13579 59480 13588
rect 63112 13628 63480 13637
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63112 13579 63480 13588
rect 67112 13628 67480 13637
rect 67152 13588 67194 13628
rect 67234 13588 67276 13628
rect 67316 13588 67358 13628
rect 67398 13588 67440 13628
rect 67112 13579 67480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 8352 12872 8720 12881
rect 8392 12832 8434 12872
rect 8474 12832 8516 12872
rect 8556 12832 8598 12872
rect 8638 12832 8680 12872
rect 8352 12823 8720 12832
rect 12352 12872 12720 12881
rect 12392 12832 12434 12872
rect 12474 12832 12516 12872
rect 12556 12832 12598 12872
rect 12638 12832 12680 12872
rect 12352 12823 12720 12832
rect 16352 12872 16720 12881
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16352 12823 16720 12832
rect 20352 12872 20720 12881
rect 20392 12832 20434 12872
rect 20474 12832 20516 12872
rect 20556 12832 20598 12872
rect 20638 12832 20680 12872
rect 20352 12823 20720 12832
rect 24352 12872 24720 12881
rect 24392 12832 24434 12872
rect 24474 12832 24516 12872
rect 24556 12832 24598 12872
rect 24638 12832 24680 12872
rect 24352 12823 24720 12832
rect 28352 12872 28720 12881
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28352 12823 28720 12832
rect 32352 12872 32720 12881
rect 32392 12832 32434 12872
rect 32474 12832 32516 12872
rect 32556 12832 32598 12872
rect 32638 12832 32680 12872
rect 32352 12823 32720 12832
rect 36352 12872 36720 12881
rect 36392 12832 36434 12872
rect 36474 12832 36516 12872
rect 36556 12832 36598 12872
rect 36638 12832 36680 12872
rect 36352 12823 36720 12832
rect 40352 12872 40720 12881
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40352 12823 40720 12832
rect 44352 12872 44720 12881
rect 44392 12832 44434 12872
rect 44474 12832 44516 12872
rect 44556 12832 44598 12872
rect 44638 12832 44680 12872
rect 44352 12823 44720 12832
rect 48352 12872 48720 12881
rect 48392 12832 48434 12872
rect 48474 12832 48516 12872
rect 48556 12832 48598 12872
rect 48638 12832 48680 12872
rect 48352 12823 48720 12832
rect 52352 12872 52720 12881
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52352 12823 52720 12832
rect 56352 12872 56720 12881
rect 56392 12832 56434 12872
rect 56474 12832 56516 12872
rect 56556 12832 56598 12872
rect 56638 12832 56680 12872
rect 56352 12823 56720 12832
rect 60352 12872 60720 12881
rect 60392 12832 60434 12872
rect 60474 12832 60516 12872
rect 60556 12832 60598 12872
rect 60638 12832 60680 12872
rect 60352 12823 60720 12832
rect 64352 12872 64720 12881
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64352 12823 64720 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 7112 12116 7480 12125
rect 7152 12076 7194 12116
rect 7234 12076 7276 12116
rect 7316 12076 7358 12116
rect 7398 12076 7440 12116
rect 7112 12067 7480 12076
rect 11112 12116 11480 12125
rect 11152 12076 11194 12116
rect 11234 12076 11276 12116
rect 11316 12076 11358 12116
rect 11398 12076 11440 12116
rect 11112 12067 11480 12076
rect 15112 12116 15480 12125
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15112 12067 15480 12076
rect 19112 12116 19480 12125
rect 19152 12076 19194 12116
rect 19234 12076 19276 12116
rect 19316 12076 19358 12116
rect 19398 12076 19440 12116
rect 19112 12067 19480 12076
rect 23112 12116 23480 12125
rect 23152 12076 23194 12116
rect 23234 12076 23276 12116
rect 23316 12076 23358 12116
rect 23398 12076 23440 12116
rect 23112 12067 23480 12076
rect 27112 12116 27480 12125
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27112 12067 27480 12076
rect 31112 12116 31480 12125
rect 31152 12076 31194 12116
rect 31234 12076 31276 12116
rect 31316 12076 31358 12116
rect 31398 12076 31440 12116
rect 31112 12067 31480 12076
rect 35112 12116 35480 12125
rect 35152 12076 35194 12116
rect 35234 12076 35276 12116
rect 35316 12076 35358 12116
rect 35398 12076 35440 12116
rect 35112 12067 35480 12076
rect 39112 12116 39480 12125
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39112 12067 39480 12076
rect 43112 12116 43480 12125
rect 43152 12076 43194 12116
rect 43234 12076 43276 12116
rect 43316 12076 43358 12116
rect 43398 12076 43440 12116
rect 43112 12067 43480 12076
rect 47112 12116 47480 12125
rect 47152 12076 47194 12116
rect 47234 12076 47276 12116
rect 47316 12076 47358 12116
rect 47398 12076 47440 12116
rect 47112 12067 47480 12076
rect 51112 12116 51480 12125
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51112 12067 51480 12076
rect 55112 12116 55480 12125
rect 55152 12076 55194 12116
rect 55234 12076 55276 12116
rect 55316 12076 55358 12116
rect 55398 12076 55440 12116
rect 55112 12067 55480 12076
rect 59112 12116 59480 12125
rect 59152 12076 59194 12116
rect 59234 12076 59276 12116
rect 59316 12076 59358 12116
rect 59398 12076 59440 12116
rect 59112 12067 59480 12076
rect 63112 12116 63480 12125
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63112 12067 63480 12076
rect 67112 12116 67480 12125
rect 67152 12076 67194 12116
rect 67234 12076 67276 12116
rect 67316 12076 67358 12116
rect 67398 12076 67440 12116
rect 67112 12067 67480 12076
rect 2188 11780 2228 11789
rect 2188 10949 2228 11740
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 8352 11360 8720 11369
rect 8392 11320 8434 11360
rect 8474 11320 8516 11360
rect 8556 11320 8598 11360
rect 8638 11320 8680 11360
rect 8352 11311 8720 11320
rect 12352 11360 12720 11369
rect 12392 11320 12434 11360
rect 12474 11320 12516 11360
rect 12556 11320 12598 11360
rect 12638 11320 12680 11360
rect 12352 11311 12720 11320
rect 16352 11360 16720 11369
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16352 11311 16720 11320
rect 20352 11360 20720 11369
rect 20392 11320 20434 11360
rect 20474 11320 20516 11360
rect 20556 11320 20598 11360
rect 20638 11320 20680 11360
rect 20352 11311 20720 11320
rect 24352 11360 24720 11369
rect 24392 11320 24434 11360
rect 24474 11320 24516 11360
rect 24556 11320 24598 11360
rect 24638 11320 24680 11360
rect 24352 11311 24720 11320
rect 28352 11360 28720 11369
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28352 11311 28720 11320
rect 32352 11360 32720 11369
rect 32392 11320 32434 11360
rect 32474 11320 32516 11360
rect 32556 11320 32598 11360
rect 32638 11320 32680 11360
rect 32352 11311 32720 11320
rect 36352 11360 36720 11369
rect 36392 11320 36434 11360
rect 36474 11320 36516 11360
rect 36556 11320 36598 11360
rect 36638 11320 36680 11360
rect 36352 11311 36720 11320
rect 40352 11360 40720 11369
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40352 11311 40720 11320
rect 44352 11360 44720 11369
rect 44392 11320 44434 11360
rect 44474 11320 44516 11360
rect 44556 11320 44598 11360
rect 44638 11320 44680 11360
rect 44352 11311 44720 11320
rect 48352 11360 48720 11369
rect 48392 11320 48434 11360
rect 48474 11320 48516 11360
rect 48556 11320 48598 11360
rect 48638 11320 48680 11360
rect 48352 11311 48720 11320
rect 52352 11360 52720 11369
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52352 11311 52720 11320
rect 56352 11360 56720 11369
rect 56392 11320 56434 11360
rect 56474 11320 56516 11360
rect 56556 11320 56598 11360
rect 56638 11320 56680 11360
rect 56352 11311 56720 11320
rect 60352 11360 60720 11369
rect 60392 11320 60434 11360
rect 60474 11320 60516 11360
rect 60556 11320 60598 11360
rect 60638 11320 60680 11360
rect 60352 11311 60720 11320
rect 64352 11360 64720 11369
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64352 11311 64720 11320
rect 2187 10940 2229 10949
rect 2187 10900 2188 10940
rect 2228 10900 2229 10940
rect 2187 10891 2229 10900
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 7112 10604 7480 10613
rect 7152 10564 7194 10604
rect 7234 10564 7276 10604
rect 7316 10564 7358 10604
rect 7398 10564 7440 10604
rect 7112 10555 7480 10564
rect 11112 10604 11480 10613
rect 11152 10564 11194 10604
rect 11234 10564 11276 10604
rect 11316 10564 11358 10604
rect 11398 10564 11440 10604
rect 11112 10555 11480 10564
rect 15112 10604 15480 10613
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15112 10555 15480 10564
rect 19112 10604 19480 10613
rect 19152 10564 19194 10604
rect 19234 10564 19276 10604
rect 19316 10564 19358 10604
rect 19398 10564 19440 10604
rect 19112 10555 19480 10564
rect 23112 10604 23480 10613
rect 23152 10564 23194 10604
rect 23234 10564 23276 10604
rect 23316 10564 23358 10604
rect 23398 10564 23440 10604
rect 23112 10555 23480 10564
rect 27112 10604 27480 10613
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27112 10555 27480 10564
rect 31112 10604 31480 10613
rect 31152 10564 31194 10604
rect 31234 10564 31276 10604
rect 31316 10564 31358 10604
rect 31398 10564 31440 10604
rect 31112 10555 31480 10564
rect 35112 10604 35480 10613
rect 35152 10564 35194 10604
rect 35234 10564 35276 10604
rect 35316 10564 35358 10604
rect 35398 10564 35440 10604
rect 35112 10555 35480 10564
rect 39112 10604 39480 10613
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39112 10555 39480 10564
rect 43112 10604 43480 10613
rect 43152 10564 43194 10604
rect 43234 10564 43276 10604
rect 43316 10564 43358 10604
rect 43398 10564 43440 10604
rect 43112 10555 43480 10564
rect 47112 10604 47480 10613
rect 47152 10564 47194 10604
rect 47234 10564 47276 10604
rect 47316 10564 47358 10604
rect 47398 10564 47440 10604
rect 47112 10555 47480 10564
rect 51112 10604 51480 10613
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51112 10555 51480 10564
rect 55112 10604 55480 10613
rect 55152 10564 55194 10604
rect 55234 10564 55276 10604
rect 55316 10564 55358 10604
rect 55398 10564 55440 10604
rect 55112 10555 55480 10564
rect 59112 10604 59480 10613
rect 59152 10564 59194 10604
rect 59234 10564 59276 10604
rect 59316 10564 59358 10604
rect 59398 10564 59440 10604
rect 59112 10555 59480 10564
rect 63112 10604 63480 10613
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63112 10555 63480 10564
rect 67112 10604 67480 10613
rect 67152 10564 67194 10604
rect 67234 10564 67276 10604
rect 67316 10564 67358 10604
rect 67398 10564 67440 10604
rect 67112 10555 67480 10564
rect 67564 10436 67604 15352
rect 67756 15342 67796 15427
rect 68236 15140 68276 15520
rect 68427 15560 68469 15569
rect 68427 15520 68428 15560
rect 68468 15520 68469 15560
rect 68427 15511 68469 15520
rect 68428 15426 68468 15511
rect 68140 15100 68276 15140
rect 68043 14804 68085 14813
rect 68043 14764 68044 14804
rect 68084 14764 68085 14804
rect 68043 14755 68085 14764
rect 68044 14670 68084 14755
rect 68140 14729 68180 15100
rect 68716 14972 68756 14981
rect 68812 14972 68852 15847
rect 69100 15569 69140 16276
rect 69292 16064 69332 16073
rect 69099 15560 69141 15569
rect 69099 15520 69100 15560
rect 69140 15520 69141 15560
rect 69099 15511 69141 15520
rect 69292 15065 69332 16024
rect 71691 16064 71733 16073
rect 71691 16024 71692 16064
rect 71732 16024 71733 16064
rect 71691 16015 71733 16024
rect 69963 15812 70005 15821
rect 69963 15772 69964 15812
rect 70004 15772 70005 15812
rect 69963 15763 70005 15772
rect 69867 15728 69909 15737
rect 69867 15688 69868 15728
rect 69908 15688 69909 15728
rect 69867 15679 69909 15688
rect 69483 15644 69525 15653
rect 69483 15604 69484 15644
rect 69524 15604 69525 15644
rect 69483 15595 69525 15604
rect 69291 15056 69333 15065
rect 69291 15016 69292 15056
rect 69332 15016 69333 15056
rect 69291 15007 69333 15016
rect 68756 14932 68852 14972
rect 69099 14972 69141 14981
rect 69099 14932 69100 14972
rect 69140 14932 69141 14972
rect 68716 14923 68756 14932
rect 69099 14923 69141 14932
rect 69484 14972 69524 15595
rect 69484 14923 69524 14932
rect 69868 14972 69908 15679
rect 69868 14923 69908 14932
rect 69100 14838 69140 14923
rect 69291 14888 69333 14897
rect 69291 14848 69292 14888
rect 69332 14848 69333 14888
rect 69291 14839 69333 14848
rect 68139 14720 68181 14729
rect 68139 14680 68140 14720
rect 68180 14680 68181 14720
rect 68139 14671 68181 14680
rect 68619 14720 68661 14729
rect 68619 14680 68620 14720
rect 68660 14680 68661 14720
rect 68619 14671 68661 14680
rect 69004 14720 69044 14729
rect 68140 14586 68180 14671
rect 68620 14586 68660 14671
rect 68352 14384 68720 14393
rect 68392 14344 68434 14384
rect 68474 14344 68516 14384
rect 68556 14344 68598 14384
rect 68638 14344 68680 14384
rect 68352 14335 68720 14344
rect 69004 13973 69044 14680
rect 69292 14216 69332 14839
rect 69676 14804 69716 14813
rect 69484 14764 69676 14804
rect 69716 14764 69812 14804
rect 69387 14720 69429 14729
rect 69484 14720 69524 14764
rect 69676 14755 69716 14764
rect 69387 14680 69388 14720
rect 69428 14680 69524 14720
rect 69387 14671 69429 14680
rect 69388 14586 69428 14671
rect 69388 14216 69428 14225
rect 69292 14176 69388 14216
rect 69388 14167 69428 14176
rect 69772 14048 69812 14764
rect 69868 14216 69908 14225
rect 69964 14216 70004 15763
rect 71692 15485 71732 16015
rect 71691 15476 71733 15485
rect 71691 15436 71692 15476
rect 71732 15436 71733 15476
rect 71691 15427 71733 15436
rect 71691 15140 71733 15149
rect 71691 15100 71692 15140
rect 71732 15100 71733 15140
rect 71691 15091 71733 15100
rect 71692 14813 71732 15091
rect 71691 14804 71733 14813
rect 71691 14764 71692 14804
rect 71732 14764 71733 14804
rect 71691 14755 71733 14764
rect 69908 14176 70004 14216
rect 69868 14167 69908 14176
rect 69772 13999 69812 14008
rect 69003 13964 69045 13973
rect 69003 13924 69004 13964
rect 69044 13924 69045 13964
rect 69003 13915 69045 13924
rect 69195 13964 69237 13973
rect 69195 13924 69196 13964
rect 69236 13924 69237 13964
rect 69195 13915 69237 13924
rect 70059 13964 70101 13973
rect 70059 13924 70060 13964
rect 70100 13924 70101 13964
rect 70059 13915 70101 13924
rect 69196 13830 69236 13915
rect 68352 12872 68720 12881
rect 68392 12832 68434 12872
rect 68474 12832 68516 12872
rect 68556 12832 68598 12872
rect 68638 12832 68680 12872
rect 68352 12823 68720 12832
rect 68352 11360 68720 11369
rect 68392 11320 68434 11360
rect 68474 11320 68516 11360
rect 68556 11320 68598 11360
rect 68638 11320 68680 11360
rect 68352 11311 68720 11320
rect 68523 11024 68565 11033
rect 68523 10984 68524 11024
rect 68564 10984 68565 11024
rect 68523 10975 68565 10984
rect 69771 11024 69813 11033
rect 69771 10984 69772 11024
rect 69812 10984 69813 11024
rect 69771 10975 69813 10984
rect 67468 10396 67604 10436
rect 67468 10268 67508 10396
rect 67468 10193 67508 10228
rect 67660 10352 67700 10361
rect 67467 10184 67509 10193
rect 67467 10144 67468 10184
rect 67508 10144 67509 10184
rect 67467 10135 67509 10144
rect 67468 10104 67508 10135
rect 67660 10109 67700 10312
rect 68524 10193 68564 10975
rect 69292 10940 69332 10949
rect 69196 10352 69236 10361
rect 69004 10268 69044 10277
rect 68332 10184 68372 10193
rect 67659 10100 67701 10109
rect 67659 10060 67660 10100
rect 67700 10060 67701 10100
rect 67659 10051 67701 10060
rect 68236 10100 68276 10109
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 8352 9848 8720 9857
rect 8392 9808 8434 9848
rect 8474 9808 8516 9848
rect 8556 9808 8598 9848
rect 8638 9808 8680 9848
rect 8352 9799 8720 9808
rect 12352 9848 12720 9857
rect 12392 9808 12434 9848
rect 12474 9808 12516 9848
rect 12556 9808 12598 9848
rect 12638 9808 12680 9848
rect 12352 9799 12720 9808
rect 16352 9848 16720 9857
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16352 9799 16720 9808
rect 20352 9848 20720 9857
rect 20392 9808 20434 9848
rect 20474 9808 20516 9848
rect 20556 9808 20598 9848
rect 20638 9808 20680 9848
rect 20352 9799 20720 9808
rect 24352 9848 24720 9857
rect 24392 9808 24434 9848
rect 24474 9808 24516 9848
rect 24556 9808 24598 9848
rect 24638 9808 24680 9848
rect 24352 9799 24720 9808
rect 28352 9848 28720 9857
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28352 9799 28720 9808
rect 32352 9848 32720 9857
rect 32392 9808 32434 9848
rect 32474 9808 32516 9848
rect 32556 9808 32598 9848
rect 32638 9808 32680 9848
rect 32352 9799 32720 9808
rect 36352 9848 36720 9857
rect 36392 9808 36434 9848
rect 36474 9808 36516 9848
rect 36556 9808 36598 9848
rect 36638 9808 36680 9848
rect 36352 9799 36720 9808
rect 40352 9848 40720 9857
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40352 9799 40720 9808
rect 44352 9848 44720 9857
rect 44392 9808 44434 9848
rect 44474 9808 44516 9848
rect 44556 9808 44598 9848
rect 44638 9808 44680 9848
rect 44352 9799 44720 9808
rect 48352 9848 48720 9857
rect 48392 9808 48434 9848
rect 48474 9808 48516 9848
rect 48556 9808 48598 9848
rect 48638 9808 48680 9848
rect 48352 9799 48720 9808
rect 52352 9848 52720 9857
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52352 9799 52720 9808
rect 56352 9848 56720 9857
rect 56392 9808 56434 9848
rect 56474 9808 56516 9848
rect 56556 9808 56598 9848
rect 56638 9808 56680 9848
rect 56352 9799 56720 9808
rect 60352 9848 60720 9857
rect 60392 9808 60434 9848
rect 60474 9808 60516 9848
rect 60556 9808 60598 9848
rect 60638 9808 60680 9848
rect 60352 9799 60720 9808
rect 64352 9848 64720 9857
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64352 9799 64720 9808
rect 68236 9605 68276 10060
rect 68332 10025 68372 10144
rect 68523 10184 68565 10193
rect 68523 10144 68524 10184
rect 68564 10144 68565 10184
rect 68523 10135 68565 10144
rect 68716 10184 68756 10193
rect 68524 10050 68564 10135
rect 68716 10025 68756 10144
rect 69004 10025 69044 10228
rect 68331 10016 68373 10025
rect 68331 9976 68332 10016
rect 68372 9976 68373 10016
rect 68331 9967 68373 9976
rect 68715 10016 68757 10025
rect 68715 9976 68716 10016
rect 68756 9976 68757 10016
rect 68715 9967 68757 9976
rect 69003 10016 69045 10025
rect 69003 9976 69004 10016
rect 69044 9976 69045 10016
rect 69003 9967 69045 9976
rect 68352 9848 68720 9857
rect 68392 9808 68434 9848
rect 68474 9808 68516 9848
rect 68556 9808 68598 9848
rect 68638 9808 68680 9848
rect 68352 9799 68720 9808
rect 68235 9596 68277 9605
rect 68235 9556 68236 9596
rect 68276 9556 68277 9596
rect 68235 9547 68277 9556
rect 69004 9428 69044 9967
rect 69196 9521 69236 10312
rect 69292 10184 69332 10900
rect 69772 10890 69812 10975
rect 69484 10772 69524 10781
rect 69484 10268 69524 10732
rect 69868 10772 69908 10781
rect 69908 10732 70004 10772
rect 69868 10723 69908 10732
rect 69484 10228 69620 10268
rect 69387 10184 69429 10193
rect 69292 10144 69388 10184
rect 69428 10144 69429 10184
rect 69387 10135 69429 10144
rect 69388 10025 69428 10135
rect 69484 10100 69524 10109
rect 69387 10016 69429 10025
rect 69387 9976 69388 10016
rect 69428 9976 69429 10016
rect 69387 9967 69429 9976
rect 69195 9512 69237 9521
rect 69195 9472 69196 9512
rect 69236 9472 69237 9512
rect 69195 9463 69237 9472
rect 69484 9437 69524 10060
rect 69580 10016 69620 10228
rect 69676 10193 69716 10278
rect 69675 10184 69717 10193
rect 69675 10144 69676 10184
rect 69716 10144 69717 10184
rect 69675 10135 69717 10144
rect 69772 10100 69812 10109
rect 69580 9976 69716 10016
rect 69579 9848 69621 9857
rect 69579 9808 69580 9848
rect 69620 9808 69621 9848
rect 69579 9799 69621 9808
rect 69580 9680 69620 9799
rect 69580 9631 69620 9640
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 7112 9092 7480 9101
rect 7152 9052 7194 9092
rect 7234 9052 7276 9092
rect 7316 9052 7358 9092
rect 7398 9052 7440 9092
rect 7112 9043 7480 9052
rect 11112 9092 11480 9101
rect 11152 9052 11194 9092
rect 11234 9052 11276 9092
rect 11316 9052 11358 9092
rect 11398 9052 11440 9092
rect 11112 9043 11480 9052
rect 15112 9092 15480 9101
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15112 9043 15480 9052
rect 19112 9092 19480 9101
rect 19152 9052 19194 9092
rect 19234 9052 19276 9092
rect 19316 9052 19358 9092
rect 19398 9052 19440 9092
rect 19112 9043 19480 9052
rect 23112 9092 23480 9101
rect 23152 9052 23194 9092
rect 23234 9052 23276 9092
rect 23316 9052 23358 9092
rect 23398 9052 23440 9092
rect 23112 9043 23480 9052
rect 27112 9092 27480 9101
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27112 9043 27480 9052
rect 31112 9092 31480 9101
rect 31152 9052 31194 9092
rect 31234 9052 31276 9092
rect 31316 9052 31358 9092
rect 31398 9052 31440 9092
rect 31112 9043 31480 9052
rect 35112 9092 35480 9101
rect 35152 9052 35194 9092
rect 35234 9052 35276 9092
rect 35316 9052 35358 9092
rect 35398 9052 35440 9092
rect 35112 9043 35480 9052
rect 39112 9092 39480 9101
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39112 9043 39480 9052
rect 43112 9092 43480 9101
rect 43152 9052 43194 9092
rect 43234 9052 43276 9092
rect 43316 9052 43358 9092
rect 43398 9052 43440 9092
rect 43112 9043 43480 9052
rect 47112 9092 47480 9101
rect 47152 9052 47194 9092
rect 47234 9052 47276 9092
rect 47316 9052 47358 9092
rect 47398 9052 47440 9092
rect 47112 9043 47480 9052
rect 51112 9092 51480 9101
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51112 9043 51480 9052
rect 55112 9092 55480 9101
rect 55152 9052 55194 9092
rect 55234 9052 55276 9092
rect 55316 9052 55358 9092
rect 55398 9052 55440 9092
rect 55112 9043 55480 9052
rect 59112 9092 59480 9101
rect 59152 9052 59194 9092
rect 59234 9052 59276 9092
rect 59316 9052 59358 9092
rect 59398 9052 59440 9092
rect 59112 9043 59480 9052
rect 63112 9092 63480 9101
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63112 9043 63480 9052
rect 67112 9092 67480 9101
rect 67152 9052 67194 9092
rect 67234 9052 67276 9092
rect 67316 9052 67358 9092
rect 67398 9052 67440 9092
rect 67112 9043 67480 9052
rect 69004 8849 69044 9388
rect 69388 9428 69428 9437
rect 69195 9344 69237 9353
rect 69195 9304 69196 9344
rect 69236 9304 69237 9344
rect 69195 9295 69237 9304
rect 69196 9210 69236 9295
rect 69388 9092 69428 9388
rect 69483 9428 69525 9437
rect 69483 9388 69484 9428
rect 69524 9388 69525 9428
rect 69483 9379 69525 9388
rect 69676 9269 69716 9976
rect 69772 9941 69812 10060
rect 69771 9932 69813 9941
rect 69771 9892 69772 9932
rect 69812 9892 69813 9932
rect 69771 9883 69813 9892
rect 69867 9764 69909 9773
rect 69867 9724 69868 9764
rect 69908 9724 69909 9764
rect 69867 9715 69909 9724
rect 69868 9680 69908 9715
rect 69868 9629 69908 9640
rect 69772 9512 69812 9521
rect 69675 9260 69717 9269
rect 69675 9220 69676 9260
rect 69716 9220 69717 9260
rect 69675 9211 69717 9220
rect 69772 9092 69812 9472
rect 69964 9185 70004 10732
rect 69963 9176 70005 9185
rect 69963 9136 69964 9176
rect 70004 9136 70005 9176
rect 69963 9127 70005 9136
rect 69388 9052 69812 9092
rect 69772 9008 69812 9052
rect 70060 9008 70100 13915
rect 70731 10100 70773 10109
rect 70731 10060 70732 10100
rect 70772 10060 70773 10100
rect 70731 10051 70773 10060
rect 70732 9689 70772 10051
rect 70731 9680 70773 9689
rect 70731 9640 70732 9680
rect 70772 9640 70773 9680
rect 70731 9631 70773 9640
rect 69772 8968 70100 9008
rect 69003 8840 69045 8849
rect 69003 8800 69004 8840
rect 69044 8800 69045 8840
rect 69003 8791 69045 8800
rect 1652 8716 1748 8756
rect 1612 8707 1652 8716
rect 652 8504 692 8513
rect 652 8177 692 8464
rect 1708 8504 1748 8716
rect 2036 8716 2132 8756
rect 1996 8707 2036 8716
rect 1804 8504 1844 8513
rect 1708 8464 1804 8504
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 844 7916 884 7927
rect 844 7841 884 7876
rect 1708 7916 1748 8464
rect 1804 8455 1844 8464
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 8352 8336 8720 8345
rect 8392 8296 8434 8336
rect 8474 8296 8516 8336
rect 8556 8296 8598 8336
rect 8638 8296 8680 8336
rect 8352 8287 8720 8296
rect 12352 8336 12720 8345
rect 12392 8296 12434 8336
rect 12474 8296 12516 8336
rect 12556 8296 12598 8336
rect 12638 8296 12680 8336
rect 12352 8287 12720 8296
rect 16352 8336 16720 8345
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16352 8287 16720 8296
rect 20352 8336 20720 8345
rect 20392 8296 20434 8336
rect 20474 8296 20516 8336
rect 20556 8296 20598 8336
rect 20638 8296 20680 8336
rect 20352 8287 20720 8296
rect 24352 8336 24720 8345
rect 24392 8296 24434 8336
rect 24474 8296 24516 8336
rect 24556 8296 24598 8336
rect 24638 8296 24680 8336
rect 24352 8287 24720 8296
rect 28352 8336 28720 8345
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28352 8287 28720 8296
rect 32352 8336 32720 8345
rect 32392 8296 32434 8336
rect 32474 8296 32516 8336
rect 32556 8296 32598 8336
rect 32638 8296 32680 8336
rect 32352 8287 32720 8296
rect 36352 8336 36720 8345
rect 36392 8296 36434 8336
rect 36474 8296 36516 8336
rect 36556 8296 36598 8336
rect 36638 8296 36680 8336
rect 36352 8287 36720 8296
rect 40352 8336 40720 8345
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40352 8287 40720 8296
rect 44352 8336 44720 8345
rect 44392 8296 44434 8336
rect 44474 8296 44516 8336
rect 44556 8296 44598 8336
rect 44638 8296 44680 8336
rect 44352 8287 44720 8296
rect 48352 8336 48720 8345
rect 48392 8296 48434 8336
rect 48474 8296 48516 8336
rect 48556 8296 48598 8336
rect 48638 8296 48680 8336
rect 48352 8287 48720 8296
rect 52352 8336 52720 8345
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52352 8287 52720 8296
rect 56352 8336 56720 8345
rect 56392 8296 56434 8336
rect 56474 8296 56516 8336
rect 56556 8296 56598 8336
rect 56638 8296 56680 8336
rect 56352 8287 56720 8296
rect 60352 8336 60720 8345
rect 60392 8296 60434 8336
rect 60474 8296 60516 8336
rect 60556 8296 60598 8336
rect 60638 8296 60680 8336
rect 60352 8287 60720 8296
rect 64352 8336 64720 8345
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64352 8287 64720 8296
rect 68352 8336 68720 8345
rect 68392 8296 68434 8336
rect 68474 8296 68516 8336
rect 68556 8296 68598 8336
rect 68638 8296 68680 8336
rect 68352 8287 68720 8296
rect 69772 8177 69812 8968
rect 69771 8168 69813 8177
rect 69771 8128 69772 8168
rect 69812 8128 69813 8168
rect 69771 8119 69813 8128
rect 843 7832 885 7841
rect 843 7792 844 7832
rect 884 7792 885 7832
rect 843 7783 885 7792
rect 1515 7832 1557 7841
rect 1515 7792 1516 7832
rect 1556 7792 1557 7832
rect 1515 7783 1557 7792
rect 652 7748 692 7757
rect 652 7337 692 7708
rect 1516 7698 1556 7783
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 844 7244 884 7253
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 844 6665 884 7204
rect 843 6656 885 6665
rect 843 6616 844 6656
rect 884 6616 885 6656
rect 843 6607 885 6616
rect 1323 6656 1365 6665
rect 1323 6616 1324 6656
rect 1364 6616 1365 6656
rect 1323 6607 1365 6616
rect 1324 6522 1364 6607
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 1516 6404 1556 6413
rect 1708 6404 1748 7876
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 7112 7580 7480 7589
rect 7152 7540 7194 7580
rect 7234 7540 7276 7580
rect 7316 7540 7358 7580
rect 7398 7540 7440 7580
rect 7112 7531 7480 7540
rect 11112 7580 11480 7589
rect 11152 7540 11194 7580
rect 11234 7540 11276 7580
rect 11316 7540 11358 7580
rect 11398 7540 11440 7580
rect 11112 7531 11480 7540
rect 15112 7580 15480 7589
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15112 7531 15480 7540
rect 19112 7580 19480 7589
rect 19152 7540 19194 7580
rect 19234 7540 19276 7580
rect 19316 7540 19358 7580
rect 19398 7540 19440 7580
rect 19112 7531 19480 7540
rect 23112 7580 23480 7589
rect 23152 7540 23194 7580
rect 23234 7540 23276 7580
rect 23316 7540 23358 7580
rect 23398 7540 23440 7580
rect 23112 7531 23480 7540
rect 27112 7580 27480 7589
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27112 7531 27480 7540
rect 31112 7580 31480 7589
rect 31152 7540 31194 7580
rect 31234 7540 31276 7580
rect 31316 7540 31358 7580
rect 31398 7540 31440 7580
rect 31112 7531 31480 7540
rect 35112 7580 35480 7589
rect 35152 7540 35194 7580
rect 35234 7540 35276 7580
rect 35316 7540 35358 7580
rect 35398 7540 35440 7580
rect 35112 7531 35480 7540
rect 39112 7580 39480 7589
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39112 7531 39480 7540
rect 43112 7580 43480 7589
rect 43152 7540 43194 7580
rect 43234 7540 43276 7580
rect 43316 7540 43358 7580
rect 43398 7540 43440 7580
rect 43112 7531 43480 7540
rect 47112 7580 47480 7589
rect 47152 7540 47194 7580
rect 47234 7540 47276 7580
rect 47316 7540 47358 7580
rect 47398 7540 47440 7580
rect 47112 7531 47480 7540
rect 51112 7580 51480 7589
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51112 7531 51480 7540
rect 55112 7580 55480 7589
rect 55152 7540 55194 7580
rect 55234 7540 55276 7580
rect 55316 7540 55358 7580
rect 55398 7540 55440 7580
rect 55112 7531 55480 7540
rect 59112 7580 59480 7589
rect 59152 7540 59194 7580
rect 59234 7540 59276 7580
rect 59316 7540 59358 7580
rect 59398 7540 59440 7580
rect 59112 7531 59480 7540
rect 63112 7580 63480 7589
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63112 7531 63480 7540
rect 67112 7580 67480 7589
rect 67152 7540 67194 7580
rect 67234 7540 67276 7580
rect 67316 7540 67358 7580
rect 67398 7540 67440 7580
rect 67112 7531 67480 7540
rect 71112 7580 71480 7589
rect 71152 7540 71194 7580
rect 71234 7540 71276 7580
rect 71316 7540 71358 7580
rect 71398 7540 71440 7580
rect 71112 7531 71480 7540
rect 71788 7253 71828 19207
rect 74956 19088 74996 19097
rect 74996 19048 75188 19088
rect 74956 19039 74996 19048
rect 75148 18929 75188 19048
rect 72352 18920 72720 18929
rect 72392 18880 72434 18920
rect 72474 18880 72516 18920
rect 72556 18880 72598 18920
rect 72638 18880 72680 18920
rect 72352 18871 72720 18880
rect 75147 18920 75189 18929
rect 75147 18880 75148 18920
rect 75188 18880 75189 18920
rect 75147 18871 75189 18880
rect 74571 18836 74613 18845
rect 74571 18796 74572 18836
rect 74612 18796 74613 18836
rect 74571 18787 74613 18796
rect 74955 18836 74997 18845
rect 74955 18796 74956 18836
rect 74996 18796 74997 18836
rect 74955 18787 74997 18796
rect 72939 18584 72981 18593
rect 72939 18544 72940 18584
rect 72980 18544 72981 18584
rect 72939 18535 72981 18544
rect 73707 18584 73749 18593
rect 73707 18544 73708 18584
rect 73748 18544 73749 18584
rect 73707 18535 73749 18544
rect 74283 18584 74325 18593
rect 74283 18544 74284 18584
rect 74324 18544 74325 18584
rect 74283 18535 74325 18544
rect 72940 18450 72980 18535
rect 73036 18332 73076 18341
rect 72352 17408 72720 17417
rect 72392 17368 72434 17408
rect 72474 17368 72516 17408
rect 72556 17368 72598 17408
rect 72638 17368 72680 17408
rect 72352 17359 72720 17368
rect 73036 15569 73076 18292
rect 73708 17837 73748 18535
rect 74284 18450 74324 18535
rect 74572 18500 74612 18787
rect 74956 18752 74996 18787
rect 74956 18701 74996 18712
rect 74476 18460 74572 18500
rect 74188 18332 74228 18341
rect 73707 17828 73749 17837
rect 73707 17788 73708 17828
rect 73748 17788 73749 17828
rect 73707 17779 73749 17788
rect 74091 17828 74133 17837
rect 74091 17788 74092 17828
rect 74132 17788 74133 17828
rect 74091 17779 74133 17788
rect 73708 17694 73748 17779
rect 74092 17694 74132 17779
rect 73900 17576 73940 17585
rect 73940 17536 74036 17576
rect 73900 17527 73940 17536
rect 73227 15980 73269 15989
rect 73227 15940 73228 15980
rect 73268 15940 73269 15980
rect 73227 15931 73269 15940
rect 73131 15644 73173 15653
rect 73228 15644 73268 15931
rect 73899 15896 73941 15905
rect 73899 15856 73900 15896
rect 73940 15856 73941 15896
rect 73899 15847 73941 15856
rect 73131 15604 73132 15644
rect 73172 15604 73173 15644
rect 73131 15595 73173 15604
rect 73215 15604 73268 15644
rect 73611 15644 73653 15653
rect 73900 15644 73940 15847
rect 73996 15644 74036 17536
rect 74188 16577 74228 18292
rect 74476 17828 74516 18460
rect 74572 18451 74612 18460
rect 75148 18500 75188 18871
rect 75244 18593 75284 19216
rect 75435 19256 75477 19265
rect 75435 19216 75436 19256
rect 75476 19216 75477 19256
rect 75435 19207 75477 19216
rect 75436 19122 75476 19207
rect 75243 18584 75285 18593
rect 75243 18544 75244 18584
rect 75284 18544 75285 18584
rect 75243 18535 75285 18544
rect 75148 18451 75188 18460
rect 74764 18332 74804 18341
rect 74956 18332 74996 18341
rect 74804 18292 74900 18332
rect 74764 18283 74804 18292
rect 74476 17779 74516 17788
rect 74860 17660 74900 18292
rect 74956 17744 74996 18292
rect 75112 18164 75480 18173
rect 75152 18124 75194 18164
rect 75234 18124 75276 18164
rect 75316 18124 75358 18164
rect 75398 18124 75440 18164
rect 75112 18115 75480 18124
rect 75340 17828 75380 17837
rect 75052 17744 75092 17753
rect 75340 17744 75380 17788
rect 75532 17744 75572 19972
rect 80619 20012 80661 20021
rect 80619 19972 80620 20012
rect 80660 19972 80661 20012
rect 80619 19963 80661 19972
rect 86859 20012 86901 20021
rect 86859 19972 86860 20012
rect 86900 19972 86901 20012
rect 86859 19963 86901 19972
rect 93196 20012 93236 20021
rect 75723 19928 75765 19937
rect 75723 19888 75724 19928
rect 75764 19888 75765 19928
rect 75723 19879 75765 19888
rect 75724 19265 75764 19879
rect 80620 19878 80660 19963
rect 86860 19878 86900 19963
rect 80428 19844 80468 19853
rect 87052 19844 87092 19853
rect 80468 19804 80564 19844
rect 80428 19795 80468 19804
rect 79112 19676 79480 19685
rect 79152 19636 79194 19676
rect 79234 19636 79276 19676
rect 79316 19636 79358 19676
rect 79398 19636 79440 19676
rect 79112 19627 79480 19636
rect 76588 19265 76628 19350
rect 80524 19349 80564 19804
rect 86956 19804 87052 19844
rect 83112 19676 83480 19685
rect 83152 19636 83194 19676
rect 83234 19636 83276 19676
rect 83316 19636 83358 19676
rect 83398 19636 83440 19676
rect 83112 19627 83480 19636
rect 77644 19340 77684 19349
rect 75628 19256 75668 19265
rect 75628 18845 75668 19216
rect 75723 19256 75765 19265
rect 75723 19216 75724 19256
rect 75764 19216 75765 19256
rect 75723 19207 75765 19216
rect 76587 19256 76629 19265
rect 76587 19216 76588 19256
rect 76628 19216 76629 19256
rect 76587 19207 76629 19216
rect 77068 19256 77108 19265
rect 77644 19256 77684 19300
rect 78220 19340 78260 19349
rect 77644 19216 78068 19256
rect 77068 19172 77108 19216
rect 76972 19132 77108 19172
rect 75724 19088 75764 19097
rect 76684 19088 76724 19097
rect 75764 19048 75956 19088
rect 75724 19039 75764 19048
rect 75819 18920 75861 18929
rect 75819 18880 75820 18920
rect 75860 18880 75861 18920
rect 75819 18871 75861 18880
rect 75627 18836 75669 18845
rect 75627 18796 75628 18836
rect 75668 18796 75669 18836
rect 75627 18787 75669 18796
rect 75820 18500 75860 18871
rect 75820 18451 75860 18460
rect 74956 17704 75052 17744
rect 75092 17704 75380 17744
rect 75436 17704 75572 17744
rect 75819 17744 75861 17753
rect 75819 17704 75820 17744
rect 75860 17704 75861 17744
rect 75052 17695 75092 17704
rect 75436 17660 75476 17704
rect 75819 17695 75861 17704
rect 74860 17620 74996 17660
rect 74284 17576 74324 17585
rect 74668 17576 74708 17585
rect 74324 17536 74420 17576
rect 74284 17527 74324 17536
rect 74187 16568 74229 16577
rect 74187 16528 74188 16568
rect 74228 16528 74229 16568
rect 74187 16519 74229 16528
rect 74283 15812 74325 15821
rect 74283 15772 74284 15812
rect 74324 15772 74325 15812
rect 74283 15763 74325 15772
rect 73611 15604 73612 15644
rect 73652 15604 73655 15644
rect 73900 15604 73945 15644
rect 73996 15604 74055 15644
rect 72814 15560 72856 15569
rect 72814 15520 72815 15560
rect 72855 15520 72856 15560
rect 72814 15511 72856 15520
rect 73035 15560 73077 15569
rect 73035 15520 73036 15560
rect 73076 15520 73077 15560
rect 73035 15511 73077 15520
rect 72704 15476 72746 15485
rect 72704 15436 72705 15476
rect 72745 15436 72746 15476
rect 72704 15427 72746 15436
rect 72414 15392 72456 15401
rect 71884 15352 72345 15392
rect 71884 14981 71924 15352
rect 72305 15204 72345 15352
rect 72414 15352 72415 15392
rect 72455 15352 72456 15392
rect 72414 15343 72456 15352
rect 72415 15204 72455 15343
rect 72705 15204 72745 15427
rect 72815 15204 72855 15511
rect 73132 15476 73172 15595
rect 73105 15436 73172 15476
rect 73105 15204 73145 15436
rect 73215 15204 73255 15604
rect 73611 15595 73655 15604
rect 73504 15560 73546 15569
rect 73504 15520 73505 15560
rect 73545 15520 73546 15560
rect 73504 15511 73546 15520
rect 73505 15204 73545 15511
rect 73615 15204 73655 15595
rect 73905 15204 73945 15604
rect 74015 15204 74055 15604
rect 74284 15560 74324 15763
rect 74380 15644 74420 17536
rect 74708 17536 74804 17576
rect 74668 17527 74708 17536
rect 74667 16568 74709 16577
rect 74667 16528 74668 16568
rect 74708 16528 74709 16568
rect 74667 16519 74709 16528
rect 74380 15604 74455 15644
rect 74284 15520 74345 15560
rect 74305 15204 74345 15520
rect 74415 15204 74455 15604
rect 74668 15560 74708 16519
rect 74764 15644 74804 17536
rect 74956 15644 74996 17620
rect 75340 17620 75476 17660
rect 75148 17576 75188 17585
rect 75148 15728 75188 17536
rect 75340 16073 75380 17620
rect 75820 17610 75860 17695
rect 75532 17576 75572 17585
rect 75724 17576 75764 17585
rect 75572 17536 75668 17576
rect 75532 17527 75572 17536
rect 75339 16064 75381 16073
rect 75339 16024 75340 16064
rect 75380 16024 75381 16064
rect 75339 16015 75381 16024
rect 75148 15688 75476 15728
rect 75436 15644 75476 15688
rect 75628 15644 75668 17536
rect 74764 15604 74855 15644
rect 74956 15604 75255 15644
rect 75436 15604 75545 15644
rect 74668 15520 74745 15560
rect 74705 15204 74745 15520
rect 74815 15204 74855 15604
rect 75104 15392 75146 15401
rect 75104 15352 75105 15392
rect 75145 15352 75146 15392
rect 75104 15343 75146 15352
rect 75105 15204 75145 15343
rect 75215 15204 75255 15604
rect 75505 15204 75545 15604
rect 75615 15604 75668 15644
rect 75615 15204 75655 15604
rect 75724 15401 75764 17536
rect 75916 15644 75956 19048
rect 76108 19048 76684 19088
rect 75905 15604 75956 15644
rect 76012 18332 76052 18341
rect 76012 15644 76052 18292
rect 76012 15604 76055 15644
rect 75723 15392 75765 15401
rect 75723 15352 75724 15392
rect 75764 15352 75765 15392
rect 75723 15343 75765 15352
rect 75905 15204 75945 15604
rect 76015 15204 76055 15604
rect 76108 15476 76148 19048
rect 76684 19039 76724 19048
rect 76203 18920 76245 18929
rect 76203 18880 76204 18920
rect 76244 18880 76245 18920
rect 76203 18871 76245 18880
rect 76352 18920 76720 18929
rect 76392 18880 76434 18920
rect 76474 18880 76516 18920
rect 76556 18880 76598 18920
rect 76638 18880 76680 18920
rect 76352 18871 76720 18880
rect 76204 17828 76244 18871
rect 76972 18845 77012 19132
rect 77164 19088 77204 19097
rect 77068 19048 77164 19088
rect 76971 18836 77013 18845
rect 76971 18796 76972 18836
rect 77012 18796 77013 18836
rect 76971 18787 77013 18796
rect 76491 18584 76533 18593
rect 76491 18544 76492 18584
rect 76532 18544 76533 18584
rect 76491 18535 76533 18544
rect 76204 17779 76244 17788
rect 76492 17753 76532 18535
rect 76588 18332 76628 18341
rect 76628 18292 76724 18332
rect 76588 18283 76628 18292
rect 76587 17828 76629 17837
rect 76587 17788 76588 17828
rect 76628 17788 76629 17828
rect 76587 17779 76629 17788
rect 76491 17744 76533 17753
rect 76491 17704 76492 17744
rect 76532 17704 76533 17744
rect 76491 17695 76533 17704
rect 76588 17694 76628 17779
rect 76684 17585 76724 18292
rect 76972 17837 77012 18787
rect 76971 17828 77013 17837
rect 76971 17788 76972 17828
rect 77012 17788 77013 17828
rect 76971 17779 77013 17788
rect 76972 17694 77012 17779
rect 76396 17576 76436 17585
rect 76204 17536 76396 17576
rect 76204 15560 76244 17536
rect 76396 17527 76436 17536
rect 76683 17576 76725 17585
rect 76683 17536 76684 17576
rect 76724 17536 76725 17576
rect 76683 17527 76725 17536
rect 76780 17576 76820 17585
rect 76352 17408 76720 17417
rect 76392 17368 76434 17408
rect 76474 17368 76516 17408
rect 76556 17368 76598 17408
rect 76638 17368 76680 17408
rect 76352 17359 76720 17368
rect 76683 17240 76725 17249
rect 76683 17200 76684 17240
rect 76724 17200 76725 17240
rect 76683 17191 76725 17200
rect 76204 15520 76455 15560
rect 76108 15436 76345 15476
rect 76305 15204 76345 15436
rect 76415 15204 76455 15520
rect 76684 15392 76724 17191
rect 76780 15476 76820 17536
rect 77068 15644 77108 19048
rect 77164 19039 77204 19048
rect 77836 19088 77876 19097
rect 78028 19088 78068 19216
rect 77876 19048 77972 19088
rect 77836 19039 77876 19048
rect 77451 18836 77493 18845
rect 77451 18796 77452 18836
rect 77492 18796 77493 18836
rect 77451 18787 77493 18796
rect 77452 18593 77492 18787
rect 77451 18584 77493 18593
rect 77451 18544 77452 18584
rect 77492 18544 77493 18584
rect 77451 18535 77493 18544
rect 77452 18450 77492 18535
rect 77548 18332 77588 18341
rect 77452 18292 77548 18332
rect 77355 17828 77397 17837
rect 77355 17788 77356 17828
rect 77396 17788 77397 17828
rect 77355 17779 77397 17788
rect 77356 17694 77396 17779
rect 77164 17576 77204 17585
rect 77204 17536 77300 17576
rect 77164 17527 77204 17536
rect 77260 15644 77300 17536
rect 77068 15604 77145 15644
rect 76780 15436 76855 15476
rect 76684 15352 76745 15392
rect 76705 15204 76745 15352
rect 76815 15204 76855 15436
rect 77105 15204 77145 15604
rect 77215 15604 77300 15644
rect 77452 15644 77492 18292
rect 77548 18283 77588 18292
rect 77739 17828 77781 17837
rect 77739 17788 77740 17828
rect 77780 17788 77781 17828
rect 77739 17779 77781 17788
rect 77740 17744 77780 17779
rect 77740 17693 77780 17704
rect 77548 17576 77588 17585
rect 77836 17576 77876 17585
rect 77588 17536 77684 17576
rect 77548 17527 77588 17536
rect 77644 15644 77684 17536
rect 77452 15604 77545 15644
rect 77215 15204 77255 15604
rect 77505 15204 77545 15604
rect 77615 15604 77684 15644
rect 77615 15204 77655 15604
rect 77836 15569 77876 17536
rect 77932 15644 77972 19048
rect 78068 19048 78164 19088
rect 78028 19039 78068 19048
rect 78124 18929 78164 19048
rect 78123 18920 78165 18929
rect 78123 18880 78124 18920
rect 78164 18880 78165 18920
rect 78123 18871 78165 18880
rect 78124 18584 78164 18871
rect 78220 18845 78260 19300
rect 80523 19340 80565 19349
rect 80523 19300 80524 19340
rect 80564 19300 80565 19340
rect 80523 19291 80565 19300
rect 82059 19340 82101 19349
rect 82059 19300 82060 19340
rect 82100 19300 82101 19340
rect 82059 19291 82101 19300
rect 82347 19340 82389 19349
rect 82347 19300 82348 19340
rect 82388 19300 82389 19340
rect 82347 19291 82389 19300
rect 84075 19340 84117 19349
rect 84075 19300 84076 19340
rect 84116 19300 84117 19340
rect 84075 19291 84117 19300
rect 85611 19340 85653 19349
rect 85611 19300 85612 19340
rect 85652 19300 85653 19340
rect 85611 19291 85653 19300
rect 86572 19340 86612 19351
rect 86956 19349 86996 19804
rect 87052 19795 87092 19804
rect 93004 19844 93044 19853
rect 93044 19804 93140 19844
rect 93004 19795 93044 19804
rect 87112 19676 87480 19685
rect 87152 19636 87194 19676
rect 87234 19636 87276 19676
rect 87316 19636 87358 19676
rect 87398 19636 87440 19676
rect 87112 19627 87480 19636
rect 91112 19676 91480 19685
rect 91152 19636 91194 19676
rect 91234 19636 91276 19676
rect 91316 19636 91358 19676
rect 91398 19636 91440 19676
rect 91112 19627 91480 19636
rect 90124 19508 90164 19517
rect 89740 19468 90124 19508
rect 88204 19349 88244 19434
rect 78604 19256 78644 19265
rect 78604 18929 78644 19216
rect 80044 19256 80084 19265
rect 80084 19216 80372 19256
rect 78700 19088 78740 19097
rect 78603 18920 78645 18929
rect 78603 18880 78604 18920
rect 78644 18880 78645 18920
rect 78603 18871 78645 18880
rect 78219 18836 78261 18845
rect 78219 18796 78220 18836
rect 78260 18796 78261 18836
rect 78219 18787 78261 18796
rect 78124 17828 78164 18544
rect 78411 18500 78453 18509
rect 78411 18460 78412 18500
rect 78452 18460 78453 18500
rect 78411 18451 78453 18460
rect 78412 18366 78452 18451
rect 78220 18332 78260 18341
rect 78604 18332 78644 18341
rect 78260 18292 78356 18332
rect 78220 18283 78260 18292
rect 78219 17828 78261 17837
rect 78124 17788 78220 17828
rect 78260 17788 78261 17828
rect 78219 17779 78261 17788
rect 78220 17694 78260 17779
rect 78316 15644 78356 18292
rect 78508 18292 78604 18332
rect 77932 15604 78055 15644
rect 77835 15560 77877 15569
rect 77835 15520 77836 15560
rect 77876 15520 77877 15560
rect 77835 15511 77877 15520
rect 77904 15392 77946 15401
rect 77904 15352 77905 15392
rect 77945 15352 77946 15392
rect 77904 15343 77946 15352
rect 77905 15204 77945 15343
rect 78015 15204 78055 15604
rect 78305 15604 78356 15644
rect 78412 17576 78452 17585
rect 78305 15204 78345 15604
rect 78412 15476 78452 17536
rect 78508 15569 78548 18292
rect 78604 18283 78644 18292
rect 78700 17996 78740 19048
rect 79371 18920 79413 18929
rect 79371 18880 79372 18920
rect 79412 18880 79413 18920
rect 79371 18871 79413 18880
rect 78987 18836 79029 18845
rect 78987 18796 78988 18836
rect 79028 18796 79029 18836
rect 78987 18787 79029 18796
rect 78795 18500 78837 18509
rect 78795 18460 78796 18500
rect 78836 18460 78837 18500
rect 78795 18451 78837 18460
rect 78988 18500 79028 18787
rect 79372 18509 79412 18871
rect 80044 18509 80084 19216
rect 80140 19088 80180 19097
rect 80332 19088 80372 19216
rect 80524 19206 80564 19291
rect 81868 19181 81908 19212
rect 82060 19206 82100 19291
rect 81867 19172 81909 19181
rect 81867 19132 81868 19172
rect 81908 19132 81909 19172
rect 81867 19123 81909 19132
rect 80180 19048 80276 19088
rect 80140 19039 80180 19048
rect 78604 17956 78740 17996
rect 78796 18416 78836 18451
rect 78604 15644 78644 17956
rect 78796 17921 78836 18376
rect 78988 18257 79028 18460
rect 79371 18500 79413 18509
rect 79371 18460 79372 18500
rect 79412 18460 79413 18500
rect 79371 18451 79413 18460
rect 79851 18500 79893 18509
rect 79851 18460 79852 18500
rect 79892 18460 79893 18500
rect 79851 18451 79893 18460
rect 80043 18500 80085 18509
rect 80043 18460 80044 18500
rect 80084 18460 80180 18500
rect 80043 18451 80085 18460
rect 79372 18366 79412 18451
rect 79852 18366 79892 18451
rect 79564 18332 79604 18341
rect 80044 18332 80084 18341
rect 79604 18292 79700 18332
rect 79564 18283 79604 18292
rect 78987 18248 79029 18257
rect 78987 18208 78988 18248
rect 79028 18208 79029 18248
rect 78987 18199 79029 18208
rect 79112 18164 79480 18173
rect 79152 18124 79194 18164
rect 79234 18124 79276 18164
rect 79316 18124 79358 18164
rect 79398 18124 79440 18164
rect 79112 18115 79480 18124
rect 78795 17912 78837 17921
rect 78700 17872 78796 17912
rect 78836 17872 78837 17912
rect 78700 17828 78740 17872
rect 78795 17863 78837 17872
rect 79179 17912 79221 17921
rect 79179 17872 79180 17912
rect 79220 17872 79221 17912
rect 79179 17863 79221 17872
rect 79467 17912 79509 17921
rect 79467 17872 79468 17912
rect 79508 17872 79509 17912
rect 79467 17863 79509 17872
rect 78700 17779 78740 17788
rect 79180 17744 79220 17863
rect 79180 17695 79220 17704
rect 79468 17744 79508 17863
rect 79468 17695 79508 17704
rect 78892 17576 78932 17585
rect 79084 17576 79124 17585
rect 79564 17576 79604 17585
rect 78932 17536 79028 17576
rect 78892 17527 78932 17536
rect 78604 15604 78745 15644
rect 78507 15560 78549 15569
rect 78507 15520 78508 15560
rect 78548 15520 78549 15560
rect 78507 15511 78549 15520
rect 78412 15436 78455 15476
rect 78415 15204 78455 15436
rect 78705 15204 78745 15604
rect 78988 15401 79028 17536
rect 79084 15644 79124 17536
rect 79468 17536 79564 17576
rect 79468 15644 79508 17536
rect 79564 17527 79604 17536
rect 79660 15644 79700 18292
rect 79851 18248 79893 18257
rect 79851 18208 79852 18248
rect 79892 18208 79893 18248
rect 79851 18199 79893 18208
rect 79852 17744 79892 18199
rect 79852 17695 79892 17704
rect 79948 17576 79988 17585
rect 79084 15604 79145 15644
rect 79468 15604 79545 15644
rect 78814 15392 78856 15401
rect 78814 15352 78815 15392
rect 78855 15352 78856 15392
rect 78814 15343 78856 15352
rect 78987 15392 79029 15401
rect 78987 15352 78988 15392
rect 79028 15352 79029 15392
rect 78987 15343 79029 15352
rect 78815 15204 78855 15343
rect 79105 15204 79145 15604
rect 79214 15560 79256 15569
rect 79214 15520 79215 15560
rect 79255 15520 79256 15560
rect 79214 15511 79256 15520
rect 79215 15204 79255 15511
rect 79505 15204 79545 15604
rect 79615 15604 79700 15644
rect 79852 17536 79948 17576
rect 79852 15644 79892 17536
rect 79948 17527 79988 17536
rect 80044 15644 80084 18292
rect 80140 17828 80180 18460
rect 80140 17779 80180 17788
rect 80236 17660 80276 19048
rect 80332 19039 80372 19048
rect 81868 19088 81908 19123
rect 80352 18920 80720 18929
rect 80392 18880 80434 18920
rect 80474 18880 80516 18920
rect 80556 18880 80598 18920
rect 80638 18880 80680 18920
rect 80352 18871 80720 18880
rect 81388 18509 81428 18594
rect 80523 18500 80565 18509
rect 80523 18460 80524 18500
rect 80564 18460 80565 18500
rect 80523 18451 80565 18460
rect 81003 18500 81045 18509
rect 81003 18460 81004 18500
rect 81044 18460 81045 18500
rect 81003 18451 81045 18460
rect 81387 18500 81429 18509
rect 81387 18460 81388 18500
rect 81428 18460 81429 18500
rect 81387 18451 81429 18460
rect 81772 18500 81812 18528
rect 81868 18500 81908 19048
rect 82252 18500 82292 18509
rect 81812 18460 82252 18500
rect 81772 18451 81812 18460
rect 80524 17828 80564 18451
rect 80524 17779 80564 17788
rect 81004 17744 81044 18451
rect 81196 18332 81236 18341
rect 81580 18332 81620 18341
rect 81964 18332 82004 18341
rect 81236 18292 81428 18332
rect 81196 18283 81236 18292
rect 81291 17744 81333 17753
rect 81044 17704 81292 17744
rect 81332 17704 81333 17744
rect 81004 17695 81044 17704
rect 81291 17695 81333 17704
rect 79852 15604 79945 15644
rect 79615 15204 79655 15604
rect 79905 15204 79945 15604
rect 80015 15604 80084 15644
rect 80140 17620 80276 17660
rect 80015 15204 80055 15604
rect 80140 15476 80180 17620
rect 80716 17585 80756 17670
rect 81292 17610 81332 17695
rect 80332 17576 80372 17585
rect 80236 17536 80332 17576
rect 80236 15560 80276 17536
rect 80332 17527 80372 17536
rect 80715 17576 80757 17585
rect 80715 17536 80716 17576
rect 80756 17536 80757 17576
rect 80715 17527 80757 17536
rect 80908 17576 80948 17585
rect 80352 17408 80720 17417
rect 80392 17368 80434 17408
rect 80474 17368 80516 17408
rect 80556 17368 80598 17408
rect 80638 17368 80680 17408
rect 80352 17359 80720 17368
rect 80908 15728 80948 17536
rect 81003 17576 81045 17585
rect 81003 17536 81004 17576
rect 81044 17536 81045 17576
rect 81003 17527 81045 17536
rect 81196 17576 81236 17585
rect 80716 15688 80948 15728
rect 80716 15644 80756 15688
rect 80705 15604 80756 15644
rect 80236 15520 80455 15560
rect 80140 15436 80345 15476
rect 80305 15204 80345 15436
rect 80415 15204 80455 15520
rect 80705 15204 80745 15604
rect 81004 15392 81044 17527
rect 81196 15644 81236 17536
rect 80815 15352 81044 15392
rect 81105 15604 81236 15644
rect 80815 15204 80855 15352
rect 81105 15204 81145 15604
rect 81388 15560 81428 18292
rect 81620 18292 81716 18332
rect 81580 18283 81620 18292
rect 81484 17753 81524 17838
rect 81483 17744 81525 17753
rect 81483 17704 81484 17744
rect 81524 17704 81525 17744
rect 81483 17695 81525 17704
rect 81580 17576 81620 17585
rect 81484 17536 81580 17576
rect 81484 15644 81524 17536
rect 81580 17527 81620 17536
rect 81676 15644 81716 18292
rect 82004 18292 82100 18332
rect 81964 18283 82004 18292
rect 81964 17753 82004 17838
rect 81963 17744 82005 17753
rect 81963 17704 81964 17744
rect 82004 17704 82005 17744
rect 81963 17695 82005 17704
rect 81868 17660 81908 17669
rect 81868 17576 81908 17620
rect 81868 17536 82004 17576
rect 81964 15644 82004 17536
rect 81484 15604 81545 15644
rect 81215 15520 81428 15560
rect 81215 15204 81255 15520
rect 81505 15204 81545 15604
rect 81615 15604 81716 15644
rect 81905 15604 82004 15644
rect 81615 15204 81655 15604
rect 81905 15204 81945 15604
rect 82060 15560 82100 18292
rect 82252 17744 82292 18460
rect 82348 17753 82388 19291
rect 82636 19256 82676 19267
rect 82636 19181 82676 19216
rect 84076 19206 84116 19291
rect 85612 19206 85652 19291
rect 86572 19265 86612 19300
rect 86763 19340 86805 19349
rect 86763 19300 86764 19340
rect 86804 19300 86805 19340
rect 86763 19291 86805 19300
rect 86955 19340 86997 19349
rect 86955 19300 86956 19340
rect 86996 19300 86997 19340
rect 86955 19291 86997 19300
rect 87436 19340 87476 19349
rect 86571 19256 86613 19265
rect 86571 19216 86572 19256
rect 86612 19216 86613 19256
rect 86571 19207 86613 19216
rect 86764 19206 86804 19291
rect 82635 19172 82677 19181
rect 82635 19132 82636 19172
rect 82676 19132 82677 19172
rect 82635 19123 82677 19132
rect 83019 19172 83061 19181
rect 83019 19132 83020 19172
rect 83060 19132 83061 19172
rect 83019 19123 83061 19132
rect 86955 19172 86997 19181
rect 86955 19132 86956 19172
rect 86996 19132 86997 19172
rect 86955 19123 86997 19132
rect 82444 18332 82484 18341
rect 82252 17695 82292 17704
rect 82347 17744 82389 17753
rect 82347 17704 82348 17744
rect 82388 17704 82389 17744
rect 82347 17695 82389 17704
rect 82348 17576 82388 17585
rect 82252 17536 82348 17576
rect 82252 15644 82292 17536
rect 82348 17527 82388 17536
rect 82444 15644 82484 18292
rect 82636 17828 82676 19123
rect 82636 17779 82676 17788
rect 82732 19088 82772 19097
rect 82732 15644 82772 19048
rect 83020 18500 83060 19123
rect 83884 19088 83924 19097
rect 82924 18460 83020 18500
rect 82924 17744 82964 18460
rect 83020 18451 83060 18460
rect 83403 18500 83445 18509
rect 83403 18460 83404 18500
rect 83444 18460 83445 18500
rect 83403 18451 83445 18460
rect 83787 18500 83829 18509
rect 83884 18500 83924 19048
rect 85804 19088 85844 19097
rect 86380 19088 86420 19097
rect 85844 19048 85940 19088
rect 85804 19039 85844 19048
rect 84352 18920 84720 18929
rect 84392 18880 84434 18920
rect 84474 18880 84516 18920
rect 84556 18880 84598 18920
rect 84638 18880 84680 18920
rect 84352 18871 84720 18880
rect 85036 18584 85076 18595
rect 85036 18509 85076 18544
rect 85900 18509 85940 19048
rect 86284 18584 86324 18595
rect 86380 18584 86420 19048
rect 86956 19088 86996 19123
rect 86956 19037 86996 19048
rect 87436 18593 87476 19300
rect 88203 19340 88245 19349
rect 88203 19300 88204 19340
rect 88244 19300 88245 19340
rect 88203 19291 88245 19300
rect 89740 19340 89780 19468
rect 90124 19459 90164 19468
rect 92908 19424 92948 19433
rect 89740 19291 89780 19300
rect 89932 19340 89972 19351
rect 89932 19265 89972 19300
rect 91372 19340 91412 19349
rect 88492 19256 88532 19265
rect 88300 19216 88492 19256
rect 88300 19172 88340 19216
rect 88492 19207 88532 19216
rect 89931 19256 89973 19265
rect 89931 19216 89932 19256
rect 89972 19216 89973 19256
rect 89931 19207 89973 19216
rect 88108 19132 88340 19172
rect 87628 19088 87668 19097
rect 86571 18584 86613 18593
rect 86380 18544 86572 18584
rect 86612 18544 86613 18584
rect 86284 18509 86324 18544
rect 86571 18535 86613 18544
rect 87051 18584 87093 18593
rect 87051 18544 87052 18584
rect 87092 18544 87093 18584
rect 87051 18535 87093 18544
rect 87435 18584 87477 18593
rect 87435 18544 87436 18584
rect 87476 18544 87477 18584
rect 87435 18535 87477 18544
rect 83787 18460 83788 18500
rect 83828 18460 83924 18500
rect 84267 18500 84309 18509
rect 84267 18460 84268 18500
rect 84308 18460 84309 18500
rect 83787 18451 83829 18460
rect 84267 18451 84309 18460
rect 84651 18500 84693 18509
rect 84651 18460 84652 18500
rect 84692 18460 84693 18500
rect 84651 18451 84693 18460
rect 85035 18500 85077 18509
rect 85515 18500 85557 18509
rect 85899 18500 85941 18509
rect 85035 18460 85036 18500
rect 85076 18460 85077 18500
rect 85035 18451 85077 18460
rect 85420 18460 85516 18500
rect 85556 18460 85557 18500
rect 83404 18366 83444 18451
rect 83212 18332 83252 18341
rect 83020 18292 83212 18332
rect 83020 17996 83060 18292
rect 83212 18283 83252 18292
rect 83596 18332 83636 18341
rect 83112 18164 83480 18173
rect 83152 18124 83194 18164
rect 83234 18124 83276 18164
rect 83316 18124 83358 18164
rect 83398 18124 83440 18164
rect 83112 18115 83480 18124
rect 83020 17956 83252 17996
rect 83020 17744 83060 17753
rect 82924 17704 83020 17744
rect 83020 17695 83060 17704
rect 82252 15604 82345 15644
rect 82015 15520 82100 15560
rect 82015 15204 82055 15520
rect 82305 15204 82345 15604
rect 82415 15604 82484 15644
rect 82705 15604 82772 15644
rect 82828 17576 82868 17585
rect 82415 15204 82455 15604
rect 82705 15204 82745 15604
rect 82828 15476 82868 17536
rect 83116 17576 83156 17585
rect 83116 15644 83156 17536
rect 82815 15436 82868 15476
rect 83105 15604 83156 15644
rect 83212 15644 83252 17956
rect 83403 17744 83445 17753
rect 83403 17704 83404 17744
rect 83444 17704 83445 17744
rect 83403 17695 83445 17704
rect 83404 17610 83444 17695
rect 83500 17576 83540 17585
rect 83500 15644 83540 17536
rect 83596 15644 83636 18292
rect 83788 17753 83828 18451
rect 84268 18366 84308 18451
rect 84652 18366 84692 18451
rect 83980 18332 84020 18341
rect 83787 17744 83829 17753
rect 83787 17704 83788 17744
rect 83828 17704 83829 17744
rect 83787 17695 83829 17704
rect 83788 17610 83828 17695
rect 83884 17576 83924 17585
rect 83884 15644 83924 17536
rect 83980 15728 84020 18292
rect 84460 18332 84500 18341
rect 84171 17744 84213 17753
rect 84171 17704 84172 17744
rect 84212 17704 84213 17744
rect 84171 17695 84213 17704
rect 84172 17610 84212 17695
rect 84460 17585 84500 18292
rect 84844 18332 84884 18341
rect 85132 18332 85172 18341
rect 84747 17828 84789 17837
rect 84747 17788 84748 17828
rect 84788 17788 84789 17828
rect 84747 17779 84789 17788
rect 84748 17744 84788 17779
rect 84748 17693 84788 17704
rect 84651 17660 84693 17669
rect 84651 17620 84652 17660
rect 84692 17620 84693 17660
rect 84651 17611 84693 17620
rect 84268 17576 84308 17585
rect 83980 15688 84055 15728
rect 83212 15604 83255 15644
rect 83500 15604 83545 15644
rect 83596 15604 83655 15644
rect 83884 15604 83945 15644
rect 82815 15204 82855 15436
rect 83105 15204 83145 15604
rect 83215 15204 83255 15604
rect 83505 15204 83545 15604
rect 83615 15204 83655 15604
rect 83905 15204 83945 15604
rect 84015 15204 84055 15688
rect 84268 15644 84308 17536
rect 84459 17576 84501 17585
rect 84459 17536 84460 17576
rect 84500 17536 84501 17576
rect 84459 17527 84501 17536
rect 84652 17526 84692 17611
rect 84352 17408 84720 17417
rect 84392 17368 84434 17408
rect 84474 17368 84516 17408
rect 84556 17368 84598 17408
rect 84638 17368 84680 17408
rect 84352 17359 84720 17368
rect 84844 15644 84884 18292
rect 85036 18292 85132 18332
rect 84940 17837 84980 17922
rect 84939 17828 84981 17837
rect 84939 17788 84940 17828
rect 84980 17788 84981 17828
rect 84939 17779 84981 17788
rect 85036 17660 85076 18292
rect 85132 18283 85172 18292
rect 85420 17837 85460 18460
rect 85515 18451 85557 18460
rect 85804 18460 85900 18500
rect 85940 18460 85941 18500
rect 85516 18366 85556 18451
rect 85708 18332 85748 18341
rect 85419 17828 85461 17837
rect 85419 17788 85420 17828
rect 85460 17788 85461 17828
rect 85419 17779 85461 17788
rect 85420 17744 85460 17779
rect 85420 17694 85460 17704
rect 84268 15604 84345 15644
rect 84305 15204 84345 15604
rect 84815 15604 84884 15644
rect 84940 17620 85076 17660
rect 84414 15560 84456 15569
rect 84414 15520 84415 15560
rect 84455 15520 84456 15560
rect 84414 15511 84456 15520
rect 84704 15560 84746 15569
rect 84704 15520 84705 15560
rect 84745 15520 84746 15560
rect 84704 15511 84746 15520
rect 84415 15204 84455 15511
rect 84705 15204 84745 15511
rect 84815 15204 84855 15604
rect 84940 15569 84980 17620
rect 85132 17576 85172 17585
rect 85035 17492 85077 17501
rect 85035 17452 85036 17492
rect 85076 17452 85077 17492
rect 85035 17443 85077 17452
rect 84939 15560 84981 15569
rect 84939 15520 84940 15560
rect 84980 15520 84981 15560
rect 84939 15511 84981 15520
rect 85036 15392 85076 17443
rect 85132 15644 85172 17536
rect 85516 17576 85556 17585
rect 85516 15644 85556 17536
rect 85708 16400 85748 18292
rect 85804 17744 85844 18460
rect 85899 18451 85941 18460
rect 86283 18500 86325 18509
rect 86283 18460 86284 18500
rect 86324 18460 86325 18500
rect 86283 18451 86325 18460
rect 86572 18500 86612 18535
rect 85900 18366 85940 18451
rect 85804 17695 85844 17704
rect 86092 18332 86132 18341
rect 86380 18332 86420 18341
rect 85132 15604 85255 15644
rect 85036 15352 85145 15392
rect 85105 15204 85145 15352
rect 85215 15204 85255 15604
rect 85505 15604 85556 15644
rect 85612 16360 85748 16400
rect 85900 17576 85940 17585
rect 85612 15644 85652 16360
rect 85900 15644 85940 17536
rect 86092 15644 86132 18292
rect 86284 18292 86380 18332
rect 86188 17828 86228 17839
rect 86188 17753 86228 17788
rect 86187 17744 86229 17753
rect 86187 17704 86188 17744
rect 86228 17704 86229 17744
rect 86187 17695 86229 17704
rect 85612 15604 85655 15644
rect 85900 15604 85945 15644
rect 85505 15204 85545 15604
rect 85615 15204 85655 15604
rect 85905 15204 85945 15604
rect 86015 15604 86132 15644
rect 86015 15204 86055 15604
rect 86284 15392 86324 18292
rect 86380 18283 86420 18292
rect 86572 17753 86612 18460
rect 87052 18500 87092 18535
rect 87052 18449 87092 18460
rect 86764 18332 86804 18341
rect 87244 18332 87284 18341
rect 86804 18292 86900 18332
rect 86764 18283 86804 18292
rect 86571 17744 86613 17753
rect 86571 17704 86572 17744
rect 86612 17704 86613 17744
rect 86571 17695 86613 17704
rect 86572 17610 86612 17695
rect 86380 17576 86420 17585
rect 86380 15476 86420 17536
rect 86668 17576 86708 17585
rect 86668 15644 86708 17536
rect 86860 15644 86900 18292
rect 86956 18292 87244 18332
rect 86956 17912 86996 18292
rect 87244 18283 87284 18292
rect 87112 18164 87480 18173
rect 87152 18124 87194 18164
rect 87234 18124 87276 18164
rect 87316 18124 87358 18164
rect 87398 18124 87440 18164
rect 87112 18115 87480 18124
rect 86956 17872 87284 17912
rect 87051 17744 87093 17753
rect 87051 17704 87052 17744
rect 87092 17704 87093 17744
rect 87051 17695 87093 17704
rect 87052 17610 87092 17695
rect 87148 17576 87188 17585
rect 87148 15728 87188 17536
rect 86668 15604 86745 15644
rect 86380 15436 86455 15476
rect 86284 15352 86345 15392
rect 86305 15204 86345 15352
rect 86415 15204 86455 15436
rect 86705 15204 86745 15604
rect 86815 15604 86900 15644
rect 87052 15688 87188 15728
rect 86815 15204 86855 15604
rect 87052 15560 87092 15688
rect 87244 15644 87284 17872
rect 87435 17744 87477 17753
rect 87435 17704 87436 17744
rect 87476 17704 87477 17744
rect 87435 17695 87477 17704
rect 87436 17610 87476 17695
rect 87532 17576 87572 17585
rect 87532 15644 87572 17536
rect 87628 15644 87668 19048
rect 88012 19088 88052 19097
rect 88108 19088 88148 19132
rect 88396 19088 88436 19097
rect 88052 19048 88148 19088
rect 88204 19048 88396 19088
rect 88012 18509 88052 19048
rect 88204 18668 88244 19048
rect 88396 19039 88436 19048
rect 89548 19088 89588 19097
rect 88352 18920 88720 18929
rect 88392 18880 88434 18920
rect 88474 18880 88516 18920
rect 88556 18880 88598 18920
rect 88638 18880 88680 18920
rect 88352 18871 88720 18880
rect 89548 18668 89588 19048
rect 90124 19088 90164 19097
rect 90124 18929 90164 19048
rect 91372 18929 91412 19300
rect 92524 19340 92564 19349
rect 92908 19340 92948 19384
rect 93100 19349 93140 19804
rect 93099 19340 93141 19349
rect 92564 19300 93044 19340
rect 92524 19291 92564 19300
rect 91564 19088 91604 19097
rect 91468 19048 91564 19088
rect 90123 18920 90165 18929
rect 90123 18880 90124 18920
rect 90164 18880 90165 18920
rect 90123 18871 90165 18880
rect 90507 18920 90549 18929
rect 90507 18880 90508 18920
rect 90548 18880 90549 18920
rect 90507 18871 90549 18880
rect 91371 18920 91413 18929
rect 91371 18880 91372 18920
rect 91412 18880 91413 18920
rect 91371 18871 91413 18880
rect 88108 18628 88244 18668
rect 89452 18628 89588 18668
rect 87723 18500 87765 18509
rect 87723 18460 87724 18500
rect 87764 18460 87765 18500
rect 87723 18451 87765 18460
rect 88011 18500 88053 18509
rect 88011 18460 88012 18500
rect 88052 18460 88053 18500
rect 88011 18451 88053 18460
rect 87724 18366 87764 18451
rect 87916 18332 87956 18341
rect 87956 18292 88052 18332
rect 87916 18283 87956 18292
rect 87915 17660 87957 17669
rect 87915 17620 87916 17660
rect 87956 17620 87957 17660
rect 87915 17611 87957 17620
rect 87916 15644 87956 17611
rect 87215 15604 87284 15644
rect 87505 15604 87572 15644
rect 87615 15604 87668 15644
rect 87905 15604 87956 15644
rect 88012 15644 88052 18292
rect 88108 17669 88148 18628
rect 89452 18595 89492 18628
rect 89452 18546 89492 18555
rect 89548 18509 89588 18628
rect 89740 18509 89780 18594
rect 88203 18500 88245 18509
rect 88203 18460 88204 18500
rect 88244 18460 88245 18500
rect 88203 18451 88245 18460
rect 88587 18500 88629 18509
rect 88587 18460 88588 18500
rect 88628 18460 88629 18500
rect 88587 18451 88629 18460
rect 88971 18500 89013 18509
rect 88971 18460 88972 18500
rect 89012 18460 89013 18500
rect 89547 18500 89589 18509
rect 89547 18497 89548 18500
rect 88971 18451 89013 18460
rect 89454 18460 89548 18497
rect 89588 18460 89589 18500
rect 89454 18457 89589 18460
rect 88204 17744 88244 18451
rect 88204 17695 88244 17704
rect 88396 18332 88436 18341
rect 88107 17660 88149 17669
rect 88107 17620 88108 17660
rect 88148 17620 88149 17660
rect 88107 17611 88149 17620
rect 88396 17585 88436 18292
rect 88588 17753 88628 18451
rect 88972 18366 89012 18451
rect 89454 18416 89494 18457
rect 89547 18451 89589 18457
rect 89739 18500 89781 18509
rect 89739 18460 89740 18500
rect 89780 18460 89781 18500
rect 89739 18451 89781 18460
rect 90123 18500 90165 18509
rect 90123 18460 90124 18500
rect 90164 18460 90165 18500
rect 90123 18451 90165 18460
rect 89452 18376 89494 18416
rect 88780 18332 88820 18341
rect 89164 18332 89204 18341
rect 88820 18292 88916 18332
rect 88780 18283 88820 18292
rect 88587 17744 88629 17753
rect 88587 17704 88588 17744
rect 88628 17704 88629 17744
rect 88587 17695 88629 17704
rect 88588 17610 88628 17695
rect 88300 17576 88340 17585
rect 88204 17536 88300 17576
rect 88204 15644 88244 17536
rect 88300 17527 88340 17536
rect 88395 17576 88437 17585
rect 88395 17536 88396 17576
rect 88436 17536 88437 17576
rect 88395 17527 88437 17536
rect 88684 17576 88724 17585
rect 88724 17536 88820 17576
rect 88684 17527 88724 17536
rect 88352 17408 88720 17417
rect 88392 17368 88434 17408
rect 88474 17368 88516 17408
rect 88556 17368 88598 17408
rect 88638 17368 88680 17408
rect 88352 17359 88720 17368
rect 88395 17240 88437 17249
rect 88395 17200 88396 17240
rect 88436 17200 88437 17240
rect 88395 17191 88437 17200
rect 88396 15644 88436 17191
rect 88780 15644 88820 17536
rect 88012 15604 88055 15644
rect 88204 15604 88345 15644
rect 88396 15604 88455 15644
rect 87052 15520 87145 15560
rect 87105 15204 87145 15520
rect 87215 15204 87255 15604
rect 87505 15204 87545 15604
rect 87615 15204 87655 15604
rect 87905 15204 87945 15604
rect 88015 15204 88055 15604
rect 88305 15204 88345 15604
rect 88415 15204 88455 15604
rect 88705 15604 88820 15644
rect 88705 15204 88745 15604
rect 88876 15560 88916 18292
rect 89204 18292 89300 18332
rect 89164 18283 89204 18292
rect 89068 17753 89108 17838
rect 89067 17744 89109 17753
rect 89067 17704 89068 17744
rect 89108 17704 89109 17744
rect 89067 17695 89109 17704
rect 89164 17576 89204 17585
rect 89068 17536 89164 17576
rect 89068 15644 89108 17536
rect 89164 17527 89204 17536
rect 89260 15644 89300 18292
rect 89452 17828 89492 18376
rect 90124 18366 90164 18451
rect 89548 18332 89588 18341
rect 89932 18332 89972 18341
rect 90316 18332 90356 18341
rect 89588 18292 89780 18332
rect 89548 18283 89588 18292
rect 89452 17753 89492 17788
rect 89451 17744 89493 17753
rect 89451 17704 89452 17744
rect 89492 17704 89493 17744
rect 89451 17695 89493 17704
rect 89452 17664 89492 17695
rect 89068 15604 89145 15644
rect 88815 15520 88916 15560
rect 88815 15204 88855 15520
rect 89105 15204 89145 15604
rect 89215 15604 89300 15644
rect 89644 17576 89684 17585
rect 89215 15204 89255 15604
rect 89504 15476 89546 15485
rect 89644 15476 89684 17536
rect 89740 15560 89780 18292
rect 89972 18292 90068 18332
rect 89932 18283 89972 18292
rect 89932 17753 89972 17838
rect 89931 17744 89973 17753
rect 89931 17704 89932 17744
rect 89972 17704 89973 17744
rect 89931 17695 89973 17704
rect 89836 17576 89876 17585
rect 89836 15737 89876 17536
rect 89835 15728 89877 15737
rect 89835 15688 89836 15728
rect 89876 15688 89877 15728
rect 89835 15679 89877 15688
rect 90028 15644 90068 18292
rect 90356 18292 90452 18332
rect 90316 18283 90356 18292
rect 90220 17753 90260 17838
rect 90219 17744 90261 17753
rect 90219 17704 90220 17744
rect 90260 17704 90261 17744
rect 90219 17695 90261 17704
rect 90316 17576 90356 17585
rect 90316 15644 90356 17536
rect 90015 15604 90068 15644
rect 90305 15604 90356 15644
rect 90412 15644 90452 18292
rect 90508 17744 90548 18871
rect 91468 18593 91508 19048
rect 91564 19039 91604 19048
rect 92716 19088 92756 19097
rect 92756 19048 92852 19088
rect 92716 19039 92756 19048
rect 92352 18920 92720 18929
rect 92392 18880 92434 18920
rect 92474 18880 92516 18920
rect 92556 18880 92598 18920
rect 92638 18880 92680 18920
rect 92352 18871 92720 18880
rect 92812 18836 92852 19048
rect 93004 18836 93044 19300
rect 93099 19300 93100 19340
rect 93140 19300 93141 19340
rect 93099 19291 93141 19300
rect 93100 19206 93140 19291
rect 93196 19265 93236 19972
rect 95112 19676 95480 19685
rect 95152 19636 95194 19676
rect 95234 19636 95276 19676
rect 95316 19636 95358 19676
rect 95398 19636 95440 19676
rect 95112 19627 95480 19636
rect 99112 19676 99480 19685
rect 99152 19636 99194 19676
rect 99234 19636 99276 19676
rect 99316 19636 99358 19676
rect 99398 19636 99440 19676
rect 99112 19627 99480 19636
rect 94155 19340 94197 19349
rect 94155 19300 94156 19340
rect 94196 19300 94197 19340
rect 94155 19291 94197 19300
rect 95787 19340 95829 19349
rect 95787 19300 95788 19340
rect 95828 19300 95829 19340
rect 95787 19291 95829 19300
rect 97131 19340 97173 19349
rect 97131 19300 97132 19340
rect 97172 19300 97173 19340
rect 97131 19291 97173 19300
rect 93195 19256 93237 19265
rect 93195 19216 93196 19256
rect 93236 19216 93237 19256
rect 93195 19207 93237 19216
rect 92812 18796 92961 18836
rect 93004 18796 93140 18836
rect 92921 18752 92961 18796
rect 92921 18712 93044 18752
rect 91467 18584 91509 18593
rect 91276 18544 91468 18584
rect 91508 18544 91509 18584
rect 90603 18500 90645 18509
rect 90603 18460 90604 18500
rect 90644 18460 90645 18500
rect 90603 18451 90645 18460
rect 91276 18500 91316 18544
rect 91467 18535 91509 18544
rect 91851 18584 91893 18593
rect 91851 18544 91852 18584
rect 91892 18544 91893 18584
rect 91851 18535 91893 18544
rect 92235 18584 92277 18593
rect 92235 18544 92236 18584
rect 92276 18544 92277 18584
rect 92235 18535 92277 18544
rect 92908 18584 92948 18595
rect 91276 18451 91316 18460
rect 91852 18500 91892 18535
rect 90604 18366 90644 18451
rect 90796 18332 90836 18341
rect 90603 17744 90645 17753
rect 90508 17704 90604 17744
rect 90644 17704 90645 17744
rect 90603 17695 90645 17704
rect 90604 17610 90644 17695
rect 90700 17576 90740 17585
rect 90700 17156 90740 17536
rect 90604 17116 90740 17156
rect 90604 15644 90644 17116
rect 90796 15644 90836 18292
rect 91468 18332 91508 18341
rect 91660 18332 91700 18341
rect 91508 18292 91604 18332
rect 91468 18283 91508 18292
rect 91112 18164 91480 18173
rect 91152 18124 91194 18164
rect 91234 18124 91276 18164
rect 91316 18124 91358 18164
rect 91398 18124 91440 18164
rect 91112 18115 91480 18124
rect 90987 17744 91029 17753
rect 90987 17704 90988 17744
rect 91028 17704 91029 17744
rect 90987 17695 91029 17704
rect 91371 17744 91413 17753
rect 91371 17704 91372 17744
rect 91412 17704 91413 17744
rect 91371 17695 91413 17704
rect 90988 17610 91028 17695
rect 91372 17610 91412 17695
rect 91084 17576 91124 17585
rect 91084 15644 91124 17536
rect 91468 17576 91508 17585
rect 91179 16568 91221 16577
rect 91179 16528 91180 16568
rect 91220 16528 91221 16568
rect 91179 16519 91221 16528
rect 91180 15728 91220 16519
rect 91180 15688 91255 15728
rect 90412 15604 90455 15644
rect 90604 15604 90745 15644
rect 90796 15604 90855 15644
rect 91084 15604 91145 15644
rect 89740 15520 89945 15560
rect 89504 15436 89505 15476
rect 89545 15436 89546 15476
rect 89504 15427 89546 15436
rect 89615 15436 89684 15476
rect 89505 15204 89545 15427
rect 89615 15204 89655 15436
rect 89905 15204 89945 15520
rect 90015 15204 90055 15604
rect 90305 15204 90345 15604
rect 90415 15204 90455 15604
rect 90705 15204 90745 15604
rect 90815 15204 90855 15604
rect 91105 15204 91145 15604
rect 91215 15204 91255 15688
rect 91468 15644 91508 17536
rect 91564 15728 91604 18292
rect 91660 16577 91700 18292
rect 91852 17753 91892 18460
rect 92236 18500 92276 18535
rect 92908 18509 92948 18544
rect 92236 18449 92276 18460
rect 92619 18500 92661 18509
rect 92619 18460 92620 18500
rect 92660 18460 92661 18500
rect 92619 18451 92661 18460
rect 92907 18500 92949 18509
rect 92907 18460 92908 18500
rect 92948 18460 92949 18500
rect 92907 18451 92949 18460
rect 92620 18366 92660 18451
rect 92044 18332 92084 18341
rect 92428 18332 92468 18341
rect 92812 18332 92852 18341
rect 91851 17744 91893 17753
rect 91851 17704 91852 17744
rect 91892 17704 91893 17744
rect 91851 17695 91893 17704
rect 91948 17576 91988 17585
rect 91852 17536 91948 17576
rect 91659 16568 91701 16577
rect 91659 16528 91660 16568
rect 91700 16528 91701 16568
rect 91659 16519 91701 16528
rect 91564 15688 91655 15728
rect 91468 15604 91545 15644
rect 91505 15204 91545 15604
rect 91615 15204 91655 15688
rect 91852 15644 91892 17536
rect 91948 17527 91988 17536
rect 92044 15644 92084 18292
rect 91852 15604 91945 15644
rect 91905 15204 91945 15604
rect 92015 15604 92084 15644
rect 92140 18292 92428 18332
rect 92015 15204 92055 15604
rect 92140 15569 92180 18292
rect 92428 18283 92468 18292
rect 92716 18292 92812 18332
rect 92236 17753 92276 17838
rect 92235 17744 92277 17753
rect 92235 17704 92236 17744
rect 92276 17704 92277 17744
rect 92235 17695 92277 17704
rect 92332 17576 92372 17585
rect 92236 17536 92332 17576
rect 92716 17576 92756 18292
rect 92812 18283 92852 18292
rect 92811 17996 92853 18005
rect 92811 17956 92812 17996
rect 92852 17956 92853 17996
rect 92811 17947 92853 17956
rect 92812 17744 92852 17947
rect 92812 17695 92852 17704
rect 92907 17660 92949 17669
rect 92907 17620 92908 17660
rect 92948 17620 92949 17660
rect 92907 17611 92949 17620
rect 92716 17536 92852 17576
rect 92139 15560 92181 15569
rect 92139 15520 92140 15560
rect 92180 15520 92181 15560
rect 92236 15560 92276 17536
rect 92332 17527 92372 17536
rect 92352 17408 92720 17417
rect 92392 17368 92434 17408
rect 92474 17368 92516 17408
rect 92556 17368 92598 17408
rect 92638 17368 92680 17408
rect 92352 17359 92720 17368
rect 92812 15644 92852 17536
rect 92908 17526 92948 17611
rect 92705 15604 92852 15644
rect 92414 15560 92456 15569
rect 92236 15520 92345 15560
rect 92139 15511 92181 15520
rect 92305 15204 92345 15520
rect 92414 15520 92415 15560
rect 92455 15520 92456 15560
rect 92414 15511 92456 15520
rect 92415 15204 92455 15511
rect 92705 15204 92745 15604
rect 93004 15560 93044 18712
rect 93100 18509 93140 18796
rect 93196 18593 93236 19207
rect 94156 19206 94196 19291
rect 95788 19206 95828 19291
rect 93964 19088 94004 19097
rect 95596 19088 95636 19097
rect 93195 18584 93237 18593
rect 93195 18544 93196 18584
rect 93236 18544 93237 18584
rect 93195 18535 93237 18544
rect 93099 18500 93141 18509
rect 93099 18460 93100 18500
rect 93140 18460 93141 18500
rect 93099 18451 93141 18460
rect 93100 17828 93140 18451
rect 93196 18005 93236 18535
rect 93868 18500 93908 18509
rect 93964 18500 94004 19048
rect 95500 19048 95596 19088
rect 95115 18584 95157 18593
rect 95115 18544 95116 18584
rect 95156 18544 95157 18584
rect 95115 18535 95157 18544
rect 94252 18500 94292 18509
rect 93908 18460 94252 18500
rect 93868 18451 93908 18460
rect 93292 18332 93332 18341
rect 93195 17996 93237 18005
rect 93195 17956 93196 17996
rect 93236 17956 93237 17996
rect 93195 17947 93237 17956
rect 93195 17828 93237 17837
rect 93100 17788 93196 17828
rect 93236 17788 93237 17828
rect 93188 17779 93237 17788
rect 93188 17749 93228 17779
rect 93188 17672 93228 17709
rect 93100 17576 93140 17585
rect 93100 15644 93140 17536
rect 93100 15604 93145 15644
rect 92815 15520 93044 15560
rect 92815 15204 92855 15520
rect 93105 15204 93145 15604
rect 93292 15392 93332 18292
rect 93771 17828 93813 17837
rect 93771 17788 93772 17828
rect 93812 17788 93813 17828
rect 93771 17779 93813 17788
rect 93772 17694 93812 17779
rect 93964 17744 94004 18460
rect 94060 18332 94100 18341
rect 94100 18292 94196 18332
rect 94060 18283 94100 18292
rect 94060 17744 94100 17753
rect 93964 17704 94060 17744
rect 94060 17695 94100 17704
rect 93483 17660 93525 17669
rect 93483 17620 93484 17660
rect 93524 17620 93525 17660
rect 93483 17611 93525 17620
rect 93215 15352 93332 15392
rect 93484 15392 93524 17611
rect 93580 17576 93620 17585
rect 93964 17576 94004 17585
rect 93580 15476 93620 17536
rect 93868 17536 93964 17576
rect 93868 15644 93908 17536
rect 93964 17527 94004 17536
rect 94156 15644 94196 18292
rect 94252 17744 94292 18460
rect 94924 18500 94964 18509
rect 94252 17695 94292 17704
rect 94444 18332 94484 18341
rect 94348 17576 94388 17585
rect 93868 15604 93945 15644
rect 93580 15436 93655 15476
rect 93484 15352 93545 15392
rect 93215 15204 93255 15352
rect 93505 15204 93545 15352
rect 93615 15204 93655 15436
rect 93905 15204 93945 15604
rect 94015 15604 94196 15644
rect 94252 17536 94348 17576
rect 94252 15644 94292 17536
rect 94348 17527 94388 17536
rect 94444 15644 94484 18292
rect 94539 18332 94581 18341
rect 94732 18332 94772 18341
rect 94539 18292 94540 18332
rect 94580 18292 94581 18332
rect 94539 18283 94581 18292
rect 94636 18292 94732 18332
rect 94252 15604 94345 15644
rect 94015 15204 94055 15604
rect 94305 15204 94345 15604
rect 94415 15604 94484 15644
rect 94415 15204 94455 15604
rect 94540 15560 94580 18283
rect 94636 15644 94676 18292
rect 94732 18283 94772 18292
rect 94924 17837 94964 18460
rect 95116 18450 95156 18535
rect 95500 18500 95540 19048
rect 95596 19039 95636 19048
rect 96352 18920 96720 18929
rect 96392 18880 96434 18920
rect 96474 18880 96516 18920
rect 96556 18880 96598 18920
rect 96638 18880 96680 18920
rect 96352 18871 96720 18880
rect 95980 18584 96020 18593
rect 96940 18584 96980 18593
rect 96020 18544 96116 18584
rect 95980 18535 96020 18544
rect 95212 18341 95252 18426
rect 95500 18341 95540 18460
rect 96076 18500 96116 18544
rect 96980 18544 97076 18584
rect 96940 18535 96980 18544
rect 96268 18500 96308 18509
rect 96076 18460 96268 18500
rect 95211 18332 95253 18341
rect 95211 18292 95212 18332
rect 95252 18292 95253 18332
rect 95211 18283 95253 18292
rect 95499 18332 95541 18341
rect 95499 18292 95500 18332
rect 95540 18292 95541 18332
rect 95499 18283 95541 18292
rect 95692 18332 95732 18341
rect 95112 18164 95480 18173
rect 95152 18124 95194 18164
rect 95234 18124 95276 18164
rect 95316 18124 95358 18164
rect 95398 18124 95440 18164
rect 95112 18115 95480 18124
rect 95403 17996 95445 18005
rect 95403 17956 95404 17996
rect 95444 17956 95445 17996
rect 95403 17947 95445 17956
rect 94731 17828 94773 17837
rect 94731 17788 94732 17828
rect 94772 17788 94773 17828
rect 94731 17779 94773 17788
rect 94923 17828 94965 17837
rect 95020 17828 95060 17856
rect 94923 17788 94924 17828
rect 94964 17788 95020 17828
rect 94923 17779 94965 17788
rect 95020 17779 95060 17788
rect 94732 17744 94772 17779
rect 94732 17693 94772 17704
rect 95404 17744 95444 17947
rect 95404 17695 95444 17704
rect 94828 17576 94868 17585
rect 95212 17576 95252 17585
rect 94868 17536 95060 17576
rect 94828 17527 94868 17536
rect 95020 15644 95060 17536
rect 94636 15604 94855 15644
rect 95020 15604 95145 15644
rect 94540 15520 94745 15560
rect 94705 15204 94745 15520
rect 94815 15204 94855 15604
rect 95105 15204 95145 15604
rect 95212 15476 95252 17536
rect 95500 17576 95540 17585
rect 95500 15644 95540 17536
rect 95500 15604 95545 15644
rect 95212 15436 95255 15476
rect 95215 15204 95255 15436
rect 95505 15204 95545 15604
rect 95692 15392 95732 18292
rect 95884 18332 95924 18341
rect 95924 18292 96020 18332
rect 95884 18283 95924 18292
rect 95883 17996 95925 18005
rect 95883 17956 95884 17996
rect 95924 17956 95925 17996
rect 95883 17947 95925 17956
rect 95884 17828 95924 17947
rect 95884 17779 95924 17788
rect 95980 17660 96020 18292
rect 96076 18005 96116 18460
rect 96268 18451 96308 18460
rect 96460 18332 96500 18341
rect 96172 18292 96460 18332
rect 96075 17996 96117 18005
rect 96075 17956 96076 17996
rect 96116 17956 96117 17996
rect 96075 17947 96117 17956
rect 95615 15352 95732 15392
rect 95884 17620 96020 17660
rect 95884 15392 95924 17620
rect 96076 17576 96116 17585
rect 96076 15653 96116 17536
rect 96075 15644 96117 15653
rect 96075 15604 96076 15644
rect 96116 15604 96117 15644
rect 96075 15595 96117 15604
rect 96172 15569 96212 18292
rect 96460 18283 96500 18292
rect 96844 18332 96884 18341
rect 96884 18292 96980 18332
rect 96844 18283 96884 18292
rect 96363 17996 96405 18005
rect 96363 17956 96364 17996
rect 96404 17956 96405 17996
rect 96363 17947 96405 17956
rect 96651 17996 96693 18005
rect 96651 17956 96652 17996
rect 96692 17956 96693 17996
rect 96651 17947 96693 17956
rect 96364 17744 96404 17947
rect 96652 17828 96692 17947
rect 96652 17779 96692 17788
rect 96364 17695 96404 17704
rect 96940 17660 96980 18292
rect 97036 17837 97076 18544
rect 97132 18500 97172 19291
rect 97612 18584 97652 18593
rect 97612 18500 97652 18544
rect 97035 17828 97077 17837
rect 97035 17788 97036 17828
rect 97076 17788 97077 17828
rect 97035 17779 97077 17788
rect 97132 17744 97172 18460
rect 97420 18460 97652 18500
rect 97324 18332 97364 18341
rect 97420 18332 97460 18460
rect 97364 18292 97460 18332
rect 97516 18332 97556 18341
rect 97556 18292 97652 18332
rect 97324 17921 97364 18292
rect 97516 18283 97556 18292
rect 97323 17912 97365 17921
rect 97323 17872 97324 17912
rect 97364 17872 97365 17912
rect 97323 17863 97365 17872
rect 97420 17744 97460 17753
rect 97132 17704 97364 17744
rect 97324 17660 97364 17704
rect 97420 17660 97460 17704
rect 96940 17620 97076 17660
rect 97324 17620 97460 17660
rect 96268 17576 96308 17585
rect 96268 15644 96308 17536
rect 96844 17576 96884 17585
rect 96352 17408 96720 17417
rect 96392 17368 96434 17408
rect 96474 17368 96516 17408
rect 96556 17368 96598 17408
rect 96638 17368 96680 17408
rect 96352 17359 96720 17368
rect 96747 16400 96789 16409
rect 96747 16360 96748 16400
rect 96788 16360 96789 16400
rect 96747 16351 96789 16360
rect 96748 15644 96788 16351
rect 96268 15604 96345 15644
rect 96171 15560 96213 15569
rect 96171 15520 96172 15560
rect 96212 15520 96213 15560
rect 96171 15511 96213 15520
rect 96014 15392 96056 15401
rect 95884 15352 95945 15392
rect 95615 15204 95655 15352
rect 95905 15204 95945 15352
rect 96014 15352 96015 15392
rect 96055 15352 96056 15392
rect 96014 15343 96056 15352
rect 96015 15204 96055 15343
rect 96305 15204 96345 15604
rect 96705 15604 96788 15644
rect 96414 15560 96456 15569
rect 96414 15520 96415 15560
rect 96455 15520 96456 15560
rect 96414 15511 96456 15520
rect 96415 15204 96455 15511
rect 96705 15204 96745 15604
rect 96844 15476 96884 17536
rect 97036 15644 97076 17620
rect 97228 17576 97268 17585
rect 97036 15604 97145 15644
rect 96815 15436 96884 15476
rect 96815 15204 96855 15436
rect 97105 15204 97145 15604
rect 97228 15476 97268 17536
rect 97516 17576 97556 17585
rect 97516 16409 97556 17536
rect 97515 16400 97557 16409
rect 97515 16360 97516 16400
rect 97556 16360 97557 16400
rect 97515 16351 97557 16360
rect 97612 15728 97652 18292
rect 99112 18164 99480 18173
rect 99152 18124 99194 18164
rect 99234 18124 99276 18164
rect 99316 18124 99358 18164
rect 99398 18124 99440 18164
rect 99112 18115 99480 18124
rect 98475 17996 98517 18005
rect 98475 17956 98476 17996
rect 98516 17956 98517 17996
rect 98475 17947 98517 17956
rect 97900 17837 97940 17922
rect 98284 17912 98324 17921
rect 98092 17872 98284 17912
rect 97899 17828 97941 17837
rect 97899 17788 97900 17828
rect 97940 17788 97941 17828
rect 97899 17779 97941 17788
rect 97899 17660 97941 17669
rect 97899 17620 97900 17660
rect 97940 17620 97941 17660
rect 97899 17611 97941 17620
rect 97516 15688 97652 15728
rect 97708 17576 97748 17585
rect 97516 15644 97556 15688
rect 97708 15644 97748 17536
rect 97215 15436 97268 15476
rect 97505 15604 97556 15644
rect 97615 15604 97748 15644
rect 97900 15644 97940 17611
rect 98092 15644 98132 17872
rect 98284 17863 98324 17872
rect 98476 17828 98516 17947
rect 98476 17779 98516 17788
rect 98667 17744 98709 17753
rect 98667 17704 98668 17744
rect 98708 17704 98709 17744
rect 98667 17695 98709 17704
rect 98668 17610 98708 17695
rect 98763 17660 98805 17669
rect 98763 17620 98764 17660
rect 98804 17620 98805 17660
rect 98763 17611 98805 17620
rect 98764 17526 98804 17611
rect 97900 15604 97945 15644
rect 97215 15204 97255 15436
rect 97505 15204 97545 15604
rect 97615 15204 97655 15604
rect 97905 15204 97945 15604
rect 98015 15604 98132 15644
rect 98015 15204 98055 15604
rect 98414 15476 98456 15485
rect 98414 15436 98415 15476
rect 98455 15436 98456 15476
rect 98414 15427 98456 15436
rect 98304 15392 98346 15401
rect 98304 15352 98305 15392
rect 98345 15352 98346 15392
rect 98304 15343 98346 15352
rect 98305 15204 98345 15343
rect 98415 15204 98455 15427
rect 98955 15392 98997 15401
rect 98955 15352 98956 15392
rect 98996 15352 98997 15392
rect 98955 15343 98997 15352
rect 71883 14972 71925 14981
rect 71883 14932 71884 14972
rect 71924 14932 71925 14972
rect 71883 14923 71925 14932
rect 98956 11528 98996 15343
rect 98860 11488 98996 11528
rect 72305 9857 72345 10080
rect 72304 9848 72346 9857
rect 72304 9808 72305 9848
rect 72345 9808 72346 9848
rect 72304 9799 72346 9808
rect 72415 9773 72455 10080
rect 72414 9764 72456 9773
rect 72705 9764 72745 10080
rect 72414 9724 72415 9764
rect 72455 9724 72456 9764
rect 72414 9715 72456 9724
rect 72652 9724 72745 9764
rect 72815 9764 72855 10080
rect 72815 9724 72884 9764
rect 72652 9353 72692 9724
rect 72844 9605 72884 9724
rect 73105 9680 73145 10080
rect 73215 9941 73255 10080
rect 73214 9932 73256 9941
rect 73214 9892 73215 9932
rect 73255 9892 73256 9932
rect 73214 9883 73256 9892
rect 73505 9848 73545 10080
rect 73324 9808 73545 9848
rect 73227 9764 73269 9773
rect 73227 9724 73228 9764
rect 73268 9724 73269 9764
rect 73227 9715 73269 9724
rect 73105 9640 73172 9680
rect 72843 9596 72885 9605
rect 72843 9556 72844 9596
rect 72884 9556 72885 9596
rect 72843 9547 72885 9556
rect 73132 9521 73172 9640
rect 73131 9512 73173 9521
rect 73131 9472 73132 9512
rect 73172 9472 73173 9512
rect 73131 9463 73173 9472
rect 72651 9344 72693 9353
rect 72651 9304 72652 9344
rect 72692 9304 72693 9344
rect 72651 9295 72693 9304
rect 73228 9269 73268 9715
rect 73324 9689 73364 9808
rect 73323 9680 73365 9689
rect 73615 9680 73655 10080
rect 73905 9941 73945 10080
rect 73904 9932 73946 9941
rect 73904 9892 73905 9932
rect 73945 9892 73946 9932
rect 73904 9883 73946 9892
rect 74015 9764 74055 10080
rect 73323 9640 73324 9680
rect 73364 9640 73365 9680
rect 73323 9631 73365 9640
rect 73612 9640 73655 9680
rect 73708 9724 74055 9764
rect 73612 9437 73652 9640
rect 73611 9428 73653 9437
rect 73611 9388 73612 9428
rect 73652 9388 73653 9428
rect 73611 9379 73653 9388
rect 73227 9260 73269 9269
rect 73227 9220 73228 9260
rect 73268 9220 73269 9260
rect 73227 9211 73269 9220
rect 73323 8840 73365 8849
rect 73323 8800 73324 8840
rect 73364 8800 73365 8840
rect 73323 8791 73365 8800
rect 71787 7244 71829 7253
rect 71787 7204 71788 7244
rect 71828 7204 71829 7244
rect 71787 7195 71829 7204
rect 73324 7244 73364 8791
rect 73420 7412 73460 7421
rect 73708 7412 73748 9724
rect 74305 9680 74345 10080
rect 73460 7372 73748 7412
rect 73804 9640 74345 9680
rect 73804 7412 73844 9640
rect 74415 9596 74455 10080
rect 74571 9764 74613 9773
rect 74571 9724 74572 9764
rect 74612 9724 74613 9764
rect 74571 9715 74613 9724
rect 74380 9556 74455 9596
rect 74380 9185 74420 9556
rect 74379 9176 74421 9185
rect 74379 9136 74380 9176
rect 74420 9136 74421 9176
rect 74379 9127 74421 9136
rect 74187 7580 74229 7589
rect 74187 7540 74188 7580
rect 74228 7540 74229 7580
rect 74187 7531 74229 7540
rect 73420 7363 73460 7372
rect 73804 7363 73844 7372
rect 73612 7244 73652 7253
rect 73324 7204 73612 7244
rect 73324 7160 73364 7204
rect 73612 7195 73652 7204
rect 73324 7111 73364 7120
rect 74091 7076 74133 7085
rect 74091 7036 74092 7076
rect 74132 7036 74133 7076
rect 74091 7027 74133 7036
rect 74092 6992 74132 7027
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 8352 6824 8720 6833
rect 8392 6784 8434 6824
rect 8474 6784 8516 6824
rect 8556 6784 8598 6824
rect 8638 6784 8680 6824
rect 8352 6775 8720 6784
rect 12352 6824 12720 6833
rect 12392 6784 12434 6824
rect 12474 6784 12516 6824
rect 12556 6784 12598 6824
rect 12638 6784 12680 6824
rect 12352 6775 12720 6784
rect 16352 6824 16720 6833
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16352 6775 16720 6784
rect 20352 6824 20720 6833
rect 20392 6784 20434 6824
rect 20474 6784 20516 6824
rect 20556 6784 20598 6824
rect 20638 6784 20680 6824
rect 20352 6775 20720 6784
rect 24352 6824 24720 6833
rect 24392 6784 24434 6824
rect 24474 6784 24516 6824
rect 24556 6784 24598 6824
rect 24638 6784 24680 6824
rect 24352 6775 24720 6784
rect 28352 6824 28720 6833
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28352 6775 28720 6784
rect 32352 6824 32720 6833
rect 32392 6784 32434 6824
rect 32474 6784 32516 6824
rect 32556 6784 32598 6824
rect 32638 6784 32680 6824
rect 32352 6775 32720 6784
rect 36352 6824 36720 6833
rect 36392 6784 36434 6824
rect 36474 6784 36516 6824
rect 36556 6784 36598 6824
rect 36638 6784 36680 6824
rect 36352 6775 36720 6784
rect 40352 6824 40720 6833
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40352 6775 40720 6784
rect 44352 6824 44720 6833
rect 44392 6784 44434 6824
rect 44474 6784 44516 6824
rect 44556 6784 44598 6824
rect 44638 6784 44680 6824
rect 44352 6775 44720 6784
rect 48352 6824 48720 6833
rect 48392 6784 48434 6824
rect 48474 6784 48516 6824
rect 48556 6784 48598 6824
rect 48638 6784 48680 6824
rect 48352 6775 48720 6784
rect 52352 6824 52720 6833
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52352 6775 52720 6784
rect 56352 6824 56720 6833
rect 56392 6784 56434 6824
rect 56474 6784 56516 6824
rect 56556 6784 56598 6824
rect 56638 6784 56680 6824
rect 56352 6775 56720 6784
rect 60352 6824 60720 6833
rect 60392 6784 60434 6824
rect 60474 6784 60516 6824
rect 60556 6784 60598 6824
rect 60638 6784 60680 6824
rect 60352 6775 60720 6784
rect 64352 6824 64720 6833
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64352 6775 64720 6784
rect 68352 6824 68720 6833
rect 68392 6784 68434 6824
rect 68474 6784 68516 6824
rect 68556 6784 68598 6824
rect 68638 6784 68680 6824
rect 68352 6775 68720 6784
rect 72352 6824 72720 6833
rect 72392 6784 72434 6824
rect 72474 6784 72516 6824
rect 72556 6784 72598 6824
rect 72638 6784 72680 6824
rect 72352 6775 72720 6784
rect 74092 6488 74132 6952
rect 74188 6656 74228 7531
rect 74283 7328 74325 7337
rect 74283 7288 74284 7328
rect 74324 7288 74325 7328
rect 74283 7279 74325 7288
rect 74475 7328 74517 7337
rect 74475 7288 74476 7328
rect 74516 7288 74517 7328
rect 74475 7279 74517 7288
rect 74284 7244 74324 7279
rect 74284 7193 74324 7204
rect 74476 7194 74516 7279
rect 74572 7076 74612 9715
rect 74705 9680 74745 10080
rect 74815 9848 74855 10080
rect 74955 9848 74997 9857
rect 74815 9808 74900 9848
rect 74668 9640 74745 9680
rect 74668 7505 74708 9640
rect 74763 7748 74805 7757
rect 74763 7708 74764 7748
rect 74804 7708 74805 7748
rect 74763 7699 74805 7708
rect 74667 7496 74709 7505
rect 74667 7456 74668 7496
rect 74708 7456 74709 7496
rect 74667 7447 74709 7456
rect 74668 7253 74708 7338
rect 74667 7244 74709 7253
rect 74667 7204 74668 7244
rect 74708 7204 74709 7244
rect 74667 7195 74709 7204
rect 74572 7036 74708 7076
rect 74379 6824 74421 6833
rect 74379 6784 74380 6824
rect 74420 6784 74421 6824
rect 74379 6775 74421 6784
rect 74188 6607 74228 6616
rect 74092 6439 74132 6448
rect 1556 6364 1748 6404
rect 74380 6404 74420 6775
rect 1516 6355 1556 6364
rect 1612 5984 1652 6364
rect 74380 6355 74420 6364
rect 74571 6404 74613 6413
rect 74571 6364 74572 6404
rect 74612 6364 74613 6404
rect 74571 6355 74613 6364
rect 74572 6236 74612 6355
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 7112 6068 7480 6077
rect 7152 6028 7194 6068
rect 7234 6028 7276 6068
rect 7316 6028 7358 6068
rect 7398 6028 7440 6068
rect 7112 6019 7480 6028
rect 11112 6068 11480 6077
rect 11152 6028 11194 6068
rect 11234 6028 11276 6068
rect 11316 6028 11358 6068
rect 11398 6028 11440 6068
rect 11112 6019 11480 6028
rect 15112 6068 15480 6077
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15112 6019 15480 6028
rect 19112 6068 19480 6077
rect 19152 6028 19194 6068
rect 19234 6028 19276 6068
rect 19316 6028 19358 6068
rect 19398 6028 19440 6068
rect 19112 6019 19480 6028
rect 23112 6068 23480 6077
rect 23152 6028 23194 6068
rect 23234 6028 23276 6068
rect 23316 6028 23358 6068
rect 23398 6028 23440 6068
rect 23112 6019 23480 6028
rect 27112 6068 27480 6077
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27112 6019 27480 6028
rect 31112 6068 31480 6077
rect 31152 6028 31194 6068
rect 31234 6028 31276 6068
rect 31316 6028 31358 6068
rect 31398 6028 31440 6068
rect 31112 6019 31480 6028
rect 35112 6068 35480 6077
rect 35152 6028 35194 6068
rect 35234 6028 35276 6068
rect 35316 6028 35358 6068
rect 35398 6028 35440 6068
rect 35112 6019 35480 6028
rect 39112 6068 39480 6077
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39112 6019 39480 6028
rect 43112 6068 43480 6077
rect 43152 6028 43194 6068
rect 43234 6028 43276 6068
rect 43316 6028 43358 6068
rect 43398 6028 43440 6068
rect 43112 6019 43480 6028
rect 47112 6068 47480 6077
rect 47152 6028 47194 6068
rect 47234 6028 47276 6068
rect 47316 6028 47358 6068
rect 47398 6028 47440 6068
rect 47112 6019 47480 6028
rect 51112 6068 51480 6077
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51112 6019 51480 6028
rect 55112 6068 55480 6077
rect 55152 6028 55194 6068
rect 55234 6028 55276 6068
rect 55316 6028 55358 6068
rect 55398 6028 55440 6068
rect 55112 6019 55480 6028
rect 59112 6068 59480 6077
rect 59152 6028 59194 6068
rect 59234 6028 59276 6068
rect 59316 6028 59358 6068
rect 59398 6028 59440 6068
rect 59112 6019 59480 6028
rect 63112 6068 63480 6077
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63112 6019 63480 6028
rect 67112 6068 67480 6077
rect 67152 6028 67194 6068
rect 67234 6028 67276 6068
rect 67316 6028 67358 6068
rect 67398 6028 67440 6068
rect 67112 6019 67480 6028
rect 71112 6068 71480 6077
rect 71152 6028 71194 6068
rect 71234 6028 71276 6068
rect 71316 6028 71358 6068
rect 71398 6028 71440 6068
rect 71112 6019 71480 6028
rect 1612 5944 2036 5984
rect 843 5816 885 5825
rect 843 5776 844 5816
rect 884 5776 885 5816
rect 843 5767 885 5776
rect 844 5732 884 5767
rect 844 5681 884 5692
rect 1612 5732 1652 5944
rect 1612 5683 1652 5692
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5480 692 5599
rect 652 5431 692 5440
rect 843 5480 885 5489
rect 843 5440 844 5480
rect 884 5440 885 5480
rect 843 5431 885 5440
rect 1419 5480 1461 5489
rect 1419 5440 1420 5480
rect 1460 5440 1461 5480
rect 1419 5431 1461 5440
rect 844 4892 884 5431
rect 1420 5346 1460 5431
rect 844 4843 884 4852
rect 1420 4892 1460 4901
rect 1708 4892 1748 5944
rect 1803 5816 1845 5825
rect 1803 5776 1804 5816
rect 1844 5776 1845 5816
rect 1803 5767 1845 5776
rect 1804 5682 1844 5767
rect 1996 5732 2036 5944
rect 74572 5732 74612 6196
rect 74668 5984 74708 7036
rect 74764 6740 74804 7699
rect 74860 7589 74900 9808
rect 74955 9808 74956 9848
rect 74996 9808 74997 9848
rect 74955 9799 74997 9808
rect 74859 7580 74901 7589
rect 74859 7540 74860 7580
rect 74900 7540 74901 7580
rect 74859 7531 74901 7540
rect 74859 6992 74901 7001
rect 74859 6952 74860 6992
rect 74900 6952 74901 6992
rect 74859 6943 74901 6952
rect 74860 6858 74900 6943
rect 74764 6700 74900 6740
rect 74764 6413 74804 6498
rect 74763 6404 74805 6413
rect 74763 6364 74764 6404
rect 74804 6364 74805 6404
rect 74763 6355 74805 6364
rect 74860 6320 74900 6700
rect 74956 6656 74996 9799
rect 75105 9764 75145 10080
rect 75215 9857 75255 10080
rect 75214 9848 75256 9857
rect 75214 9808 75215 9848
rect 75255 9808 75256 9848
rect 75214 9799 75256 9808
rect 75505 9773 75545 10080
rect 75052 9724 75145 9764
rect 75504 9764 75546 9773
rect 75504 9724 75505 9764
rect 75545 9724 75546 9764
rect 75052 7757 75092 9724
rect 75504 9715 75546 9724
rect 75615 9680 75655 10080
rect 75905 9680 75945 10080
rect 76015 9680 76055 10080
rect 76305 9680 76345 10080
rect 76415 9680 76455 10080
rect 76705 9764 76745 10080
rect 75615 9640 75668 9680
rect 75905 9640 75956 9680
rect 75628 8168 75668 9640
rect 75532 8128 75668 8168
rect 75051 7748 75093 7757
rect 75051 7708 75052 7748
rect 75092 7708 75093 7748
rect 75051 7699 75093 7708
rect 75112 7580 75480 7589
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75112 7531 75480 7540
rect 75243 7412 75285 7421
rect 75243 7372 75244 7412
rect 75284 7372 75285 7412
rect 75243 7363 75285 7372
rect 75147 7328 75189 7337
rect 75147 7288 75148 7328
rect 75188 7288 75189 7328
rect 75147 7279 75189 7288
rect 75052 7244 75092 7253
rect 75052 7085 75092 7204
rect 75051 7076 75093 7085
rect 75051 7036 75052 7076
rect 75092 7036 75093 7076
rect 75051 7027 75093 7036
rect 75148 6917 75188 7279
rect 75244 7278 75284 7363
rect 75436 7253 75476 7338
rect 75435 7244 75477 7253
rect 75340 7204 75436 7244
rect 75476 7204 75477 7244
rect 75147 6908 75189 6917
rect 75147 6868 75148 6908
rect 75188 6868 75189 6908
rect 75147 6859 75189 6868
rect 75340 6665 75380 7204
rect 75435 7195 75477 7204
rect 75435 6992 75477 7001
rect 75435 6952 75436 6992
rect 75476 6952 75477 6992
rect 75435 6943 75477 6952
rect 75244 6656 75284 6665
rect 74956 6616 75244 6656
rect 75244 6607 75284 6616
rect 75339 6656 75381 6665
rect 75339 6616 75340 6656
rect 75380 6616 75381 6656
rect 75339 6607 75381 6616
rect 75436 6497 75476 6943
rect 75532 6656 75572 8128
rect 75916 7412 75956 9640
rect 75916 7363 75956 7372
rect 76012 9640 76055 9680
rect 76300 9640 76345 9680
rect 76396 9640 76455 9680
rect 76588 9724 76745 9764
rect 75724 7253 75764 7338
rect 75723 7244 75765 7253
rect 75723 7204 75724 7244
rect 75764 7204 75765 7244
rect 75723 7195 75765 7204
rect 75723 6992 75765 7001
rect 75723 6952 75724 6992
rect 75764 6952 75765 6992
rect 75723 6943 75765 6952
rect 75532 6607 75572 6616
rect 75145 6475 75185 6496
rect 75435 6488 75477 6497
rect 75435 6448 75436 6488
rect 75476 6448 75477 6488
rect 75435 6439 75477 6448
rect 75724 6488 75764 6943
rect 75820 6656 75860 6665
rect 76012 6656 76052 9640
rect 76300 7412 76340 9640
rect 76300 7363 76340 7372
rect 75860 6616 76052 6656
rect 76108 7244 76148 7253
rect 75820 6607 75860 6616
rect 76108 6497 76148 7204
rect 76396 6992 76436 9640
rect 76588 7421 76628 9724
rect 76815 9680 76855 10080
rect 76780 9640 76855 9680
rect 77105 9680 77145 10080
rect 77215 9764 77255 10080
rect 77215 9724 77300 9764
rect 77105 9640 77204 9680
rect 76587 7412 76629 7421
rect 76587 7372 76588 7412
rect 76628 7372 76629 7412
rect 76587 7363 76629 7372
rect 76588 7085 76628 7170
rect 76683 7160 76725 7169
rect 76683 7120 76684 7160
rect 76724 7120 76725 7160
rect 76683 7111 76725 7120
rect 76587 7076 76629 7085
rect 76587 7036 76588 7076
rect 76628 7036 76629 7076
rect 76587 7027 76629 7036
rect 76684 7026 76724 7111
rect 76204 6952 76436 6992
rect 76204 6656 76244 6952
rect 76352 6824 76720 6833
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76352 6775 76720 6784
rect 76396 6656 76436 6665
rect 76204 6616 76396 6656
rect 76396 6607 76436 6616
rect 76587 6656 76629 6665
rect 76587 6616 76588 6656
rect 76628 6616 76629 6656
rect 76587 6607 76629 6616
rect 76780 6656 76820 9640
rect 77067 7412 77109 7421
rect 77067 7372 77068 7412
rect 77108 7372 77109 7412
rect 77067 7363 77109 7372
rect 77068 7278 77108 7363
rect 76875 7244 76917 7253
rect 76875 7204 76876 7244
rect 76916 7204 76917 7244
rect 76875 7195 76917 7204
rect 76876 7110 76916 7195
rect 76780 6607 76820 6616
rect 77164 6656 77204 9640
rect 77260 7337 77300 9724
rect 77505 9680 77545 10080
rect 77452 9640 77545 9680
rect 77615 9680 77655 10080
rect 77905 9680 77945 10080
rect 78015 9680 78055 10080
rect 78305 9680 78345 10080
rect 77615 9640 77684 9680
rect 77905 9640 77972 9680
rect 78015 9640 78068 9680
rect 77452 7421 77492 9640
rect 77644 7421 77684 9640
rect 77451 7412 77493 7421
rect 77451 7372 77452 7412
rect 77492 7372 77493 7412
rect 77451 7363 77493 7372
rect 77643 7412 77685 7421
rect 77643 7372 77644 7412
rect 77684 7372 77685 7412
rect 77643 7363 77685 7372
rect 77259 7328 77301 7337
rect 77259 7288 77260 7328
rect 77300 7288 77301 7328
rect 77259 7279 77301 7288
rect 77452 7244 77492 7253
rect 77259 7160 77301 7169
rect 77259 7120 77260 7160
rect 77300 7120 77301 7160
rect 77259 7111 77301 7120
rect 77260 6992 77300 7111
rect 77452 7001 77492 7204
rect 77643 7244 77685 7253
rect 77643 7204 77644 7244
rect 77684 7204 77685 7244
rect 77643 7195 77685 7204
rect 77835 7244 77877 7253
rect 77835 7204 77836 7244
rect 77876 7204 77877 7244
rect 77835 7195 77877 7204
rect 77644 7085 77684 7195
rect 77836 7110 77876 7195
rect 77643 7076 77685 7085
rect 77643 7036 77644 7076
rect 77684 7036 77685 7076
rect 77643 7027 77685 7036
rect 77260 6943 77300 6952
rect 77451 6992 77493 7001
rect 77451 6952 77452 6992
rect 77492 6952 77493 6992
rect 77451 6943 77493 6952
rect 77644 6992 77684 7027
rect 77164 6607 77204 6616
rect 75724 6439 75764 6448
rect 76107 6488 76149 6497
rect 76107 6448 76108 6488
rect 76148 6448 76149 6488
rect 76107 6439 76149 6448
rect 76299 6488 76341 6497
rect 76299 6448 76300 6488
rect 76340 6448 76341 6488
rect 76588 6488 76628 6607
rect 76684 6488 76724 6497
rect 76588 6448 76684 6488
rect 76299 6439 76341 6448
rect 75145 6413 75185 6435
rect 75145 6404 75189 6413
rect 75145 6364 75148 6404
rect 75188 6364 75189 6404
rect 75147 6355 75189 6364
rect 75436 6354 75476 6439
rect 76300 6354 76340 6439
rect 76684 6404 76724 6448
rect 76972 6404 77012 6413
rect 76684 6364 76972 6404
rect 77644 6404 77684 6952
rect 77932 6656 77972 9640
rect 78028 7589 78068 9640
rect 78220 9640 78345 9680
rect 78415 9680 78455 10080
rect 78705 9680 78745 10080
rect 78815 9764 78855 10080
rect 79105 9764 79145 10080
rect 78415 9640 78548 9680
rect 78027 7580 78069 7589
rect 78027 7540 78028 7580
rect 78068 7540 78069 7580
rect 78027 7531 78069 7540
rect 78027 7412 78069 7421
rect 78027 7372 78028 7412
rect 78068 7372 78069 7412
rect 78027 7363 78069 7372
rect 78028 7278 78068 7363
rect 78124 7160 78164 7169
rect 78124 7001 78164 7120
rect 78123 6992 78165 7001
rect 78123 6952 78124 6992
rect 78164 6952 78165 6992
rect 78123 6943 78165 6952
rect 78220 6656 78260 9640
rect 78315 7580 78357 7589
rect 78315 7540 78316 7580
rect 78356 7540 78357 7580
rect 78315 7531 78357 7540
rect 78316 7412 78356 7531
rect 78316 7363 78356 7372
rect 78412 7160 78452 7171
rect 78412 7085 78452 7120
rect 78411 7076 78453 7085
rect 78411 7036 78412 7076
rect 78452 7036 78453 7076
rect 78411 7027 78453 7036
rect 78316 6656 78356 6665
rect 78220 6616 78316 6656
rect 77932 6607 77972 6616
rect 78316 6607 78356 6616
rect 77740 6413 77780 6498
rect 78124 6413 78164 6498
rect 77739 6404 77781 6413
rect 77644 6364 77740 6404
rect 77780 6364 77781 6404
rect 74956 6320 74996 6329
rect 74860 6280 74956 6320
rect 74956 6271 74996 6280
rect 75112 6068 75480 6077
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75112 6019 75480 6028
rect 74668 5944 74996 5984
rect 74956 5900 74996 5944
rect 76684 5909 76724 5994
rect 75340 5900 75380 5909
rect 74956 5860 75340 5900
rect 75340 5851 75380 5860
rect 76683 5900 76725 5909
rect 76683 5860 76684 5900
rect 76724 5860 76725 5900
rect 76683 5851 76725 5860
rect 75148 5732 75188 5741
rect 74572 5692 75148 5732
rect 1996 5683 2036 5692
rect 75148 5683 75188 5692
rect 76492 5732 76532 5741
rect 76780 5732 76820 6364
rect 76972 6355 77012 6364
rect 77739 6355 77781 6364
rect 78123 6404 78165 6413
rect 78123 6364 78124 6404
rect 78164 6364 78165 6404
rect 78123 6355 78165 6364
rect 76532 5692 76820 5732
rect 76492 5683 76532 5692
rect 78124 5648 78164 6355
rect 78508 6320 78548 9640
rect 78700 9640 78745 9680
rect 78796 9724 78855 9764
rect 78903 9724 79145 9764
rect 78700 7244 78740 9640
rect 78796 7412 78836 9724
rect 78903 9680 78943 9724
rect 79215 9680 79255 10080
rect 79505 9857 79545 10080
rect 79504 9848 79546 9857
rect 79504 9808 79505 9848
rect 79545 9808 79546 9848
rect 79504 9799 79546 9808
rect 79615 9680 79655 10080
rect 79755 9848 79797 9857
rect 79755 9808 79756 9848
rect 79796 9808 79797 9848
rect 79755 9799 79797 9808
rect 78796 7363 78836 7372
rect 78892 9640 78943 9680
rect 78988 9640 79255 9680
rect 79564 9640 79655 9680
rect 78700 7204 78836 7244
rect 78700 7149 78740 7158
rect 78700 7085 78740 7109
rect 78699 7076 78741 7085
rect 78699 7036 78700 7076
rect 78740 7036 78741 7076
rect 78699 7027 78741 7036
rect 78700 7014 78740 7027
rect 78603 6404 78645 6413
rect 78603 6364 78604 6404
rect 78644 6364 78645 6404
rect 78603 6355 78645 6364
rect 78316 6280 78548 6320
rect 78316 5900 78356 6280
rect 78316 5851 78356 5860
rect 78604 5732 78644 6355
rect 78796 5900 78836 7204
rect 78892 6992 78932 9640
rect 78988 7412 79028 9640
rect 79112 7580 79480 7589
rect 79152 7540 79194 7580
rect 79234 7540 79276 7580
rect 79316 7540 79358 7580
rect 79398 7540 79440 7580
rect 79112 7531 79480 7540
rect 79180 7412 79220 7421
rect 78988 7372 79180 7412
rect 79180 7363 79220 7372
rect 79468 7412 79508 7421
rect 79564 7412 79604 9640
rect 79508 7372 79604 7412
rect 79468 7363 79508 7372
rect 79659 7328 79701 7337
rect 79659 7288 79660 7328
rect 79700 7288 79701 7328
rect 79659 7279 79701 7288
rect 79083 7244 79125 7253
rect 79083 7204 79084 7244
rect 79124 7204 79125 7244
rect 79083 7195 79125 7204
rect 79660 7244 79700 7279
rect 79084 7160 79124 7195
rect 79660 7193 79700 7204
rect 79084 7109 79124 7120
rect 79372 7160 79412 7169
rect 79372 7001 79412 7120
rect 79371 6992 79413 7001
rect 78892 6952 79124 6992
rect 79084 6656 79124 6952
rect 79371 6952 79372 6992
rect 79412 6952 79413 6992
rect 79371 6943 79413 6952
rect 79084 6607 79124 6616
rect 79756 6572 79796 9799
rect 79905 9680 79945 10080
rect 79852 9640 79945 9680
rect 79852 7412 79892 9640
rect 80015 9596 80055 10080
rect 80305 9773 80345 10080
rect 80304 9764 80346 9773
rect 80304 9724 80305 9764
rect 80345 9724 80346 9764
rect 80304 9715 80346 9724
rect 80415 9680 80455 10080
rect 80705 9680 80745 10080
rect 80815 9764 80855 10080
rect 80815 9724 80948 9764
rect 80415 9640 80468 9680
rect 80705 9640 80852 9680
rect 79852 7363 79892 7372
rect 79948 9556 80055 9596
rect 79948 6656 79988 9556
rect 80043 7328 80085 7337
rect 80043 7288 80044 7328
rect 80084 7288 80180 7328
rect 80043 7279 80085 7288
rect 80044 7194 80084 7279
rect 80044 6656 80084 6665
rect 79948 6616 80044 6656
rect 80044 6607 80084 6616
rect 79372 6532 79796 6572
rect 78892 6413 78932 6498
rect 78891 6404 78933 6413
rect 78891 6364 78892 6404
rect 78932 6364 78933 6404
rect 78891 6355 78933 6364
rect 79372 6320 79412 6532
rect 79948 6488 79988 6497
rect 80140 6488 80180 7288
rect 80236 7253 80276 7338
rect 80235 7244 80277 7253
rect 80235 7204 80236 7244
rect 80276 7204 80277 7244
rect 80235 7195 80277 7204
rect 80428 7076 80468 9640
rect 80716 7328 80756 7339
rect 80716 7253 80756 7288
rect 79988 6448 80180 6488
rect 80236 7036 80468 7076
rect 80524 7244 80564 7253
rect 79564 6404 79604 6413
rect 79948 6404 79988 6448
rect 79604 6364 79988 6404
rect 79564 6355 79604 6364
rect 79372 6271 79412 6280
rect 79112 6068 79480 6077
rect 79152 6028 79194 6068
rect 79234 6028 79276 6068
rect 79316 6028 79358 6068
rect 79398 6028 79440 6068
rect 79112 6019 79480 6028
rect 78796 5851 78836 5860
rect 78604 5683 78644 5692
rect 79948 5732 79988 6364
rect 80139 5900 80181 5909
rect 80139 5860 80140 5900
rect 80180 5860 80181 5900
rect 80236 5900 80276 7036
rect 80524 7001 80564 7204
rect 80715 7244 80757 7253
rect 80715 7204 80716 7244
rect 80756 7204 80757 7244
rect 80715 7195 80757 7204
rect 80523 6992 80565 7001
rect 80523 6952 80524 6992
rect 80564 6952 80565 6992
rect 80523 6943 80565 6952
rect 80352 6824 80720 6833
rect 80392 6784 80434 6824
rect 80474 6784 80516 6824
rect 80556 6784 80598 6824
rect 80638 6784 80680 6824
rect 80352 6775 80720 6784
rect 80620 6656 80660 6665
rect 80812 6656 80852 9640
rect 80908 7421 80948 9724
rect 81105 9680 81145 10080
rect 81215 9680 81255 10080
rect 81505 9680 81545 10080
rect 81004 9640 81145 9680
rect 81196 9640 81255 9680
rect 81484 9640 81545 9680
rect 81615 9680 81655 10080
rect 81905 9932 81945 10080
rect 81880 9892 81945 9932
rect 81615 9640 81716 9680
rect 80907 7412 80949 7421
rect 80907 7372 80908 7412
rect 80948 7372 80949 7412
rect 80907 7363 80949 7372
rect 80907 7160 80949 7169
rect 80907 7120 80908 7160
rect 80948 7120 80949 7160
rect 80907 7111 80949 7120
rect 80660 6616 80852 6656
rect 80908 6992 80948 7111
rect 80620 6607 80660 6616
rect 80428 6404 80468 6413
rect 80332 5900 80372 5909
rect 80236 5860 80332 5900
rect 80139 5851 80181 5860
rect 80332 5851 80372 5860
rect 80140 5766 80180 5851
rect 79948 5683 79988 5692
rect 78220 5648 78260 5657
rect 78124 5608 78220 5648
rect 78220 5599 78260 5608
rect 80428 5648 80468 6364
rect 80908 6404 80948 6952
rect 81004 6656 81044 9640
rect 81099 7244 81141 7253
rect 81099 7204 81100 7244
rect 81140 7204 81141 7244
rect 81099 7195 81141 7204
rect 81100 7110 81140 7195
rect 81100 6656 81140 6665
rect 81004 6616 81100 6656
rect 81100 6607 81140 6616
rect 80908 5648 80948 6364
rect 81196 5900 81236 9640
rect 81484 7412 81524 9640
rect 81579 8252 81621 8261
rect 81579 8212 81580 8252
rect 81620 8212 81621 8252
rect 81579 8203 81621 8212
rect 81484 7363 81524 7372
rect 81292 7244 81332 7255
rect 81292 7169 81332 7204
rect 81291 7160 81333 7169
rect 81291 7120 81292 7160
rect 81332 7120 81333 7160
rect 81291 7111 81333 7120
rect 81292 6488 81332 7111
rect 81484 6656 81524 6665
rect 81580 6656 81620 8203
rect 81676 7589 81716 9640
rect 81880 9512 81920 9892
rect 82015 9848 82055 10080
rect 82305 9857 82345 10080
rect 82304 9848 82346 9857
rect 82015 9808 82100 9848
rect 82060 9680 82100 9808
rect 82304 9808 82305 9848
rect 82345 9808 82346 9848
rect 82304 9799 82346 9808
rect 82415 9680 82455 10080
rect 82539 9848 82581 9857
rect 82539 9808 82540 9848
rect 82580 9808 82581 9848
rect 82539 9799 82581 9808
rect 82060 9640 82292 9680
rect 81880 9472 82004 9512
rect 81964 7748 82004 9472
rect 82252 8261 82292 9640
rect 82348 9640 82455 9680
rect 82251 8252 82293 8261
rect 82251 8212 82252 8252
rect 82292 8212 82293 8252
rect 82251 8203 82293 8212
rect 81880 7708 82004 7748
rect 81675 7580 81717 7589
rect 81675 7540 81676 7580
rect 81716 7540 81717 7580
rect 81675 7531 81717 7540
rect 81675 7412 81717 7421
rect 81675 7372 81676 7412
rect 81716 7372 81717 7412
rect 81675 7363 81717 7372
rect 81676 7278 81716 7363
rect 81880 7328 81920 7708
rect 81963 7580 82005 7589
rect 81963 7540 81964 7580
rect 82004 7540 82005 7580
rect 81963 7531 82005 7540
rect 81868 7288 81920 7328
rect 81772 7160 81812 7169
rect 81772 7001 81812 7120
rect 81771 6992 81813 7001
rect 81771 6952 81772 6992
rect 81812 6952 81813 6992
rect 81771 6943 81813 6952
rect 81524 6616 81620 6656
rect 81868 6656 81908 7288
rect 81964 7244 82004 7531
rect 82348 7412 82388 9640
rect 82348 7363 82388 7372
rect 82251 7244 82293 7253
rect 81964 7204 82100 7244
rect 82060 7160 82100 7204
rect 82251 7204 82252 7244
rect 82292 7204 82293 7244
rect 82251 7195 82293 7204
rect 81964 7149 82004 7158
rect 82060 7111 82100 7120
rect 82252 7160 82292 7195
rect 82540 7160 82580 9799
rect 82705 9680 82745 10080
rect 82815 9680 82855 10080
rect 83105 9680 83145 10080
rect 83215 9680 83255 10080
rect 83505 9680 83545 10080
rect 83615 9773 83655 10080
rect 83614 9764 83656 9773
rect 83614 9724 83615 9764
rect 83655 9724 83656 9764
rect 83614 9715 83656 9724
rect 82705 9640 82772 9680
rect 82815 9640 82964 9680
rect 83105 9640 83156 9680
rect 82252 7109 82292 7120
rect 82348 7120 82580 7160
rect 82635 7160 82677 7169
rect 82635 7120 82636 7160
rect 82676 7120 82677 7160
rect 81964 7085 82004 7109
rect 81960 7076 82004 7085
rect 81960 7036 81961 7076
rect 82001 7036 82004 7076
rect 81960 7027 82002 7036
rect 81961 7017 82001 7027
rect 81484 6607 81524 6616
rect 81868 6607 81908 6616
rect 82252 6656 82292 6665
rect 82348 6656 82388 7120
rect 82635 7111 82677 7120
rect 82636 6992 82676 7111
rect 82292 6616 82388 6656
rect 82540 6952 82636 6992
rect 82252 6607 82292 6616
rect 81388 6488 81428 6497
rect 81292 6448 81388 6488
rect 81428 6448 81716 6488
rect 81388 6439 81428 6448
rect 81676 6404 81716 6448
rect 82540 6413 82580 6952
rect 82636 6943 82676 6952
rect 82732 6824 82772 9640
rect 82827 7244 82869 7253
rect 82827 7204 82828 7244
rect 82868 7204 82869 7244
rect 82924 7244 82964 9640
rect 83116 7925 83156 9640
rect 83212 9640 83255 9680
rect 83500 9640 83545 9680
rect 83905 9680 83945 10080
rect 84015 9764 84055 10080
rect 84015 9724 84116 9764
rect 83905 9640 84020 9680
rect 83115 7916 83157 7925
rect 83115 7876 83116 7916
rect 83156 7876 83157 7916
rect 83115 7867 83157 7876
rect 83212 7748 83252 9640
rect 83020 7708 83252 7748
rect 83500 7748 83540 9640
rect 83500 7708 83636 7748
rect 83020 7412 83060 7708
rect 83112 7580 83480 7589
rect 83152 7540 83194 7580
rect 83234 7540 83276 7580
rect 83316 7540 83358 7580
rect 83398 7540 83440 7580
rect 83112 7531 83480 7540
rect 83404 7412 83444 7421
rect 83020 7372 83404 7412
rect 83404 7363 83444 7372
rect 83020 7244 83060 7253
rect 82924 7204 83020 7244
rect 82827 7195 82869 7204
rect 83020 7195 83060 7204
rect 82828 7110 82868 7195
rect 83115 7160 83157 7169
rect 83115 7120 83116 7160
rect 83156 7120 83157 7160
rect 83115 7111 83157 7120
rect 83307 7160 83349 7169
rect 83307 7120 83308 7160
rect 83348 7120 83349 7160
rect 83307 7111 83349 7120
rect 82923 7076 82965 7085
rect 82923 7036 82924 7076
rect 82964 7036 82965 7076
rect 82923 7027 82965 7036
rect 82636 6784 82772 6824
rect 81676 6355 81716 6364
rect 82059 6404 82101 6413
rect 82059 6364 82060 6404
rect 82100 6364 82101 6404
rect 82059 6355 82101 6364
rect 82539 6404 82581 6413
rect 82539 6364 82540 6404
rect 82580 6364 82581 6404
rect 82539 6355 82581 6364
rect 82060 6270 82100 6355
rect 81196 5851 81236 5860
rect 82636 5900 82676 6784
rect 82924 6656 82964 7027
rect 83116 7026 83156 7111
rect 83308 7026 83348 7111
rect 82924 6607 82964 6616
rect 83404 6656 83444 6665
rect 83596 6656 83636 7708
rect 83883 7412 83925 7421
rect 83883 7372 83884 7412
rect 83924 7372 83925 7412
rect 83883 7363 83925 7372
rect 83884 7278 83924 7363
rect 83787 7160 83829 7169
rect 83787 7120 83788 7160
rect 83828 7120 83829 7160
rect 83787 7111 83829 7120
rect 83788 7026 83828 7111
rect 83444 6616 83636 6656
rect 83884 6656 83924 6665
rect 83980 6656 84020 9640
rect 84076 7421 84116 9724
rect 84305 9680 84345 10080
rect 84415 9764 84455 10080
rect 84415 9724 84500 9764
rect 84305 9640 84404 9680
rect 84075 7412 84117 7421
rect 84075 7372 84076 7412
rect 84116 7372 84117 7412
rect 84075 7363 84117 7372
rect 84267 7244 84309 7253
rect 84267 7204 84268 7244
rect 84308 7204 84309 7244
rect 84267 7195 84309 7204
rect 84075 7160 84117 7169
rect 84075 7120 84076 7160
rect 84116 7120 84117 7160
rect 84075 7111 84117 7120
rect 83924 6616 84020 6656
rect 84076 6992 84116 7111
rect 84268 7110 84308 7195
rect 84364 6992 84404 9640
rect 84460 7589 84500 9724
rect 84705 9680 84745 10080
rect 84815 9764 84855 10080
rect 84815 9724 84884 9764
rect 84705 9640 84788 9680
rect 84459 7580 84501 7589
rect 84459 7540 84460 7580
rect 84500 7540 84501 7580
rect 84459 7531 84501 7540
rect 84651 7412 84693 7421
rect 84651 7372 84652 7412
rect 84692 7372 84693 7412
rect 84651 7363 84693 7372
rect 84652 7278 84692 7363
rect 84556 7160 84596 7169
rect 84556 7001 84596 7120
rect 83404 6607 83444 6616
rect 83884 6607 83924 6616
rect 82731 6404 82773 6413
rect 82731 6364 82732 6404
rect 82772 6364 82773 6404
rect 82731 6355 82773 6364
rect 83211 6404 83253 6413
rect 83211 6364 83212 6404
rect 83252 6364 83253 6404
rect 83211 6355 83253 6364
rect 83691 6404 83733 6413
rect 83691 6364 83692 6404
rect 83732 6364 83733 6404
rect 84076 6404 84116 6952
rect 84268 6952 84404 6992
rect 84555 6992 84597 7001
rect 84555 6952 84556 6992
rect 84596 6952 84597 6992
rect 84268 6656 84308 6952
rect 84555 6943 84597 6952
rect 84748 6908 84788 9640
rect 84844 7421 84884 9724
rect 85105 9680 85145 10080
rect 85036 9640 85145 9680
rect 85215 9680 85255 10080
rect 85505 9680 85545 10080
rect 85615 9680 85655 10080
rect 85905 9680 85945 10080
rect 86015 9680 86055 10080
rect 85215 9640 85268 9680
rect 85505 9640 85556 9680
rect 84843 7412 84885 7421
rect 84843 7372 84844 7412
rect 84884 7372 84885 7412
rect 84843 7363 84885 7372
rect 85036 7412 85076 9640
rect 85228 7412 85268 9640
rect 85036 7363 85076 7372
rect 85132 7372 85268 7412
rect 84844 7244 84884 7255
rect 84844 7169 84884 7204
rect 84843 7160 84885 7169
rect 84843 7120 84844 7160
rect 84884 7120 84885 7160
rect 84843 7111 84885 7120
rect 84748 6868 84884 6908
rect 84352 6824 84720 6833
rect 84392 6784 84434 6824
rect 84474 6784 84516 6824
rect 84556 6784 84598 6824
rect 84638 6784 84680 6824
rect 84352 6775 84720 6784
rect 84364 6656 84404 6665
rect 84268 6616 84364 6656
rect 84364 6607 84404 6616
rect 84748 6656 84788 6665
rect 84844 6656 84884 6868
rect 84788 6616 84884 6656
rect 84940 6656 84980 6665
rect 85132 6656 85172 7372
rect 85227 7244 85269 7253
rect 85227 7204 85228 7244
rect 85268 7204 85269 7244
rect 85227 7195 85269 7204
rect 85228 7110 85268 7195
rect 85420 6992 85460 7001
rect 84980 6616 85172 6656
rect 85324 6952 85420 6992
rect 84748 6607 84788 6616
rect 84940 6607 84980 6616
rect 85036 6488 85076 6499
rect 85036 6413 85076 6448
rect 84171 6404 84213 6413
rect 84076 6364 84172 6404
rect 84212 6364 84213 6404
rect 83691 6355 83733 6364
rect 84171 6355 84213 6364
rect 84555 6404 84597 6413
rect 84555 6364 84556 6404
rect 84596 6364 84597 6404
rect 84555 6355 84597 6364
rect 85035 6404 85077 6413
rect 85035 6364 85036 6404
rect 85076 6364 85077 6404
rect 85035 6355 85077 6364
rect 85227 6404 85269 6413
rect 85324 6404 85364 6952
rect 85420 6943 85460 6952
rect 85420 6656 85460 6665
rect 85516 6656 85556 9640
rect 85612 9640 85655 9680
rect 85804 9640 85945 9680
rect 85996 9640 86055 9680
rect 86305 9680 86345 10080
rect 86415 9764 86455 10080
rect 86415 9724 86516 9764
rect 86305 9640 86420 9680
rect 85612 8849 85652 9640
rect 85611 8840 85653 8849
rect 85611 8800 85612 8840
rect 85652 8800 85653 8840
rect 85611 8791 85653 8800
rect 85707 7580 85749 7589
rect 85707 7540 85708 7580
rect 85748 7540 85749 7580
rect 85707 7531 85749 7540
rect 85708 7412 85748 7531
rect 85708 7363 85748 7372
rect 85612 7169 85652 7254
rect 85611 7160 85653 7169
rect 85611 7120 85612 7160
rect 85652 7120 85653 7160
rect 85611 7111 85653 7120
rect 85460 6616 85556 6656
rect 85804 6656 85844 9640
rect 85996 7001 86036 9640
rect 86187 8168 86229 8177
rect 86187 8128 86188 8168
rect 86228 8128 86229 8168
rect 86187 8119 86229 8128
rect 86091 7244 86133 7253
rect 86091 7204 86092 7244
rect 86132 7204 86133 7244
rect 86091 7195 86133 7204
rect 86092 7110 86132 7195
rect 85995 6992 86037 7001
rect 85995 6952 85996 6992
rect 86036 6952 86037 6992
rect 85995 6943 86037 6952
rect 85420 6607 85460 6616
rect 85804 6607 85844 6616
rect 86091 6572 86133 6581
rect 86091 6532 86092 6572
rect 86132 6532 86133 6572
rect 86091 6523 86133 6532
rect 86092 6413 86132 6523
rect 85227 6364 85228 6404
rect 85268 6364 85364 6404
rect 85227 6355 85269 6364
rect 82636 5851 82676 5860
rect 82444 5732 82484 5741
rect 82732 5732 82772 6355
rect 83212 6270 83252 6355
rect 83112 6068 83480 6077
rect 83152 6028 83194 6068
rect 83234 6028 83276 6068
rect 83316 6028 83358 6068
rect 83398 6028 83440 6068
rect 83112 6019 83480 6028
rect 83595 5900 83637 5909
rect 83595 5860 83596 5900
rect 83636 5860 83637 5900
rect 83595 5851 83637 5860
rect 83596 5766 83636 5851
rect 82484 5692 82772 5732
rect 82444 5683 82484 5692
rect 81100 5648 81140 5657
rect 80468 5608 81100 5648
rect 80428 5599 80468 5608
rect 81100 5599 81140 5608
rect 83500 5648 83540 5657
rect 83692 5648 83732 6355
rect 84172 6270 84212 6355
rect 84556 6270 84596 6355
rect 85228 6270 85268 6355
rect 83540 5608 83732 5648
rect 85324 5648 85364 6364
rect 85611 6404 85653 6413
rect 85611 6364 85612 6404
rect 85652 6364 85653 6404
rect 85611 6355 85653 6364
rect 86091 6404 86133 6413
rect 86091 6364 86092 6404
rect 86132 6364 86133 6404
rect 86091 6355 86133 6364
rect 85612 6270 85652 6355
rect 86092 6270 86132 6355
rect 85515 5900 85557 5909
rect 85515 5860 85516 5900
rect 85556 5860 85557 5900
rect 85515 5851 85557 5860
rect 85516 5766 85556 5851
rect 86188 5825 86228 8119
rect 86283 7328 86325 7337
rect 86283 7288 86284 7328
rect 86324 7288 86325 7328
rect 86283 7279 86325 7288
rect 86284 7194 86324 7279
rect 86284 6656 86324 6665
rect 86380 6656 86420 9640
rect 86476 7589 86516 9724
rect 86705 9680 86745 10080
rect 86815 9764 86855 10080
rect 86815 9724 86900 9764
rect 86705 9640 86804 9680
rect 86475 7580 86517 7589
rect 86475 7540 86476 7580
rect 86516 7540 86517 7580
rect 86475 7531 86517 7540
rect 86667 7412 86709 7421
rect 86667 7372 86668 7412
rect 86708 7372 86709 7412
rect 86667 7363 86709 7372
rect 86476 7328 86516 7339
rect 86476 7253 86516 7288
rect 86475 7244 86517 7253
rect 86475 7204 86476 7244
rect 86516 7204 86517 7244
rect 86475 7195 86517 7204
rect 86668 7244 86708 7363
rect 86668 6917 86708 7204
rect 86667 6908 86709 6917
rect 86667 6868 86668 6908
rect 86708 6868 86709 6908
rect 86667 6859 86709 6868
rect 86324 6616 86420 6656
rect 86284 6607 86324 6616
rect 86764 5900 86804 9640
rect 86860 7328 86900 9724
rect 87105 9680 87145 10080
rect 87215 9773 87255 10080
rect 87214 9764 87256 9773
rect 87214 9724 87215 9764
rect 87255 9724 87256 9764
rect 87214 9715 87256 9724
rect 86956 9640 87145 9680
rect 87505 9680 87545 10080
rect 87615 9680 87655 10080
rect 87723 9764 87765 9773
rect 87723 9724 87724 9764
rect 87764 9724 87765 9764
rect 87723 9715 87765 9724
rect 87505 9640 87572 9680
rect 87615 9640 87668 9680
rect 86956 7412 86996 9640
rect 87112 7580 87480 7589
rect 87152 7540 87194 7580
rect 87234 7540 87276 7580
rect 87316 7540 87358 7580
rect 87398 7540 87440 7580
rect 87112 7531 87480 7540
rect 87147 7412 87189 7421
rect 86956 7372 87092 7412
rect 86860 7288 86996 7328
rect 86956 7169 86996 7288
rect 86860 7160 86900 7169
rect 86860 6581 86900 7120
rect 86955 7160 86997 7169
rect 86955 7120 86956 7160
rect 86996 7120 86997 7160
rect 86955 7111 86997 7120
rect 86955 6992 86997 7001
rect 86955 6952 86956 6992
rect 86996 6952 86997 6992
rect 86955 6943 86997 6952
rect 86956 6858 86996 6943
rect 87052 6656 87092 7372
rect 87147 7372 87148 7412
rect 87188 7372 87189 7412
rect 87147 7363 87189 7372
rect 87148 7278 87188 7363
rect 87243 7328 87285 7337
rect 87532 7328 87572 9640
rect 87243 7288 87244 7328
rect 87284 7288 87285 7328
rect 87243 7279 87285 7288
rect 87340 7288 87572 7328
rect 87244 7160 87284 7279
rect 87244 7085 87284 7120
rect 87243 7076 87285 7085
rect 87243 7036 87244 7076
rect 87284 7036 87285 7076
rect 87243 7027 87285 7036
rect 87052 6607 87092 6616
rect 86859 6572 86901 6581
rect 86859 6532 86860 6572
rect 86900 6532 86901 6572
rect 86859 6523 86901 6532
rect 86764 5851 86804 5860
rect 86860 6404 86900 6413
rect 87244 6404 87284 7027
rect 87340 6656 87380 7288
rect 87435 7160 87477 7169
rect 87435 7120 87436 7160
rect 87476 7120 87477 7160
rect 87435 7111 87477 7120
rect 87532 7160 87572 7171
rect 87436 7026 87476 7111
rect 87532 7085 87572 7120
rect 87531 7076 87573 7085
rect 87531 7036 87532 7076
rect 87572 7036 87573 7076
rect 87531 7027 87573 7036
rect 87532 6656 87572 6665
rect 87340 6616 87532 6656
rect 87532 6607 87572 6616
rect 87340 6404 87380 6413
rect 86900 6364 87340 6404
rect 86187 5816 86229 5825
rect 86187 5776 86188 5816
rect 86228 5776 86229 5816
rect 86187 5767 86229 5776
rect 86572 5732 86612 5741
rect 86860 5732 86900 6364
rect 87340 6355 87380 6364
rect 87112 6068 87480 6077
rect 87152 6028 87194 6068
rect 87234 6028 87276 6068
rect 87316 6028 87358 6068
rect 87398 6028 87440 6068
rect 87112 6019 87480 6028
rect 87628 5900 87668 9640
rect 87724 7412 87764 9715
rect 87905 9680 87945 10080
rect 88015 9680 88055 10080
rect 88305 9680 88345 10080
rect 88415 9680 88455 10080
rect 87905 9640 87956 9680
rect 87724 7363 87764 7372
rect 87820 7160 87860 7171
rect 87820 7085 87860 7120
rect 87819 7076 87861 7085
rect 87628 5851 87668 5860
rect 87724 7036 87820 7076
rect 87860 7036 87861 7076
rect 87724 6404 87764 7036
rect 87819 7027 87861 7036
rect 87916 6656 87956 9640
rect 88012 9640 88055 9680
rect 88204 9640 88345 9680
rect 88396 9640 88455 9680
rect 88705 9680 88745 10080
rect 88815 9764 88855 10080
rect 89105 9773 89145 10080
rect 89104 9764 89146 9773
rect 88815 9724 88916 9764
rect 88705 9640 88820 9680
rect 88012 7589 88052 9640
rect 88011 7580 88053 7589
rect 88011 7540 88012 7580
rect 88052 7540 88053 7580
rect 88011 7531 88053 7540
rect 88011 7244 88053 7253
rect 88011 7204 88012 7244
rect 88052 7204 88053 7244
rect 88011 7195 88053 7204
rect 88012 7085 88052 7195
rect 88204 7160 88244 9640
rect 88299 7244 88341 7253
rect 88299 7204 88300 7244
rect 88340 7204 88341 7244
rect 88299 7195 88341 7204
rect 88108 7120 88244 7160
rect 88011 7076 88053 7085
rect 88011 7036 88012 7076
rect 88052 7036 88053 7076
rect 88011 7027 88053 7036
rect 88108 6824 88148 7120
rect 88204 6992 88244 7001
rect 88300 6992 88340 7195
rect 88396 7001 88436 9640
rect 88780 7412 88820 9640
rect 88780 7363 88820 7372
rect 88587 7244 88629 7253
rect 88587 7204 88588 7244
rect 88628 7204 88629 7244
rect 88587 7195 88629 7204
rect 88588 7110 88628 7195
rect 88244 6952 88340 6992
rect 88395 6992 88437 7001
rect 88395 6952 88396 6992
rect 88436 6952 88437 6992
rect 88204 6943 88244 6952
rect 88395 6943 88437 6952
rect 88352 6824 88720 6833
rect 88108 6784 88244 6824
rect 88204 6656 88244 6784
rect 88392 6784 88434 6824
rect 88474 6784 88516 6824
rect 88556 6784 88598 6824
rect 88638 6784 88680 6824
rect 88352 6775 88720 6784
rect 88300 6656 88340 6665
rect 88204 6616 88300 6656
rect 87916 6607 87956 6616
rect 88300 6607 88340 6616
rect 88491 6656 88533 6665
rect 88876 6656 88916 9724
rect 89104 9724 89105 9764
rect 89145 9724 89146 9764
rect 89104 9715 89146 9724
rect 89215 9680 89255 10080
rect 89505 9680 89545 10080
rect 89615 9848 89655 10080
rect 89615 9808 89780 9848
rect 89215 9640 89300 9680
rect 89505 9640 89588 9680
rect 88971 7580 89013 7589
rect 88971 7540 88972 7580
rect 89012 7540 89013 7580
rect 88971 7531 89013 7540
rect 88972 7412 89012 7531
rect 88972 7363 89012 7372
rect 89067 7244 89109 7253
rect 89067 7204 89068 7244
rect 89108 7204 89109 7244
rect 89067 7195 89109 7204
rect 88491 6616 88492 6656
rect 88532 6616 88533 6656
rect 88491 6607 88533 6616
rect 88780 6616 88916 6656
rect 89068 7160 89108 7195
rect 88492 6522 88532 6607
rect 88107 6488 88149 6497
rect 88107 6448 88108 6488
rect 88148 6448 88149 6488
rect 88107 6439 88149 6448
rect 88587 6488 88629 6497
rect 88587 6448 88588 6488
rect 88628 6448 88629 6488
rect 88587 6439 88629 6448
rect 88780 6488 88820 6616
rect 88780 6439 88820 6448
rect 88875 6488 88917 6497
rect 89068 6488 89108 7120
rect 89260 6656 89300 9640
rect 89452 7244 89492 7255
rect 89452 7169 89492 7204
rect 89451 7160 89493 7169
rect 89451 7120 89452 7160
rect 89492 7120 89493 7160
rect 89451 7111 89493 7120
rect 89260 6607 89300 6616
rect 89164 6488 89204 6497
rect 88875 6448 88876 6488
rect 88916 6448 89164 6488
rect 88875 6439 88917 6448
rect 89164 6439 89204 6448
rect 86612 5692 86900 5732
rect 86572 5683 86612 5692
rect 85420 5648 85460 5657
rect 85324 5608 85420 5648
rect 83500 5599 83540 5608
rect 85420 5599 85460 5608
rect 87532 5648 87572 5657
rect 87724 5648 87764 6364
rect 88108 6404 88148 6439
rect 88108 6353 88148 6364
rect 88588 6354 88628 6439
rect 88876 5732 88916 6439
rect 89452 6320 89492 6329
rect 89548 6320 89588 9640
rect 89643 7412 89685 7421
rect 89643 7372 89644 7412
rect 89684 7372 89685 7412
rect 89643 7363 89685 7372
rect 89644 7278 89684 7363
rect 89643 6404 89685 6413
rect 89643 6364 89644 6404
rect 89684 6364 89685 6404
rect 89643 6355 89685 6364
rect 89492 6280 89588 6320
rect 89452 6271 89492 6280
rect 89644 6152 89684 6355
rect 89548 6112 89684 6152
rect 89067 5900 89109 5909
rect 89067 5860 89068 5900
rect 89108 5860 89109 5900
rect 89067 5851 89109 5860
rect 89068 5766 89108 5851
rect 88876 5683 88916 5692
rect 87572 5608 87764 5648
rect 89548 5648 89588 6112
rect 89644 5900 89684 5909
rect 89740 5900 89780 9808
rect 89905 9680 89945 10080
rect 89836 9640 89945 9680
rect 90015 9680 90055 10080
rect 90305 9680 90345 10080
rect 90415 9680 90455 10080
rect 90705 9680 90745 10080
rect 90015 9640 90068 9680
rect 89836 7421 89876 9640
rect 90028 7421 90068 9640
rect 90220 9640 90345 9680
rect 90412 9640 90455 9680
rect 90508 9640 90745 9680
rect 90815 9680 90855 10080
rect 91105 9680 91145 10080
rect 90815 9640 90932 9680
rect 89835 7412 89877 7421
rect 89835 7372 89836 7412
rect 89876 7372 89877 7412
rect 89835 7363 89877 7372
rect 90027 7412 90069 7421
rect 90027 7372 90028 7412
rect 90068 7372 90069 7412
rect 90027 7363 90069 7372
rect 90028 7244 90068 7253
rect 89835 7160 89877 7169
rect 89835 7120 89836 7160
rect 89876 7120 89877 7160
rect 89835 7111 89877 7120
rect 89836 6992 89876 7111
rect 90028 7085 90068 7204
rect 90027 7076 90069 7085
rect 90027 7036 90028 7076
rect 90068 7036 90069 7076
rect 90027 7027 90069 7036
rect 89836 6943 89876 6952
rect 89684 5860 89780 5900
rect 90220 5900 90260 9640
rect 90412 7412 90452 9640
rect 90412 7363 90452 7372
rect 90316 7160 90356 7169
rect 90316 6917 90356 7120
rect 90315 6908 90357 6917
rect 90315 6868 90316 6908
rect 90356 6868 90357 6908
rect 90315 6859 90357 6868
rect 90508 6656 90548 9640
rect 90892 7421 90932 9640
rect 90988 9640 91145 9680
rect 91215 9680 91255 10080
rect 91505 9857 91545 10080
rect 91504 9848 91546 9857
rect 91504 9808 91505 9848
rect 91545 9808 91546 9848
rect 91504 9799 91546 9808
rect 91615 9764 91655 10080
rect 91755 9848 91797 9857
rect 91755 9808 91756 9848
rect 91796 9808 91797 9848
rect 91755 9799 91797 9808
rect 91615 9724 91700 9764
rect 91215 9640 91604 9680
rect 90603 7412 90645 7421
rect 90603 7372 90604 7412
rect 90644 7372 90645 7412
rect 90603 7363 90645 7372
rect 90891 7412 90933 7421
rect 90891 7372 90892 7412
rect 90932 7372 90933 7412
rect 90988 7412 91028 9640
rect 91112 7580 91480 7589
rect 91152 7540 91194 7580
rect 91234 7540 91276 7580
rect 91316 7540 91358 7580
rect 91398 7540 91440 7580
rect 91112 7531 91480 7540
rect 91564 7412 91604 9640
rect 90988 7372 91124 7412
rect 90891 7363 90933 7372
rect 90604 7278 90644 7363
rect 90987 7244 91029 7253
rect 90987 7204 90988 7244
rect 91028 7204 91029 7244
rect 90987 7195 91029 7204
rect 90712 7160 90754 7169
rect 90712 7120 90713 7160
rect 90753 7120 90754 7160
rect 90712 7111 90754 7120
rect 90891 7160 90933 7169
rect 90891 7120 90892 7160
rect 90932 7120 90933 7160
rect 90891 7111 90933 7120
rect 90713 7026 90753 7111
rect 90604 6656 90644 6665
rect 90508 6616 90604 6656
rect 90604 6607 90644 6616
rect 90892 6413 90932 7111
rect 90988 7110 91028 7195
rect 91084 6656 91124 7372
rect 91276 7372 91604 7412
rect 91179 7328 91221 7337
rect 91179 7288 91180 7328
rect 91220 7288 91221 7328
rect 91179 7279 91221 7288
rect 91180 7194 91220 7279
rect 91084 6607 91124 6616
rect 91276 6656 91316 7372
rect 91372 7244 91412 7253
rect 91372 7085 91412 7204
rect 91563 7244 91605 7253
rect 91563 7204 91564 7244
rect 91604 7204 91605 7244
rect 91563 7195 91605 7204
rect 91371 7076 91413 7085
rect 91371 7036 91372 7076
rect 91412 7036 91413 7076
rect 91371 7027 91413 7036
rect 91564 6992 91604 7195
rect 91276 6607 91316 6616
rect 91468 6952 91564 6992
rect 91468 6572 91508 6952
rect 91564 6943 91604 6952
rect 91660 6572 91700 9724
rect 91756 7337 91796 9799
rect 91905 9680 91945 10080
rect 92015 9764 92055 10080
rect 92015 9724 92084 9764
rect 91905 9640 91988 9680
rect 91851 7412 91893 7421
rect 91851 7372 91852 7412
rect 91892 7372 91893 7412
rect 91851 7363 91893 7372
rect 91755 7328 91797 7337
rect 91755 7288 91756 7328
rect 91796 7288 91797 7328
rect 91755 7279 91797 7288
rect 91852 7278 91892 7363
rect 91755 7160 91797 7169
rect 91755 7120 91756 7160
rect 91796 7120 91797 7160
rect 91755 7111 91797 7120
rect 91756 7026 91796 7111
rect 91852 6656 91892 6665
rect 91948 6656 91988 9640
rect 91892 6616 91988 6656
rect 91852 6607 91892 6616
rect 91372 6532 91508 6572
rect 91564 6532 91700 6572
rect 92044 6572 92084 9724
rect 92305 9680 92345 10080
rect 92236 9640 92345 9680
rect 92415 9680 92455 10080
rect 92705 9773 92745 10080
rect 92704 9764 92746 9773
rect 92704 9724 92705 9764
rect 92745 9724 92746 9764
rect 92704 9715 92746 9724
rect 92815 9680 92855 10080
rect 93003 9848 93045 9857
rect 93003 9808 93004 9848
rect 93044 9808 93045 9848
rect 93003 9799 93045 9808
rect 92907 9764 92949 9773
rect 92907 9724 92908 9764
rect 92948 9724 92949 9764
rect 92907 9715 92949 9724
rect 92415 9640 92468 9680
rect 92139 7244 92181 7253
rect 92139 7204 92140 7244
rect 92180 7204 92181 7244
rect 92139 7195 92181 7204
rect 92140 7110 92180 7195
rect 92236 6656 92276 9640
rect 92428 7589 92468 9640
rect 92812 9640 92855 9680
rect 92427 7580 92469 7589
rect 92427 7540 92428 7580
rect 92468 7540 92469 7580
rect 92427 7531 92469 7540
rect 92331 7328 92373 7337
rect 92331 7288 92332 7328
rect 92372 7288 92373 7328
rect 92331 7279 92373 7288
rect 92524 7328 92564 7339
rect 92332 7194 92372 7279
rect 92524 7253 92564 7288
rect 92523 7244 92565 7253
rect 92523 7204 92524 7244
rect 92564 7204 92565 7244
rect 92523 7195 92565 7204
rect 92716 7244 92756 7253
rect 92716 7085 92756 7204
rect 92715 7076 92757 7085
rect 92715 7036 92716 7076
rect 92756 7036 92757 7076
rect 92715 7027 92757 7036
rect 92352 6824 92720 6833
rect 92392 6784 92434 6824
rect 92474 6784 92516 6824
rect 92556 6784 92598 6824
rect 92638 6784 92680 6824
rect 92352 6775 92720 6784
rect 92332 6656 92372 6665
rect 92620 6656 92660 6665
rect 92236 6616 92332 6656
rect 92332 6607 92372 6616
rect 92428 6616 92620 6656
rect 92044 6532 92276 6572
rect 91372 6488 91412 6532
rect 91372 6413 91412 6448
rect 90411 6404 90453 6413
rect 90411 6364 90412 6404
rect 90452 6364 90453 6404
rect 90411 6355 90453 6364
rect 90891 6404 90933 6413
rect 90891 6364 90892 6404
rect 90932 6364 90933 6404
rect 90891 6355 90933 6364
rect 91371 6404 91413 6413
rect 91371 6364 91372 6404
rect 91412 6364 91413 6404
rect 91371 6355 91413 6364
rect 89644 5851 89684 5860
rect 90220 5851 90260 5860
rect 90412 5732 90452 6355
rect 90892 6270 90932 6355
rect 91372 6324 91412 6355
rect 91112 6068 91480 6077
rect 91152 6028 91194 6068
rect 91234 6028 91276 6068
rect 91316 6028 91358 6068
rect 91398 6028 91440 6068
rect 91112 6019 91480 6028
rect 91564 5900 91604 6532
rect 92236 6488 92276 6532
rect 92428 6488 92468 6616
rect 92620 6607 92660 6616
rect 92236 6448 92468 6488
rect 92524 6488 92564 6499
rect 92524 6413 92564 6448
rect 91659 6404 91701 6413
rect 92139 6404 92181 6413
rect 91659 6364 91660 6404
rect 91700 6364 91796 6404
rect 91659 6355 91701 6364
rect 91660 6270 91700 6355
rect 91660 5900 91700 5909
rect 91564 5860 91660 5900
rect 91660 5851 91700 5860
rect 90412 5683 90452 5692
rect 87532 5599 87572 5608
rect 89548 5599 89588 5608
rect 91564 5648 91604 5657
rect 91756 5648 91796 6364
rect 92139 6364 92140 6404
rect 92180 6364 92181 6404
rect 92139 6355 92181 6364
rect 92523 6404 92565 6413
rect 92523 6364 92524 6404
rect 92564 6364 92565 6404
rect 92523 6355 92565 6364
rect 92140 6270 92180 6355
rect 92812 5900 92852 9640
rect 92908 7412 92948 9715
rect 92908 7363 92948 7372
rect 93004 6572 93044 9799
rect 93105 9680 93145 10080
rect 93215 9857 93255 10080
rect 93214 9848 93256 9857
rect 93214 9808 93215 9848
rect 93255 9808 93256 9848
rect 93214 9799 93256 9808
rect 93505 9680 93545 10080
rect 93615 9764 93655 10080
rect 93905 9848 93945 10080
rect 93772 9808 93945 9848
rect 93615 9724 93716 9764
rect 93105 9640 93236 9680
rect 93505 9640 93620 9680
rect 93099 7328 93141 7337
rect 93099 7288 93100 7328
rect 93140 7288 93141 7328
rect 93099 7279 93141 7288
rect 93100 7244 93140 7279
rect 93100 7193 93140 7204
rect 93196 6656 93236 9640
rect 93291 7580 93333 7589
rect 93291 7540 93292 7580
rect 93332 7540 93333 7580
rect 93291 7531 93333 7540
rect 93292 7412 93332 7531
rect 93292 7363 93332 7372
rect 93483 7412 93525 7421
rect 93483 7372 93484 7412
rect 93524 7372 93525 7412
rect 93483 7363 93525 7372
rect 93387 7328 93429 7337
rect 93387 7288 93388 7328
rect 93428 7288 93429 7328
rect 93387 7279 93429 7288
rect 93196 6607 93236 6616
rect 93388 7160 93428 7279
rect 93004 6532 93140 6572
rect 93004 6404 93044 6415
rect 93004 6329 93044 6364
rect 93003 6320 93045 6329
rect 93003 6280 93004 6320
rect 93044 6280 93045 6320
rect 93003 6271 93045 6280
rect 92812 5851 92852 5860
rect 91604 5608 91796 5648
rect 92908 5648 92948 5657
rect 93004 5648 93044 6271
rect 93100 5900 93140 6532
rect 93388 6404 93428 7120
rect 93388 6329 93428 6364
rect 93387 6320 93429 6329
rect 93387 6280 93388 6320
rect 93428 6280 93429 6320
rect 93387 6271 93429 6280
rect 93388 6240 93428 6271
rect 93196 5900 93236 5909
rect 93100 5860 93196 5900
rect 93484 5900 93524 7363
rect 93580 6656 93620 9640
rect 93676 7421 93716 9724
rect 93675 7412 93717 7421
rect 93675 7372 93676 7412
rect 93716 7372 93717 7412
rect 93675 7363 93717 7372
rect 93772 7169 93812 9808
rect 94015 9680 94055 10080
rect 94305 9680 94345 10080
rect 94015 9640 94100 9680
rect 93963 7328 94005 7337
rect 93963 7288 93964 7328
rect 94004 7288 94005 7328
rect 93963 7279 94005 7288
rect 93964 7194 94004 7279
rect 93676 7160 93716 7169
rect 93676 7085 93716 7120
rect 93771 7160 93813 7169
rect 93771 7120 93772 7160
rect 93812 7120 93813 7160
rect 93771 7111 93813 7120
rect 93675 7076 93717 7085
rect 93675 7036 93676 7076
rect 93716 7036 93717 7076
rect 93675 7027 93717 7036
rect 93676 6665 93716 7027
rect 93771 6992 93813 7001
rect 93771 6952 93772 6992
rect 93812 6952 93813 6992
rect 93771 6943 93813 6952
rect 93772 6858 93812 6943
rect 94060 6824 94100 9640
rect 94252 9640 94345 9680
rect 94415 9680 94455 10080
rect 94705 9680 94745 10080
rect 94815 9680 94855 10080
rect 95105 9680 95145 10080
rect 95215 9680 95255 10080
rect 95505 9680 95545 10080
rect 95615 9680 95655 10080
rect 95905 9932 95945 10080
rect 94415 9640 94484 9680
rect 94705 9640 94772 9680
rect 94815 9640 94868 9680
rect 94156 7253 94196 7338
rect 94155 7244 94197 7253
rect 94155 7204 94156 7244
rect 94196 7204 94197 7244
rect 94155 7195 94197 7204
rect 94155 7076 94197 7085
rect 94155 7036 94156 7076
rect 94196 7036 94197 7076
rect 94155 7027 94197 7036
rect 93964 6784 94100 6824
rect 93580 6607 93620 6616
rect 93675 6656 93717 6665
rect 93675 6616 93676 6656
rect 93716 6616 93717 6656
rect 93675 6607 93717 6616
rect 93868 6404 93908 6415
rect 93868 6329 93908 6364
rect 93867 6320 93909 6329
rect 93867 6280 93868 6320
rect 93908 6280 93909 6320
rect 93867 6271 93909 6280
rect 93580 5900 93620 5909
rect 93484 5860 93580 5900
rect 93196 5851 93236 5860
rect 93580 5851 93620 5860
rect 93964 5900 94004 6784
rect 94060 6656 94100 6665
rect 94156 6656 94196 7027
rect 94100 6616 94196 6656
rect 94252 6656 94292 9640
rect 94348 7244 94388 7253
rect 94348 6917 94388 7204
rect 94444 7001 94484 9640
rect 94732 7412 94772 9640
rect 94732 7363 94772 7372
rect 94731 7160 94773 7169
rect 94731 7120 94732 7160
rect 94772 7120 94773 7160
rect 94731 7111 94773 7120
rect 94443 6992 94485 7001
rect 94443 6952 94444 6992
rect 94484 6952 94485 6992
rect 94443 6943 94485 6952
rect 94540 6992 94580 7001
rect 94347 6908 94389 6917
rect 94347 6868 94348 6908
rect 94388 6868 94389 6908
rect 94347 6859 94389 6868
rect 94540 6665 94580 6952
rect 94060 6607 94100 6616
rect 94252 6607 94292 6616
rect 94539 6656 94581 6665
rect 94539 6616 94540 6656
rect 94580 6616 94581 6656
rect 94539 6607 94581 6616
rect 94732 6488 94772 7111
rect 94828 6656 94868 9640
rect 95020 9640 95145 9680
rect 95212 9640 95255 9680
rect 95404 9640 95545 9680
rect 95596 9640 95655 9680
rect 95788 9892 95945 9932
rect 95020 7412 95060 9640
rect 95212 7757 95252 9640
rect 95404 7841 95444 9640
rect 95403 7832 95445 7841
rect 95403 7792 95404 7832
rect 95444 7792 95445 7832
rect 95403 7783 95445 7792
rect 95211 7748 95253 7757
rect 95211 7708 95212 7748
rect 95252 7708 95253 7748
rect 95211 7699 95253 7708
rect 95112 7580 95480 7589
rect 95152 7540 95194 7580
rect 95234 7540 95276 7580
rect 95316 7540 95358 7580
rect 95398 7540 95440 7580
rect 95112 7531 95480 7540
rect 95116 7412 95156 7421
rect 95020 7372 95116 7412
rect 94924 7337 94964 7368
rect 95116 7363 95156 7372
rect 94923 7328 94965 7337
rect 94923 7288 94924 7328
rect 94964 7288 94965 7328
rect 94923 7279 94965 7288
rect 95307 7328 95349 7337
rect 95307 7288 95308 7328
rect 95348 7288 95349 7328
rect 95307 7279 95349 7288
rect 94828 6607 94868 6616
rect 94924 7244 94964 7279
rect 94732 6439 94772 6448
rect 94924 6413 94964 7204
rect 95308 7244 95348 7279
rect 95308 7193 95348 7204
rect 95307 6740 95349 6749
rect 95307 6700 95308 6740
rect 95348 6700 95349 6740
rect 95307 6691 95349 6700
rect 95308 6656 95348 6691
rect 95308 6605 95348 6616
rect 95596 6656 95636 9640
rect 95691 7244 95733 7253
rect 95691 7204 95692 7244
rect 95732 7204 95733 7244
rect 95691 7195 95733 7204
rect 95692 7110 95732 7195
rect 95596 6607 95636 6616
rect 95691 6656 95733 6665
rect 95691 6616 95692 6656
rect 95732 6616 95733 6656
rect 95691 6607 95733 6616
rect 95692 6488 95732 6607
rect 95692 6439 95732 6448
rect 94059 6404 94101 6413
rect 94059 6364 94060 6404
rect 94100 6364 94101 6404
rect 94059 6355 94101 6364
rect 94443 6404 94485 6413
rect 94443 6364 94444 6404
rect 94484 6364 94485 6404
rect 94443 6355 94485 6364
rect 94923 6404 94965 6413
rect 94923 6364 94924 6404
rect 94964 6364 94965 6404
rect 94923 6355 94965 6364
rect 95115 6404 95157 6413
rect 95115 6364 95116 6404
rect 95156 6364 95157 6404
rect 95115 6355 95157 6364
rect 93964 5851 94004 5860
rect 93291 5648 93333 5657
rect 92948 5608 93292 5648
rect 93332 5608 93333 5648
rect 91564 5599 91604 5608
rect 92908 5599 92948 5608
rect 93291 5599 93333 5608
rect 93675 5648 93717 5657
rect 93675 5608 93676 5648
rect 93716 5608 93717 5648
rect 93675 5599 93717 5608
rect 93868 5648 93908 5657
rect 94060 5648 94100 6355
rect 94444 6270 94484 6355
rect 95116 6270 95156 6355
rect 95112 6068 95480 6077
rect 95152 6028 95194 6068
rect 95234 6028 95276 6068
rect 95316 6028 95358 6068
rect 95398 6028 95440 6068
rect 95112 6019 95480 6028
rect 95692 5900 95732 5909
rect 95788 5900 95828 9892
rect 95883 9764 95925 9773
rect 95883 9724 95884 9764
rect 95924 9724 95925 9764
rect 95883 9715 95925 9724
rect 95884 7412 95924 9715
rect 96015 9680 96055 10080
rect 96305 9773 96345 10080
rect 96304 9764 96346 9773
rect 96304 9724 96305 9764
rect 96345 9724 96346 9764
rect 96304 9715 96346 9724
rect 95884 7363 95924 7372
rect 95980 9640 96055 9680
rect 96415 9680 96455 10080
rect 96705 9680 96745 10080
rect 96815 9764 96855 10080
rect 96815 9724 96884 9764
rect 96415 9640 96500 9680
rect 96705 9640 96788 9680
rect 95884 6497 95924 6582
rect 95883 6488 95925 6497
rect 95883 6448 95884 6488
rect 95924 6448 95925 6488
rect 95883 6439 95925 6448
rect 95980 6404 96020 9640
rect 96171 7748 96213 7757
rect 96171 7708 96172 7748
rect 96212 7708 96213 7748
rect 96171 7699 96213 7708
rect 96075 7244 96117 7253
rect 96075 7204 96076 7244
rect 96116 7204 96117 7244
rect 96075 7195 96117 7204
rect 96076 6992 96116 7195
rect 96076 6581 96116 6952
rect 96075 6572 96117 6581
rect 96075 6532 96076 6572
rect 96116 6532 96117 6572
rect 96075 6523 96117 6532
rect 95980 6364 96116 6404
rect 95883 6320 95925 6329
rect 95883 6280 95884 6320
rect 95924 6280 95925 6320
rect 95883 6271 95925 6280
rect 95732 5860 95828 5900
rect 95692 5851 95732 5860
rect 95500 5732 95540 5741
rect 95884 5732 95924 6271
rect 95979 6236 96021 6245
rect 95979 6196 95980 6236
rect 96020 6196 96021 6236
rect 95979 6187 96021 6196
rect 95980 6102 96020 6187
rect 95980 5900 96020 5909
rect 96076 5900 96116 6364
rect 96172 6245 96212 7699
rect 96460 7421 96500 9640
rect 96459 7412 96501 7421
rect 96459 7372 96460 7412
rect 96500 7372 96501 7412
rect 96459 7363 96501 7372
rect 96652 7328 96692 7339
rect 96652 7253 96692 7288
rect 96267 7244 96309 7253
rect 96267 7204 96268 7244
rect 96308 7204 96309 7244
rect 96267 7195 96309 7204
rect 96460 7244 96500 7253
rect 96268 7110 96308 7195
rect 96460 7085 96500 7204
rect 96651 7244 96693 7253
rect 96651 7204 96652 7244
rect 96692 7204 96693 7244
rect 96651 7195 96693 7204
rect 96459 7076 96501 7085
rect 96459 7036 96460 7076
rect 96500 7036 96501 7076
rect 96459 7027 96501 7036
rect 96748 6908 96788 9640
rect 96844 7589 96884 9724
rect 97105 9680 97145 10080
rect 97036 9640 97145 9680
rect 97215 9680 97255 10080
rect 97505 9680 97545 10080
rect 97215 9640 97364 9680
rect 96843 7580 96885 7589
rect 96843 7540 96844 7580
rect 96884 7540 96885 7580
rect 96843 7531 96885 7540
rect 96843 7412 96885 7421
rect 96843 7372 96844 7412
rect 96884 7372 96885 7412
rect 96843 7363 96885 7372
rect 96844 7278 96884 7363
rect 96939 7160 96981 7169
rect 96939 7120 96940 7160
rect 96980 7120 96981 7160
rect 96939 7111 96981 7120
rect 96748 6868 96884 6908
rect 96352 6824 96720 6833
rect 96392 6784 96434 6824
rect 96474 6784 96516 6824
rect 96556 6784 96598 6824
rect 96638 6784 96680 6824
rect 96352 6775 96720 6784
rect 96844 6740 96884 6868
rect 96748 6700 96884 6740
rect 96556 6656 96596 6665
rect 96748 6656 96788 6700
rect 96596 6616 96788 6656
rect 96556 6607 96596 6616
rect 96364 6404 96404 6415
rect 96364 6329 96404 6364
rect 96940 6404 96980 7111
rect 97036 6656 97076 9640
rect 97131 7580 97173 7589
rect 97131 7540 97132 7580
rect 97172 7540 97173 7580
rect 97131 7531 97173 7540
rect 97132 7412 97172 7531
rect 97132 7363 97172 7372
rect 97227 7160 97269 7169
rect 97227 7120 97228 7160
rect 97268 7120 97269 7160
rect 97227 7111 97269 7120
rect 97228 7026 97268 7111
rect 97132 6656 97172 6665
rect 97036 6616 97132 6656
rect 97324 6656 97364 9640
rect 97420 9640 97545 9680
rect 97615 9680 97655 10080
rect 97905 9680 97945 10080
rect 98015 9764 98055 10080
rect 98015 9724 98132 9764
rect 97615 9640 97748 9680
rect 97905 9640 98036 9680
rect 97420 7412 97460 9640
rect 97515 9512 97557 9521
rect 97515 9472 97516 9512
rect 97556 9472 97557 9512
rect 97515 9463 97557 9472
rect 97420 7363 97460 7372
rect 97420 6656 97460 6665
rect 97324 6616 97420 6656
rect 97132 6607 97172 6616
rect 97420 6607 97460 6616
rect 96940 6329 96980 6364
rect 97324 6488 97364 6497
rect 97324 6329 97364 6448
rect 96363 6320 96405 6329
rect 96363 6280 96364 6320
rect 96404 6280 96405 6320
rect 96363 6271 96405 6280
rect 96939 6320 96981 6329
rect 96939 6280 96940 6320
rect 96980 6280 96981 6320
rect 96939 6271 96981 6280
rect 97323 6320 97365 6329
rect 97323 6280 97324 6320
rect 97364 6280 97365 6320
rect 97323 6271 97365 6280
rect 96171 6236 96213 6245
rect 96171 6196 96172 6236
rect 96212 6196 96213 6236
rect 96171 6187 96213 6196
rect 96020 5860 96116 5900
rect 95980 5851 96020 5860
rect 96939 5816 96981 5825
rect 96939 5776 96940 5816
rect 96980 5776 96981 5816
rect 96939 5767 96981 5776
rect 95540 5692 95924 5732
rect 95500 5683 95540 5692
rect 93908 5608 94100 5648
rect 95884 5648 95924 5692
rect 93868 5599 93908 5608
rect 95884 5599 95924 5608
rect 93292 5514 93332 5599
rect 93676 5514 93716 5599
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 8352 5312 8720 5321
rect 8392 5272 8434 5312
rect 8474 5272 8516 5312
rect 8556 5272 8598 5312
rect 8638 5272 8680 5312
rect 8352 5263 8720 5272
rect 12352 5312 12720 5321
rect 12392 5272 12434 5312
rect 12474 5272 12516 5312
rect 12556 5272 12598 5312
rect 12638 5272 12680 5312
rect 12352 5263 12720 5272
rect 16352 5312 16720 5321
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16352 5263 16720 5272
rect 20352 5312 20720 5321
rect 20392 5272 20434 5312
rect 20474 5272 20516 5312
rect 20556 5272 20598 5312
rect 20638 5272 20680 5312
rect 20352 5263 20720 5272
rect 24352 5312 24720 5321
rect 24392 5272 24434 5312
rect 24474 5272 24516 5312
rect 24556 5272 24598 5312
rect 24638 5272 24680 5312
rect 24352 5263 24720 5272
rect 28352 5312 28720 5321
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28352 5263 28720 5272
rect 32352 5312 32720 5321
rect 32392 5272 32434 5312
rect 32474 5272 32516 5312
rect 32556 5272 32598 5312
rect 32638 5272 32680 5312
rect 32352 5263 32720 5272
rect 36352 5312 36720 5321
rect 36392 5272 36434 5312
rect 36474 5272 36516 5312
rect 36556 5272 36598 5312
rect 36638 5272 36680 5312
rect 36352 5263 36720 5272
rect 40352 5312 40720 5321
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40352 5263 40720 5272
rect 44352 5312 44720 5321
rect 44392 5272 44434 5312
rect 44474 5272 44516 5312
rect 44556 5272 44598 5312
rect 44638 5272 44680 5312
rect 44352 5263 44720 5272
rect 48352 5312 48720 5321
rect 48392 5272 48434 5312
rect 48474 5272 48516 5312
rect 48556 5272 48598 5312
rect 48638 5272 48680 5312
rect 48352 5263 48720 5272
rect 52352 5312 52720 5321
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52352 5263 52720 5272
rect 56352 5312 56720 5321
rect 56392 5272 56434 5312
rect 56474 5272 56516 5312
rect 56556 5272 56598 5312
rect 56638 5272 56680 5312
rect 56352 5263 56720 5272
rect 60352 5312 60720 5321
rect 60392 5272 60434 5312
rect 60474 5272 60516 5312
rect 60556 5272 60598 5312
rect 60638 5272 60680 5312
rect 60352 5263 60720 5272
rect 64352 5312 64720 5321
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64352 5263 64720 5272
rect 68352 5312 68720 5321
rect 68392 5272 68434 5312
rect 68474 5272 68516 5312
rect 68556 5272 68598 5312
rect 68638 5272 68680 5312
rect 68352 5263 68720 5272
rect 72352 5312 72720 5321
rect 72392 5272 72434 5312
rect 72474 5272 72516 5312
rect 72556 5272 72598 5312
rect 72638 5272 72680 5312
rect 72352 5263 72720 5272
rect 76352 5312 76720 5321
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76352 5263 76720 5272
rect 80352 5312 80720 5321
rect 80392 5272 80434 5312
rect 80474 5272 80516 5312
rect 80556 5272 80598 5312
rect 80638 5272 80680 5312
rect 80352 5263 80720 5272
rect 84352 5312 84720 5321
rect 84392 5272 84434 5312
rect 84474 5272 84516 5312
rect 84556 5272 84598 5312
rect 84638 5272 84680 5312
rect 84352 5263 84720 5272
rect 88352 5312 88720 5321
rect 88392 5272 88434 5312
rect 88474 5272 88516 5312
rect 88556 5272 88598 5312
rect 88638 5272 88680 5312
rect 88352 5263 88720 5272
rect 92352 5312 92720 5321
rect 92392 5272 92434 5312
rect 92474 5272 92516 5312
rect 92556 5272 92598 5312
rect 92638 5272 92680 5312
rect 92352 5263 92720 5272
rect 96352 5312 96720 5321
rect 96392 5272 96434 5312
rect 96474 5272 96516 5312
rect 96556 5272 96598 5312
rect 96638 5272 96680 5312
rect 96352 5263 96720 5272
rect 1804 4892 1844 4901
rect 2188 4892 2228 4901
rect 1460 4852 1804 4892
rect 1844 4852 2188 4892
rect 1420 4843 1460 4852
rect 1804 4843 1844 4852
rect 2188 4843 2228 4852
rect 96940 4892 96980 5767
rect 97516 4976 97556 9463
rect 97611 7244 97653 7253
rect 97611 7204 97612 7244
rect 97652 7204 97653 7244
rect 97611 7195 97653 7204
rect 97612 7110 97652 7195
rect 97708 6656 97748 9640
rect 97996 7412 98036 9640
rect 97996 7363 98036 7372
rect 97803 7244 97845 7253
rect 97803 7204 97804 7244
rect 97844 7204 97845 7244
rect 97803 7195 97845 7204
rect 97708 6607 97748 6616
rect 97804 6488 97844 7195
rect 97995 6656 98037 6665
rect 97995 6616 97996 6656
rect 98036 6616 98037 6656
rect 97995 6607 98037 6616
rect 98092 6656 98132 9724
rect 98305 9680 98345 10080
rect 98415 9764 98455 10080
rect 98415 9724 98804 9764
rect 98305 9640 98516 9680
rect 98476 7412 98516 9640
rect 98476 7363 98516 7372
rect 98187 7244 98229 7253
rect 98187 7204 98188 7244
rect 98228 7204 98229 7244
rect 98187 7195 98229 7204
rect 98668 7244 98708 7253
rect 98188 7110 98228 7195
rect 98092 6607 98132 6616
rect 97804 6439 97844 6448
rect 97996 6488 98036 6607
rect 97996 6439 98036 6448
rect 98668 5825 98708 7204
rect 98764 5900 98804 9724
rect 98764 5851 98804 5860
rect 98379 5816 98421 5825
rect 98379 5776 98380 5816
rect 98420 5776 98421 5816
rect 98379 5767 98421 5776
rect 98667 5816 98709 5825
rect 98667 5776 98668 5816
rect 98708 5776 98709 5816
rect 98667 5767 98709 5776
rect 98380 5648 98420 5767
rect 98380 5599 98420 5608
rect 98668 5648 98708 5767
rect 98668 5599 98708 5608
rect 98284 5480 98324 5489
rect 98860 5480 98900 11488
rect 99112 7580 99480 7589
rect 99152 7540 99194 7580
rect 99234 7540 99276 7580
rect 99316 7540 99358 7580
rect 99398 7540 99440 7580
rect 99112 7531 99480 7540
rect 99112 6068 99480 6077
rect 99152 6028 99194 6068
rect 99234 6028 99276 6068
rect 99316 6028 99358 6068
rect 99398 6028 99440 6068
rect 99112 6019 99480 6028
rect 98324 5440 98900 5480
rect 98284 5431 98324 5440
rect 96940 4843 96980 4852
rect 97132 4936 97556 4976
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 97132 4808 97172 4936
rect 97132 4759 97172 4768
rect 652 4674 692 4759
rect 747 4724 789 4733
rect 1228 4724 1268 4733
rect 747 4684 748 4724
rect 788 4684 789 4724
rect 747 4675 789 4684
rect 940 4684 1228 4724
rect 651 3968 693 3977
rect 651 3928 652 3968
rect 692 3928 693 3968
rect 651 3919 693 3928
rect 652 3834 692 3919
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 652 3078 692 3163
rect 748 2708 788 4675
rect 843 4220 885 4229
rect 843 4180 844 4220
rect 884 4180 885 4220
rect 843 4171 885 4180
rect 844 4086 884 4171
rect 844 3380 884 3389
rect 940 3380 980 4684
rect 1228 4675 1268 4684
rect 1612 4724 1652 4733
rect 1612 4229 1652 4684
rect 1995 4724 2037 4733
rect 1995 4684 1996 4724
rect 2036 4684 2037 4724
rect 1995 4675 2037 4684
rect 1996 4590 2036 4675
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 7112 4556 7480 4565
rect 7152 4516 7194 4556
rect 7234 4516 7276 4556
rect 7316 4516 7358 4556
rect 7398 4516 7440 4556
rect 7112 4507 7480 4516
rect 11112 4556 11480 4565
rect 11152 4516 11194 4556
rect 11234 4516 11276 4556
rect 11316 4516 11358 4556
rect 11398 4516 11440 4556
rect 11112 4507 11480 4516
rect 15112 4556 15480 4565
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15112 4507 15480 4516
rect 19112 4556 19480 4565
rect 19152 4516 19194 4556
rect 19234 4516 19276 4556
rect 19316 4516 19358 4556
rect 19398 4516 19440 4556
rect 19112 4507 19480 4516
rect 23112 4556 23480 4565
rect 23152 4516 23194 4556
rect 23234 4516 23276 4556
rect 23316 4516 23358 4556
rect 23398 4516 23440 4556
rect 23112 4507 23480 4516
rect 27112 4556 27480 4565
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27112 4507 27480 4516
rect 31112 4556 31480 4565
rect 31152 4516 31194 4556
rect 31234 4516 31276 4556
rect 31316 4516 31358 4556
rect 31398 4516 31440 4556
rect 31112 4507 31480 4516
rect 35112 4556 35480 4565
rect 35152 4516 35194 4556
rect 35234 4516 35276 4556
rect 35316 4516 35358 4556
rect 35398 4516 35440 4556
rect 35112 4507 35480 4516
rect 39112 4556 39480 4565
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39112 4507 39480 4516
rect 43112 4556 43480 4565
rect 43152 4516 43194 4556
rect 43234 4516 43276 4556
rect 43316 4516 43358 4556
rect 43398 4516 43440 4556
rect 43112 4507 43480 4516
rect 47112 4556 47480 4565
rect 47152 4516 47194 4556
rect 47234 4516 47276 4556
rect 47316 4516 47358 4556
rect 47398 4516 47440 4556
rect 47112 4507 47480 4516
rect 51112 4556 51480 4565
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51112 4507 51480 4516
rect 55112 4556 55480 4565
rect 55152 4516 55194 4556
rect 55234 4516 55276 4556
rect 55316 4516 55358 4556
rect 55398 4516 55440 4556
rect 55112 4507 55480 4516
rect 59112 4556 59480 4565
rect 59152 4516 59194 4556
rect 59234 4516 59276 4556
rect 59316 4516 59358 4556
rect 59398 4516 59440 4556
rect 59112 4507 59480 4516
rect 63112 4556 63480 4565
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63112 4507 63480 4516
rect 67112 4556 67480 4565
rect 67152 4516 67194 4556
rect 67234 4516 67276 4556
rect 67316 4516 67358 4556
rect 67398 4516 67440 4556
rect 67112 4507 67480 4516
rect 71112 4556 71480 4565
rect 71152 4516 71194 4556
rect 71234 4516 71276 4556
rect 71316 4516 71358 4556
rect 71398 4516 71440 4556
rect 71112 4507 71480 4516
rect 75112 4556 75480 4565
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75112 4507 75480 4516
rect 79112 4556 79480 4565
rect 79152 4516 79194 4556
rect 79234 4516 79276 4556
rect 79316 4516 79358 4556
rect 79398 4516 79440 4556
rect 79112 4507 79480 4516
rect 83112 4556 83480 4565
rect 83152 4516 83194 4556
rect 83234 4516 83276 4556
rect 83316 4516 83358 4556
rect 83398 4516 83440 4556
rect 83112 4507 83480 4516
rect 87112 4556 87480 4565
rect 87152 4516 87194 4556
rect 87234 4516 87276 4556
rect 87316 4516 87358 4556
rect 87398 4516 87440 4556
rect 87112 4507 87480 4516
rect 91112 4556 91480 4565
rect 91152 4516 91194 4556
rect 91234 4516 91276 4556
rect 91316 4516 91358 4556
rect 91398 4516 91440 4556
rect 91112 4507 91480 4516
rect 95112 4556 95480 4565
rect 95152 4516 95194 4556
rect 95234 4516 95276 4556
rect 95316 4516 95358 4556
rect 95398 4516 95440 4556
rect 95112 4507 95480 4516
rect 99112 4556 99480 4565
rect 99152 4516 99194 4556
rect 99234 4516 99276 4556
rect 99316 4516 99358 4556
rect 99398 4516 99440 4556
rect 99112 4507 99480 4516
rect 1611 4220 1653 4229
rect 1611 4180 1612 4220
rect 1652 4180 1653 4220
rect 1611 4171 1653 4180
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 8352 3800 8720 3809
rect 8392 3760 8434 3800
rect 8474 3760 8516 3800
rect 8556 3760 8598 3800
rect 8638 3760 8680 3800
rect 8352 3751 8720 3760
rect 12352 3800 12720 3809
rect 12392 3760 12434 3800
rect 12474 3760 12516 3800
rect 12556 3760 12598 3800
rect 12638 3760 12680 3800
rect 12352 3751 12720 3760
rect 16352 3800 16720 3809
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16352 3751 16720 3760
rect 20352 3800 20720 3809
rect 20392 3760 20434 3800
rect 20474 3760 20516 3800
rect 20556 3760 20598 3800
rect 20638 3760 20680 3800
rect 20352 3751 20720 3760
rect 24352 3800 24720 3809
rect 24392 3760 24434 3800
rect 24474 3760 24516 3800
rect 24556 3760 24598 3800
rect 24638 3760 24680 3800
rect 24352 3751 24720 3760
rect 28352 3800 28720 3809
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28352 3751 28720 3760
rect 32352 3800 32720 3809
rect 32392 3760 32434 3800
rect 32474 3760 32516 3800
rect 32556 3760 32598 3800
rect 32638 3760 32680 3800
rect 32352 3751 32720 3760
rect 36352 3800 36720 3809
rect 36392 3760 36434 3800
rect 36474 3760 36516 3800
rect 36556 3760 36598 3800
rect 36638 3760 36680 3800
rect 36352 3751 36720 3760
rect 40352 3800 40720 3809
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40352 3751 40720 3760
rect 44352 3800 44720 3809
rect 44392 3760 44434 3800
rect 44474 3760 44516 3800
rect 44556 3760 44598 3800
rect 44638 3760 44680 3800
rect 44352 3751 44720 3760
rect 48352 3800 48720 3809
rect 48392 3760 48434 3800
rect 48474 3760 48516 3800
rect 48556 3760 48598 3800
rect 48638 3760 48680 3800
rect 48352 3751 48720 3760
rect 52352 3800 52720 3809
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52352 3751 52720 3760
rect 56352 3800 56720 3809
rect 56392 3760 56434 3800
rect 56474 3760 56516 3800
rect 56556 3760 56598 3800
rect 56638 3760 56680 3800
rect 56352 3751 56720 3760
rect 60352 3800 60720 3809
rect 60392 3760 60434 3800
rect 60474 3760 60516 3800
rect 60556 3760 60598 3800
rect 60638 3760 60680 3800
rect 60352 3751 60720 3760
rect 64352 3800 64720 3809
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64352 3751 64720 3760
rect 68352 3800 68720 3809
rect 68392 3760 68434 3800
rect 68474 3760 68516 3800
rect 68556 3760 68598 3800
rect 68638 3760 68680 3800
rect 68352 3751 68720 3760
rect 72352 3800 72720 3809
rect 72392 3760 72434 3800
rect 72474 3760 72516 3800
rect 72556 3760 72598 3800
rect 72638 3760 72680 3800
rect 72352 3751 72720 3760
rect 76352 3800 76720 3809
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76352 3751 76720 3760
rect 80352 3800 80720 3809
rect 80392 3760 80434 3800
rect 80474 3760 80516 3800
rect 80556 3760 80598 3800
rect 80638 3760 80680 3800
rect 80352 3751 80720 3760
rect 84352 3800 84720 3809
rect 84392 3760 84434 3800
rect 84474 3760 84516 3800
rect 84556 3760 84598 3800
rect 84638 3760 84680 3800
rect 84352 3751 84720 3760
rect 88352 3800 88720 3809
rect 88392 3760 88434 3800
rect 88474 3760 88516 3800
rect 88556 3760 88598 3800
rect 88638 3760 88680 3800
rect 88352 3751 88720 3760
rect 92352 3800 92720 3809
rect 92392 3760 92434 3800
rect 92474 3760 92516 3800
rect 92556 3760 92598 3800
rect 92638 3760 92680 3800
rect 92352 3751 92720 3760
rect 96352 3800 96720 3809
rect 96392 3760 96434 3800
rect 96474 3760 96516 3800
rect 96556 3760 96598 3800
rect 96638 3760 96680 3800
rect 96352 3751 96720 3760
rect 884 3340 980 3380
rect 844 3331 884 3340
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 7112 3044 7480 3053
rect 7152 3004 7194 3044
rect 7234 3004 7276 3044
rect 7316 3004 7358 3044
rect 7398 3004 7440 3044
rect 7112 2995 7480 3004
rect 11112 3044 11480 3053
rect 11152 3004 11194 3044
rect 11234 3004 11276 3044
rect 11316 3004 11358 3044
rect 11398 3004 11440 3044
rect 11112 2995 11480 3004
rect 15112 3044 15480 3053
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15112 2995 15480 3004
rect 19112 3044 19480 3053
rect 19152 3004 19194 3044
rect 19234 3004 19276 3044
rect 19316 3004 19358 3044
rect 19398 3004 19440 3044
rect 19112 2995 19480 3004
rect 23112 3044 23480 3053
rect 23152 3004 23194 3044
rect 23234 3004 23276 3044
rect 23316 3004 23358 3044
rect 23398 3004 23440 3044
rect 23112 2995 23480 3004
rect 27112 3044 27480 3053
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27112 2995 27480 3004
rect 31112 3044 31480 3053
rect 31152 3004 31194 3044
rect 31234 3004 31276 3044
rect 31316 3004 31358 3044
rect 31398 3004 31440 3044
rect 31112 2995 31480 3004
rect 35112 3044 35480 3053
rect 35152 3004 35194 3044
rect 35234 3004 35276 3044
rect 35316 3004 35358 3044
rect 35398 3004 35440 3044
rect 35112 2995 35480 3004
rect 39112 3044 39480 3053
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39112 2995 39480 3004
rect 43112 3044 43480 3053
rect 43152 3004 43194 3044
rect 43234 3004 43276 3044
rect 43316 3004 43358 3044
rect 43398 3004 43440 3044
rect 43112 2995 43480 3004
rect 47112 3044 47480 3053
rect 47152 3004 47194 3044
rect 47234 3004 47276 3044
rect 47316 3004 47358 3044
rect 47398 3004 47440 3044
rect 47112 2995 47480 3004
rect 51112 3044 51480 3053
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51112 2995 51480 3004
rect 55112 3044 55480 3053
rect 55152 3004 55194 3044
rect 55234 3004 55276 3044
rect 55316 3004 55358 3044
rect 55398 3004 55440 3044
rect 55112 2995 55480 3004
rect 59112 3044 59480 3053
rect 59152 3004 59194 3044
rect 59234 3004 59276 3044
rect 59316 3004 59358 3044
rect 59398 3004 59440 3044
rect 59112 2995 59480 3004
rect 63112 3044 63480 3053
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63112 2995 63480 3004
rect 67112 3044 67480 3053
rect 67152 3004 67194 3044
rect 67234 3004 67276 3044
rect 67316 3004 67358 3044
rect 67398 3004 67440 3044
rect 67112 2995 67480 3004
rect 71112 3044 71480 3053
rect 71152 3004 71194 3044
rect 71234 3004 71276 3044
rect 71316 3004 71358 3044
rect 71398 3004 71440 3044
rect 71112 2995 71480 3004
rect 75112 3044 75480 3053
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75112 2995 75480 3004
rect 79112 3044 79480 3053
rect 79152 3004 79194 3044
rect 79234 3004 79276 3044
rect 79316 3004 79358 3044
rect 79398 3004 79440 3044
rect 79112 2995 79480 3004
rect 83112 3044 83480 3053
rect 83152 3004 83194 3044
rect 83234 3004 83276 3044
rect 83316 3004 83358 3044
rect 83398 3004 83440 3044
rect 83112 2995 83480 3004
rect 87112 3044 87480 3053
rect 87152 3004 87194 3044
rect 87234 3004 87276 3044
rect 87316 3004 87358 3044
rect 87398 3004 87440 3044
rect 87112 2995 87480 3004
rect 91112 3044 91480 3053
rect 91152 3004 91194 3044
rect 91234 3004 91276 3044
rect 91316 3004 91358 3044
rect 91398 3004 91440 3044
rect 91112 2995 91480 3004
rect 95112 3044 95480 3053
rect 95152 3004 95194 3044
rect 95234 3004 95276 3044
rect 95316 3004 95358 3044
rect 95398 3004 95440 3044
rect 95112 2995 95480 3004
rect 99112 3044 99480 3053
rect 99152 3004 99194 3044
rect 99234 3004 99276 3044
rect 99316 3004 99358 3044
rect 99398 3004 99440 3044
rect 99112 2995 99480 3004
rect 844 2708 884 2717
rect 748 2668 844 2708
rect 844 2659 884 2668
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 8352 2288 8720 2297
rect 8392 2248 8434 2288
rect 8474 2248 8516 2288
rect 8556 2248 8598 2288
rect 8638 2248 8680 2288
rect 8352 2239 8720 2248
rect 12352 2288 12720 2297
rect 12392 2248 12434 2288
rect 12474 2248 12516 2288
rect 12556 2248 12598 2288
rect 12638 2248 12680 2288
rect 12352 2239 12720 2248
rect 16352 2288 16720 2297
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16352 2239 16720 2248
rect 20352 2288 20720 2297
rect 20392 2248 20434 2288
rect 20474 2248 20516 2288
rect 20556 2248 20598 2288
rect 20638 2248 20680 2288
rect 20352 2239 20720 2248
rect 24352 2288 24720 2297
rect 24392 2248 24434 2288
rect 24474 2248 24516 2288
rect 24556 2248 24598 2288
rect 24638 2248 24680 2288
rect 24352 2239 24720 2248
rect 28352 2288 28720 2297
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28352 2239 28720 2248
rect 32352 2288 32720 2297
rect 32392 2248 32434 2288
rect 32474 2248 32516 2288
rect 32556 2248 32598 2288
rect 32638 2248 32680 2288
rect 32352 2239 32720 2248
rect 36352 2288 36720 2297
rect 36392 2248 36434 2288
rect 36474 2248 36516 2288
rect 36556 2248 36598 2288
rect 36638 2248 36680 2288
rect 36352 2239 36720 2248
rect 40352 2288 40720 2297
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40352 2239 40720 2248
rect 44352 2288 44720 2297
rect 44392 2248 44434 2288
rect 44474 2248 44516 2288
rect 44556 2248 44598 2288
rect 44638 2248 44680 2288
rect 44352 2239 44720 2248
rect 48352 2288 48720 2297
rect 48392 2248 48434 2288
rect 48474 2248 48516 2288
rect 48556 2248 48598 2288
rect 48638 2248 48680 2288
rect 48352 2239 48720 2248
rect 52352 2288 52720 2297
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52352 2239 52720 2248
rect 56352 2288 56720 2297
rect 56392 2248 56434 2288
rect 56474 2248 56516 2288
rect 56556 2248 56598 2288
rect 56638 2248 56680 2288
rect 56352 2239 56720 2248
rect 60352 2288 60720 2297
rect 60392 2248 60434 2288
rect 60474 2248 60516 2288
rect 60556 2248 60598 2288
rect 60638 2248 60680 2288
rect 60352 2239 60720 2248
rect 64352 2288 64720 2297
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64352 2239 64720 2248
rect 68352 2288 68720 2297
rect 68392 2248 68434 2288
rect 68474 2248 68516 2288
rect 68556 2248 68598 2288
rect 68638 2248 68680 2288
rect 68352 2239 68720 2248
rect 72352 2288 72720 2297
rect 72392 2248 72434 2288
rect 72474 2248 72516 2288
rect 72556 2248 72598 2288
rect 72638 2248 72680 2288
rect 72352 2239 72720 2248
rect 76352 2288 76720 2297
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76352 2239 76720 2248
rect 80352 2288 80720 2297
rect 80392 2248 80434 2288
rect 80474 2248 80516 2288
rect 80556 2248 80598 2288
rect 80638 2248 80680 2288
rect 80352 2239 80720 2248
rect 84352 2288 84720 2297
rect 84392 2248 84434 2288
rect 84474 2248 84516 2288
rect 84556 2248 84598 2288
rect 84638 2248 84680 2288
rect 84352 2239 84720 2248
rect 88352 2288 88720 2297
rect 88392 2248 88434 2288
rect 88474 2248 88516 2288
rect 88556 2248 88598 2288
rect 88638 2248 88680 2288
rect 88352 2239 88720 2248
rect 92352 2288 92720 2297
rect 92392 2248 92434 2288
rect 92474 2248 92516 2288
rect 92556 2248 92598 2288
rect 92638 2248 92680 2288
rect 92352 2239 92720 2248
rect 96352 2288 96720 2297
rect 96392 2248 96434 2288
rect 96474 2248 96516 2288
rect 96556 2248 96598 2288
rect 96638 2248 96680 2288
rect 96352 2239 96720 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 7112 1532 7480 1541
rect 7152 1492 7194 1532
rect 7234 1492 7276 1532
rect 7316 1492 7358 1532
rect 7398 1492 7440 1532
rect 7112 1483 7480 1492
rect 11112 1532 11480 1541
rect 11152 1492 11194 1532
rect 11234 1492 11276 1532
rect 11316 1492 11358 1532
rect 11398 1492 11440 1532
rect 11112 1483 11480 1492
rect 15112 1532 15480 1541
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15112 1483 15480 1492
rect 19112 1532 19480 1541
rect 19152 1492 19194 1532
rect 19234 1492 19276 1532
rect 19316 1492 19358 1532
rect 19398 1492 19440 1532
rect 19112 1483 19480 1492
rect 23112 1532 23480 1541
rect 23152 1492 23194 1532
rect 23234 1492 23276 1532
rect 23316 1492 23358 1532
rect 23398 1492 23440 1532
rect 23112 1483 23480 1492
rect 27112 1532 27480 1541
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27112 1483 27480 1492
rect 31112 1532 31480 1541
rect 31152 1492 31194 1532
rect 31234 1492 31276 1532
rect 31316 1492 31358 1532
rect 31398 1492 31440 1532
rect 31112 1483 31480 1492
rect 35112 1532 35480 1541
rect 35152 1492 35194 1532
rect 35234 1492 35276 1532
rect 35316 1492 35358 1532
rect 35398 1492 35440 1532
rect 35112 1483 35480 1492
rect 39112 1532 39480 1541
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39112 1483 39480 1492
rect 43112 1532 43480 1541
rect 43152 1492 43194 1532
rect 43234 1492 43276 1532
rect 43316 1492 43358 1532
rect 43398 1492 43440 1532
rect 43112 1483 43480 1492
rect 47112 1532 47480 1541
rect 47152 1492 47194 1532
rect 47234 1492 47276 1532
rect 47316 1492 47358 1532
rect 47398 1492 47440 1532
rect 47112 1483 47480 1492
rect 51112 1532 51480 1541
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51112 1483 51480 1492
rect 55112 1532 55480 1541
rect 55152 1492 55194 1532
rect 55234 1492 55276 1532
rect 55316 1492 55358 1532
rect 55398 1492 55440 1532
rect 55112 1483 55480 1492
rect 59112 1532 59480 1541
rect 59152 1492 59194 1532
rect 59234 1492 59276 1532
rect 59316 1492 59358 1532
rect 59398 1492 59440 1532
rect 59112 1483 59480 1492
rect 63112 1532 63480 1541
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63112 1483 63480 1492
rect 67112 1532 67480 1541
rect 67152 1492 67194 1532
rect 67234 1492 67276 1532
rect 67316 1492 67358 1532
rect 67398 1492 67440 1532
rect 67112 1483 67480 1492
rect 71112 1532 71480 1541
rect 71152 1492 71194 1532
rect 71234 1492 71276 1532
rect 71316 1492 71358 1532
rect 71398 1492 71440 1532
rect 71112 1483 71480 1492
rect 75112 1532 75480 1541
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75112 1483 75480 1492
rect 79112 1532 79480 1541
rect 79152 1492 79194 1532
rect 79234 1492 79276 1532
rect 79316 1492 79358 1532
rect 79398 1492 79440 1532
rect 79112 1483 79480 1492
rect 83112 1532 83480 1541
rect 83152 1492 83194 1532
rect 83234 1492 83276 1532
rect 83316 1492 83358 1532
rect 83398 1492 83440 1532
rect 83112 1483 83480 1492
rect 87112 1532 87480 1541
rect 87152 1492 87194 1532
rect 87234 1492 87276 1532
rect 87316 1492 87358 1532
rect 87398 1492 87440 1532
rect 87112 1483 87480 1492
rect 91112 1532 91480 1541
rect 91152 1492 91194 1532
rect 91234 1492 91276 1532
rect 91316 1492 91358 1532
rect 91398 1492 91440 1532
rect 91112 1483 91480 1492
rect 95112 1532 95480 1541
rect 95152 1492 95194 1532
rect 95234 1492 95276 1532
rect 95316 1492 95358 1532
rect 95398 1492 95440 1532
rect 95112 1483 95480 1492
rect 99112 1532 99480 1541
rect 99152 1492 99194 1532
rect 99234 1492 99276 1532
rect 99316 1492 99358 1532
rect 99398 1492 99440 1532
rect 99112 1483 99480 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 8352 776 8720 785
rect 8392 736 8434 776
rect 8474 736 8516 776
rect 8556 736 8598 776
rect 8638 736 8680 776
rect 8352 727 8720 736
rect 12352 776 12720 785
rect 12392 736 12434 776
rect 12474 736 12516 776
rect 12556 736 12598 776
rect 12638 736 12680 776
rect 12352 727 12720 736
rect 16352 776 16720 785
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16352 727 16720 736
rect 20352 776 20720 785
rect 20392 736 20434 776
rect 20474 736 20516 776
rect 20556 736 20598 776
rect 20638 736 20680 776
rect 20352 727 20720 736
rect 24352 776 24720 785
rect 24392 736 24434 776
rect 24474 736 24516 776
rect 24556 736 24598 776
rect 24638 736 24680 776
rect 24352 727 24720 736
rect 28352 776 28720 785
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28352 727 28720 736
rect 32352 776 32720 785
rect 32392 736 32434 776
rect 32474 736 32516 776
rect 32556 736 32598 776
rect 32638 736 32680 776
rect 32352 727 32720 736
rect 36352 776 36720 785
rect 36392 736 36434 776
rect 36474 736 36516 776
rect 36556 736 36598 776
rect 36638 736 36680 776
rect 36352 727 36720 736
rect 40352 776 40720 785
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40352 727 40720 736
rect 44352 776 44720 785
rect 44392 736 44434 776
rect 44474 736 44516 776
rect 44556 736 44598 776
rect 44638 736 44680 776
rect 44352 727 44720 736
rect 48352 776 48720 785
rect 48392 736 48434 776
rect 48474 736 48516 776
rect 48556 736 48598 776
rect 48638 736 48680 776
rect 48352 727 48720 736
rect 52352 776 52720 785
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52352 727 52720 736
rect 56352 776 56720 785
rect 56392 736 56434 776
rect 56474 736 56516 776
rect 56556 736 56598 776
rect 56638 736 56680 776
rect 56352 727 56720 736
rect 60352 776 60720 785
rect 60392 736 60434 776
rect 60474 736 60516 776
rect 60556 736 60598 776
rect 60638 736 60680 776
rect 60352 727 60720 736
rect 64352 776 64720 785
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64352 727 64720 736
rect 68352 776 68720 785
rect 68392 736 68434 776
rect 68474 736 68516 776
rect 68556 736 68598 776
rect 68638 736 68680 776
rect 68352 727 68720 736
rect 72352 776 72720 785
rect 72392 736 72434 776
rect 72474 736 72516 776
rect 72556 736 72598 776
rect 72638 736 72680 776
rect 72352 727 72720 736
rect 76352 776 76720 785
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76352 727 76720 736
rect 80352 776 80720 785
rect 80392 736 80434 776
rect 80474 736 80516 776
rect 80556 736 80598 776
rect 80638 736 80680 776
rect 80352 727 80720 736
rect 84352 776 84720 785
rect 84392 736 84434 776
rect 84474 736 84516 776
rect 84556 736 84598 776
rect 84638 736 84680 776
rect 84352 727 84720 736
rect 88352 776 88720 785
rect 88392 736 88434 776
rect 88474 736 88516 776
rect 88556 736 88598 776
rect 88638 736 88680 776
rect 88352 727 88720 736
rect 92352 776 92720 785
rect 92392 736 92434 776
rect 92474 736 92516 776
rect 92556 736 92598 776
rect 92638 736 92680 776
rect 92352 727 92720 736
rect 96352 776 96720 785
rect 96392 736 96434 776
rect 96474 736 96516 776
rect 96556 736 96598 776
rect 96638 736 96680 776
rect 96352 727 96720 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 8352 38536 8392 38576
rect 8434 38536 8474 38576
rect 8516 38536 8556 38576
rect 8598 38536 8638 38576
rect 8680 38536 8720 38576
rect 12352 38536 12392 38576
rect 12434 38536 12474 38576
rect 12516 38536 12556 38576
rect 12598 38536 12638 38576
rect 12680 38536 12720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 20352 38536 20392 38576
rect 20434 38536 20474 38576
rect 20516 38536 20556 38576
rect 20598 38536 20638 38576
rect 20680 38536 20720 38576
rect 24352 38536 24392 38576
rect 24434 38536 24474 38576
rect 24516 38536 24556 38576
rect 24598 38536 24638 38576
rect 24680 38536 24720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 32352 38536 32392 38576
rect 32434 38536 32474 38576
rect 32516 38536 32556 38576
rect 32598 38536 32638 38576
rect 32680 38536 32720 38576
rect 36352 38536 36392 38576
rect 36434 38536 36474 38576
rect 36516 38536 36556 38576
rect 36598 38536 36638 38576
rect 36680 38536 36720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 44352 38536 44392 38576
rect 44434 38536 44474 38576
rect 44516 38536 44556 38576
rect 44598 38536 44638 38576
rect 44680 38536 44720 38576
rect 48352 38536 48392 38576
rect 48434 38536 48474 38576
rect 48516 38536 48556 38576
rect 48598 38536 48638 38576
rect 48680 38536 48720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 56352 38536 56392 38576
rect 56434 38536 56474 38576
rect 56516 38536 56556 38576
rect 56598 38536 56638 38576
rect 56680 38536 56720 38576
rect 60352 38536 60392 38576
rect 60434 38536 60474 38576
rect 60516 38536 60556 38576
rect 60598 38536 60638 38576
rect 60680 38536 60720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 68352 38536 68392 38576
rect 68434 38536 68474 38576
rect 68516 38536 68556 38576
rect 68598 38536 68638 38576
rect 68680 38536 68720 38576
rect 72352 38536 72392 38576
rect 72434 38536 72474 38576
rect 72516 38536 72556 38576
rect 72598 38536 72638 38576
rect 72680 38536 72720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 80352 38536 80392 38576
rect 80434 38536 80474 38576
rect 80516 38536 80556 38576
rect 80598 38536 80638 38576
rect 80680 38536 80720 38576
rect 84352 38536 84392 38576
rect 84434 38536 84474 38576
rect 84516 38536 84556 38576
rect 84598 38536 84638 38576
rect 84680 38536 84720 38576
rect 88352 38536 88392 38576
rect 88434 38536 88474 38576
rect 88516 38536 88556 38576
rect 88598 38536 88638 38576
rect 88680 38536 88720 38576
rect 92352 38536 92392 38576
rect 92434 38536 92474 38576
rect 92516 38536 92556 38576
rect 92598 38536 92638 38576
rect 92680 38536 92720 38576
rect 96352 38536 96392 38576
rect 96434 38536 96474 38576
rect 96516 38536 96556 38576
rect 96598 38536 96638 38576
rect 96680 38536 96720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 7112 37780 7152 37820
rect 7194 37780 7234 37820
rect 7276 37780 7316 37820
rect 7358 37780 7398 37820
rect 7440 37780 7480 37820
rect 11112 37780 11152 37820
rect 11194 37780 11234 37820
rect 11276 37780 11316 37820
rect 11358 37780 11398 37820
rect 11440 37780 11480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 19112 37780 19152 37820
rect 19194 37780 19234 37820
rect 19276 37780 19316 37820
rect 19358 37780 19398 37820
rect 19440 37780 19480 37820
rect 23112 37780 23152 37820
rect 23194 37780 23234 37820
rect 23276 37780 23316 37820
rect 23358 37780 23398 37820
rect 23440 37780 23480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 31112 37780 31152 37820
rect 31194 37780 31234 37820
rect 31276 37780 31316 37820
rect 31358 37780 31398 37820
rect 31440 37780 31480 37820
rect 35112 37780 35152 37820
rect 35194 37780 35234 37820
rect 35276 37780 35316 37820
rect 35358 37780 35398 37820
rect 35440 37780 35480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 43112 37780 43152 37820
rect 43194 37780 43234 37820
rect 43276 37780 43316 37820
rect 43358 37780 43398 37820
rect 43440 37780 43480 37820
rect 47112 37780 47152 37820
rect 47194 37780 47234 37820
rect 47276 37780 47316 37820
rect 47358 37780 47398 37820
rect 47440 37780 47480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 55112 37780 55152 37820
rect 55194 37780 55234 37820
rect 55276 37780 55316 37820
rect 55358 37780 55398 37820
rect 55440 37780 55480 37820
rect 59112 37780 59152 37820
rect 59194 37780 59234 37820
rect 59276 37780 59316 37820
rect 59358 37780 59398 37820
rect 59440 37780 59480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 67112 37780 67152 37820
rect 67194 37780 67234 37820
rect 67276 37780 67316 37820
rect 67358 37780 67398 37820
rect 67440 37780 67480 37820
rect 71112 37780 71152 37820
rect 71194 37780 71234 37820
rect 71276 37780 71316 37820
rect 71358 37780 71398 37820
rect 71440 37780 71480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 79112 37780 79152 37820
rect 79194 37780 79234 37820
rect 79276 37780 79316 37820
rect 79358 37780 79398 37820
rect 79440 37780 79480 37820
rect 83112 37780 83152 37820
rect 83194 37780 83234 37820
rect 83276 37780 83316 37820
rect 83358 37780 83398 37820
rect 83440 37780 83480 37820
rect 87112 37780 87152 37820
rect 87194 37780 87234 37820
rect 87276 37780 87316 37820
rect 87358 37780 87398 37820
rect 87440 37780 87480 37820
rect 91112 37780 91152 37820
rect 91194 37780 91234 37820
rect 91276 37780 91316 37820
rect 91358 37780 91398 37820
rect 91440 37780 91480 37820
rect 95112 37780 95152 37820
rect 95194 37780 95234 37820
rect 95276 37780 95316 37820
rect 95358 37780 95398 37820
rect 95440 37780 95480 37820
rect 99112 37780 99152 37820
rect 99194 37780 99234 37820
rect 99276 37780 99316 37820
rect 99358 37780 99398 37820
rect 99440 37780 99480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 8352 37024 8392 37064
rect 8434 37024 8474 37064
rect 8516 37024 8556 37064
rect 8598 37024 8638 37064
rect 8680 37024 8720 37064
rect 12352 37024 12392 37064
rect 12434 37024 12474 37064
rect 12516 37024 12556 37064
rect 12598 37024 12638 37064
rect 12680 37024 12720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 20352 37024 20392 37064
rect 20434 37024 20474 37064
rect 20516 37024 20556 37064
rect 20598 37024 20638 37064
rect 20680 37024 20720 37064
rect 24352 37024 24392 37064
rect 24434 37024 24474 37064
rect 24516 37024 24556 37064
rect 24598 37024 24638 37064
rect 24680 37024 24720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 32352 37024 32392 37064
rect 32434 37024 32474 37064
rect 32516 37024 32556 37064
rect 32598 37024 32638 37064
rect 32680 37024 32720 37064
rect 36352 37024 36392 37064
rect 36434 37024 36474 37064
rect 36516 37024 36556 37064
rect 36598 37024 36638 37064
rect 36680 37024 36720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 44352 37024 44392 37064
rect 44434 37024 44474 37064
rect 44516 37024 44556 37064
rect 44598 37024 44638 37064
rect 44680 37024 44720 37064
rect 48352 37024 48392 37064
rect 48434 37024 48474 37064
rect 48516 37024 48556 37064
rect 48598 37024 48638 37064
rect 48680 37024 48720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 56352 37024 56392 37064
rect 56434 37024 56474 37064
rect 56516 37024 56556 37064
rect 56598 37024 56638 37064
rect 56680 37024 56720 37064
rect 60352 37024 60392 37064
rect 60434 37024 60474 37064
rect 60516 37024 60556 37064
rect 60598 37024 60638 37064
rect 60680 37024 60720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 68352 37024 68392 37064
rect 68434 37024 68474 37064
rect 68516 37024 68556 37064
rect 68598 37024 68638 37064
rect 68680 37024 68720 37064
rect 72352 37024 72392 37064
rect 72434 37024 72474 37064
rect 72516 37024 72556 37064
rect 72598 37024 72638 37064
rect 72680 37024 72720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 80352 37024 80392 37064
rect 80434 37024 80474 37064
rect 80516 37024 80556 37064
rect 80598 37024 80638 37064
rect 80680 37024 80720 37064
rect 84352 37024 84392 37064
rect 84434 37024 84474 37064
rect 84516 37024 84556 37064
rect 84598 37024 84638 37064
rect 84680 37024 84720 37064
rect 88352 37024 88392 37064
rect 88434 37024 88474 37064
rect 88516 37024 88556 37064
rect 88598 37024 88638 37064
rect 88680 37024 88720 37064
rect 92352 37024 92392 37064
rect 92434 37024 92474 37064
rect 92516 37024 92556 37064
rect 92598 37024 92638 37064
rect 92680 37024 92720 37064
rect 96352 37024 96392 37064
rect 96434 37024 96474 37064
rect 96516 37024 96556 37064
rect 96598 37024 96638 37064
rect 96680 37024 96720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 7112 36268 7152 36308
rect 7194 36268 7234 36308
rect 7276 36268 7316 36308
rect 7358 36268 7398 36308
rect 7440 36268 7480 36308
rect 11112 36268 11152 36308
rect 11194 36268 11234 36308
rect 11276 36268 11316 36308
rect 11358 36268 11398 36308
rect 11440 36268 11480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 19112 36268 19152 36308
rect 19194 36268 19234 36308
rect 19276 36268 19316 36308
rect 19358 36268 19398 36308
rect 19440 36268 19480 36308
rect 23112 36268 23152 36308
rect 23194 36268 23234 36308
rect 23276 36268 23316 36308
rect 23358 36268 23398 36308
rect 23440 36268 23480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 31112 36268 31152 36308
rect 31194 36268 31234 36308
rect 31276 36268 31316 36308
rect 31358 36268 31398 36308
rect 31440 36268 31480 36308
rect 35112 36268 35152 36308
rect 35194 36268 35234 36308
rect 35276 36268 35316 36308
rect 35358 36268 35398 36308
rect 35440 36268 35480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 43112 36268 43152 36308
rect 43194 36268 43234 36308
rect 43276 36268 43316 36308
rect 43358 36268 43398 36308
rect 43440 36268 43480 36308
rect 47112 36268 47152 36308
rect 47194 36268 47234 36308
rect 47276 36268 47316 36308
rect 47358 36268 47398 36308
rect 47440 36268 47480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 55112 36268 55152 36308
rect 55194 36268 55234 36308
rect 55276 36268 55316 36308
rect 55358 36268 55398 36308
rect 55440 36268 55480 36308
rect 59112 36268 59152 36308
rect 59194 36268 59234 36308
rect 59276 36268 59316 36308
rect 59358 36268 59398 36308
rect 59440 36268 59480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 67112 36268 67152 36308
rect 67194 36268 67234 36308
rect 67276 36268 67316 36308
rect 67358 36268 67398 36308
rect 67440 36268 67480 36308
rect 71112 36268 71152 36308
rect 71194 36268 71234 36308
rect 71276 36268 71316 36308
rect 71358 36268 71398 36308
rect 71440 36268 71480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 79112 36268 79152 36308
rect 79194 36268 79234 36308
rect 79276 36268 79316 36308
rect 79358 36268 79398 36308
rect 79440 36268 79480 36308
rect 83112 36268 83152 36308
rect 83194 36268 83234 36308
rect 83276 36268 83316 36308
rect 83358 36268 83398 36308
rect 83440 36268 83480 36308
rect 87112 36268 87152 36308
rect 87194 36268 87234 36308
rect 87276 36268 87316 36308
rect 87358 36268 87398 36308
rect 87440 36268 87480 36308
rect 91112 36268 91152 36308
rect 91194 36268 91234 36308
rect 91276 36268 91316 36308
rect 91358 36268 91398 36308
rect 91440 36268 91480 36308
rect 95112 36268 95152 36308
rect 95194 36268 95234 36308
rect 95276 36268 95316 36308
rect 95358 36268 95398 36308
rect 95440 36268 95480 36308
rect 99112 36268 99152 36308
rect 99194 36268 99234 36308
rect 99276 36268 99316 36308
rect 99358 36268 99398 36308
rect 99440 36268 99480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 8352 35512 8392 35552
rect 8434 35512 8474 35552
rect 8516 35512 8556 35552
rect 8598 35512 8638 35552
rect 8680 35512 8720 35552
rect 12352 35512 12392 35552
rect 12434 35512 12474 35552
rect 12516 35512 12556 35552
rect 12598 35512 12638 35552
rect 12680 35512 12720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 20352 35512 20392 35552
rect 20434 35512 20474 35552
rect 20516 35512 20556 35552
rect 20598 35512 20638 35552
rect 20680 35512 20720 35552
rect 24352 35512 24392 35552
rect 24434 35512 24474 35552
rect 24516 35512 24556 35552
rect 24598 35512 24638 35552
rect 24680 35512 24720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 32352 35512 32392 35552
rect 32434 35512 32474 35552
rect 32516 35512 32556 35552
rect 32598 35512 32638 35552
rect 32680 35512 32720 35552
rect 36352 35512 36392 35552
rect 36434 35512 36474 35552
rect 36516 35512 36556 35552
rect 36598 35512 36638 35552
rect 36680 35512 36720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 44352 35512 44392 35552
rect 44434 35512 44474 35552
rect 44516 35512 44556 35552
rect 44598 35512 44638 35552
rect 44680 35512 44720 35552
rect 48352 35512 48392 35552
rect 48434 35512 48474 35552
rect 48516 35512 48556 35552
rect 48598 35512 48638 35552
rect 48680 35512 48720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 56352 35512 56392 35552
rect 56434 35512 56474 35552
rect 56516 35512 56556 35552
rect 56598 35512 56638 35552
rect 56680 35512 56720 35552
rect 60352 35512 60392 35552
rect 60434 35512 60474 35552
rect 60516 35512 60556 35552
rect 60598 35512 60638 35552
rect 60680 35512 60720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 68352 35512 68392 35552
rect 68434 35512 68474 35552
rect 68516 35512 68556 35552
rect 68598 35512 68638 35552
rect 68680 35512 68720 35552
rect 72352 35512 72392 35552
rect 72434 35512 72474 35552
rect 72516 35512 72556 35552
rect 72598 35512 72638 35552
rect 72680 35512 72720 35552
rect 73900 35092 73940 35132
rect 74092 35092 74132 35132
rect 73708 35008 73748 35048
rect 74476 35008 74516 35048
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 7112 34756 7152 34796
rect 7194 34756 7234 34796
rect 7276 34756 7316 34796
rect 7358 34756 7398 34796
rect 7440 34756 7480 34796
rect 11112 34756 11152 34796
rect 11194 34756 11234 34796
rect 11276 34756 11316 34796
rect 11358 34756 11398 34796
rect 11440 34756 11480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 19112 34756 19152 34796
rect 19194 34756 19234 34796
rect 19276 34756 19316 34796
rect 19358 34756 19398 34796
rect 19440 34756 19480 34796
rect 23112 34756 23152 34796
rect 23194 34756 23234 34796
rect 23276 34756 23316 34796
rect 23358 34756 23398 34796
rect 23440 34756 23480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 31112 34756 31152 34796
rect 31194 34756 31234 34796
rect 31276 34756 31316 34796
rect 31358 34756 31398 34796
rect 31440 34756 31480 34796
rect 35112 34756 35152 34796
rect 35194 34756 35234 34796
rect 35276 34756 35316 34796
rect 35358 34756 35398 34796
rect 35440 34756 35480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 43112 34756 43152 34796
rect 43194 34756 43234 34796
rect 43276 34756 43316 34796
rect 43358 34756 43398 34796
rect 43440 34756 43480 34796
rect 47112 34756 47152 34796
rect 47194 34756 47234 34796
rect 47276 34756 47316 34796
rect 47358 34756 47398 34796
rect 47440 34756 47480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 55112 34756 55152 34796
rect 55194 34756 55234 34796
rect 55276 34756 55316 34796
rect 55358 34756 55398 34796
rect 55440 34756 55480 34796
rect 59112 34756 59152 34796
rect 59194 34756 59234 34796
rect 59276 34756 59316 34796
rect 59358 34756 59398 34796
rect 59440 34756 59480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 67112 34756 67152 34796
rect 67194 34756 67234 34796
rect 67276 34756 67316 34796
rect 67358 34756 67398 34796
rect 67440 34756 67480 34796
rect 71112 34756 71152 34796
rect 71194 34756 71234 34796
rect 71276 34756 71316 34796
rect 71358 34756 71398 34796
rect 71440 34756 71480 34796
rect 69772 34420 69812 34460
rect 73420 34420 73460 34460
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 8352 34000 8392 34040
rect 8434 34000 8474 34040
rect 8516 34000 8556 34040
rect 8598 34000 8638 34040
rect 8680 34000 8720 34040
rect 12352 34000 12392 34040
rect 12434 34000 12474 34040
rect 12516 34000 12556 34040
rect 12598 34000 12638 34040
rect 12680 34000 12720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 20352 34000 20392 34040
rect 20434 34000 20474 34040
rect 20516 34000 20556 34040
rect 20598 34000 20638 34040
rect 20680 34000 20720 34040
rect 24352 34000 24392 34040
rect 24434 34000 24474 34040
rect 24516 34000 24556 34040
rect 24598 34000 24638 34040
rect 24680 34000 24720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 32352 34000 32392 34040
rect 32434 34000 32474 34040
rect 32516 34000 32556 34040
rect 32598 34000 32638 34040
rect 32680 34000 32720 34040
rect 36352 34000 36392 34040
rect 36434 34000 36474 34040
rect 36516 34000 36556 34040
rect 36598 34000 36638 34040
rect 36680 34000 36720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 44352 34000 44392 34040
rect 44434 34000 44474 34040
rect 44516 34000 44556 34040
rect 44598 34000 44638 34040
rect 44680 34000 44720 34040
rect 48352 34000 48392 34040
rect 48434 34000 48474 34040
rect 48516 34000 48556 34040
rect 48598 34000 48638 34040
rect 48680 34000 48720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 56352 34000 56392 34040
rect 56434 34000 56474 34040
rect 56516 34000 56556 34040
rect 56598 34000 56638 34040
rect 56680 34000 56720 34040
rect 60352 34000 60392 34040
rect 60434 34000 60474 34040
rect 60516 34000 60556 34040
rect 60598 34000 60638 34040
rect 60680 34000 60720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 68352 34000 68392 34040
rect 68434 34000 68474 34040
rect 68516 34000 68556 34040
rect 68598 34000 68638 34040
rect 68680 34000 68720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 7112 33244 7152 33284
rect 7194 33244 7234 33284
rect 7276 33244 7316 33284
rect 7358 33244 7398 33284
rect 7440 33244 7480 33284
rect 11112 33244 11152 33284
rect 11194 33244 11234 33284
rect 11276 33244 11316 33284
rect 11358 33244 11398 33284
rect 11440 33244 11480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 19112 33244 19152 33284
rect 19194 33244 19234 33284
rect 19276 33244 19316 33284
rect 19358 33244 19398 33284
rect 19440 33244 19480 33284
rect 23112 33244 23152 33284
rect 23194 33244 23234 33284
rect 23276 33244 23316 33284
rect 23358 33244 23398 33284
rect 23440 33244 23480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 31112 33244 31152 33284
rect 31194 33244 31234 33284
rect 31276 33244 31316 33284
rect 31358 33244 31398 33284
rect 31440 33244 31480 33284
rect 35112 33244 35152 33284
rect 35194 33244 35234 33284
rect 35276 33244 35316 33284
rect 35358 33244 35398 33284
rect 35440 33244 35480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 43112 33244 43152 33284
rect 43194 33244 43234 33284
rect 43276 33244 43316 33284
rect 43358 33244 43398 33284
rect 43440 33244 43480 33284
rect 47112 33244 47152 33284
rect 47194 33244 47234 33284
rect 47276 33244 47316 33284
rect 47358 33244 47398 33284
rect 47440 33244 47480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 55112 33244 55152 33284
rect 55194 33244 55234 33284
rect 55276 33244 55316 33284
rect 55358 33244 55398 33284
rect 55440 33244 55480 33284
rect 59112 33244 59152 33284
rect 59194 33244 59234 33284
rect 59276 33244 59316 33284
rect 59358 33244 59398 33284
rect 59440 33244 59480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 67112 33244 67152 33284
rect 67194 33244 67234 33284
rect 67276 33244 67316 33284
rect 67358 33244 67398 33284
rect 67440 33244 67480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 8352 32488 8392 32528
rect 8434 32488 8474 32528
rect 8516 32488 8556 32528
rect 8598 32488 8638 32528
rect 8680 32488 8720 32528
rect 12352 32488 12392 32528
rect 12434 32488 12474 32528
rect 12516 32488 12556 32528
rect 12598 32488 12638 32528
rect 12680 32488 12720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 20352 32488 20392 32528
rect 20434 32488 20474 32528
rect 20516 32488 20556 32528
rect 20598 32488 20638 32528
rect 20680 32488 20720 32528
rect 24352 32488 24392 32528
rect 24434 32488 24474 32528
rect 24516 32488 24556 32528
rect 24598 32488 24638 32528
rect 24680 32488 24720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 32352 32488 32392 32528
rect 32434 32488 32474 32528
rect 32516 32488 32556 32528
rect 32598 32488 32638 32528
rect 32680 32488 32720 32528
rect 36352 32488 36392 32528
rect 36434 32488 36474 32528
rect 36516 32488 36556 32528
rect 36598 32488 36638 32528
rect 36680 32488 36720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 44352 32488 44392 32528
rect 44434 32488 44474 32528
rect 44516 32488 44556 32528
rect 44598 32488 44638 32528
rect 44680 32488 44720 32528
rect 48352 32488 48392 32528
rect 48434 32488 48474 32528
rect 48516 32488 48556 32528
rect 48598 32488 48638 32528
rect 48680 32488 48720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 56352 32488 56392 32528
rect 56434 32488 56474 32528
rect 56516 32488 56556 32528
rect 56598 32488 56638 32528
rect 56680 32488 56720 32528
rect 60352 32488 60392 32528
rect 60434 32488 60474 32528
rect 60516 32488 60556 32528
rect 60598 32488 60638 32528
rect 60680 32488 60720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 68352 32488 68392 32528
rect 68434 32488 68474 32528
rect 68516 32488 68556 32528
rect 68598 32488 68638 32528
rect 68680 32488 68720 32528
rect 72352 34000 72392 34040
rect 72434 34000 72474 34040
rect 72516 34000 72556 34040
rect 72598 34000 72638 34040
rect 72680 34000 72720 34040
rect 71788 32740 71828 32780
rect 67564 32068 67604 32108
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 7112 31732 7152 31772
rect 7194 31732 7234 31772
rect 7276 31732 7316 31772
rect 7358 31732 7398 31772
rect 7440 31732 7480 31772
rect 11112 31732 11152 31772
rect 11194 31732 11234 31772
rect 11276 31732 11316 31772
rect 11358 31732 11398 31772
rect 11440 31732 11480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 19112 31732 19152 31772
rect 19194 31732 19234 31772
rect 19276 31732 19316 31772
rect 19358 31732 19398 31772
rect 19440 31732 19480 31772
rect 23112 31732 23152 31772
rect 23194 31732 23234 31772
rect 23276 31732 23316 31772
rect 23358 31732 23398 31772
rect 23440 31732 23480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 31112 31732 31152 31772
rect 31194 31732 31234 31772
rect 31276 31732 31316 31772
rect 31358 31732 31398 31772
rect 31440 31732 31480 31772
rect 35112 31732 35152 31772
rect 35194 31732 35234 31772
rect 35276 31732 35316 31772
rect 35358 31732 35398 31772
rect 35440 31732 35480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 43112 31732 43152 31772
rect 43194 31732 43234 31772
rect 43276 31732 43316 31772
rect 43358 31732 43398 31772
rect 43440 31732 43480 31772
rect 47112 31732 47152 31772
rect 47194 31732 47234 31772
rect 47276 31732 47316 31772
rect 47358 31732 47398 31772
rect 47440 31732 47480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 55112 31732 55152 31772
rect 55194 31732 55234 31772
rect 55276 31732 55316 31772
rect 55358 31732 55398 31772
rect 55440 31732 55480 31772
rect 59112 31732 59152 31772
rect 59194 31732 59234 31772
rect 59276 31732 59316 31772
rect 59358 31732 59398 31772
rect 59440 31732 59480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 67112 31732 67152 31772
rect 67194 31732 67234 31772
rect 67276 31732 67316 31772
rect 67358 31732 67398 31772
rect 67440 31732 67480 31772
rect 68908 31816 68948 31856
rect 67180 31564 67220 31604
rect 67564 31564 67604 31604
rect 68812 31564 68852 31604
rect 67660 31480 67700 31520
rect 67276 31228 67316 31268
rect 67564 31228 67604 31268
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 8352 30976 8392 31016
rect 8434 30976 8474 31016
rect 8516 30976 8556 31016
rect 8598 30976 8638 31016
rect 8680 30976 8720 31016
rect 12352 30976 12392 31016
rect 12434 30976 12474 31016
rect 12516 30976 12556 31016
rect 12598 30976 12638 31016
rect 12680 30976 12720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 20352 30976 20392 31016
rect 20434 30976 20474 31016
rect 20516 30976 20556 31016
rect 20598 30976 20638 31016
rect 20680 30976 20720 31016
rect 24352 30976 24392 31016
rect 24434 30976 24474 31016
rect 24516 30976 24556 31016
rect 24598 30976 24638 31016
rect 24680 30976 24720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 32352 30976 32392 31016
rect 32434 30976 32474 31016
rect 32516 30976 32556 31016
rect 32598 30976 32638 31016
rect 32680 30976 32720 31016
rect 36352 30976 36392 31016
rect 36434 30976 36474 31016
rect 36516 30976 36556 31016
rect 36598 30976 36638 31016
rect 36680 30976 36720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 44352 30976 44392 31016
rect 44434 30976 44474 31016
rect 44516 30976 44556 31016
rect 44598 30976 44638 31016
rect 44680 30976 44720 31016
rect 48352 30976 48392 31016
rect 48434 30976 48474 31016
rect 48516 30976 48556 31016
rect 48598 30976 48638 31016
rect 48680 30976 48720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 56352 30976 56392 31016
rect 56434 30976 56474 31016
rect 56516 30976 56556 31016
rect 56598 30976 56638 31016
rect 56680 30976 56720 31016
rect 60352 30976 60392 31016
rect 60434 30976 60474 31016
rect 60516 30976 60556 31016
rect 60598 30976 60638 31016
rect 60680 30976 60720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 68620 31228 68660 31268
rect 68352 30976 68392 31016
rect 68434 30976 68474 31016
rect 68516 30976 68556 31016
rect 68598 30976 68638 31016
rect 68680 30976 68720 31016
rect 69484 31732 69524 31772
rect 69196 31480 69236 31520
rect 68524 30724 68564 30764
rect 67756 30640 67796 30680
rect 68044 30640 68084 30680
rect 69292 31228 69332 31268
rect 69100 30808 69140 30848
rect 69388 31144 69428 31184
rect 69580 31480 69620 31520
rect 69676 31312 69716 31352
rect 69868 31900 69908 31940
rect 69868 31564 69908 31604
rect 69580 31144 69620 31184
rect 69292 30724 69332 30764
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 7112 30220 7152 30260
rect 7194 30220 7234 30260
rect 7276 30220 7316 30260
rect 7358 30220 7398 30260
rect 7440 30220 7480 30260
rect 11112 30220 11152 30260
rect 11194 30220 11234 30260
rect 11276 30220 11316 30260
rect 11358 30220 11398 30260
rect 11440 30220 11480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 19112 30220 19152 30260
rect 19194 30220 19234 30260
rect 19276 30220 19316 30260
rect 19358 30220 19398 30260
rect 19440 30220 19480 30260
rect 23112 30220 23152 30260
rect 23194 30220 23234 30260
rect 23276 30220 23316 30260
rect 23358 30220 23398 30260
rect 23440 30220 23480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 31112 30220 31152 30260
rect 31194 30220 31234 30260
rect 31276 30220 31316 30260
rect 31358 30220 31398 30260
rect 31440 30220 31480 30260
rect 35112 30220 35152 30260
rect 35194 30220 35234 30260
rect 35276 30220 35316 30260
rect 35358 30220 35398 30260
rect 35440 30220 35480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 43112 30220 43152 30260
rect 43194 30220 43234 30260
rect 43276 30220 43316 30260
rect 43358 30220 43398 30260
rect 43440 30220 43480 30260
rect 47112 30220 47152 30260
rect 47194 30220 47234 30260
rect 47276 30220 47316 30260
rect 47358 30220 47398 30260
rect 47440 30220 47480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 55112 30220 55152 30260
rect 55194 30220 55234 30260
rect 55276 30220 55316 30260
rect 55358 30220 55398 30260
rect 55440 30220 55480 30260
rect 59112 30220 59152 30260
rect 59194 30220 59234 30260
rect 59276 30220 59316 30260
rect 59358 30220 59398 30260
rect 59440 30220 59480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 67112 30220 67152 30260
rect 67194 30220 67234 30260
rect 67276 30220 67316 30260
rect 67358 30220 67398 30260
rect 67440 30220 67480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 8352 29464 8392 29504
rect 8434 29464 8474 29504
rect 8516 29464 8556 29504
rect 8598 29464 8638 29504
rect 8680 29464 8720 29504
rect 12352 29464 12392 29504
rect 12434 29464 12474 29504
rect 12516 29464 12556 29504
rect 12598 29464 12638 29504
rect 12680 29464 12720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 20352 29464 20392 29504
rect 20434 29464 20474 29504
rect 20516 29464 20556 29504
rect 20598 29464 20638 29504
rect 20680 29464 20720 29504
rect 24352 29464 24392 29504
rect 24434 29464 24474 29504
rect 24516 29464 24556 29504
rect 24598 29464 24638 29504
rect 24680 29464 24720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 32352 29464 32392 29504
rect 32434 29464 32474 29504
rect 32516 29464 32556 29504
rect 32598 29464 32638 29504
rect 32680 29464 32720 29504
rect 36352 29464 36392 29504
rect 36434 29464 36474 29504
rect 36516 29464 36556 29504
rect 36598 29464 36638 29504
rect 36680 29464 36720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 44352 29464 44392 29504
rect 44434 29464 44474 29504
rect 44516 29464 44556 29504
rect 44598 29464 44638 29504
rect 44680 29464 44720 29504
rect 48352 29464 48392 29504
rect 48434 29464 48474 29504
rect 48516 29464 48556 29504
rect 48598 29464 48638 29504
rect 48680 29464 48720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 56352 29464 56392 29504
rect 56434 29464 56474 29504
rect 56516 29464 56556 29504
rect 56598 29464 56638 29504
rect 56680 29464 56720 29504
rect 60352 29464 60392 29504
rect 60434 29464 60474 29504
rect 60516 29464 60556 29504
rect 60598 29464 60638 29504
rect 60680 29464 60720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 7112 28708 7152 28748
rect 7194 28708 7234 28748
rect 7276 28708 7316 28748
rect 7358 28708 7398 28748
rect 7440 28708 7480 28748
rect 11112 28708 11152 28748
rect 11194 28708 11234 28748
rect 11276 28708 11316 28748
rect 11358 28708 11398 28748
rect 11440 28708 11480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 19112 28708 19152 28748
rect 19194 28708 19234 28748
rect 19276 28708 19316 28748
rect 19358 28708 19398 28748
rect 19440 28708 19480 28748
rect 23112 28708 23152 28748
rect 23194 28708 23234 28748
rect 23276 28708 23316 28748
rect 23358 28708 23398 28748
rect 23440 28708 23480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 31112 28708 31152 28748
rect 31194 28708 31234 28748
rect 31276 28708 31316 28748
rect 31358 28708 31398 28748
rect 31440 28708 31480 28748
rect 35112 28708 35152 28748
rect 35194 28708 35234 28748
rect 35276 28708 35316 28748
rect 35358 28708 35398 28748
rect 35440 28708 35480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 43112 28708 43152 28748
rect 43194 28708 43234 28748
rect 43276 28708 43316 28748
rect 43358 28708 43398 28748
rect 43440 28708 43480 28748
rect 47112 28708 47152 28748
rect 47194 28708 47234 28748
rect 47276 28708 47316 28748
rect 47358 28708 47398 28748
rect 47440 28708 47480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 55112 28708 55152 28748
rect 55194 28708 55234 28748
rect 55276 28708 55316 28748
rect 55358 28708 55398 28748
rect 55440 28708 55480 28748
rect 59112 28708 59152 28748
rect 59194 28708 59234 28748
rect 59276 28708 59316 28748
rect 59358 28708 59398 28748
rect 59440 28708 59480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 67112 28708 67152 28748
rect 67194 28708 67234 28748
rect 67276 28708 67316 28748
rect 67358 28708 67398 28748
rect 67440 28708 67480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 8352 27952 8392 27992
rect 8434 27952 8474 27992
rect 8516 27952 8556 27992
rect 8598 27952 8638 27992
rect 8680 27952 8720 27992
rect 12352 27952 12392 27992
rect 12434 27952 12474 27992
rect 12516 27952 12556 27992
rect 12598 27952 12638 27992
rect 12680 27952 12720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 20352 27952 20392 27992
rect 20434 27952 20474 27992
rect 20516 27952 20556 27992
rect 20598 27952 20638 27992
rect 20680 27952 20720 27992
rect 24352 27952 24392 27992
rect 24434 27952 24474 27992
rect 24516 27952 24556 27992
rect 24598 27952 24638 27992
rect 24680 27952 24720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 32352 27952 32392 27992
rect 32434 27952 32474 27992
rect 32516 27952 32556 27992
rect 32598 27952 32638 27992
rect 32680 27952 32720 27992
rect 36352 27952 36392 27992
rect 36434 27952 36474 27992
rect 36516 27952 36556 27992
rect 36598 27952 36638 27992
rect 36680 27952 36720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 44352 27952 44392 27992
rect 44434 27952 44474 27992
rect 44516 27952 44556 27992
rect 44598 27952 44638 27992
rect 44680 27952 44720 27992
rect 48352 27952 48392 27992
rect 48434 27952 48474 27992
rect 48516 27952 48556 27992
rect 48598 27952 48638 27992
rect 48680 27952 48720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 56352 27952 56392 27992
rect 56434 27952 56474 27992
rect 56516 27952 56556 27992
rect 56598 27952 56638 27992
rect 56680 27952 56720 27992
rect 60352 27952 60392 27992
rect 60434 27952 60474 27992
rect 60516 27952 60556 27992
rect 60598 27952 60638 27992
rect 60680 27952 60720 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 7112 27196 7152 27236
rect 7194 27196 7234 27236
rect 7276 27196 7316 27236
rect 7358 27196 7398 27236
rect 7440 27196 7480 27236
rect 11112 27196 11152 27236
rect 11194 27196 11234 27236
rect 11276 27196 11316 27236
rect 11358 27196 11398 27236
rect 11440 27196 11480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 19112 27196 19152 27236
rect 19194 27196 19234 27236
rect 19276 27196 19316 27236
rect 19358 27196 19398 27236
rect 19440 27196 19480 27236
rect 23112 27196 23152 27236
rect 23194 27196 23234 27236
rect 23276 27196 23316 27236
rect 23358 27196 23398 27236
rect 23440 27196 23480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 31112 27196 31152 27236
rect 31194 27196 31234 27236
rect 31276 27196 31316 27236
rect 31358 27196 31398 27236
rect 31440 27196 31480 27236
rect 35112 27196 35152 27236
rect 35194 27196 35234 27236
rect 35276 27196 35316 27236
rect 35358 27196 35398 27236
rect 35440 27196 35480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 43112 27196 43152 27236
rect 43194 27196 43234 27236
rect 43276 27196 43316 27236
rect 43358 27196 43398 27236
rect 43440 27196 43480 27236
rect 47112 27196 47152 27236
rect 47194 27196 47234 27236
rect 47276 27196 47316 27236
rect 47358 27196 47398 27236
rect 47440 27196 47480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 55112 27196 55152 27236
rect 55194 27196 55234 27236
rect 55276 27196 55316 27236
rect 55358 27196 55398 27236
rect 55440 27196 55480 27236
rect 59112 27196 59152 27236
rect 59194 27196 59234 27236
rect 59276 27196 59316 27236
rect 59358 27196 59398 27236
rect 59440 27196 59480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 67112 27196 67152 27236
rect 67194 27196 67234 27236
rect 67276 27196 67316 27236
rect 67358 27196 67398 27236
rect 67440 27196 67480 27236
rect 69004 30640 69044 30680
rect 69772 31228 69812 31268
rect 68352 29464 68392 29504
rect 68434 29464 68474 29504
rect 68516 29464 68556 29504
rect 68598 29464 68638 29504
rect 68680 29464 68720 29504
rect 68352 27952 68392 27992
rect 68434 27952 68474 27992
rect 68516 27952 68556 27992
rect 68598 27952 68638 27992
rect 68680 27952 68720 27992
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 8352 26440 8392 26480
rect 8434 26440 8474 26480
rect 8516 26440 8556 26480
rect 8598 26440 8638 26480
rect 8680 26440 8720 26480
rect 12352 26440 12392 26480
rect 12434 26440 12474 26480
rect 12516 26440 12556 26480
rect 12598 26440 12638 26480
rect 12680 26440 12720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 20352 26440 20392 26480
rect 20434 26440 20474 26480
rect 20516 26440 20556 26480
rect 20598 26440 20638 26480
rect 20680 26440 20720 26480
rect 24352 26440 24392 26480
rect 24434 26440 24474 26480
rect 24516 26440 24556 26480
rect 24598 26440 24638 26480
rect 24680 26440 24720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 32352 26440 32392 26480
rect 32434 26440 32474 26480
rect 32516 26440 32556 26480
rect 32598 26440 32638 26480
rect 32680 26440 32720 26480
rect 36352 26440 36392 26480
rect 36434 26440 36474 26480
rect 36516 26440 36556 26480
rect 36598 26440 36638 26480
rect 36680 26440 36720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 44352 26440 44392 26480
rect 44434 26440 44474 26480
rect 44516 26440 44556 26480
rect 44598 26440 44638 26480
rect 44680 26440 44720 26480
rect 48352 26440 48392 26480
rect 48434 26440 48474 26480
rect 48516 26440 48556 26480
rect 48598 26440 48638 26480
rect 48680 26440 48720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 56352 26440 56392 26480
rect 56434 26440 56474 26480
rect 56516 26440 56556 26480
rect 56598 26440 56638 26480
rect 56680 26440 56720 26480
rect 60352 26440 60392 26480
rect 60434 26440 60474 26480
rect 60516 26440 60556 26480
rect 60598 26440 60638 26480
rect 60680 26440 60720 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 7112 25684 7152 25724
rect 7194 25684 7234 25724
rect 7276 25684 7316 25724
rect 7358 25684 7398 25724
rect 7440 25684 7480 25724
rect 11112 25684 11152 25724
rect 11194 25684 11234 25724
rect 11276 25684 11316 25724
rect 11358 25684 11398 25724
rect 11440 25684 11480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 19112 25684 19152 25724
rect 19194 25684 19234 25724
rect 19276 25684 19316 25724
rect 19358 25684 19398 25724
rect 19440 25684 19480 25724
rect 23112 25684 23152 25724
rect 23194 25684 23234 25724
rect 23276 25684 23316 25724
rect 23358 25684 23398 25724
rect 23440 25684 23480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 31112 25684 31152 25724
rect 31194 25684 31234 25724
rect 31276 25684 31316 25724
rect 31358 25684 31398 25724
rect 31440 25684 31480 25724
rect 35112 25684 35152 25724
rect 35194 25684 35234 25724
rect 35276 25684 35316 25724
rect 35358 25684 35398 25724
rect 35440 25684 35480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 43112 25684 43152 25724
rect 43194 25684 43234 25724
rect 43276 25684 43316 25724
rect 43358 25684 43398 25724
rect 43440 25684 43480 25724
rect 47112 25684 47152 25724
rect 47194 25684 47234 25724
rect 47276 25684 47316 25724
rect 47358 25684 47398 25724
rect 47440 25684 47480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 55112 25684 55152 25724
rect 55194 25684 55234 25724
rect 55276 25684 55316 25724
rect 55358 25684 55398 25724
rect 55440 25684 55480 25724
rect 59112 25684 59152 25724
rect 59194 25684 59234 25724
rect 59276 25684 59316 25724
rect 59358 25684 59398 25724
rect 59440 25684 59480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 67112 25684 67152 25724
rect 67194 25684 67234 25724
rect 67276 25684 67316 25724
rect 67358 25684 67398 25724
rect 67440 25684 67480 25724
rect 844 25264 884 25304
rect 652 24928 692 24968
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 8352 24928 8392 24968
rect 8434 24928 8474 24968
rect 8516 24928 8556 24968
rect 8598 24928 8638 24968
rect 8680 24928 8720 24968
rect 12352 24928 12392 24968
rect 12434 24928 12474 24968
rect 12516 24928 12556 24968
rect 12598 24928 12638 24968
rect 12680 24928 12720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 20352 24928 20392 24968
rect 20434 24928 20474 24968
rect 20516 24928 20556 24968
rect 20598 24928 20638 24968
rect 20680 24928 20720 24968
rect 24352 24928 24392 24968
rect 24434 24928 24474 24968
rect 24516 24928 24556 24968
rect 24598 24928 24638 24968
rect 24680 24928 24720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 32352 24928 32392 24968
rect 32434 24928 32474 24968
rect 32516 24928 32556 24968
rect 32598 24928 32638 24968
rect 32680 24928 32720 24968
rect 36352 24928 36392 24968
rect 36434 24928 36474 24968
rect 36516 24928 36556 24968
rect 36598 24928 36638 24968
rect 36680 24928 36720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 44352 24928 44392 24968
rect 44434 24928 44474 24968
rect 44516 24928 44556 24968
rect 44598 24928 44638 24968
rect 44680 24928 44720 24968
rect 48352 24928 48392 24968
rect 48434 24928 48474 24968
rect 48516 24928 48556 24968
rect 48598 24928 48638 24968
rect 48680 24928 48720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 56352 24928 56392 24968
rect 56434 24928 56474 24968
rect 56516 24928 56556 24968
rect 56598 24928 56638 24968
rect 56680 24928 56720 24968
rect 60352 24928 60392 24968
rect 60434 24928 60474 24968
rect 60516 24928 60556 24968
rect 60598 24928 60638 24968
rect 60680 24928 60720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 67948 25600 67988 25640
rect 67756 25264 67796 25304
rect 67564 24844 67604 24884
rect 652 24088 692 24128
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 7112 24172 7152 24212
rect 7194 24172 7234 24212
rect 7276 24172 7316 24212
rect 7358 24172 7398 24212
rect 7440 24172 7480 24212
rect 11112 24172 11152 24212
rect 11194 24172 11234 24212
rect 11276 24172 11316 24212
rect 11358 24172 11398 24212
rect 11440 24172 11480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 19112 24172 19152 24212
rect 19194 24172 19234 24212
rect 19276 24172 19316 24212
rect 19358 24172 19398 24212
rect 19440 24172 19480 24212
rect 23112 24172 23152 24212
rect 23194 24172 23234 24212
rect 23276 24172 23316 24212
rect 23358 24172 23398 24212
rect 23440 24172 23480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 31112 24172 31152 24212
rect 31194 24172 31234 24212
rect 31276 24172 31316 24212
rect 31358 24172 31398 24212
rect 31440 24172 31480 24212
rect 35112 24172 35152 24212
rect 35194 24172 35234 24212
rect 35276 24172 35316 24212
rect 35358 24172 35398 24212
rect 35440 24172 35480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 43112 24172 43152 24212
rect 43194 24172 43234 24212
rect 43276 24172 43316 24212
rect 43358 24172 43398 24212
rect 43440 24172 43480 24212
rect 47112 24172 47152 24212
rect 47194 24172 47234 24212
rect 47276 24172 47316 24212
rect 47358 24172 47398 24212
rect 47440 24172 47480 24212
rect 51112 24172 51152 24212
rect 51194 24172 51234 24212
rect 51276 24172 51316 24212
rect 51358 24172 51398 24212
rect 51440 24172 51480 24212
rect 55112 24172 55152 24212
rect 55194 24172 55234 24212
rect 55276 24172 55316 24212
rect 55358 24172 55398 24212
rect 55440 24172 55480 24212
rect 59112 24172 59152 24212
rect 59194 24172 59234 24212
rect 59276 24172 59316 24212
rect 59358 24172 59398 24212
rect 59440 24172 59480 24212
rect 63112 24172 63152 24212
rect 63194 24172 63234 24212
rect 63276 24172 63316 24212
rect 63358 24172 63398 24212
rect 63440 24172 63480 24212
rect 67112 24172 67152 24212
rect 67194 24172 67234 24212
rect 67276 24172 67316 24212
rect 67358 24172 67398 24212
rect 67440 24172 67480 24212
rect 844 23752 884 23792
rect 652 23248 692 23288
rect 844 23080 884 23120
rect 556 22408 596 22448
rect 2092 23752 2132 23792
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 8352 23416 8392 23456
rect 8434 23416 8474 23456
rect 8516 23416 8556 23456
rect 8598 23416 8638 23456
rect 8680 23416 8720 23456
rect 12352 23416 12392 23456
rect 12434 23416 12474 23456
rect 12516 23416 12556 23456
rect 12598 23416 12638 23456
rect 12680 23416 12720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 20352 23416 20392 23456
rect 20434 23416 20474 23456
rect 20516 23416 20556 23456
rect 20598 23416 20638 23456
rect 20680 23416 20720 23456
rect 24352 23416 24392 23456
rect 24434 23416 24474 23456
rect 24516 23416 24556 23456
rect 24598 23416 24638 23456
rect 24680 23416 24720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 32352 23416 32392 23456
rect 32434 23416 32474 23456
rect 32516 23416 32556 23456
rect 32598 23416 32638 23456
rect 32680 23416 32720 23456
rect 36352 23416 36392 23456
rect 36434 23416 36474 23456
rect 36516 23416 36556 23456
rect 36598 23416 36638 23456
rect 36680 23416 36720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 44352 23416 44392 23456
rect 44434 23416 44474 23456
rect 44516 23416 44556 23456
rect 44598 23416 44638 23456
rect 44680 23416 44720 23456
rect 48352 23416 48392 23456
rect 48434 23416 48474 23456
rect 48516 23416 48556 23456
rect 48598 23416 48638 23456
rect 48680 23416 48720 23456
rect 52352 23416 52392 23456
rect 52434 23416 52474 23456
rect 52516 23416 52556 23456
rect 52598 23416 52638 23456
rect 52680 23416 52720 23456
rect 56352 23416 56392 23456
rect 56434 23416 56474 23456
rect 56516 23416 56556 23456
rect 56598 23416 56638 23456
rect 56680 23416 56720 23456
rect 60352 23416 60392 23456
rect 60434 23416 60474 23456
rect 60516 23416 60556 23456
rect 60598 23416 60638 23456
rect 60680 23416 60720 23456
rect 64352 23416 64392 23456
rect 64434 23416 64474 23456
rect 64516 23416 64556 23456
rect 64598 23416 64638 23456
rect 64680 23416 64720 23456
rect 68352 26440 68392 26480
rect 68434 26440 68474 26480
rect 68516 26440 68556 26480
rect 68598 26440 68638 26480
rect 68680 26440 68720 26480
rect 68620 26104 68660 26144
rect 68812 26104 68852 26144
rect 68332 26020 68372 26060
rect 68812 25936 68852 25976
rect 68524 25600 68564 25640
rect 68332 25348 68372 25388
rect 68620 25264 68660 25304
rect 69292 26104 69332 26144
rect 69484 26104 69524 26144
rect 69100 26020 69140 26060
rect 69196 25768 69236 25808
rect 69004 25684 69044 25724
rect 69388 26020 69428 26060
rect 69580 26020 69620 26060
rect 69580 25852 69620 25892
rect 69772 26104 69812 26144
rect 68908 25096 68948 25136
rect 69484 25264 69524 25304
rect 69868 25516 69908 25556
rect 69964 25432 70004 25472
rect 69772 25180 69812 25220
rect 69292 25012 69332 25052
rect 69676 25012 69716 25052
rect 68352 24928 68392 24968
rect 68434 24928 68474 24968
rect 68516 24928 68556 24968
rect 68598 24928 68638 24968
rect 68680 24928 68720 24968
rect 68352 23416 68392 23456
rect 68434 23416 68474 23456
rect 68516 23416 68556 23456
rect 68598 23416 68638 23456
rect 68680 23416 68720 23456
rect 73900 32068 73940 32108
rect 73612 31984 73652 32024
rect 73228 31732 73268 31772
rect 72415 31480 72455 31520
rect 74668 34588 74708 34628
rect 74476 34252 74516 34292
rect 74284 32908 74324 32948
rect 74860 35092 74900 35132
rect 74860 34504 74900 34544
rect 76780 35680 76820 35720
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 76204 35176 76244 35216
rect 76684 35176 76724 35216
rect 77260 35176 77300 35216
rect 77548 35176 77588 35216
rect 75628 35092 75668 35132
rect 76108 35092 76148 35132
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 75148 34420 75188 34460
rect 74860 34252 74900 34292
rect 75628 34336 75668 34376
rect 74764 32908 74804 32948
rect 74284 31816 74324 31856
rect 72305 31312 72345 31352
rect 72815 31396 72855 31436
rect 73215 31564 73255 31604
rect 73505 31480 73545 31520
rect 74668 32740 74708 32780
rect 74668 31900 74708 31940
rect 75340 32740 75380 32780
rect 75628 32740 75668 32780
rect 76588 35092 76628 35132
rect 76204 34336 76244 34376
rect 77068 35092 77108 35132
rect 75916 34252 75956 34292
rect 75724 31312 75764 31352
rect 76780 34168 76820 34208
rect 77836 35176 77876 35216
rect 76972 34336 77012 34376
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 76684 33832 76724 33872
rect 76684 32488 76724 32528
rect 76015 31312 76055 31352
rect 76815 31480 76855 31520
rect 77356 32488 77396 32528
rect 77836 34336 77876 34376
rect 78220 34336 78260 34376
rect 77548 34252 77588 34292
rect 78316 34168 78356 34208
rect 78700 34336 78740 34376
rect 78604 34168 78644 34208
rect 78988 35092 79028 35132
rect 79112 34756 79152 34796
rect 79194 34756 79234 34796
rect 79276 34756 79316 34796
rect 79358 34756 79398 34796
rect 79440 34756 79480 34796
rect 79276 34252 79316 34292
rect 80140 35008 80180 35048
rect 79756 34336 79796 34376
rect 80352 35512 80392 35552
rect 80434 35512 80474 35552
rect 80516 35512 80556 35552
rect 80598 35512 80638 35552
rect 80680 35512 80720 35552
rect 81580 35092 81620 35132
rect 80428 35008 80468 35048
rect 80620 35008 80660 35048
rect 80908 35008 80948 35048
rect 81388 35008 81428 35048
rect 80236 34672 80276 34712
rect 80716 34672 80756 34712
rect 80332 34168 80372 34208
rect 80352 34000 80392 34040
rect 80434 34000 80474 34040
rect 80516 34000 80556 34040
rect 80598 34000 80638 34040
rect 80680 34000 80720 34040
rect 80428 33832 80468 33872
rect 80332 33748 80372 33788
rect 80236 32740 80276 32780
rect 80716 32740 80756 32780
rect 81004 34420 81044 34460
rect 81004 34252 81044 34292
rect 81196 34420 81236 34460
rect 81484 34420 81524 34460
rect 81292 32740 81332 32780
rect 84352 35512 84392 35552
rect 84434 35512 84474 35552
rect 84516 35512 84556 35552
rect 84598 35512 84638 35552
rect 84680 35512 84720 35552
rect 83884 35176 83924 35216
rect 84268 35176 84308 35216
rect 84652 35176 84692 35216
rect 85228 35680 85268 35720
rect 81772 35092 81812 35132
rect 82348 35092 82388 35132
rect 82636 35092 82676 35132
rect 83308 35092 83348 35132
rect 83500 35092 83540 35132
rect 81676 34336 81716 34376
rect 81868 34420 81908 34460
rect 82252 34504 82292 34544
rect 82156 34336 82196 34376
rect 82060 34084 82100 34124
rect 81868 32740 81908 32780
rect 82305 31564 82345 31604
rect 82636 34504 82676 34544
rect 82732 31732 82772 31772
rect 83112 34756 83152 34796
rect 83194 34756 83234 34796
rect 83276 34756 83316 34796
rect 83358 34756 83398 34796
rect 83440 34756 83480 34796
rect 83308 34588 83348 34628
rect 83596 34588 83636 34628
rect 83116 34420 83156 34460
rect 83116 33832 83156 33872
rect 83500 34000 83540 34040
rect 83505 31564 83545 31604
rect 83884 34588 83924 34628
rect 83884 34168 83924 34208
rect 83788 31564 83828 31604
rect 84172 34588 84212 34628
rect 84652 34504 84692 34544
rect 84076 34168 84116 34208
rect 84172 34084 84212 34124
rect 85036 34588 85076 34628
rect 85036 34420 85076 34460
rect 84748 34336 84788 34376
rect 84364 34168 84404 34208
rect 84352 34000 84392 34040
rect 84434 34000 84474 34040
rect 84516 34000 84556 34040
rect 84598 34000 84638 34040
rect 84680 34000 84720 34040
rect 84940 34168 84980 34208
rect 84705 31564 84745 31604
rect 85228 34504 85268 34544
rect 85420 34504 85460 34544
rect 86092 35092 86132 35132
rect 86380 35092 86420 35132
rect 86572 35092 86612 35132
rect 85804 34504 85844 34544
rect 86188 34168 86228 34208
rect 84940 31564 84980 31604
rect 85215 31480 85255 31520
rect 86476 35008 86516 35048
rect 86668 34924 86708 34964
rect 87628 35176 87668 35216
rect 87052 35092 87092 35132
rect 86860 34588 86900 34628
rect 87436 35092 87476 35132
rect 87916 35008 87956 35048
rect 87244 34924 87284 34964
rect 87112 34756 87152 34796
rect 87194 34756 87234 34796
rect 87276 34756 87316 34796
rect 87358 34756 87398 34796
rect 87440 34756 87480 34796
rect 86764 34168 86804 34208
rect 86815 31480 86855 31520
rect 87215 31564 87255 31604
rect 87724 34924 87764 34964
rect 87628 34000 87668 34040
rect 87820 34420 87860 34460
rect 88352 35512 88392 35552
rect 88434 35512 88474 35552
rect 88516 35512 88556 35552
rect 88598 35512 88638 35552
rect 88680 35512 88720 35552
rect 88108 35176 88148 35216
rect 88492 35176 88532 35216
rect 88684 35092 88724 35132
rect 88300 34924 88340 34964
rect 88108 34420 88148 34460
rect 88300 34420 88340 34460
rect 88684 34420 88724 34460
rect 88352 34000 88392 34040
rect 88434 34000 88474 34040
rect 88516 34000 88556 34040
rect 88598 34000 88638 34040
rect 88680 34000 88720 34040
rect 88300 33832 88340 33872
rect 88204 31564 88244 31604
rect 88415 31564 88455 31604
rect 89356 35008 89396 35048
rect 89164 34336 89204 34376
rect 89068 34168 89108 34208
rect 89932 35260 89972 35300
rect 89932 35092 89972 35132
rect 89452 34336 89492 34376
rect 89644 34336 89684 34376
rect 89356 34252 89396 34292
rect 89548 34168 89588 34208
rect 89932 34337 89972 34376
rect 89932 34336 89972 34337
rect 89505 31396 89545 31436
rect 92428 35680 92468 35720
rect 92352 35512 92392 35552
rect 92434 35512 92474 35552
rect 92516 35512 92556 35552
rect 92598 35512 92638 35552
rect 92680 35512 92720 35552
rect 90220 35092 90260 35132
rect 90682 35129 90722 35132
rect 90682 35092 90722 35129
rect 91084 35092 91124 35132
rect 91468 35092 91508 35132
rect 91756 35092 91796 35132
rect 92236 35092 92276 35132
rect 92428 35092 92468 35132
rect 92620 35092 92660 35132
rect 93100 35092 93140 35132
rect 90220 34840 90260 34880
rect 90220 34504 90260 34544
rect 90316 34168 90356 34208
rect 90604 34420 90644 34460
rect 90604 34168 90644 34208
rect 91112 34756 91152 34796
rect 91194 34756 91234 34796
rect 91276 34756 91316 34796
rect 91358 34756 91398 34796
rect 91440 34756 91480 34796
rect 90988 34252 91028 34292
rect 89905 31480 89945 31520
rect 89740 31396 89780 31436
rect 91180 34420 91220 34460
rect 91468 34420 91508 34460
rect 91756 34420 91796 34460
rect 91105 31480 91145 31520
rect 90988 31396 91028 31436
rect 92044 34336 92084 34376
rect 91948 34168 91988 34208
rect 92236 34336 92276 34376
rect 92620 34504 92660 34544
rect 92812 34336 92852 34376
rect 92812 34168 92852 34208
rect 91372 31480 91412 31520
rect 91615 31396 91655 31436
rect 92352 34000 92392 34040
rect 92434 34000 92474 34040
rect 92516 34000 92556 34040
rect 92598 34000 92638 34040
rect 92680 34000 92720 34040
rect 93100 34420 93140 34460
rect 93100 34168 93140 34208
rect 93580 34420 93620 34460
rect 93580 34252 93620 34292
rect 93484 34168 93524 34208
rect 93868 34420 93908 34460
rect 94060 34420 94100 34460
rect 94252 34336 94292 34376
rect 92415 31480 92455 31520
rect 94636 34420 94676 34460
rect 96352 35512 96392 35552
rect 96434 35512 96474 35552
rect 96516 35512 96556 35552
rect 96598 35512 96638 35552
rect 96680 35512 96720 35552
rect 95212 35092 95252 35132
rect 95404 35092 95444 35132
rect 95884 35092 95924 35132
rect 96172 35092 96212 35132
rect 95116 34924 95156 34964
rect 95112 34756 95152 34796
rect 95194 34756 95234 34796
rect 95276 34756 95316 34796
rect 95358 34756 95398 34796
rect 95440 34756 95480 34796
rect 95020 34252 95060 34292
rect 95596 34336 95636 34376
rect 95788 34924 95828 34964
rect 96172 34924 96212 34964
rect 96076 34420 96116 34460
rect 96268 34336 96308 34376
rect 96460 34420 96500 34460
rect 96940 34924 96980 34964
rect 96844 34504 96884 34544
rect 97804 35092 97844 35132
rect 97132 34504 97172 34544
rect 96748 34336 96788 34376
rect 97036 34336 97076 34376
rect 96652 34168 96692 34208
rect 96940 34084 96980 34124
rect 96352 34000 96392 34040
rect 96434 34000 96474 34040
rect 96516 34000 96556 34040
rect 96598 34000 96638 34040
rect 96680 34000 96720 34040
rect 96844 34000 96884 34040
rect 97516 34420 97556 34460
rect 97804 34420 97844 34460
rect 97900 34336 97940 34376
rect 97900 34168 97940 34208
rect 97996 34000 98036 34040
rect 97505 31564 97545 31604
rect 99112 34756 99152 34796
rect 99194 34756 99234 34796
rect 99276 34756 99316 34796
rect 99358 34756 99398 34796
rect 99440 34756 99480 34796
rect 98284 34336 98324 34376
rect 98860 34336 98900 34376
rect 98956 34168 98996 34208
rect 98188 31564 98228 31604
rect 98305 31564 98345 31604
rect 71884 30808 71924 30848
rect 72305 25852 72345 25892
rect 72415 25768 72455 25808
rect 72705 25768 72745 25808
rect 72844 25684 72884 25724
rect 73228 25516 73268 25556
rect 73036 25264 73076 25304
rect 72352 23416 72392 23456
rect 72434 23416 72474 23456
rect 72516 23416 72556 23456
rect 72598 23416 72638 23456
rect 72680 23416 72720 23456
rect 71788 23332 71828 23372
rect 2092 23248 2132 23288
rect 68236 23248 68276 23288
rect 1996 23080 2036 23120
rect 940 21988 980 22028
rect 652 21568 692 21608
rect 652 20728 692 20768
rect 652 19888 692 19928
rect 652 19048 692 19088
rect 652 18208 692 18248
rect 652 17368 692 17408
rect 652 16528 692 16568
rect 652 15688 692 15728
rect 1996 15436 2036 15476
rect 844 14932 884 14972
rect 1708 14932 1748 14972
rect 652 14848 692 14888
rect 844 14176 884 14216
rect 1324 14176 1364 14216
rect 652 14008 692 14048
rect 844 13336 884 13376
rect 1708 13336 1748 13376
rect 652 13168 692 13208
rect 652 12328 692 12368
rect 844 11908 884 11948
rect 844 11740 884 11780
rect 1612 11740 1652 11780
rect 652 11488 692 11528
rect 1996 11908 2036 11948
rect 1612 10900 1652 10940
rect 844 10816 884 10856
rect 1420 10816 1460 10856
rect 652 10732 692 10772
rect 844 10312 884 10352
rect 1324 10312 1364 10352
rect 1804 10900 1844 10940
rect 652 9808 692 9848
rect 844 9304 884 9344
rect 1324 9304 1364 9344
rect 652 8968 692 9008
rect 844 8800 884 8840
rect 1420 8800 1460 8840
rect 73324 25180 73364 25220
rect 73516 25180 73556 25220
rect 73324 25012 73364 25052
rect 73132 24088 73172 24128
rect 74305 25852 74345 25892
rect 73900 25684 73940 25724
rect 73804 25348 73844 25388
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 7112 22660 7152 22700
rect 7194 22660 7234 22700
rect 7276 22660 7316 22700
rect 7358 22660 7398 22700
rect 7440 22660 7480 22700
rect 11112 22660 11152 22700
rect 11194 22660 11234 22700
rect 11276 22660 11316 22700
rect 11358 22660 11398 22700
rect 11440 22660 11480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 19112 22660 19152 22700
rect 19194 22660 19234 22700
rect 19276 22660 19316 22700
rect 19358 22660 19398 22700
rect 19440 22660 19480 22700
rect 23112 22660 23152 22700
rect 23194 22660 23234 22700
rect 23276 22660 23316 22700
rect 23358 22660 23398 22700
rect 23440 22660 23480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 31112 22660 31152 22700
rect 31194 22660 31234 22700
rect 31276 22660 31316 22700
rect 31358 22660 31398 22700
rect 31440 22660 31480 22700
rect 35112 22660 35152 22700
rect 35194 22660 35234 22700
rect 35276 22660 35316 22700
rect 35358 22660 35398 22700
rect 35440 22660 35480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 43112 22660 43152 22700
rect 43194 22660 43234 22700
rect 43276 22660 43316 22700
rect 43358 22660 43398 22700
rect 43440 22660 43480 22700
rect 47112 22660 47152 22700
rect 47194 22660 47234 22700
rect 47276 22660 47316 22700
rect 47358 22660 47398 22700
rect 47440 22660 47480 22700
rect 51112 22660 51152 22700
rect 51194 22660 51234 22700
rect 51276 22660 51316 22700
rect 51358 22660 51398 22700
rect 51440 22660 51480 22700
rect 55112 22660 55152 22700
rect 55194 22660 55234 22700
rect 55276 22660 55316 22700
rect 55358 22660 55398 22700
rect 55440 22660 55480 22700
rect 59112 22660 59152 22700
rect 59194 22660 59234 22700
rect 59276 22660 59316 22700
rect 59358 22660 59398 22700
rect 59440 22660 59480 22700
rect 63112 22660 63152 22700
rect 63194 22660 63234 22700
rect 63276 22660 63316 22700
rect 63358 22660 63398 22700
rect 63440 22660 63480 22700
rect 67112 22660 67152 22700
rect 67194 22660 67234 22700
rect 67276 22660 67316 22700
rect 67358 22660 67398 22700
rect 67440 22660 67480 22700
rect 71112 22660 71152 22700
rect 71194 22660 71234 22700
rect 71276 22660 71316 22700
rect 71358 22660 71398 22700
rect 71440 22660 71480 22700
rect 74415 25684 74455 25724
rect 73996 25432 74036 25472
rect 74092 25180 74132 25220
rect 74572 22828 74612 22868
rect 75820 25684 75860 25724
rect 74860 24088 74900 24128
rect 75244 24844 75284 24884
rect 75628 25180 75668 25220
rect 75628 23332 75668 23372
rect 74764 22996 74804 23036
rect 75148 22996 75188 23036
rect 75724 22996 75764 23036
rect 75628 22912 75668 22952
rect 75340 22828 75380 22868
rect 75112 22660 75152 22700
rect 75194 22660 75234 22700
rect 75276 22660 75316 22700
rect 75358 22660 75398 22700
rect 75440 22660 75480 22700
rect 75244 22492 75284 22532
rect 75436 22492 75476 22532
rect 74380 22240 74420 22280
rect 75052 22240 75092 22280
rect 76588 25768 76628 25808
rect 76415 25684 76455 25724
rect 75820 22240 75860 22280
rect 75724 22072 75764 22112
rect 9388 21988 9428 22028
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 8352 21904 8392 21944
rect 8434 21904 8474 21944
rect 8516 21904 8556 21944
rect 8598 21904 8638 21944
rect 8680 21904 8720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 7112 21148 7152 21188
rect 7194 21148 7234 21188
rect 7276 21148 7316 21188
rect 7358 21148 7398 21188
rect 7440 21148 7480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 8352 20392 8392 20432
rect 8434 20392 8474 20432
rect 8516 20392 8556 20432
rect 8598 20392 8638 20432
rect 8680 20392 8720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 7112 19636 7152 19676
rect 7194 19636 7234 19676
rect 7276 19636 7316 19676
rect 7358 19636 7398 19676
rect 7440 19636 7480 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 8352 18880 8392 18920
rect 8434 18880 8474 18920
rect 8516 18880 8556 18920
rect 8598 18880 8638 18920
rect 8680 18880 8720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 7112 18124 7152 18164
rect 7194 18124 7234 18164
rect 7276 18124 7316 18164
rect 7358 18124 7398 18164
rect 7440 18124 7480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 8352 17368 8392 17408
rect 8434 17368 8474 17408
rect 8516 17368 8556 17408
rect 8598 17368 8638 17408
rect 8680 17368 8720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 7112 16612 7152 16652
rect 7194 16612 7234 16652
rect 7276 16612 7316 16652
rect 7358 16612 7398 16652
rect 7440 16612 7480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 8352 15856 8392 15896
rect 8434 15856 8474 15896
rect 8516 15856 8556 15896
rect 8598 15856 8638 15896
rect 8680 15856 8720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 7112 15100 7152 15140
rect 7194 15100 7234 15140
rect 7276 15100 7316 15140
rect 7358 15100 7398 15140
rect 7440 15100 7480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 8352 14344 8392 14384
rect 8434 14344 8474 14384
rect 8516 14344 8556 14384
rect 8598 14344 8638 14384
rect 8680 14344 8720 14384
rect 12352 21904 12392 21944
rect 12434 21904 12474 21944
rect 12516 21904 12556 21944
rect 12598 21904 12638 21944
rect 12680 21904 12720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 20352 21904 20392 21944
rect 20434 21904 20474 21944
rect 20516 21904 20556 21944
rect 20598 21904 20638 21944
rect 20680 21904 20720 21944
rect 24352 21904 24392 21944
rect 24434 21904 24474 21944
rect 24516 21904 24556 21944
rect 24598 21904 24638 21944
rect 24680 21904 24720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 32352 21904 32392 21944
rect 32434 21904 32474 21944
rect 32516 21904 32556 21944
rect 32598 21904 32638 21944
rect 32680 21904 32720 21944
rect 36352 21904 36392 21944
rect 36434 21904 36474 21944
rect 36516 21904 36556 21944
rect 36598 21904 36638 21944
rect 36680 21904 36720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 44352 21904 44392 21944
rect 44434 21904 44474 21944
rect 44516 21904 44556 21944
rect 44598 21904 44638 21944
rect 44680 21904 44720 21944
rect 48352 21904 48392 21944
rect 48434 21904 48474 21944
rect 48516 21904 48556 21944
rect 48598 21904 48638 21944
rect 48680 21904 48720 21944
rect 52352 21904 52392 21944
rect 52434 21904 52474 21944
rect 52516 21904 52556 21944
rect 52598 21904 52638 21944
rect 52680 21904 52720 21944
rect 56352 21904 56392 21944
rect 56434 21904 56474 21944
rect 56516 21904 56556 21944
rect 56598 21904 56638 21944
rect 56680 21904 56720 21944
rect 60352 21904 60392 21944
rect 60434 21904 60474 21944
rect 60516 21904 60556 21944
rect 60598 21904 60638 21944
rect 60680 21904 60720 21944
rect 64352 21904 64392 21944
rect 64434 21904 64474 21944
rect 64516 21904 64556 21944
rect 64598 21904 64638 21944
rect 64680 21904 64720 21944
rect 68352 21904 68392 21944
rect 68434 21904 68474 21944
rect 68516 21904 68556 21944
rect 68598 21904 68638 21944
rect 68680 21904 68720 21944
rect 72352 21904 72392 21944
rect 72434 21904 72474 21944
rect 72516 21904 72556 21944
rect 72598 21904 72638 21944
rect 72680 21904 72720 21944
rect 76108 22828 76148 22868
rect 76815 25768 76855 25808
rect 76588 23584 76628 23624
rect 76352 23416 76392 23456
rect 76434 23416 76474 23456
rect 76516 23416 76556 23456
rect 76598 23416 76638 23456
rect 76680 23416 76720 23456
rect 76300 23248 76340 23288
rect 76684 23248 76724 23288
rect 76492 22912 76532 22952
rect 76108 22072 76148 22112
rect 76588 22072 76628 22112
rect 76352 21904 76392 21944
rect 76434 21904 76474 21944
rect 76516 21904 76556 21944
rect 76598 21904 76638 21944
rect 76680 21904 76720 21944
rect 76588 21736 76628 21776
rect 76876 22996 76916 23036
rect 77260 22660 77300 22700
rect 77164 22240 77204 22280
rect 77836 22828 77876 22868
rect 77740 22660 77780 22700
rect 78124 22660 78164 22700
rect 78412 23248 78452 23288
rect 78412 22996 78452 23036
rect 77740 22324 77780 22364
rect 78124 22324 78164 22364
rect 78796 22828 78836 22868
rect 79180 23248 79220 23288
rect 78988 22996 79028 23036
rect 79564 22996 79604 23036
rect 79276 22828 79316 22868
rect 79112 22660 79152 22700
rect 79194 22660 79234 22700
rect 79276 22660 79316 22700
rect 79358 22660 79398 22700
rect 79440 22660 79480 22700
rect 78796 22240 78836 22280
rect 79756 22996 79796 23036
rect 80044 24424 80084 24464
rect 80428 24340 80468 24380
rect 80716 23584 80756 23624
rect 80352 23416 80392 23456
rect 80434 23416 80474 23456
rect 80516 23416 80556 23456
rect 80598 23416 80638 23456
rect 80680 23416 80720 23456
rect 80620 23248 80660 23288
rect 80236 23080 80276 23120
rect 80716 23164 80756 23204
rect 80716 22492 80756 22532
rect 80908 24424 80948 24464
rect 81004 23080 81044 23120
rect 79948 22324 79988 22364
rect 80428 22324 80468 22364
rect 80352 21904 80392 21944
rect 80434 21904 80474 21944
rect 80516 21904 80556 21944
rect 80598 21904 80638 21944
rect 80680 21904 80720 21944
rect 81196 24340 81236 24380
rect 81292 23080 81332 23120
rect 81580 23080 81620 23120
rect 81868 23080 81908 23120
rect 82156 23080 82196 23120
rect 81676 22324 81716 22364
rect 82444 23080 82484 23120
rect 82924 23080 82964 23120
rect 82636 22324 82676 22364
rect 83212 23080 83252 23120
rect 83500 23248 83540 23288
rect 83308 22828 83348 22868
rect 83112 22660 83152 22700
rect 83194 22660 83234 22700
rect 83276 22660 83316 22700
rect 83358 22660 83398 22700
rect 83440 22660 83480 22700
rect 83596 22660 83636 22700
rect 83788 23164 83828 23204
rect 83788 22660 83828 22700
rect 84705 25684 84745 25724
rect 84940 25684 84980 25724
rect 84268 23752 84308 23792
rect 84352 23416 84392 23456
rect 84434 23416 84474 23456
rect 84516 23416 84556 23456
rect 84598 23416 84638 23456
rect 84680 23416 84720 23456
rect 84076 23080 84116 23120
rect 83980 22996 84020 23036
rect 83980 22828 84020 22868
rect 83596 22324 83636 22364
rect 83788 22324 83828 22364
rect 84364 23080 84404 23120
rect 84748 23080 84788 23120
rect 84268 22996 84308 23036
rect 85420 23920 85460 23960
rect 85804 23164 85844 23204
rect 85132 23080 85172 23120
rect 85420 23080 85460 23120
rect 85708 22996 85748 23036
rect 85420 22492 85460 22532
rect 85900 22660 85940 22700
rect 86092 22660 86132 22700
rect 84556 22324 84596 22364
rect 84940 22324 84980 22364
rect 85612 22324 85652 22364
rect 85804 22324 85844 22364
rect 84352 21904 84392 21944
rect 84434 21904 84474 21944
rect 84516 21904 84556 21944
rect 84598 21904 84638 21944
rect 84680 21904 84720 21944
rect 84364 21736 84404 21776
rect 86284 22996 86324 23036
rect 87215 25684 87255 25724
rect 86668 23080 86708 23120
rect 86476 22912 86516 22952
rect 86572 22660 86612 22700
rect 86380 22324 86420 22364
rect 86284 22240 86324 22280
rect 86668 22408 86708 22448
rect 86572 22324 86612 22364
rect 87724 25684 87764 25724
rect 87340 22828 87380 22868
rect 87532 22996 87572 23036
rect 86956 22660 86996 22700
rect 87112 22660 87152 22700
rect 87194 22660 87234 22700
rect 87276 22660 87316 22700
rect 87358 22660 87398 22700
rect 87440 22660 87480 22700
rect 87052 22492 87092 22532
rect 87724 22996 87764 23036
rect 87628 22492 87668 22532
rect 86956 22240 86996 22280
rect 87628 22324 87668 22364
rect 87820 22828 87860 22868
rect 88108 22828 88148 22868
rect 88396 23584 88436 23624
rect 88352 23416 88392 23456
rect 88434 23416 88474 23456
rect 88516 23416 88556 23456
rect 88598 23416 88638 23456
rect 88680 23416 88720 23456
rect 88396 23248 88436 23288
rect 88492 22828 88532 22868
rect 88780 22828 88820 22868
rect 87724 22240 87764 22280
rect 88396 22324 88436 22364
rect 88876 22324 88916 22364
rect 87244 22156 87284 22196
rect 88012 22156 88052 22196
rect 88352 21904 88392 21944
rect 88434 21904 88474 21944
rect 88516 21904 88556 21944
rect 88598 21904 88638 21944
rect 88680 21904 88720 21944
rect 89356 23248 89396 23288
rect 89452 23080 89492 23120
rect 89356 22492 89396 22532
rect 90015 25684 90055 25724
rect 90508 25684 90548 25724
rect 89644 23248 89684 23288
rect 89836 23080 89876 23120
rect 89740 22492 89780 22532
rect 90124 22492 90164 22532
rect 90412 23920 90452 23960
rect 91905 25852 91945 25892
rect 90796 23836 90836 23876
rect 90508 23080 90548 23120
rect 90316 22996 90356 23036
rect 90316 22828 90356 22868
rect 90604 22492 90644 22532
rect 91180 23248 91220 23288
rect 90892 23080 90932 23120
rect 91180 23080 91220 23120
rect 91372 25180 91412 25220
rect 90892 22828 90932 22868
rect 91372 22828 91412 22868
rect 90508 22324 90548 22364
rect 91112 22660 91152 22700
rect 91194 22660 91234 22700
rect 91276 22660 91316 22700
rect 91358 22660 91398 22700
rect 91440 22660 91480 22700
rect 90988 22324 91028 22364
rect 91084 22240 91124 22280
rect 91276 22492 91316 22532
rect 91756 23248 91796 23288
rect 91660 23164 91700 23204
rect 91852 22996 91892 23036
rect 91852 22408 91892 22448
rect 92140 25852 92180 25892
rect 92044 25180 92084 25220
rect 92044 22996 92084 23036
rect 92428 24004 92468 24044
rect 92352 23416 92392 23456
rect 92434 23416 92474 23456
rect 92516 23416 92556 23456
rect 92598 23416 92638 23456
rect 92680 23416 92720 23456
rect 92236 22576 92276 22616
rect 92620 22660 92660 22700
rect 92524 22576 92564 22616
rect 92236 22324 92276 22364
rect 92908 22660 92948 22700
rect 93100 22660 93140 22700
rect 93292 22660 93332 22700
rect 91948 22240 91988 22280
rect 92620 22072 92660 22112
rect 92352 21904 92392 21944
rect 92434 21904 92474 21944
rect 92516 21904 92556 21944
rect 92598 21904 92638 21944
rect 92680 21904 92720 21944
rect 93580 23836 93620 23876
rect 93676 23248 93716 23288
rect 93484 22996 93524 23036
rect 93772 22660 93812 22700
rect 93484 22492 93524 22532
rect 93964 23248 94004 23288
rect 94060 22660 94100 22700
rect 94444 22660 94484 22700
rect 93772 22324 93812 22364
rect 95105 25768 95145 25808
rect 95215 25684 95255 25724
rect 95404 24676 95444 24716
rect 95308 23080 95348 23120
rect 95112 22660 95152 22700
rect 95194 22660 95234 22700
rect 95276 22660 95316 22700
rect 95358 22660 95398 22700
rect 95440 22660 95480 22700
rect 95404 22492 95444 22532
rect 95692 24676 95732 24716
rect 95692 23080 95732 23120
rect 95692 22912 95732 22952
rect 95116 22408 95156 22448
rect 95308 22408 95348 22448
rect 94924 22324 94964 22364
rect 93484 22072 93524 22112
rect 77548 21484 77588 21524
rect 77740 21484 77780 21524
rect 78892 21484 78932 21524
rect 79276 21484 79316 21524
rect 80812 21484 80852 21524
rect 82156 21484 82196 21524
rect 82636 21484 82676 21524
rect 83404 21484 83444 21524
rect 83788 21484 83828 21524
rect 84172 21484 84212 21524
rect 92716 21568 92756 21608
rect 95212 21736 95252 21776
rect 93388 21568 93428 21608
rect 95884 22660 95924 22700
rect 96076 23248 96116 23288
rect 96076 22492 96116 22532
rect 96352 23416 96392 23456
rect 96434 23416 96474 23456
rect 96516 23416 96556 23456
rect 96598 23416 96638 23456
rect 96680 23416 96720 23456
rect 96460 23248 96500 23288
rect 96556 22912 96596 22952
rect 96844 22912 96884 22952
rect 96364 22660 96404 22700
rect 95788 22408 95828 22448
rect 95692 22324 95732 22364
rect 96076 22324 96116 22364
rect 96364 22324 96404 22364
rect 97132 22912 97172 22952
rect 97420 22912 97460 22952
rect 97804 23080 97844 23120
rect 97804 22912 97844 22952
rect 97228 22324 97268 22364
rect 99244 31564 99284 31604
rect 99148 25432 99188 25472
rect 98188 23080 98228 23120
rect 99112 22660 99152 22700
rect 99194 22660 99234 22700
rect 99276 22660 99316 22700
rect 99358 22660 99398 22700
rect 99440 22660 99480 22700
rect 98188 22324 98228 22364
rect 96352 21904 96392 21944
rect 96434 21904 96474 21944
rect 96516 21904 96556 21944
rect 96598 21904 96638 21944
rect 96680 21904 96720 21944
rect 11112 21148 11152 21188
rect 11194 21148 11234 21188
rect 11276 21148 11316 21188
rect 11358 21148 11398 21188
rect 11440 21148 11480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 19112 21148 19152 21188
rect 19194 21148 19234 21188
rect 19276 21148 19316 21188
rect 19358 21148 19398 21188
rect 19440 21148 19480 21188
rect 23112 21148 23152 21188
rect 23194 21148 23234 21188
rect 23276 21148 23316 21188
rect 23358 21148 23398 21188
rect 23440 21148 23480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 31112 21148 31152 21188
rect 31194 21148 31234 21188
rect 31276 21148 31316 21188
rect 31358 21148 31398 21188
rect 31440 21148 31480 21188
rect 35112 21148 35152 21188
rect 35194 21148 35234 21188
rect 35276 21148 35316 21188
rect 35358 21148 35398 21188
rect 35440 21148 35480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 43112 21148 43152 21188
rect 43194 21148 43234 21188
rect 43276 21148 43316 21188
rect 43358 21148 43398 21188
rect 43440 21148 43480 21188
rect 47112 21148 47152 21188
rect 47194 21148 47234 21188
rect 47276 21148 47316 21188
rect 47358 21148 47398 21188
rect 47440 21148 47480 21188
rect 51112 21148 51152 21188
rect 51194 21148 51234 21188
rect 51276 21148 51316 21188
rect 51358 21148 51398 21188
rect 51440 21148 51480 21188
rect 55112 21148 55152 21188
rect 55194 21148 55234 21188
rect 55276 21148 55316 21188
rect 55358 21148 55398 21188
rect 55440 21148 55480 21188
rect 59112 21148 59152 21188
rect 59194 21148 59234 21188
rect 59276 21148 59316 21188
rect 59358 21148 59398 21188
rect 59440 21148 59480 21188
rect 63112 21148 63152 21188
rect 63194 21148 63234 21188
rect 63276 21148 63316 21188
rect 63358 21148 63398 21188
rect 63440 21148 63480 21188
rect 67112 21148 67152 21188
rect 67194 21148 67234 21188
rect 67276 21148 67316 21188
rect 67358 21148 67398 21188
rect 67440 21148 67480 21188
rect 71112 21148 71152 21188
rect 71194 21148 71234 21188
rect 71276 21148 71316 21188
rect 71358 21148 71398 21188
rect 71440 21148 71480 21188
rect 75112 21148 75152 21188
rect 75194 21148 75234 21188
rect 75276 21148 75316 21188
rect 75358 21148 75398 21188
rect 75440 21148 75480 21188
rect 79112 21148 79152 21188
rect 79194 21148 79234 21188
rect 79276 21148 79316 21188
rect 79358 21148 79398 21188
rect 79440 21148 79480 21188
rect 83112 21148 83152 21188
rect 83194 21148 83234 21188
rect 83276 21148 83316 21188
rect 83358 21148 83398 21188
rect 83440 21148 83480 21188
rect 87112 21148 87152 21188
rect 87194 21148 87234 21188
rect 87276 21148 87316 21188
rect 87358 21148 87398 21188
rect 87440 21148 87480 21188
rect 91112 21148 91152 21188
rect 91194 21148 91234 21188
rect 91276 21148 91316 21188
rect 91358 21148 91398 21188
rect 91440 21148 91480 21188
rect 95112 21148 95152 21188
rect 95194 21148 95234 21188
rect 95276 21148 95316 21188
rect 95358 21148 95398 21188
rect 95440 21148 95480 21188
rect 99112 21148 99152 21188
rect 99194 21148 99234 21188
rect 99276 21148 99316 21188
rect 99358 21148 99398 21188
rect 99440 21148 99480 21188
rect 12352 20392 12392 20432
rect 12434 20392 12474 20432
rect 12516 20392 12556 20432
rect 12598 20392 12638 20432
rect 12680 20392 12720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 20352 20392 20392 20432
rect 20434 20392 20474 20432
rect 20516 20392 20556 20432
rect 20598 20392 20638 20432
rect 20680 20392 20720 20432
rect 24352 20392 24392 20432
rect 24434 20392 24474 20432
rect 24516 20392 24556 20432
rect 24598 20392 24638 20432
rect 24680 20392 24720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 32352 20392 32392 20432
rect 32434 20392 32474 20432
rect 32516 20392 32556 20432
rect 32598 20392 32638 20432
rect 32680 20392 32720 20432
rect 36352 20392 36392 20432
rect 36434 20392 36474 20432
rect 36516 20392 36556 20432
rect 36598 20392 36638 20432
rect 36680 20392 36720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 44352 20392 44392 20432
rect 44434 20392 44474 20432
rect 44516 20392 44556 20432
rect 44598 20392 44638 20432
rect 44680 20392 44720 20432
rect 48352 20392 48392 20432
rect 48434 20392 48474 20432
rect 48516 20392 48556 20432
rect 48598 20392 48638 20432
rect 48680 20392 48720 20432
rect 52352 20392 52392 20432
rect 52434 20392 52474 20432
rect 52516 20392 52556 20432
rect 52598 20392 52638 20432
rect 52680 20392 52720 20432
rect 56352 20392 56392 20432
rect 56434 20392 56474 20432
rect 56516 20392 56556 20432
rect 56598 20392 56638 20432
rect 56680 20392 56720 20432
rect 60352 20392 60392 20432
rect 60434 20392 60474 20432
rect 60516 20392 60556 20432
rect 60598 20392 60638 20432
rect 60680 20392 60720 20432
rect 64352 20392 64392 20432
rect 64434 20392 64474 20432
rect 64516 20392 64556 20432
rect 64598 20392 64638 20432
rect 64680 20392 64720 20432
rect 68352 20392 68392 20432
rect 68434 20392 68474 20432
rect 68516 20392 68556 20432
rect 68598 20392 68638 20432
rect 68680 20392 68720 20432
rect 72352 20392 72392 20432
rect 72434 20392 72474 20432
rect 72516 20392 72556 20432
rect 72598 20392 72638 20432
rect 72680 20392 72720 20432
rect 76352 20392 76392 20432
rect 76434 20392 76474 20432
rect 76516 20392 76556 20432
rect 76598 20392 76638 20432
rect 76680 20392 76720 20432
rect 80352 20392 80392 20432
rect 80434 20392 80474 20432
rect 80516 20392 80556 20432
rect 80598 20392 80638 20432
rect 80680 20392 80720 20432
rect 84352 20392 84392 20432
rect 84434 20392 84474 20432
rect 84516 20392 84556 20432
rect 84598 20392 84638 20432
rect 84680 20392 84720 20432
rect 88352 20392 88392 20432
rect 88434 20392 88474 20432
rect 88516 20392 88556 20432
rect 88598 20392 88638 20432
rect 88680 20392 88720 20432
rect 92352 20392 92392 20432
rect 92434 20392 92474 20432
rect 92516 20392 92556 20432
rect 92598 20392 92638 20432
rect 92680 20392 92720 20432
rect 96352 20392 96392 20432
rect 96434 20392 96474 20432
rect 96516 20392 96556 20432
rect 96598 20392 96638 20432
rect 96680 20392 96720 20432
rect 11112 19636 11152 19676
rect 11194 19636 11234 19676
rect 11276 19636 11316 19676
rect 11358 19636 11398 19676
rect 11440 19636 11480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 19112 19636 19152 19676
rect 19194 19636 19234 19676
rect 19276 19636 19316 19676
rect 19358 19636 19398 19676
rect 19440 19636 19480 19676
rect 23112 19636 23152 19676
rect 23194 19636 23234 19676
rect 23276 19636 23316 19676
rect 23358 19636 23398 19676
rect 23440 19636 23480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 31112 19636 31152 19676
rect 31194 19636 31234 19676
rect 31276 19636 31316 19676
rect 31358 19636 31398 19676
rect 31440 19636 31480 19676
rect 35112 19636 35152 19676
rect 35194 19636 35234 19676
rect 35276 19636 35316 19676
rect 35358 19636 35398 19676
rect 35440 19636 35480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 43112 19636 43152 19676
rect 43194 19636 43234 19676
rect 43276 19636 43316 19676
rect 43358 19636 43398 19676
rect 43440 19636 43480 19676
rect 47112 19636 47152 19676
rect 47194 19636 47234 19676
rect 47276 19636 47316 19676
rect 47358 19636 47398 19676
rect 47440 19636 47480 19676
rect 51112 19636 51152 19676
rect 51194 19636 51234 19676
rect 51276 19636 51316 19676
rect 51358 19636 51398 19676
rect 51440 19636 51480 19676
rect 55112 19636 55152 19676
rect 55194 19636 55234 19676
rect 55276 19636 55316 19676
rect 55358 19636 55398 19676
rect 55440 19636 55480 19676
rect 59112 19636 59152 19676
rect 59194 19636 59234 19676
rect 59276 19636 59316 19676
rect 59358 19636 59398 19676
rect 59440 19636 59480 19676
rect 63112 19636 63152 19676
rect 63194 19636 63234 19676
rect 63276 19636 63316 19676
rect 63358 19636 63398 19676
rect 63440 19636 63480 19676
rect 67112 19636 67152 19676
rect 67194 19636 67234 19676
rect 67276 19636 67316 19676
rect 67358 19636 67398 19676
rect 67440 19636 67480 19676
rect 71112 19636 71152 19676
rect 71194 19636 71234 19676
rect 71276 19636 71316 19676
rect 71358 19636 71398 19676
rect 71440 19636 71480 19676
rect 75112 19636 75152 19676
rect 75194 19636 75234 19676
rect 75276 19636 75316 19676
rect 75358 19636 75398 19676
rect 75440 19636 75480 19676
rect 71788 19216 71828 19256
rect 12352 18880 12392 18920
rect 12434 18880 12474 18920
rect 12516 18880 12556 18920
rect 12598 18880 12638 18920
rect 12680 18880 12720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 20352 18880 20392 18920
rect 20434 18880 20474 18920
rect 20516 18880 20556 18920
rect 20598 18880 20638 18920
rect 20680 18880 20720 18920
rect 24352 18880 24392 18920
rect 24434 18880 24474 18920
rect 24516 18880 24556 18920
rect 24598 18880 24638 18920
rect 24680 18880 24720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 32352 18880 32392 18920
rect 32434 18880 32474 18920
rect 32516 18880 32556 18920
rect 32598 18880 32638 18920
rect 32680 18880 32720 18920
rect 36352 18880 36392 18920
rect 36434 18880 36474 18920
rect 36516 18880 36556 18920
rect 36598 18880 36638 18920
rect 36680 18880 36720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 44352 18880 44392 18920
rect 44434 18880 44474 18920
rect 44516 18880 44556 18920
rect 44598 18880 44638 18920
rect 44680 18880 44720 18920
rect 48352 18880 48392 18920
rect 48434 18880 48474 18920
rect 48516 18880 48556 18920
rect 48598 18880 48638 18920
rect 48680 18880 48720 18920
rect 52352 18880 52392 18920
rect 52434 18880 52474 18920
rect 52516 18880 52556 18920
rect 52598 18880 52638 18920
rect 52680 18880 52720 18920
rect 56352 18880 56392 18920
rect 56434 18880 56474 18920
rect 56516 18880 56556 18920
rect 56598 18880 56638 18920
rect 56680 18880 56720 18920
rect 60352 18880 60392 18920
rect 60434 18880 60474 18920
rect 60516 18880 60556 18920
rect 60598 18880 60638 18920
rect 60680 18880 60720 18920
rect 64352 18880 64392 18920
rect 64434 18880 64474 18920
rect 64516 18880 64556 18920
rect 64598 18880 64638 18920
rect 64680 18880 64720 18920
rect 68352 18880 68392 18920
rect 68434 18880 68474 18920
rect 68516 18880 68556 18920
rect 68598 18880 68638 18920
rect 68680 18880 68720 18920
rect 68236 18544 68276 18584
rect 11112 18124 11152 18164
rect 11194 18124 11234 18164
rect 11276 18124 11316 18164
rect 11358 18124 11398 18164
rect 11440 18124 11480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 19112 18124 19152 18164
rect 19194 18124 19234 18164
rect 19276 18124 19316 18164
rect 19358 18124 19398 18164
rect 19440 18124 19480 18164
rect 23112 18124 23152 18164
rect 23194 18124 23234 18164
rect 23276 18124 23316 18164
rect 23358 18124 23398 18164
rect 23440 18124 23480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 31112 18124 31152 18164
rect 31194 18124 31234 18164
rect 31276 18124 31316 18164
rect 31358 18124 31398 18164
rect 31440 18124 31480 18164
rect 35112 18124 35152 18164
rect 35194 18124 35234 18164
rect 35276 18124 35316 18164
rect 35358 18124 35398 18164
rect 35440 18124 35480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 43112 18124 43152 18164
rect 43194 18124 43234 18164
rect 43276 18124 43316 18164
rect 43358 18124 43398 18164
rect 43440 18124 43480 18164
rect 47112 18124 47152 18164
rect 47194 18124 47234 18164
rect 47276 18124 47316 18164
rect 47358 18124 47398 18164
rect 47440 18124 47480 18164
rect 51112 18124 51152 18164
rect 51194 18124 51234 18164
rect 51276 18124 51316 18164
rect 51358 18124 51398 18164
rect 51440 18124 51480 18164
rect 55112 18124 55152 18164
rect 55194 18124 55234 18164
rect 55276 18124 55316 18164
rect 55358 18124 55398 18164
rect 55440 18124 55480 18164
rect 59112 18124 59152 18164
rect 59194 18124 59234 18164
rect 59276 18124 59316 18164
rect 59358 18124 59398 18164
rect 59440 18124 59480 18164
rect 63112 18124 63152 18164
rect 63194 18124 63234 18164
rect 63276 18124 63316 18164
rect 63358 18124 63398 18164
rect 63440 18124 63480 18164
rect 67112 18124 67152 18164
rect 67194 18124 67234 18164
rect 67276 18124 67316 18164
rect 67358 18124 67398 18164
rect 67440 18124 67480 18164
rect 12352 17368 12392 17408
rect 12434 17368 12474 17408
rect 12516 17368 12556 17408
rect 12598 17368 12638 17408
rect 12680 17368 12720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 20352 17368 20392 17408
rect 20434 17368 20474 17408
rect 20516 17368 20556 17408
rect 20598 17368 20638 17408
rect 20680 17368 20720 17408
rect 24352 17368 24392 17408
rect 24434 17368 24474 17408
rect 24516 17368 24556 17408
rect 24598 17368 24638 17408
rect 24680 17368 24720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 32352 17368 32392 17408
rect 32434 17368 32474 17408
rect 32516 17368 32556 17408
rect 32598 17368 32638 17408
rect 32680 17368 32720 17408
rect 36352 17368 36392 17408
rect 36434 17368 36474 17408
rect 36516 17368 36556 17408
rect 36598 17368 36638 17408
rect 36680 17368 36720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 44352 17368 44392 17408
rect 44434 17368 44474 17408
rect 44516 17368 44556 17408
rect 44598 17368 44638 17408
rect 44680 17368 44720 17408
rect 48352 17368 48392 17408
rect 48434 17368 48474 17408
rect 48516 17368 48556 17408
rect 48598 17368 48638 17408
rect 48680 17368 48720 17408
rect 52352 17368 52392 17408
rect 52434 17368 52474 17408
rect 52516 17368 52556 17408
rect 52598 17368 52638 17408
rect 52680 17368 52720 17408
rect 56352 17368 56392 17408
rect 56434 17368 56474 17408
rect 56516 17368 56556 17408
rect 56598 17368 56638 17408
rect 56680 17368 56720 17408
rect 60352 17368 60392 17408
rect 60434 17368 60474 17408
rect 60516 17368 60556 17408
rect 60598 17368 60638 17408
rect 60680 17368 60720 17408
rect 64352 17368 64392 17408
rect 64434 17368 64474 17408
rect 64516 17368 64556 17408
rect 64598 17368 64638 17408
rect 64680 17368 64720 17408
rect 11112 16612 11152 16652
rect 11194 16612 11234 16652
rect 11276 16612 11316 16652
rect 11358 16612 11398 16652
rect 11440 16612 11480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 19112 16612 19152 16652
rect 19194 16612 19234 16652
rect 19276 16612 19316 16652
rect 19358 16612 19398 16652
rect 19440 16612 19480 16652
rect 23112 16612 23152 16652
rect 23194 16612 23234 16652
rect 23276 16612 23316 16652
rect 23358 16612 23398 16652
rect 23440 16612 23480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 31112 16612 31152 16652
rect 31194 16612 31234 16652
rect 31276 16612 31316 16652
rect 31358 16612 31398 16652
rect 31440 16612 31480 16652
rect 35112 16612 35152 16652
rect 35194 16612 35234 16652
rect 35276 16612 35316 16652
rect 35358 16612 35398 16652
rect 35440 16612 35480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 43112 16612 43152 16652
rect 43194 16612 43234 16652
rect 43276 16612 43316 16652
rect 43358 16612 43398 16652
rect 43440 16612 43480 16652
rect 47112 16612 47152 16652
rect 47194 16612 47234 16652
rect 47276 16612 47316 16652
rect 47358 16612 47398 16652
rect 47440 16612 47480 16652
rect 51112 16612 51152 16652
rect 51194 16612 51234 16652
rect 51276 16612 51316 16652
rect 51358 16612 51398 16652
rect 51440 16612 51480 16652
rect 55112 16612 55152 16652
rect 55194 16612 55234 16652
rect 55276 16612 55316 16652
rect 55358 16612 55398 16652
rect 55440 16612 55480 16652
rect 59112 16612 59152 16652
rect 59194 16612 59234 16652
rect 59276 16612 59316 16652
rect 59358 16612 59398 16652
rect 59440 16612 59480 16652
rect 63112 16612 63152 16652
rect 63194 16612 63234 16652
rect 63276 16612 63316 16652
rect 63358 16612 63398 16652
rect 63440 16612 63480 16652
rect 67112 16612 67152 16652
rect 67194 16612 67234 16652
rect 67276 16612 67316 16652
rect 67358 16612 67398 16652
rect 67440 16612 67480 16652
rect 67372 15940 67412 15980
rect 12352 15856 12392 15896
rect 12434 15856 12474 15896
rect 12516 15856 12556 15896
rect 12598 15856 12638 15896
rect 12680 15856 12720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 20352 15856 20392 15896
rect 20434 15856 20474 15896
rect 20516 15856 20556 15896
rect 20598 15856 20638 15896
rect 20680 15856 20720 15896
rect 24352 15856 24392 15896
rect 24434 15856 24474 15896
rect 24516 15856 24556 15896
rect 24598 15856 24638 15896
rect 24680 15856 24720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 32352 15856 32392 15896
rect 32434 15856 32474 15896
rect 32516 15856 32556 15896
rect 32598 15856 32638 15896
rect 32680 15856 32720 15896
rect 36352 15856 36392 15896
rect 36434 15856 36474 15896
rect 36516 15856 36556 15896
rect 36598 15856 36638 15896
rect 36680 15856 36720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 44352 15856 44392 15896
rect 44434 15856 44474 15896
rect 44516 15856 44556 15896
rect 44598 15856 44638 15896
rect 44680 15856 44720 15896
rect 48352 15856 48392 15896
rect 48434 15856 48474 15896
rect 48516 15856 48556 15896
rect 48598 15856 48638 15896
rect 48680 15856 48720 15896
rect 52352 15856 52392 15896
rect 52434 15856 52474 15896
rect 52516 15856 52556 15896
rect 52598 15856 52638 15896
rect 52680 15856 52720 15896
rect 56352 15856 56392 15896
rect 56434 15856 56474 15896
rect 56516 15856 56556 15896
rect 56598 15856 56638 15896
rect 56680 15856 56720 15896
rect 60352 15856 60392 15896
rect 60434 15856 60474 15896
rect 60516 15856 60556 15896
rect 60598 15856 60638 15896
rect 60680 15856 60720 15896
rect 64352 15856 64392 15896
rect 64434 15856 64474 15896
rect 64516 15856 64556 15896
rect 64598 15856 64638 15896
rect 64680 15856 64720 15896
rect 67180 15520 67220 15560
rect 67564 15520 67604 15560
rect 71112 18124 71152 18164
rect 71194 18124 71234 18164
rect 71276 18124 71316 18164
rect 71358 18124 71398 18164
rect 71440 18124 71480 18164
rect 68352 17368 68392 17408
rect 68434 17368 68474 17408
rect 68516 17368 68556 17408
rect 68598 17368 68638 17408
rect 68680 17368 68720 17408
rect 68352 15856 68392 15896
rect 68434 15856 68474 15896
rect 68516 15856 68556 15896
rect 68598 15856 68638 15896
rect 68680 15856 68720 15896
rect 68812 15856 68852 15896
rect 67756 15436 67796 15476
rect 11112 15100 11152 15140
rect 11194 15100 11234 15140
rect 11276 15100 11316 15140
rect 11358 15100 11398 15140
rect 11440 15100 11480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 19112 15100 19152 15140
rect 19194 15100 19234 15140
rect 19276 15100 19316 15140
rect 19358 15100 19398 15140
rect 19440 15100 19480 15140
rect 23112 15100 23152 15140
rect 23194 15100 23234 15140
rect 23276 15100 23316 15140
rect 23358 15100 23398 15140
rect 23440 15100 23480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 31112 15100 31152 15140
rect 31194 15100 31234 15140
rect 31276 15100 31316 15140
rect 31358 15100 31398 15140
rect 31440 15100 31480 15140
rect 35112 15100 35152 15140
rect 35194 15100 35234 15140
rect 35276 15100 35316 15140
rect 35358 15100 35398 15140
rect 35440 15100 35480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 43112 15100 43152 15140
rect 43194 15100 43234 15140
rect 43276 15100 43316 15140
rect 43358 15100 43398 15140
rect 43440 15100 43480 15140
rect 47112 15100 47152 15140
rect 47194 15100 47234 15140
rect 47276 15100 47316 15140
rect 47358 15100 47398 15140
rect 47440 15100 47480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 55112 15100 55152 15140
rect 55194 15100 55234 15140
rect 55276 15100 55316 15140
rect 55358 15100 55398 15140
rect 55440 15100 55480 15140
rect 59112 15100 59152 15140
rect 59194 15100 59234 15140
rect 59276 15100 59316 15140
rect 59358 15100 59398 15140
rect 59440 15100 59480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 67112 15100 67152 15140
rect 67194 15100 67234 15140
rect 67276 15100 67316 15140
rect 67358 15100 67398 15140
rect 67440 15100 67480 15140
rect 12352 14344 12392 14384
rect 12434 14344 12474 14384
rect 12516 14344 12556 14384
rect 12598 14344 12638 14384
rect 12680 14344 12720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 20352 14344 20392 14384
rect 20434 14344 20474 14384
rect 20516 14344 20556 14384
rect 20598 14344 20638 14384
rect 20680 14344 20720 14384
rect 24352 14344 24392 14384
rect 24434 14344 24474 14384
rect 24516 14344 24556 14384
rect 24598 14344 24638 14384
rect 24680 14344 24720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 32352 14344 32392 14384
rect 32434 14344 32474 14384
rect 32516 14344 32556 14384
rect 32598 14344 32638 14384
rect 32680 14344 32720 14384
rect 36352 14344 36392 14384
rect 36434 14344 36474 14384
rect 36516 14344 36556 14384
rect 36598 14344 36638 14384
rect 36680 14344 36720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 44352 14344 44392 14384
rect 44434 14344 44474 14384
rect 44516 14344 44556 14384
rect 44598 14344 44638 14384
rect 44680 14344 44720 14384
rect 48352 14344 48392 14384
rect 48434 14344 48474 14384
rect 48516 14344 48556 14384
rect 48598 14344 48638 14384
rect 48680 14344 48720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 56352 14344 56392 14384
rect 56434 14344 56474 14384
rect 56516 14344 56556 14384
rect 56598 14344 56638 14384
rect 56680 14344 56720 14384
rect 60352 14344 60392 14384
rect 60434 14344 60474 14384
rect 60516 14344 60556 14384
rect 60598 14344 60638 14384
rect 60680 14344 60720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 9388 13924 9428 13964
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 7112 13588 7152 13628
rect 7194 13588 7234 13628
rect 7276 13588 7316 13628
rect 7358 13588 7398 13628
rect 7440 13588 7480 13628
rect 11112 13588 11152 13628
rect 11194 13588 11234 13628
rect 11276 13588 11316 13628
rect 11358 13588 11398 13628
rect 11440 13588 11480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 19112 13588 19152 13628
rect 19194 13588 19234 13628
rect 19276 13588 19316 13628
rect 19358 13588 19398 13628
rect 19440 13588 19480 13628
rect 23112 13588 23152 13628
rect 23194 13588 23234 13628
rect 23276 13588 23316 13628
rect 23358 13588 23398 13628
rect 23440 13588 23480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 31112 13588 31152 13628
rect 31194 13588 31234 13628
rect 31276 13588 31316 13628
rect 31358 13588 31398 13628
rect 31440 13588 31480 13628
rect 35112 13588 35152 13628
rect 35194 13588 35234 13628
rect 35276 13588 35316 13628
rect 35358 13588 35398 13628
rect 35440 13588 35480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 43112 13588 43152 13628
rect 43194 13588 43234 13628
rect 43276 13588 43316 13628
rect 43358 13588 43398 13628
rect 43440 13588 43480 13628
rect 47112 13588 47152 13628
rect 47194 13588 47234 13628
rect 47276 13588 47316 13628
rect 47358 13588 47398 13628
rect 47440 13588 47480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 55112 13588 55152 13628
rect 55194 13588 55234 13628
rect 55276 13588 55316 13628
rect 55358 13588 55398 13628
rect 55440 13588 55480 13628
rect 59112 13588 59152 13628
rect 59194 13588 59234 13628
rect 59276 13588 59316 13628
rect 59358 13588 59398 13628
rect 59440 13588 59480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 67112 13588 67152 13628
rect 67194 13588 67234 13628
rect 67276 13588 67316 13628
rect 67358 13588 67398 13628
rect 67440 13588 67480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 8352 12832 8392 12872
rect 8434 12832 8474 12872
rect 8516 12832 8556 12872
rect 8598 12832 8638 12872
rect 8680 12832 8720 12872
rect 12352 12832 12392 12872
rect 12434 12832 12474 12872
rect 12516 12832 12556 12872
rect 12598 12832 12638 12872
rect 12680 12832 12720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 20352 12832 20392 12872
rect 20434 12832 20474 12872
rect 20516 12832 20556 12872
rect 20598 12832 20638 12872
rect 20680 12832 20720 12872
rect 24352 12832 24392 12872
rect 24434 12832 24474 12872
rect 24516 12832 24556 12872
rect 24598 12832 24638 12872
rect 24680 12832 24720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 32352 12832 32392 12872
rect 32434 12832 32474 12872
rect 32516 12832 32556 12872
rect 32598 12832 32638 12872
rect 32680 12832 32720 12872
rect 36352 12832 36392 12872
rect 36434 12832 36474 12872
rect 36516 12832 36556 12872
rect 36598 12832 36638 12872
rect 36680 12832 36720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 44352 12832 44392 12872
rect 44434 12832 44474 12872
rect 44516 12832 44556 12872
rect 44598 12832 44638 12872
rect 44680 12832 44720 12872
rect 48352 12832 48392 12872
rect 48434 12832 48474 12872
rect 48516 12832 48556 12872
rect 48598 12832 48638 12872
rect 48680 12832 48720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 56352 12832 56392 12872
rect 56434 12832 56474 12872
rect 56516 12832 56556 12872
rect 56598 12832 56638 12872
rect 56680 12832 56720 12872
rect 60352 12832 60392 12872
rect 60434 12832 60474 12872
rect 60516 12832 60556 12872
rect 60598 12832 60638 12872
rect 60680 12832 60720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 7112 12076 7152 12116
rect 7194 12076 7234 12116
rect 7276 12076 7316 12116
rect 7358 12076 7398 12116
rect 7440 12076 7480 12116
rect 11112 12076 11152 12116
rect 11194 12076 11234 12116
rect 11276 12076 11316 12116
rect 11358 12076 11398 12116
rect 11440 12076 11480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 19112 12076 19152 12116
rect 19194 12076 19234 12116
rect 19276 12076 19316 12116
rect 19358 12076 19398 12116
rect 19440 12076 19480 12116
rect 23112 12076 23152 12116
rect 23194 12076 23234 12116
rect 23276 12076 23316 12116
rect 23358 12076 23398 12116
rect 23440 12076 23480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 31112 12076 31152 12116
rect 31194 12076 31234 12116
rect 31276 12076 31316 12116
rect 31358 12076 31398 12116
rect 31440 12076 31480 12116
rect 35112 12076 35152 12116
rect 35194 12076 35234 12116
rect 35276 12076 35316 12116
rect 35358 12076 35398 12116
rect 35440 12076 35480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 43112 12076 43152 12116
rect 43194 12076 43234 12116
rect 43276 12076 43316 12116
rect 43358 12076 43398 12116
rect 43440 12076 43480 12116
rect 47112 12076 47152 12116
rect 47194 12076 47234 12116
rect 47276 12076 47316 12116
rect 47358 12076 47398 12116
rect 47440 12076 47480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 55112 12076 55152 12116
rect 55194 12076 55234 12116
rect 55276 12076 55316 12116
rect 55358 12076 55398 12116
rect 55440 12076 55480 12116
rect 59112 12076 59152 12116
rect 59194 12076 59234 12116
rect 59276 12076 59316 12116
rect 59358 12076 59398 12116
rect 59440 12076 59480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 67112 12076 67152 12116
rect 67194 12076 67234 12116
rect 67276 12076 67316 12116
rect 67358 12076 67398 12116
rect 67440 12076 67480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 8352 11320 8392 11360
rect 8434 11320 8474 11360
rect 8516 11320 8556 11360
rect 8598 11320 8638 11360
rect 8680 11320 8720 11360
rect 12352 11320 12392 11360
rect 12434 11320 12474 11360
rect 12516 11320 12556 11360
rect 12598 11320 12638 11360
rect 12680 11320 12720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 20352 11320 20392 11360
rect 20434 11320 20474 11360
rect 20516 11320 20556 11360
rect 20598 11320 20638 11360
rect 20680 11320 20720 11360
rect 24352 11320 24392 11360
rect 24434 11320 24474 11360
rect 24516 11320 24556 11360
rect 24598 11320 24638 11360
rect 24680 11320 24720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 32352 11320 32392 11360
rect 32434 11320 32474 11360
rect 32516 11320 32556 11360
rect 32598 11320 32638 11360
rect 32680 11320 32720 11360
rect 36352 11320 36392 11360
rect 36434 11320 36474 11360
rect 36516 11320 36556 11360
rect 36598 11320 36638 11360
rect 36680 11320 36720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 44352 11320 44392 11360
rect 44434 11320 44474 11360
rect 44516 11320 44556 11360
rect 44598 11320 44638 11360
rect 44680 11320 44720 11360
rect 48352 11320 48392 11360
rect 48434 11320 48474 11360
rect 48516 11320 48556 11360
rect 48598 11320 48638 11360
rect 48680 11320 48720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 56352 11320 56392 11360
rect 56434 11320 56474 11360
rect 56516 11320 56556 11360
rect 56598 11320 56638 11360
rect 56680 11320 56720 11360
rect 60352 11320 60392 11360
rect 60434 11320 60474 11360
rect 60516 11320 60556 11360
rect 60598 11320 60638 11360
rect 60680 11320 60720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 2188 10900 2228 10940
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 7112 10564 7152 10604
rect 7194 10564 7234 10604
rect 7276 10564 7316 10604
rect 7358 10564 7398 10604
rect 7440 10564 7480 10604
rect 11112 10564 11152 10604
rect 11194 10564 11234 10604
rect 11276 10564 11316 10604
rect 11358 10564 11398 10604
rect 11440 10564 11480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 19112 10564 19152 10604
rect 19194 10564 19234 10604
rect 19276 10564 19316 10604
rect 19358 10564 19398 10604
rect 19440 10564 19480 10604
rect 23112 10564 23152 10604
rect 23194 10564 23234 10604
rect 23276 10564 23316 10604
rect 23358 10564 23398 10604
rect 23440 10564 23480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 31112 10564 31152 10604
rect 31194 10564 31234 10604
rect 31276 10564 31316 10604
rect 31358 10564 31398 10604
rect 31440 10564 31480 10604
rect 35112 10564 35152 10604
rect 35194 10564 35234 10604
rect 35276 10564 35316 10604
rect 35358 10564 35398 10604
rect 35440 10564 35480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 43112 10564 43152 10604
rect 43194 10564 43234 10604
rect 43276 10564 43316 10604
rect 43358 10564 43398 10604
rect 43440 10564 43480 10604
rect 47112 10564 47152 10604
rect 47194 10564 47234 10604
rect 47276 10564 47316 10604
rect 47358 10564 47398 10604
rect 47440 10564 47480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 55112 10564 55152 10604
rect 55194 10564 55234 10604
rect 55276 10564 55316 10604
rect 55358 10564 55398 10604
rect 55440 10564 55480 10604
rect 59112 10564 59152 10604
rect 59194 10564 59234 10604
rect 59276 10564 59316 10604
rect 59358 10564 59398 10604
rect 59440 10564 59480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 67112 10564 67152 10604
rect 67194 10564 67234 10604
rect 67276 10564 67316 10604
rect 67358 10564 67398 10604
rect 67440 10564 67480 10604
rect 68428 15520 68468 15560
rect 68044 14764 68084 14804
rect 69100 15520 69140 15560
rect 71692 16024 71732 16064
rect 69964 15772 70004 15812
rect 69868 15688 69908 15728
rect 69484 15604 69524 15644
rect 69292 15016 69332 15056
rect 69100 14932 69140 14972
rect 69292 14848 69332 14888
rect 68140 14680 68180 14720
rect 68620 14680 68660 14720
rect 68352 14344 68392 14384
rect 68434 14344 68474 14384
rect 68516 14344 68556 14384
rect 68598 14344 68638 14384
rect 68680 14344 68720 14384
rect 69388 14680 69428 14720
rect 71692 15436 71732 15476
rect 71692 15100 71732 15140
rect 71692 14764 71732 14804
rect 69004 13924 69044 13964
rect 69196 13924 69236 13964
rect 70060 13924 70100 13964
rect 68352 12832 68392 12872
rect 68434 12832 68474 12872
rect 68516 12832 68556 12872
rect 68598 12832 68638 12872
rect 68680 12832 68720 12872
rect 68352 11320 68392 11360
rect 68434 11320 68474 11360
rect 68516 11320 68556 11360
rect 68598 11320 68638 11360
rect 68680 11320 68720 11360
rect 68524 10984 68564 11024
rect 69772 10984 69812 11024
rect 67468 10144 67508 10184
rect 67660 10060 67700 10100
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 8352 9808 8392 9848
rect 8434 9808 8474 9848
rect 8516 9808 8556 9848
rect 8598 9808 8638 9848
rect 8680 9808 8720 9848
rect 12352 9808 12392 9848
rect 12434 9808 12474 9848
rect 12516 9808 12556 9848
rect 12598 9808 12638 9848
rect 12680 9808 12720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 20352 9808 20392 9848
rect 20434 9808 20474 9848
rect 20516 9808 20556 9848
rect 20598 9808 20638 9848
rect 20680 9808 20720 9848
rect 24352 9808 24392 9848
rect 24434 9808 24474 9848
rect 24516 9808 24556 9848
rect 24598 9808 24638 9848
rect 24680 9808 24720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 32352 9808 32392 9848
rect 32434 9808 32474 9848
rect 32516 9808 32556 9848
rect 32598 9808 32638 9848
rect 32680 9808 32720 9848
rect 36352 9808 36392 9848
rect 36434 9808 36474 9848
rect 36516 9808 36556 9848
rect 36598 9808 36638 9848
rect 36680 9808 36720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 44352 9808 44392 9848
rect 44434 9808 44474 9848
rect 44516 9808 44556 9848
rect 44598 9808 44638 9848
rect 44680 9808 44720 9848
rect 48352 9808 48392 9848
rect 48434 9808 48474 9848
rect 48516 9808 48556 9848
rect 48598 9808 48638 9848
rect 48680 9808 48720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 56352 9808 56392 9848
rect 56434 9808 56474 9848
rect 56516 9808 56556 9848
rect 56598 9808 56638 9848
rect 56680 9808 56720 9848
rect 60352 9808 60392 9848
rect 60434 9808 60474 9848
rect 60516 9808 60556 9848
rect 60598 9808 60638 9848
rect 60680 9808 60720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 68524 10144 68564 10184
rect 68332 9976 68372 10016
rect 68716 9976 68756 10016
rect 69004 9976 69044 10016
rect 68352 9808 68392 9848
rect 68434 9808 68474 9848
rect 68516 9808 68556 9848
rect 68598 9808 68638 9848
rect 68680 9808 68720 9848
rect 68236 9556 68276 9596
rect 69388 10144 69428 10184
rect 69388 9976 69428 10016
rect 69196 9472 69236 9512
rect 69676 10144 69716 10184
rect 69580 9808 69620 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 7112 9052 7152 9092
rect 7194 9052 7234 9092
rect 7276 9052 7316 9092
rect 7358 9052 7398 9092
rect 7440 9052 7480 9092
rect 11112 9052 11152 9092
rect 11194 9052 11234 9092
rect 11276 9052 11316 9092
rect 11358 9052 11398 9092
rect 11440 9052 11480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 19112 9052 19152 9092
rect 19194 9052 19234 9092
rect 19276 9052 19316 9092
rect 19358 9052 19398 9092
rect 19440 9052 19480 9092
rect 23112 9052 23152 9092
rect 23194 9052 23234 9092
rect 23276 9052 23316 9092
rect 23358 9052 23398 9092
rect 23440 9052 23480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 31112 9052 31152 9092
rect 31194 9052 31234 9092
rect 31276 9052 31316 9092
rect 31358 9052 31398 9092
rect 31440 9052 31480 9092
rect 35112 9052 35152 9092
rect 35194 9052 35234 9092
rect 35276 9052 35316 9092
rect 35358 9052 35398 9092
rect 35440 9052 35480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 43112 9052 43152 9092
rect 43194 9052 43234 9092
rect 43276 9052 43316 9092
rect 43358 9052 43398 9092
rect 43440 9052 43480 9092
rect 47112 9052 47152 9092
rect 47194 9052 47234 9092
rect 47276 9052 47316 9092
rect 47358 9052 47398 9092
rect 47440 9052 47480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 55112 9052 55152 9092
rect 55194 9052 55234 9092
rect 55276 9052 55316 9092
rect 55358 9052 55398 9092
rect 55440 9052 55480 9092
rect 59112 9052 59152 9092
rect 59194 9052 59234 9092
rect 59276 9052 59316 9092
rect 59358 9052 59398 9092
rect 59440 9052 59480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 67112 9052 67152 9092
rect 67194 9052 67234 9092
rect 67276 9052 67316 9092
rect 67358 9052 67398 9092
rect 67440 9052 67480 9092
rect 69196 9304 69236 9344
rect 69484 9388 69524 9428
rect 69772 9892 69812 9932
rect 69868 9724 69908 9764
rect 69676 9220 69716 9260
rect 69964 9136 70004 9176
rect 70732 10060 70772 10100
rect 70732 9640 70772 9680
rect 69004 8800 69044 8840
rect 652 8128 692 8168
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 8352 8296 8392 8336
rect 8434 8296 8474 8336
rect 8516 8296 8556 8336
rect 8598 8296 8638 8336
rect 8680 8296 8720 8336
rect 12352 8296 12392 8336
rect 12434 8296 12474 8336
rect 12516 8296 12556 8336
rect 12598 8296 12638 8336
rect 12680 8296 12720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 20352 8296 20392 8336
rect 20434 8296 20474 8336
rect 20516 8296 20556 8336
rect 20598 8296 20638 8336
rect 20680 8296 20720 8336
rect 24352 8296 24392 8336
rect 24434 8296 24474 8336
rect 24516 8296 24556 8336
rect 24598 8296 24638 8336
rect 24680 8296 24720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 32352 8296 32392 8336
rect 32434 8296 32474 8336
rect 32516 8296 32556 8336
rect 32598 8296 32638 8336
rect 32680 8296 32720 8336
rect 36352 8296 36392 8336
rect 36434 8296 36474 8336
rect 36516 8296 36556 8336
rect 36598 8296 36638 8336
rect 36680 8296 36720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 44352 8296 44392 8336
rect 44434 8296 44474 8336
rect 44516 8296 44556 8336
rect 44598 8296 44638 8336
rect 44680 8296 44720 8336
rect 48352 8296 48392 8336
rect 48434 8296 48474 8336
rect 48516 8296 48556 8336
rect 48598 8296 48638 8336
rect 48680 8296 48720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 56352 8296 56392 8336
rect 56434 8296 56474 8336
rect 56516 8296 56556 8336
rect 56598 8296 56638 8336
rect 56680 8296 56720 8336
rect 60352 8296 60392 8336
rect 60434 8296 60474 8336
rect 60516 8296 60556 8336
rect 60598 8296 60638 8336
rect 60680 8296 60720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 68352 8296 68392 8336
rect 68434 8296 68474 8336
rect 68516 8296 68556 8336
rect 68598 8296 68638 8336
rect 68680 8296 68720 8336
rect 69772 8128 69812 8168
rect 844 7792 884 7832
rect 1516 7792 1556 7832
rect 652 7288 692 7328
rect 844 6616 884 6656
rect 1324 6616 1364 6656
rect 652 6448 692 6488
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 7112 7540 7152 7580
rect 7194 7540 7234 7580
rect 7276 7540 7316 7580
rect 7358 7540 7398 7580
rect 7440 7540 7480 7580
rect 11112 7540 11152 7580
rect 11194 7540 11234 7580
rect 11276 7540 11316 7580
rect 11358 7540 11398 7580
rect 11440 7540 11480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 19112 7540 19152 7580
rect 19194 7540 19234 7580
rect 19276 7540 19316 7580
rect 19358 7540 19398 7580
rect 19440 7540 19480 7580
rect 23112 7540 23152 7580
rect 23194 7540 23234 7580
rect 23276 7540 23316 7580
rect 23358 7540 23398 7580
rect 23440 7540 23480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 31112 7540 31152 7580
rect 31194 7540 31234 7580
rect 31276 7540 31316 7580
rect 31358 7540 31398 7580
rect 31440 7540 31480 7580
rect 35112 7540 35152 7580
rect 35194 7540 35234 7580
rect 35276 7540 35316 7580
rect 35358 7540 35398 7580
rect 35440 7540 35480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 43112 7540 43152 7580
rect 43194 7540 43234 7580
rect 43276 7540 43316 7580
rect 43358 7540 43398 7580
rect 43440 7540 43480 7580
rect 47112 7540 47152 7580
rect 47194 7540 47234 7580
rect 47276 7540 47316 7580
rect 47358 7540 47398 7580
rect 47440 7540 47480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 55112 7540 55152 7580
rect 55194 7540 55234 7580
rect 55276 7540 55316 7580
rect 55358 7540 55398 7580
rect 55440 7540 55480 7580
rect 59112 7540 59152 7580
rect 59194 7540 59234 7580
rect 59276 7540 59316 7580
rect 59358 7540 59398 7580
rect 59440 7540 59480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 67112 7540 67152 7580
rect 67194 7540 67234 7580
rect 67276 7540 67316 7580
rect 67358 7540 67398 7580
rect 67440 7540 67480 7580
rect 71112 7540 71152 7580
rect 71194 7540 71234 7580
rect 71276 7540 71316 7580
rect 71358 7540 71398 7580
rect 71440 7540 71480 7580
rect 72352 18880 72392 18920
rect 72434 18880 72474 18920
rect 72516 18880 72556 18920
rect 72598 18880 72638 18920
rect 72680 18880 72720 18920
rect 75148 18880 75188 18920
rect 74572 18796 74612 18836
rect 74956 18796 74996 18836
rect 72940 18544 72980 18584
rect 73708 18544 73748 18584
rect 74284 18544 74324 18584
rect 72352 17368 72392 17408
rect 72434 17368 72474 17408
rect 72516 17368 72556 17408
rect 72598 17368 72638 17408
rect 72680 17368 72720 17408
rect 73708 17788 73748 17828
rect 74092 17788 74132 17828
rect 73228 15940 73268 15980
rect 73900 15856 73940 15896
rect 73132 15604 73172 15644
rect 75436 19216 75476 19256
rect 75244 18544 75284 18584
rect 75112 18124 75152 18164
rect 75194 18124 75234 18164
rect 75276 18124 75316 18164
rect 75358 18124 75398 18164
rect 75440 18124 75480 18164
rect 80620 19972 80660 20012
rect 86860 19972 86900 20012
rect 75724 19888 75764 19928
rect 79112 19636 79152 19676
rect 79194 19636 79234 19676
rect 79276 19636 79316 19676
rect 79358 19636 79398 19676
rect 79440 19636 79480 19676
rect 83112 19636 83152 19676
rect 83194 19636 83234 19676
rect 83276 19636 83316 19676
rect 83358 19636 83398 19676
rect 83440 19636 83480 19676
rect 75724 19216 75764 19256
rect 76588 19216 76628 19256
rect 75820 18880 75860 18920
rect 75628 18796 75668 18836
rect 75820 17704 75860 17744
rect 74188 16528 74228 16568
rect 74284 15772 74324 15812
rect 73612 15604 73652 15644
rect 72815 15520 72855 15560
rect 73036 15520 73076 15560
rect 72705 15436 72745 15476
rect 72415 15352 72455 15392
rect 73505 15520 73545 15560
rect 74668 16528 74708 16568
rect 75340 16024 75380 16064
rect 75105 15352 75145 15392
rect 75724 15352 75764 15392
rect 76204 18880 76244 18920
rect 76352 18880 76392 18920
rect 76434 18880 76474 18920
rect 76516 18880 76556 18920
rect 76598 18880 76638 18920
rect 76680 18880 76720 18920
rect 76972 18796 77012 18836
rect 76492 18544 76532 18584
rect 76588 17788 76628 17828
rect 76492 17704 76532 17744
rect 76972 17788 77012 17828
rect 76684 17536 76724 17576
rect 76352 17368 76392 17408
rect 76434 17368 76474 17408
rect 76516 17368 76556 17408
rect 76598 17368 76638 17408
rect 76680 17368 76720 17408
rect 76684 17200 76724 17240
rect 77452 18796 77492 18836
rect 77452 18544 77492 18584
rect 77356 17788 77396 17828
rect 77740 17788 77780 17828
rect 78124 18880 78164 18920
rect 80524 19300 80564 19340
rect 82060 19300 82100 19340
rect 82348 19300 82388 19340
rect 84076 19300 84116 19340
rect 85612 19300 85652 19340
rect 87112 19636 87152 19676
rect 87194 19636 87234 19676
rect 87276 19636 87316 19676
rect 87358 19636 87398 19676
rect 87440 19636 87480 19676
rect 91112 19636 91152 19676
rect 91194 19636 91234 19676
rect 91276 19636 91316 19676
rect 91358 19636 91398 19676
rect 91440 19636 91480 19676
rect 78604 18880 78644 18920
rect 78220 18796 78260 18836
rect 78412 18460 78452 18500
rect 78220 17788 78260 17828
rect 77836 15520 77876 15560
rect 77905 15352 77945 15392
rect 79372 18880 79412 18920
rect 78988 18796 79028 18836
rect 78796 18460 78836 18500
rect 81868 19132 81908 19172
rect 79372 18460 79412 18500
rect 79852 18460 79892 18500
rect 80044 18460 80084 18500
rect 78988 18208 79028 18248
rect 79112 18124 79152 18164
rect 79194 18124 79234 18164
rect 79276 18124 79316 18164
rect 79358 18124 79398 18164
rect 79440 18124 79480 18164
rect 78796 17872 78836 17912
rect 79180 17872 79220 17912
rect 79468 17872 79508 17912
rect 78508 15520 78548 15560
rect 79852 18208 79892 18248
rect 78815 15352 78855 15392
rect 78988 15352 79028 15392
rect 79215 15520 79255 15560
rect 80352 18880 80392 18920
rect 80434 18880 80474 18920
rect 80516 18880 80556 18920
rect 80598 18880 80638 18920
rect 80680 18880 80720 18920
rect 80524 18460 80564 18500
rect 81004 18460 81044 18500
rect 81388 18460 81428 18500
rect 81292 17704 81332 17744
rect 80716 17536 80756 17576
rect 80352 17368 80392 17408
rect 80434 17368 80474 17408
rect 80516 17368 80556 17408
rect 80598 17368 80638 17408
rect 80680 17368 80720 17408
rect 81004 17536 81044 17576
rect 81484 17704 81524 17744
rect 81964 17704 82004 17744
rect 86764 19300 86804 19340
rect 86956 19300 86996 19340
rect 86572 19216 86612 19256
rect 82636 19132 82676 19172
rect 83020 19132 83060 19172
rect 86956 19132 86996 19172
rect 82348 17704 82388 17744
rect 83404 18460 83444 18500
rect 84352 18880 84392 18920
rect 84434 18880 84474 18920
rect 84516 18880 84556 18920
rect 84598 18880 84638 18920
rect 84680 18880 84720 18920
rect 88204 19300 88244 19340
rect 89932 19216 89972 19256
rect 86572 18544 86612 18584
rect 87052 18544 87092 18584
rect 87436 18544 87476 18584
rect 83788 18460 83828 18500
rect 84268 18460 84308 18500
rect 84652 18460 84692 18500
rect 85036 18460 85076 18500
rect 85516 18460 85556 18500
rect 83112 18124 83152 18164
rect 83194 18124 83234 18164
rect 83276 18124 83316 18164
rect 83358 18124 83398 18164
rect 83440 18124 83480 18164
rect 83404 17704 83444 17744
rect 83788 17704 83828 17744
rect 84172 17704 84212 17744
rect 84748 17788 84788 17828
rect 84652 17620 84692 17660
rect 84460 17536 84500 17576
rect 84352 17368 84392 17408
rect 84434 17368 84474 17408
rect 84516 17368 84556 17408
rect 84598 17368 84638 17408
rect 84680 17368 84720 17408
rect 84940 17788 84980 17828
rect 85900 18460 85940 18500
rect 85420 17788 85460 17828
rect 84415 15520 84455 15560
rect 84705 15520 84745 15560
rect 85036 17452 85076 17492
rect 84940 15520 84980 15560
rect 86284 18460 86324 18500
rect 86188 17704 86228 17744
rect 86572 17704 86612 17744
rect 87112 18124 87152 18164
rect 87194 18124 87234 18164
rect 87276 18124 87316 18164
rect 87358 18124 87398 18164
rect 87440 18124 87480 18164
rect 87052 17704 87092 17744
rect 87436 17704 87476 17744
rect 88352 18880 88392 18920
rect 88434 18880 88474 18920
rect 88516 18880 88556 18920
rect 88598 18880 88638 18920
rect 88680 18880 88720 18920
rect 90124 18880 90164 18920
rect 90508 18880 90548 18920
rect 91372 18880 91412 18920
rect 87724 18460 87764 18500
rect 88012 18460 88052 18500
rect 87916 17620 87956 17660
rect 88204 18460 88244 18500
rect 88588 18460 88628 18500
rect 88972 18460 89012 18500
rect 89548 18460 89588 18500
rect 88108 17620 88148 17660
rect 89740 18460 89780 18500
rect 90124 18460 90164 18500
rect 88588 17704 88628 17744
rect 88396 17536 88436 17576
rect 88352 17368 88392 17408
rect 88434 17368 88474 17408
rect 88516 17368 88556 17408
rect 88598 17368 88638 17408
rect 88680 17368 88720 17408
rect 88396 17200 88436 17240
rect 89068 17704 89108 17744
rect 89452 17704 89492 17744
rect 89932 17704 89972 17744
rect 89836 15688 89876 15728
rect 90220 17704 90260 17744
rect 92352 18880 92392 18920
rect 92434 18880 92474 18920
rect 92516 18880 92556 18920
rect 92598 18880 92638 18920
rect 92680 18880 92720 18920
rect 93100 19300 93140 19340
rect 95112 19636 95152 19676
rect 95194 19636 95234 19676
rect 95276 19636 95316 19676
rect 95358 19636 95398 19676
rect 95440 19636 95480 19676
rect 99112 19636 99152 19676
rect 99194 19636 99234 19676
rect 99276 19636 99316 19676
rect 99358 19636 99398 19676
rect 99440 19636 99480 19676
rect 94156 19300 94196 19340
rect 95788 19300 95828 19340
rect 97132 19300 97172 19340
rect 93196 19216 93236 19256
rect 91468 18544 91508 18584
rect 90604 18460 90644 18500
rect 91852 18544 91892 18584
rect 92236 18544 92276 18584
rect 90604 17704 90644 17744
rect 91112 18124 91152 18164
rect 91194 18124 91234 18164
rect 91276 18124 91316 18164
rect 91358 18124 91398 18164
rect 91440 18124 91480 18164
rect 90988 17704 91028 17744
rect 91372 17704 91412 17744
rect 91180 16528 91220 16568
rect 89505 15436 89545 15476
rect 92620 18460 92660 18500
rect 92908 18460 92948 18500
rect 91852 17704 91892 17744
rect 91660 16528 91700 16568
rect 92236 17704 92276 17744
rect 92812 17956 92852 17996
rect 92908 17620 92948 17660
rect 92140 15520 92180 15560
rect 92352 17368 92392 17408
rect 92434 17368 92474 17408
rect 92516 17368 92556 17408
rect 92598 17368 92638 17408
rect 92680 17368 92720 17408
rect 92415 15520 92455 15560
rect 93196 18544 93236 18584
rect 93100 18460 93140 18500
rect 95116 18544 95156 18584
rect 93196 17956 93236 17996
rect 93196 17788 93236 17828
rect 93772 17788 93812 17828
rect 93484 17620 93524 17660
rect 94540 18292 94580 18332
rect 96352 18880 96392 18920
rect 96434 18880 96474 18920
rect 96516 18880 96556 18920
rect 96598 18880 96638 18920
rect 96680 18880 96720 18920
rect 95212 18292 95252 18332
rect 95500 18292 95540 18332
rect 95112 18124 95152 18164
rect 95194 18124 95234 18164
rect 95276 18124 95316 18164
rect 95358 18124 95398 18164
rect 95440 18124 95480 18164
rect 95404 17956 95444 17996
rect 94732 17788 94772 17828
rect 94924 17788 94964 17828
rect 95884 17956 95924 17996
rect 96076 17956 96116 17996
rect 96076 15604 96116 15644
rect 96364 17956 96404 17996
rect 96652 17956 96692 17996
rect 97036 17788 97076 17828
rect 97324 17872 97364 17912
rect 96352 17368 96392 17408
rect 96434 17368 96474 17408
rect 96516 17368 96556 17408
rect 96598 17368 96638 17408
rect 96680 17368 96720 17408
rect 96748 16360 96788 16400
rect 96172 15520 96212 15560
rect 96015 15352 96055 15392
rect 96415 15520 96455 15560
rect 97516 16360 97556 16400
rect 99112 18124 99152 18164
rect 99194 18124 99234 18164
rect 99276 18124 99316 18164
rect 99358 18124 99398 18164
rect 99440 18124 99480 18164
rect 98476 17956 98516 17996
rect 97900 17788 97940 17828
rect 97900 17620 97940 17660
rect 98668 17704 98708 17744
rect 98764 17620 98804 17660
rect 98415 15436 98455 15476
rect 98305 15352 98345 15392
rect 98956 15352 98996 15392
rect 71884 14932 71924 14972
rect 72305 9808 72345 9848
rect 72415 9724 72455 9764
rect 73215 9892 73255 9932
rect 73228 9724 73268 9764
rect 72844 9556 72884 9596
rect 73132 9472 73172 9512
rect 72652 9304 72692 9344
rect 73905 9892 73945 9932
rect 73324 9640 73364 9680
rect 73612 9388 73652 9428
rect 73228 9220 73268 9260
rect 73324 8800 73364 8840
rect 71788 7204 71828 7244
rect 74572 9724 74612 9764
rect 74380 9136 74420 9176
rect 74188 7540 74228 7580
rect 74092 7036 74132 7076
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 8352 6784 8392 6824
rect 8434 6784 8474 6824
rect 8516 6784 8556 6824
rect 8598 6784 8638 6824
rect 8680 6784 8720 6824
rect 12352 6784 12392 6824
rect 12434 6784 12474 6824
rect 12516 6784 12556 6824
rect 12598 6784 12638 6824
rect 12680 6784 12720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 20352 6784 20392 6824
rect 20434 6784 20474 6824
rect 20516 6784 20556 6824
rect 20598 6784 20638 6824
rect 20680 6784 20720 6824
rect 24352 6784 24392 6824
rect 24434 6784 24474 6824
rect 24516 6784 24556 6824
rect 24598 6784 24638 6824
rect 24680 6784 24720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 32352 6784 32392 6824
rect 32434 6784 32474 6824
rect 32516 6784 32556 6824
rect 32598 6784 32638 6824
rect 32680 6784 32720 6824
rect 36352 6784 36392 6824
rect 36434 6784 36474 6824
rect 36516 6784 36556 6824
rect 36598 6784 36638 6824
rect 36680 6784 36720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 44352 6784 44392 6824
rect 44434 6784 44474 6824
rect 44516 6784 44556 6824
rect 44598 6784 44638 6824
rect 44680 6784 44720 6824
rect 48352 6784 48392 6824
rect 48434 6784 48474 6824
rect 48516 6784 48556 6824
rect 48598 6784 48638 6824
rect 48680 6784 48720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 56352 6784 56392 6824
rect 56434 6784 56474 6824
rect 56516 6784 56556 6824
rect 56598 6784 56638 6824
rect 56680 6784 56720 6824
rect 60352 6784 60392 6824
rect 60434 6784 60474 6824
rect 60516 6784 60556 6824
rect 60598 6784 60638 6824
rect 60680 6784 60720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 68352 6784 68392 6824
rect 68434 6784 68474 6824
rect 68516 6784 68556 6824
rect 68598 6784 68638 6824
rect 68680 6784 68720 6824
rect 72352 6784 72392 6824
rect 72434 6784 72474 6824
rect 72516 6784 72556 6824
rect 72598 6784 72638 6824
rect 72680 6784 72720 6824
rect 74284 7288 74324 7328
rect 74476 7288 74516 7328
rect 74764 7708 74804 7748
rect 74668 7456 74708 7496
rect 74668 7204 74708 7244
rect 74380 6784 74420 6824
rect 74572 6364 74612 6404
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 7112 6028 7152 6068
rect 7194 6028 7234 6068
rect 7276 6028 7316 6068
rect 7358 6028 7398 6068
rect 7440 6028 7480 6068
rect 11112 6028 11152 6068
rect 11194 6028 11234 6068
rect 11276 6028 11316 6068
rect 11358 6028 11398 6068
rect 11440 6028 11480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 19112 6028 19152 6068
rect 19194 6028 19234 6068
rect 19276 6028 19316 6068
rect 19358 6028 19398 6068
rect 19440 6028 19480 6068
rect 23112 6028 23152 6068
rect 23194 6028 23234 6068
rect 23276 6028 23316 6068
rect 23358 6028 23398 6068
rect 23440 6028 23480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 31112 6028 31152 6068
rect 31194 6028 31234 6068
rect 31276 6028 31316 6068
rect 31358 6028 31398 6068
rect 31440 6028 31480 6068
rect 35112 6028 35152 6068
rect 35194 6028 35234 6068
rect 35276 6028 35316 6068
rect 35358 6028 35398 6068
rect 35440 6028 35480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 43112 6028 43152 6068
rect 43194 6028 43234 6068
rect 43276 6028 43316 6068
rect 43358 6028 43398 6068
rect 43440 6028 43480 6068
rect 47112 6028 47152 6068
rect 47194 6028 47234 6068
rect 47276 6028 47316 6068
rect 47358 6028 47398 6068
rect 47440 6028 47480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 55112 6028 55152 6068
rect 55194 6028 55234 6068
rect 55276 6028 55316 6068
rect 55358 6028 55398 6068
rect 55440 6028 55480 6068
rect 59112 6028 59152 6068
rect 59194 6028 59234 6068
rect 59276 6028 59316 6068
rect 59358 6028 59398 6068
rect 59440 6028 59480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 67112 6028 67152 6068
rect 67194 6028 67234 6068
rect 67276 6028 67316 6068
rect 67358 6028 67398 6068
rect 67440 6028 67480 6068
rect 71112 6028 71152 6068
rect 71194 6028 71234 6068
rect 71276 6028 71316 6068
rect 71358 6028 71398 6068
rect 71440 6028 71480 6068
rect 844 5776 884 5816
rect 652 5608 692 5648
rect 844 5440 884 5480
rect 1420 5440 1460 5480
rect 1804 5776 1844 5816
rect 74956 9808 74996 9848
rect 74860 7540 74900 7580
rect 74860 6952 74900 6992
rect 74764 6364 74804 6404
rect 75215 9808 75255 9848
rect 75505 9724 75545 9764
rect 75052 7708 75092 7748
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 75244 7372 75284 7412
rect 75148 7288 75188 7328
rect 75052 7036 75092 7076
rect 75436 7204 75476 7244
rect 75148 6868 75188 6908
rect 75436 6952 75476 6992
rect 75340 6616 75380 6656
rect 75724 7204 75764 7244
rect 75724 6952 75764 6992
rect 75436 6448 75476 6488
rect 76588 7372 76628 7412
rect 76684 7120 76724 7160
rect 76588 7036 76628 7076
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 76588 6616 76628 6656
rect 77068 7372 77108 7412
rect 76876 7204 76916 7244
rect 77452 7372 77492 7412
rect 77644 7372 77684 7412
rect 77260 7288 77300 7328
rect 77260 7120 77300 7160
rect 77644 7204 77684 7244
rect 77836 7204 77876 7244
rect 77644 7036 77684 7076
rect 77452 6952 77492 6992
rect 76108 6448 76148 6488
rect 76300 6448 76340 6488
rect 75148 6364 75188 6404
rect 78028 7540 78068 7580
rect 78028 7372 78068 7412
rect 78124 6952 78164 6992
rect 78316 7540 78356 7580
rect 78412 7036 78452 7076
rect 77740 6364 77780 6404
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 76684 5860 76724 5900
rect 78124 6364 78164 6404
rect 79505 9808 79545 9848
rect 79756 9808 79796 9848
rect 78700 7036 78740 7076
rect 78604 6364 78644 6404
rect 79112 7540 79152 7580
rect 79194 7540 79234 7580
rect 79276 7540 79316 7580
rect 79358 7540 79398 7580
rect 79440 7540 79480 7580
rect 79660 7288 79700 7328
rect 79084 7204 79124 7244
rect 79372 6952 79412 6992
rect 80305 9724 80345 9764
rect 80044 7288 80084 7328
rect 78892 6364 78932 6404
rect 80236 7204 80276 7244
rect 79112 6028 79152 6068
rect 79194 6028 79234 6068
rect 79276 6028 79316 6068
rect 79358 6028 79398 6068
rect 79440 6028 79480 6068
rect 80140 5860 80180 5900
rect 80716 7204 80756 7244
rect 80524 6952 80564 6992
rect 80352 6784 80392 6824
rect 80434 6784 80474 6824
rect 80516 6784 80556 6824
rect 80598 6784 80638 6824
rect 80680 6784 80720 6824
rect 80908 7372 80948 7412
rect 80908 7120 80948 7160
rect 81100 7204 81140 7244
rect 81580 8212 81620 8252
rect 81292 7120 81332 7160
rect 82305 9808 82345 9848
rect 82540 9808 82580 9848
rect 82252 8212 82292 8252
rect 81676 7540 81716 7580
rect 81676 7372 81716 7412
rect 81964 7540 82004 7580
rect 81772 6952 81812 6992
rect 82252 7204 82292 7244
rect 83615 9724 83655 9764
rect 82636 7120 82676 7160
rect 81961 7036 82001 7076
rect 82828 7204 82868 7244
rect 83116 7876 83156 7916
rect 83112 7540 83152 7580
rect 83194 7540 83234 7580
rect 83276 7540 83316 7580
rect 83358 7540 83398 7580
rect 83440 7540 83480 7580
rect 83116 7120 83156 7160
rect 83308 7120 83348 7160
rect 82924 7036 82964 7076
rect 82060 6364 82100 6404
rect 82540 6364 82580 6404
rect 83884 7372 83924 7412
rect 83788 7120 83828 7160
rect 84076 7372 84116 7412
rect 84268 7204 84308 7244
rect 84076 7120 84116 7160
rect 84460 7540 84500 7580
rect 84652 7372 84692 7412
rect 82732 6364 82772 6404
rect 83212 6364 83252 6404
rect 83692 6364 83732 6404
rect 84556 6952 84596 6992
rect 84844 7372 84884 7412
rect 84844 7120 84884 7160
rect 84352 6784 84392 6824
rect 84434 6784 84474 6824
rect 84516 6784 84556 6824
rect 84598 6784 84638 6824
rect 84680 6784 84720 6824
rect 85228 7204 85268 7244
rect 84172 6364 84212 6404
rect 84556 6364 84596 6404
rect 85036 6364 85076 6404
rect 85612 8800 85652 8840
rect 85708 7540 85748 7580
rect 85612 7120 85652 7160
rect 86188 8128 86228 8168
rect 86092 7204 86132 7244
rect 85996 6952 86036 6992
rect 86092 6532 86132 6572
rect 85228 6364 85268 6404
rect 83112 6028 83152 6068
rect 83194 6028 83234 6068
rect 83276 6028 83316 6068
rect 83358 6028 83398 6068
rect 83440 6028 83480 6068
rect 83596 5860 83636 5900
rect 85612 6364 85652 6404
rect 86092 6364 86132 6404
rect 85516 5860 85556 5900
rect 86284 7288 86324 7328
rect 86476 7540 86516 7580
rect 86668 7372 86708 7412
rect 86476 7204 86516 7244
rect 86668 6868 86708 6908
rect 87215 9724 87255 9764
rect 87724 9724 87764 9764
rect 87112 7540 87152 7580
rect 87194 7540 87234 7580
rect 87276 7540 87316 7580
rect 87358 7540 87398 7580
rect 87440 7540 87480 7580
rect 86956 7120 86996 7160
rect 86956 6952 86996 6992
rect 87148 7372 87188 7412
rect 87244 7288 87284 7328
rect 87244 7036 87284 7076
rect 86860 6532 86900 6572
rect 87436 7120 87476 7160
rect 87532 7036 87572 7076
rect 86188 5776 86228 5816
rect 87112 6028 87152 6068
rect 87194 6028 87234 6068
rect 87276 6028 87316 6068
rect 87358 6028 87398 6068
rect 87440 6028 87480 6068
rect 87820 7036 87860 7076
rect 88012 7540 88052 7580
rect 88012 7204 88052 7244
rect 88300 7204 88340 7244
rect 88012 7036 88052 7076
rect 88588 7204 88628 7244
rect 88396 6952 88436 6992
rect 88352 6784 88392 6824
rect 88434 6784 88474 6824
rect 88516 6784 88556 6824
rect 88598 6784 88638 6824
rect 88680 6784 88720 6824
rect 89105 9724 89145 9764
rect 88972 7540 89012 7580
rect 89068 7204 89108 7244
rect 88492 6616 88532 6656
rect 88108 6448 88148 6488
rect 88588 6448 88628 6488
rect 89452 7120 89492 7160
rect 88876 6448 88916 6488
rect 89644 7372 89684 7412
rect 89644 6364 89684 6404
rect 89068 5860 89108 5900
rect 89836 7372 89876 7412
rect 90028 7372 90068 7412
rect 89836 7120 89876 7160
rect 90028 7036 90068 7076
rect 90316 6868 90356 6908
rect 91505 9808 91545 9848
rect 91756 9808 91796 9848
rect 90604 7372 90644 7412
rect 90892 7372 90932 7412
rect 91112 7540 91152 7580
rect 91194 7540 91234 7580
rect 91276 7540 91316 7580
rect 91358 7540 91398 7580
rect 91440 7540 91480 7580
rect 90988 7204 91028 7244
rect 90713 7120 90753 7160
rect 90892 7120 90932 7160
rect 91180 7288 91220 7328
rect 91564 7204 91604 7244
rect 91372 7036 91412 7076
rect 91852 7372 91892 7412
rect 91756 7288 91796 7328
rect 91756 7120 91796 7160
rect 92705 9724 92745 9764
rect 93004 9808 93044 9848
rect 92908 9724 92948 9764
rect 92140 7204 92180 7244
rect 92428 7540 92468 7580
rect 92332 7288 92372 7328
rect 92524 7204 92564 7244
rect 92716 7036 92756 7076
rect 92352 6784 92392 6824
rect 92434 6784 92474 6824
rect 92516 6784 92556 6824
rect 92598 6784 92638 6824
rect 92680 6784 92720 6824
rect 90412 6364 90452 6404
rect 90892 6364 90932 6404
rect 91372 6364 91412 6404
rect 91112 6028 91152 6068
rect 91194 6028 91234 6068
rect 91276 6028 91316 6068
rect 91358 6028 91398 6068
rect 91440 6028 91480 6068
rect 91660 6364 91700 6404
rect 92140 6364 92180 6404
rect 92524 6364 92564 6404
rect 93215 9808 93255 9848
rect 93100 7288 93140 7328
rect 93292 7540 93332 7580
rect 93484 7372 93524 7412
rect 93388 7288 93428 7328
rect 93004 6280 93044 6320
rect 93388 6280 93428 6320
rect 93676 7372 93716 7412
rect 93964 7288 94004 7328
rect 93772 7120 93812 7160
rect 93676 7036 93716 7076
rect 93772 6952 93812 6992
rect 94156 7204 94196 7244
rect 94156 7036 94196 7076
rect 93676 6616 93716 6656
rect 93868 6280 93908 6320
rect 94732 7120 94772 7160
rect 94444 6952 94484 6992
rect 94348 6868 94388 6908
rect 94540 6616 94580 6656
rect 95404 7792 95444 7832
rect 95212 7708 95252 7748
rect 95112 7540 95152 7580
rect 95194 7540 95234 7580
rect 95276 7540 95316 7580
rect 95358 7540 95398 7580
rect 95440 7540 95480 7580
rect 94924 7288 94964 7328
rect 95308 7288 95348 7328
rect 95308 6700 95348 6740
rect 95692 7204 95732 7244
rect 95692 6616 95732 6656
rect 94060 6364 94100 6404
rect 94444 6364 94484 6404
rect 94924 6364 94964 6404
rect 95116 6364 95156 6404
rect 93292 5608 93332 5648
rect 93676 5608 93716 5648
rect 95112 6028 95152 6068
rect 95194 6028 95234 6068
rect 95276 6028 95316 6068
rect 95358 6028 95398 6068
rect 95440 6028 95480 6068
rect 95884 9724 95924 9764
rect 96305 9724 96345 9764
rect 95884 6448 95924 6488
rect 96172 7708 96212 7748
rect 96076 7204 96116 7244
rect 96076 6532 96116 6572
rect 95884 6280 95924 6320
rect 95980 6196 96020 6236
rect 96460 7372 96500 7412
rect 96268 7204 96308 7244
rect 96652 7204 96692 7244
rect 96460 7036 96500 7076
rect 96844 7540 96884 7580
rect 96844 7372 96884 7412
rect 96940 7120 96980 7160
rect 96352 6784 96392 6824
rect 96434 6784 96474 6824
rect 96516 6784 96556 6824
rect 96598 6784 96638 6824
rect 96680 6784 96720 6824
rect 97132 7540 97172 7580
rect 97228 7120 97268 7160
rect 97516 9472 97556 9512
rect 96364 6280 96404 6320
rect 96940 6280 96980 6320
rect 97324 6280 97364 6320
rect 96172 6196 96212 6236
rect 96940 5776 96980 5816
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 8352 5272 8392 5312
rect 8434 5272 8474 5312
rect 8516 5272 8556 5312
rect 8598 5272 8638 5312
rect 8680 5272 8720 5312
rect 12352 5272 12392 5312
rect 12434 5272 12474 5312
rect 12516 5272 12556 5312
rect 12598 5272 12638 5312
rect 12680 5272 12720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 20352 5272 20392 5312
rect 20434 5272 20474 5312
rect 20516 5272 20556 5312
rect 20598 5272 20638 5312
rect 20680 5272 20720 5312
rect 24352 5272 24392 5312
rect 24434 5272 24474 5312
rect 24516 5272 24556 5312
rect 24598 5272 24638 5312
rect 24680 5272 24720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 32352 5272 32392 5312
rect 32434 5272 32474 5312
rect 32516 5272 32556 5312
rect 32598 5272 32638 5312
rect 32680 5272 32720 5312
rect 36352 5272 36392 5312
rect 36434 5272 36474 5312
rect 36516 5272 36556 5312
rect 36598 5272 36638 5312
rect 36680 5272 36720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 44352 5272 44392 5312
rect 44434 5272 44474 5312
rect 44516 5272 44556 5312
rect 44598 5272 44638 5312
rect 44680 5272 44720 5312
rect 48352 5272 48392 5312
rect 48434 5272 48474 5312
rect 48516 5272 48556 5312
rect 48598 5272 48638 5312
rect 48680 5272 48720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 56352 5272 56392 5312
rect 56434 5272 56474 5312
rect 56516 5272 56556 5312
rect 56598 5272 56638 5312
rect 56680 5272 56720 5312
rect 60352 5272 60392 5312
rect 60434 5272 60474 5312
rect 60516 5272 60556 5312
rect 60598 5272 60638 5312
rect 60680 5272 60720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 68352 5272 68392 5312
rect 68434 5272 68474 5312
rect 68516 5272 68556 5312
rect 68598 5272 68638 5312
rect 68680 5272 68720 5312
rect 72352 5272 72392 5312
rect 72434 5272 72474 5312
rect 72516 5272 72556 5312
rect 72598 5272 72638 5312
rect 72680 5272 72720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 80352 5272 80392 5312
rect 80434 5272 80474 5312
rect 80516 5272 80556 5312
rect 80598 5272 80638 5312
rect 80680 5272 80720 5312
rect 84352 5272 84392 5312
rect 84434 5272 84474 5312
rect 84516 5272 84556 5312
rect 84598 5272 84638 5312
rect 84680 5272 84720 5312
rect 88352 5272 88392 5312
rect 88434 5272 88474 5312
rect 88516 5272 88556 5312
rect 88598 5272 88638 5312
rect 88680 5272 88720 5312
rect 92352 5272 92392 5312
rect 92434 5272 92474 5312
rect 92516 5272 92556 5312
rect 92598 5272 92638 5312
rect 92680 5272 92720 5312
rect 96352 5272 96392 5312
rect 96434 5272 96474 5312
rect 96516 5272 96556 5312
rect 96598 5272 96638 5312
rect 96680 5272 96720 5312
rect 97612 7204 97652 7244
rect 97804 7204 97844 7244
rect 97996 6616 98036 6656
rect 98188 7204 98228 7244
rect 98380 5776 98420 5816
rect 98668 5776 98708 5816
rect 99112 7540 99152 7580
rect 99194 7540 99234 7580
rect 99276 7540 99316 7580
rect 99358 7540 99398 7580
rect 99440 7540 99480 7580
rect 99112 6028 99152 6068
rect 99194 6028 99234 6068
rect 99276 6028 99316 6068
rect 99358 6028 99398 6068
rect 99440 6028 99480 6068
rect 652 4768 692 4808
rect 748 4684 788 4724
rect 652 3928 692 3968
rect 652 3172 692 3212
rect 844 4180 884 4220
rect 1996 4684 2036 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 7112 4516 7152 4556
rect 7194 4516 7234 4556
rect 7276 4516 7316 4556
rect 7358 4516 7398 4556
rect 7440 4516 7480 4556
rect 11112 4516 11152 4556
rect 11194 4516 11234 4556
rect 11276 4516 11316 4556
rect 11358 4516 11398 4556
rect 11440 4516 11480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 19112 4516 19152 4556
rect 19194 4516 19234 4556
rect 19276 4516 19316 4556
rect 19358 4516 19398 4556
rect 19440 4516 19480 4556
rect 23112 4516 23152 4556
rect 23194 4516 23234 4556
rect 23276 4516 23316 4556
rect 23358 4516 23398 4556
rect 23440 4516 23480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 31112 4516 31152 4556
rect 31194 4516 31234 4556
rect 31276 4516 31316 4556
rect 31358 4516 31398 4556
rect 31440 4516 31480 4556
rect 35112 4516 35152 4556
rect 35194 4516 35234 4556
rect 35276 4516 35316 4556
rect 35358 4516 35398 4556
rect 35440 4516 35480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 43112 4516 43152 4556
rect 43194 4516 43234 4556
rect 43276 4516 43316 4556
rect 43358 4516 43398 4556
rect 43440 4516 43480 4556
rect 47112 4516 47152 4556
rect 47194 4516 47234 4556
rect 47276 4516 47316 4556
rect 47358 4516 47398 4556
rect 47440 4516 47480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 55112 4516 55152 4556
rect 55194 4516 55234 4556
rect 55276 4516 55316 4556
rect 55358 4516 55398 4556
rect 55440 4516 55480 4556
rect 59112 4516 59152 4556
rect 59194 4516 59234 4556
rect 59276 4516 59316 4556
rect 59358 4516 59398 4556
rect 59440 4516 59480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 67112 4516 67152 4556
rect 67194 4516 67234 4556
rect 67276 4516 67316 4556
rect 67358 4516 67398 4556
rect 67440 4516 67480 4556
rect 71112 4516 71152 4556
rect 71194 4516 71234 4556
rect 71276 4516 71316 4556
rect 71358 4516 71398 4556
rect 71440 4516 71480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 79112 4516 79152 4556
rect 79194 4516 79234 4556
rect 79276 4516 79316 4556
rect 79358 4516 79398 4556
rect 79440 4516 79480 4556
rect 83112 4516 83152 4556
rect 83194 4516 83234 4556
rect 83276 4516 83316 4556
rect 83358 4516 83398 4556
rect 83440 4516 83480 4556
rect 87112 4516 87152 4556
rect 87194 4516 87234 4556
rect 87276 4516 87316 4556
rect 87358 4516 87398 4556
rect 87440 4516 87480 4556
rect 91112 4516 91152 4556
rect 91194 4516 91234 4556
rect 91276 4516 91316 4556
rect 91358 4516 91398 4556
rect 91440 4516 91480 4556
rect 95112 4516 95152 4556
rect 95194 4516 95234 4556
rect 95276 4516 95316 4556
rect 95358 4516 95398 4556
rect 95440 4516 95480 4556
rect 99112 4516 99152 4556
rect 99194 4516 99234 4556
rect 99276 4516 99316 4556
rect 99358 4516 99398 4556
rect 99440 4516 99480 4556
rect 1612 4180 1652 4220
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 8352 3760 8392 3800
rect 8434 3760 8474 3800
rect 8516 3760 8556 3800
rect 8598 3760 8638 3800
rect 8680 3760 8720 3800
rect 12352 3760 12392 3800
rect 12434 3760 12474 3800
rect 12516 3760 12556 3800
rect 12598 3760 12638 3800
rect 12680 3760 12720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 20352 3760 20392 3800
rect 20434 3760 20474 3800
rect 20516 3760 20556 3800
rect 20598 3760 20638 3800
rect 20680 3760 20720 3800
rect 24352 3760 24392 3800
rect 24434 3760 24474 3800
rect 24516 3760 24556 3800
rect 24598 3760 24638 3800
rect 24680 3760 24720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 32352 3760 32392 3800
rect 32434 3760 32474 3800
rect 32516 3760 32556 3800
rect 32598 3760 32638 3800
rect 32680 3760 32720 3800
rect 36352 3760 36392 3800
rect 36434 3760 36474 3800
rect 36516 3760 36556 3800
rect 36598 3760 36638 3800
rect 36680 3760 36720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 44352 3760 44392 3800
rect 44434 3760 44474 3800
rect 44516 3760 44556 3800
rect 44598 3760 44638 3800
rect 44680 3760 44720 3800
rect 48352 3760 48392 3800
rect 48434 3760 48474 3800
rect 48516 3760 48556 3800
rect 48598 3760 48638 3800
rect 48680 3760 48720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 56352 3760 56392 3800
rect 56434 3760 56474 3800
rect 56516 3760 56556 3800
rect 56598 3760 56638 3800
rect 56680 3760 56720 3800
rect 60352 3760 60392 3800
rect 60434 3760 60474 3800
rect 60516 3760 60556 3800
rect 60598 3760 60638 3800
rect 60680 3760 60720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 68352 3760 68392 3800
rect 68434 3760 68474 3800
rect 68516 3760 68556 3800
rect 68598 3760 68638 3800
rect 68680 3760 68720 3800
rect 72352 3760 72392 3800
rect 72434 3760 72474 3800
rect 72516 3760 72556 3800
rect 72598 3760 72638 3800
rect 72680 3760 72720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 80352 3760 80392 3800
rect 80434 3760 80474 3800
rect 80516 3760 80556 3800
rect 80598 3760 80638 3800
rect 80680 3760 80720 3800
rect 84352 3760 84392 3800
rect 84434 3760 84474 3800
rect 84516 3760 84556 3800
rect 84598 3760 84638 3800
rect 84680 3760 84720 3800
rect 88352 3760 88392 3800
rect 88434 3760 88474 3800
rect 88516 3760 88556 3800
rect 88598 3760 88638 3800
rect 88680 3760 88720 3800
rect 92352 3760 92392 3800
rect 92434 3760 92474 3800
rect 92516 3760 92556 3800
rect 92598 3760 92638 3800
rect 92680 3760 92720 3800
rect 96352 3760 96392 3800
rect 96434 3760 96474 3800
rect 96516 3760 96556 3800
rect 96598 3760 96638 3800
rect 96680 3760 96720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 7112 3004 7152 3044
rect 7194 3004 7234 3044
rect 7276 3004 7316 3044
rect 7358 3004 7398 3044
rect 7440 3004 7480 3044
rect 11112 3004 11152 3044
rect 11194 3004 11234 3044
rect 11276 3004 11316 3044
rect 11358 3004 11398 3044
rect 11440 3004 11480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 19112 3004 19152 3044
rect 19194 3004 19234 3044
rect 19276 3004 19316 3044
rect 19358 3004 19398 3044
rect 19440 3004 19480 3044
rect 23112 3004 23152 3044
rect 23194 3004 23234 3044
rect 23276 3004 23316 3044
rect 23358 3004 23398 3044
rect 23440 3004 23480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 31112 3004 31152 3044
rect 31194 3004 31234 3044
rect 31276 3004 31316 3044
rect 31358 3004 31398 3044
rect 31440 3004 31480 3044
rect 35112 3004 35152 3044
rect 35194 3004 35234 3044
rect 35276 3004 35316 3044
rect 35358 3004 35398 3044
rect 35440 3004 35480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 43112 3004 43152 3044
rect 43194 3004 43234 3044
rect 43276 3004 43316 3044
rect 43358 3004 43398 3044
rect 43440 3004 43480 3044
rect 47112 3004 47152 3044
rect 47194 3004 47234 3044
rect 47276 3004 47316 3044
rect 47358 3004 47398 3044
rect 47440 3004 47480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 55112 3004 55152 3044
rect 55194 3004 55234 3044
rect 55276 3004 55316 3044
rect 55358 3004 55398 3044
rect 55440 3004 55480 3044
rect 59112 3004 59152 3044
rect 59194 3004 59234 3044
rect 59276 3004 59316 3044
rect 59358 3004 59398 3044
rect 59440 3004 59480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 67112 3004 67152 3044
rect 67194 3004 67234 3044
rect 67276 3004 67316 3044
rect 67358 3004 67398 3044
rect 67440 3004 67480 3044
rect 71112 3004 71152 3044
rect 71194 3004 71234 3044
rect 71276 3004 71316 3044
rect 71358 3004 71398 3044
rect 71440 3004 71480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 79112 3004 79152 3044
rect 79194 3004 79234 3044
rect 79276 3004 79316 3044
rect 79358 3004 79398 3044
rect 79440 3004 79480 3044
rect 83112 3004 83152 3044
rect 83194 3004 83234 3044
rect 83276 3004 83316 3044
rect 83358 3004 83398 3044
rect 83440 3004 83480 3044
rect 87112 3004 87152 3044
rect 87194 3004 87234 3044
rect 87276 3004 87316 3044
rect 87358 3004 87398 3044
rect 87440 3004 87480 3044
rect 91112 3004 91152 3044
rect 91194 3004 91234 3044
rect 91276 3004 91316 3044
rect 91358 3004 91398 3044
rect 91440 3004 91480 3044
rect 95112 3004 95152 3044
rect 95194 3004 95234 3044
rect 95276 3004 95316 3044
rect 95358 3004 95398 3044
rect 95440 3004 95480 3044
rect 99112 3004 99152 3044
rect 99194 3004 99234 3044
rect 99276 3004 99316 3044
rect 99358 3004 99398 3044
rect 99440 3004 99480 3044
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 8352 2248 8392 2288
rect 8434 2248 8474 2288
rect 8516 2248 8556 2288
rect 8598 2248 8638 2288
rect 8680 2248 8720 2288
rect 12352 2248 12392 2288
rect 12434 2248 12474 2288
rect 12516 2248 12556 2288
rect 12598 2248 12638 2288
rect 12680 2248 12720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 20352 2248 20392 2288
rect 20434 2248 20474 2288
rect 20516 2248 20556 2288
rect 20598 2248 20638 2288
rect 20680 2248 20720 2288
rect 24352 2248 24392 2288
rect 24434 2248 24474 2288
rect 24516 2248 24556 2288
rect 24598 2248 24638 2288
rect 24680 2248 24720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 32352 2248 32392 2288
rect 32434 2248 32474 2288
rect 32516 2248 32556 2288
rect 32598 2248 32638 2288
rect 32680 2248 32720 2288
rect 36352 2248 36392 2288
rect 36434 2248 36474 2288
rect 36516 2248 36556 2288
rect 36598 2248 36638 2288
rect 36680 2248 36720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 44352 2248 44392 2288
rect 44434 2248 44474 2288
rect 44516 2248 44556 2288
rect 44598 2248 44638 2288
rect 44680 2248 44720 2288
rect 48352 2248 48392 2288
rect 48434 2248 48474 2288
rect 48516 2248 48556 2288
rect 48598 2248 48638 2288
rect 48680 2248 48720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 56352 2248 56392 2288
rect 56434 2248 56474 2288
rect 56516 2248 56556 2288
rect 56598 2248 56638 2288
rect 56680 2248 56720 2288
rect 60352 2248 60392 2288
rect 60434 2248 60474 2288
rect 60516 2248 60556 2288
rect 60598 2248 60638 2288
rect 60680 2248 60720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 68352 2248 68392 2288
rect 68434 2248 68474 2288
rect 68516 2248 68556 2288
rect 68598 2248 68638 2288
rect 68680 2248 68720 2288
rect 72352 2248 72392 2288
rect 72434 2248 72474 2288
rect 72516 2248 72556 2288
rect 72598 2248 72638 2288
rect 72680 2248 72720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 80352 2248 80392 2288
rect 80434 2248 80474 2288
rect 80516 2248 80556 2288
rect 80598 2248 80638 2288
rect 80680 2248 80720 2288
rect 84352 2248 84392 2288
rect 84434 2248 84474 2288
rect 84516 2248 84556 2288
rect 84598 2248 84638 2288
rect 84680 2248 84720 2288
rect 88352 2248 88392 2288
rect 88434 2248 88474 2288
rect 88516 2248 88556 2288
rect 88598 2248 88638 2288
rect 88680 2248 88720 2288
rect 92352 2248 92392 2288
rect 92434 2248 92474 2288
rect 92516 2248 92556 2288
rect 92598 2248 92638 2288
rect 92680 2248 92720 2288
rect 96352 2248 96392 2288
rect 96434 2248 96474 2288
rect 96516 2248 96556 2288
rect 96598 2248 96638 2288
rect 96680 2248 96720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 7112 1492 7152 1532
rect 7194 1492 7234 1532
rect 7276 1492 7316 1532
rect 7358 1492 7398 1532
rect 7440 1492 7480 1532
rect 11112 1492 11152 1532
rect 11194 1492 11234 1532
rect 11276 1492 11316 1532
rect 11358 1492 11398 1532
rect 11440 1492 11480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 19112 1492 19152 1532
rect 19194 1492 19234 1532
rect 19276 1492 19316 1532
rect 19358 1492 19398 1532
rect 19440 1492 19480 1532
rect 23112 1492 23152 1532
rect 23194 1492 23234 1532
rect 23276 1492 23316 1532
rect 23358 1492 23398 1532
rect 23440 1492 23480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 31112 1492 31152 1532
rect 31194 1492 31234 1532
rect 31276 1492 31316 1532
rect 31358 1492 31398 1532
rect 31440 1492 31480 1532
rect 35112 1492 35152 1532
rect 35194 1492 35234 1532
rect 35276 1492 35316 1532
rect 35358 1492 35398 1532
rect 35440 1492 35480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 43112 1492 43152 1532
rect 43194 1492 43234 1532
rect 43276 1492 43316 1532
rect 43358 1492 43398 1532
rect 43440 1492 43480 1532
rect 47112 1492 47152 1532
rect 47194 1492 47234 1532
rect 47276 1492 47316 1532
rect 47358 1492 47398 1532
rect 47440 1492 47480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 55112 1492 55152 1532
rect 55194 1492 55234 1532
rect 55276 1492 55316 1532
rect 55358 1492 55398 1532
rect 55440 1492 55480 1532
rect 59112 1492 59152 1532
rect 59194 1492 59234 1532
rect 59276 1492 59316 1532
rect 59358 1492 59398 1532
rect 59440 1492 59480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 67112 1492 67152 1532
rect 67194 1492 67234 1532
rect 67276 1492 67316 1532
rect 67358 1492 67398 1532
rect 67440 1492 67480 1532
rect 71112 1492 71152 1532
rect 71194 1492 71234 1532
rect 71276 1492 71316 1532
rect 71358 1492 71398 1532
rect 71440 1492 71480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 79112 1492 79152 1532
rect 79194 1492 79234 1532
rect 79276 1492 79316 1532
rect 79358 1492 79398 1532
rect 79440 1492 79480 1532
rect 83112 1492 83152 1532
rect 83194 1492 83234 1532
rect 83276 1492 83316 1532
rect 83358 1492 83398 1532
rect 83440 1492 83480 1532
rect 87112 1492 87152 1532
rect 87194 1492 87234 1532
rect 87276 1492 87316 1532
rect 87358 1492 87398 1532
rect 87440 1492 87480 1532
rect 91112 1492 91152 1532
rect 91194 1492 91234 1532
rect 91276 1492 91316 1532
rect 91358 1492 91398 1532
rect 91440 1492 91480 1532
rect 95112 1492 95152 1532
rect 95194 1492 95234 1532
rect 95276 1492 95316 1532
rect 95358 1492 95398 1532
rect 95440 1492 95480 1532
rect 99112 1492 99152 1532
rect 99194 1492 99234 1532
rect 99276 1492 99316 1532
rect 99358 1492 99398 1532
rect 99440 1492 99480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 8352 736 8392 776
rect 8434 736 8474 776
rect 8516 736 8556 776
rect 8598 736 8638 776
rect 8680 736 8720 776
rect 12352 736 12392 776
rect 12434 736 12474 776
rect 12516 736 12556 776
rect 12598 736 12638 776
rect 12680 736 12720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 20352 736 20392 776
rect 20434 736 20474 776
rect 20516 736 20556 776
rect 20598 736 20638 776
rect 20680 736 20720 776
rect 24352 736 24392 776
rect 24434 736 24474 776
rect 24516 736 24556 776
rect 24598 736 24638 776
rect 24680 736 24720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 32352 736 32392 776
rect 32434 736 32474 776
rect 32516 736 32556 776
rect 32598 736 32638 776
rect 32680 736 32720 776
rect 36352 736 36392 776
rect 36434 736 36474 776
rect 36516 736 36556 776
rect 36598 736 36638 776
rect 36680 736 36720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 44352 736 44392 776
rect 44434 736 44474 776
rect 44516 736 44556 776
rect 44598 736 44638 776
rect 44680 736 44720 776
rect 48352 736 48392 776
rect 48434 736 48474 776
rect 48516 736 48556 776
rect 48598 736 48638 776
rect 48680 736 48720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 56352 736 56392 776
rect 56434 736 56474 776
rect 56516 736 56556 776
rect 56598 736 56638 776
rect 56680 736 56720 776
rect 60352 736 60392 776
rect 60434 736 60474 776
rect 60516 736 60556 776
rect 60598 736 60638 776
rect 60680 736 60720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 68352 736 68392 776
rect 68434 736 68474 776
rect 68516 736 68556 776
rect 68598 736 68638 776
rect 68680 736 68720 776
rect 72352 736 72392 776
rect 72434 736 72474 776
rect 72516 736 72556 776
rect 72598 736 72638 776
rect 72680 736 72720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
rect 80352 736 80392 776
rect 80434 736 80474 776
rect 80516 736 80556 776
rect 80598 736 80638 776
rect 80680 736 80720 776
rect 84352 736 84392 776
rect 84434 736 84474 776
rect 84516 736 84556 776
rect 84598 736 84638 776
rect 84680 736 84720 776
rect 88352 736 88392 776
rect 88434 736 88474 776
rect 88516 736 88556 776
rect 88598 736 88638 776
rect 88680 736 88720 776
rect 92352 736 92392 776
rect 92434 736 92474 776
rect 92516 736 92556 776
rect 92598 736 92638 776
rect 92680 736 92720 776
rect 96352 736 96392 776
rect 96434 736 96474 776
rect 96516 736 96556 776
rect 96598 736 96638 776
rect 96680 736 96720 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 8343 38536 8352 38576
rect 8392 38536 8434 38576
rect 8474 38536 8516 38576
rect 8556 38536 8598 38576
rect 8638 38536 8680 38576
rect 8720 38536 8729 38576
rect 12343 38536 12352 38576
rect 12392 38536 12434 38576
rect 12474 38536 12516 38576
rect 12556 38536 12598 38576
rect 12638 38536 12680 38576
rect 12720 38536 12729 38576
rect 16343 38536 16352 38576
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16720 38536 16729 38576
rect 20343 38536 20352 38576
rect 20392 38536 20434 38576
rect 20474 38536 20516 38576
rect 20556 38536 20598 38576
rect 20638 38536 20680 38576
rect 20720 38536 20729 38576
rect 24343 38536 24352 38576
rect 24392 38536 24434 38576
rect 24474 38536 24516 38576
rect 24556 38536 24598 38576
rect 24638 38536 24680 38576
rect 24720 38536 24729 38576
rect 28343 38536 28352 38576
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28720 38536 28729 38576
rect 32343 38536 32352 38576
rect 32392 38536 32434 38576
rect 32474 38536 32516 38576
rect 32556 38536 32598 38576
rect 32638 38536 32680 38576
rect 32720 38536 32729 38576
rect 36343 38536 36352 38576
rect 36392 38536 36434 38576
rect 36474 38536 36516 38576
rect 36556 38536 36598 38576
rect 36638 38536 36680 38576
rect 36720 38536 36729 38576
rect 40343 38536 40352 38576
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40720 38536 40729 38576
rect 44343 38536 44352 38576
rect 44392 38536 44434 38576
rect 44474 38536 44516 38576
rect 44556 38536 44598 38576
rect 44638 38536 44680 38576
rect 44720 38536 44729 38576
rect 48343 38536 48352 38576
rect 48392 38536 48434 38576
rect 48474 38536 48516 38576
rect 48556 38536 48598 38576
rect 48638 38536 48680 38576
rect 48720 38536 48729 38576
rect 52343 38536 52352 38576
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52720 38536 52729 38576
rect 56343 38536 56352 38576
rect 56392 38536 56434 38576
rect 56474 38536 56516 38576
rect 56556 38536 56598 38576
rect 56638 38536 56680 38576
rect 56720 38536 56729 38576
rect 60343 38536 60352 38576
rect 60392 38536 60434 38576
rect 60474 38536 60516 38576
rect 60556 38536 60598 38576
rect 60638 38536 60680 38576
rect 60720 38536 60729 38576
rect 64343 38536 64352 38576
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64720 38536 64729 38576
rect 68343 38536 68352 38576
rect 68392 38536 68434 38576
rect 68474 38536 68516 38576
rect 68556 38536 68598 38576
rect 68638 38536 68680 38576
rect 68720 38536 68729 38576
rect 72343 38536 72352 38576
rect 72392 38536 72434 38576
rect 72474 38536 72516 38576
rect 72556 38536 72598 38576
rect 72638 38536 72680 38576
rect 72720 38536 72729 38576
rect 76343 38536 76352 38576
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76720 38536 76729 38576
rect 80343 38536 80352 38576
rect 80392 38536 80434 38576
rect 80474 38536 80516 38576
rect 80556 38536 80598 38576
rect 80638 38536 80680 38576
rect 80720 38536 80729 38576
rect 84343 38536 84352 38576
rect 84392 38536 84434 38576
rect 84474 38536 84516 38576
rect 84556 38536 84598 38576
rect 84638 38536 84680 38576
rect 84720 38536 84729 38576
rect 88343 38536 88352 38576
rect 88392 38536 88434 38576
rect 88474 38536 88516 38576
rect 88556 38536 88598 38576
rect 88638 38536 88680 38576
rect 88720 38536 88729 38576
rect 92343 38536 92352 38576
rect 92392 38536 92434 38576
rect 92474 38536 92516 38576
rect 92556 38536 92598 38576
rect 92638 38536 92680 38576
rect 92720 38536 92729 38576
rect 96343 38536 96352 38576
rect 96392 38536 96434 38576
rect 96474 38536 96516 38576
rect 96556 38536 96598 38576
rect 96638 38536 96680 38576
rect 96720 38536 96729 38576
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 7103 37780 7112 37820
rect 7152 37780 7194 37820
rect 7234 37780 7276 37820
rect 7316 37780 7358 37820
rect 7398 37780 7440 37820
rect 7480 37780 7489 37820
rect 11103 37780 11112 37820
rect 11152 37780 11194 37820
rect 11234 37780 11276 37820
rect 11316 37780 11358 37820
rect 11398 37780 11440 37820
rect 11480 37780 11489 37820
rect 15103 37780 15112 37820
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15480 37780 15489 37820
rect 19103 37780 19112 37820
rect 19152 37780 19194 37820
rect 19234 37780 19276 37820
rect 19316 37780 19358 37820
rect 19398 37780 19440 37820
rect 19480 37780 19489 37820
rect 23103 37780 23112 37820
rect 23152 37780 23194 37820
rect 23234 37780 23276 37820
rect 23316 37780 23358 37820
rect 23398 37780 23440 37820
rect 23480 37780 23489 37820
rect 27103 37780 27112 37820
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27480 37780 27489 37820
rect 31103 37780 31112 37820
rect 31152 37780 31194 37820
rect 31234 37780 31276 37820
rect 31316 37780 31358 37820
rect 31398 37780 31440 37820
rect 31480 37780 31489 37820
rect 35103 37780 35112 37820
rect 35152 37780 35194 37820
rect 35234 37780 35276 37820
rect 35316 37780 35358 37820
rect 35398 37780 35440 37820
rect 35480 37780 35489 37820
rect 39103 37780 39112 37820
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39480 37780 39489 37820
rect 43103 37780 43112 37820
rect 43152 37780 43194 37820
rect 43234 37780 43276 37820
rect 43316 37780 43358 37820
rect 43398 37780 43440 37820
rect 43480 37780 43489 37820
rect 47103 37780 47112 37820
rect 47152 37780 47194 37820
rect 47234 37780 47276 37820
rect 47316 37780 47358 37820
rect 47398 37780 47440 37820
rect 47480 37780 47489 37820
rect 51103 37780 51112 37820
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51480 37780 51489 37820
rect 55103 37780 55112 37820
rect 55152 37780 55194 37820
rect 55234 37780 55276 37820
rect 55316 37780 55358 37820
rect 55398 37780 55440 37820
rect 55480 37780 55489 37820
rect 59103 37780 59112 37820
rect 59152 37780 59194 37820
rect 59234 37780 59276 37820
rect 59316 37780 59358 37820
rect 59398 37780 59440 37820
rect 59480 37780 59489 37820
rect 63103 37780 63112 37820
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63480 37780 63489 37820
rect 67103 37780 67112 37820
rect 67152 37780 67194 37820
rect 67234 37780 67276 37820
rect 67316 37780 67358 37820
rect 67398 37780 67440 37820
rect 67480 37780 67489 37820
rect 71103 37780 71112 37820
rect 71152 37780 71194 37820
rect 71234 37780 71276 37820
rect 71316 37780 71358 37820
rect 71398 37780 71440 37820
rect 71480 37780 71489 37820
rect 75103 37780 75112 37820
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75480 37780 75489 37820
rect 79103 37780 79112 37820
rect 79152 37780 79194 37820
rect 79234 37780 79276 37820
rect 79316 37780 79358 37820
rect 79398 37780 79440 37820
rect 79480 37780 79489 37820
rect 83103 37780 83112 37820
rect 83152 37780 83194 37820
rect 83234 37780 83276 37820
rect 83316 37780 83358 37820
rect 83398 37780 83440 37820
rect 83480 37780 83489 37820
rect 87103 37780 87112 37820
rect 87152 37780 87194 37820
rect 87234 37780 87276 37820
rect 87316 37780 87358 37820
rect 87398 37780 87440 37820
rect 87480 37780 87489 37820
rect 91103 37780 91112 37820
rect 91152 37780 91194 37820
rect 91234 37780 91276 37820
rect 91316 37780 91358 37820
rect 91398 37780 91440 37820
rect 91480 37780 91489 37820
rect 95103 37780 95112 37820
rect 95152 37780 95194 37820
rect 95234 37780 95276 37820
rect 95316 37780 95358 37820
rect 95398 37780 95440 37820
rect 95480 37780 95489 37820
rect 99103 37780 99112 37820
rect 99152 37780 99194 37820
rect 99234 37780 99276 37820
rect 99316 37780 99358 37820
rect 99398 37780 99440 37820
rect 99480 37780 99489 37820
rect 0 37508 80 37588
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 8343 37024 8352 37064
rect 8392 37024 8434 37064
rect 8474 37024 8516 37064
rect 8556 37024 8598 37064
rect 8638 37024 8680 37064
rect 8720 37024 8729 37064
rect 12343 37024 12352 37064
rect 12392 37024 12434 37064
rect 12474 37024 12516 37064
rect 12556 37024 12598 37064
rect 12638 37024 12680 37064
rect 12720 37024 12729 37064
rect 16343 37024 16352 37064
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16720 37024 16729 37064
rect 20343 37024 20352 37064
rect 20392 37024 20434 37064
rect 20474 37024 20516 37064
rect 20556 37024 20598 37064
rect 20638 37024 20680 37064
rect 20720 37024 20729 37064
rect 24343 37024 24352 37064
rect 24392 37024 24434 37064
rect 24474 37024 24516 37064
rect 24556 37024 24598 37064
rect 24638 37024 24680 37064
rect 24720 37024 24729 37064
rect 28343 37024 28352 37064
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28720 37024 28729 37064
rect 32343 37024 32352 37064
rect 32392 37024 32434 37064
rect 32474 37024 32516 37064
rect 32556 37024 32598 37064
rect 32638 37024 32680 37064
rect 32720 37024 32729 37064
rect 36343 37024 36352 37064
rect 36392 37024 36434 37064
rect 36474 37024 36516 37064
rect 36556 37024 36598 37064
rect 36638 37024 36680 37064
rect 36720 37024 36729 37064
rect 40343 37024 40352 37064
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40720 37024 40729 37064
rect 44343 37024 44352 37064
rect 44392 37024 44434 37064
rect 44474 37024 44516 37064
rect 44556 37024 44598 37064
rect 44638 37024 44680 37064
rect 44720 37024 44729 37064
rect 48343 37024 48352 37064
rect 48392 37024 48434 37064
rect 48474 37024 48516 37064
rect 48556 37024 48598 37064
rect 48638 37024 48680 37064
rect 48720 37024 48729 37064
rect 52343 37024 52352 37064
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52720 37024 52729 37064
rect 56343 37024 56352 37064
rect 56392 37024 56434 37064
rect 56474 37024 56516 37064
rect 56556 37024 56598 37064
rect 56638 37024 56680 37064
rect 56720 37024 56729 37064
rect 60343 37024 60352 37064
rect 60392 37024 60434 37064
rect 60474 37024 60516 37064
rect 60556 37024 60598 37064
rect 60638 37024 60680 37064
rect 60720 37024 60729 37064
rect 64343 37024 64352 37064
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64720 37024 64729 37064
rect 68343 37024 68352 37064
rect 68392 37024 68434 37064
rect 68474 37024 68516 37064
rect 68556 37024 68598 37064
rect 68638 37024 68680 37064
rect 68720 37024 68729 37064
rect 72343 37024 72352 37064
rect 72392 37024 72434 37064
rect 72474 37024 72516 37064
rect 72556 37024 72598 37064
rect 72638 37024 72680 37064
rect 72720 37024 72729 37064
rect 76343 37024 76352 37064
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76720 37024 76729 37064
rect 80343 37024 80352 37064
rect 80392 37024 80434 37064
rect 80474 37024 80516 37064
rect 80556 37024 80598 37064
rect 80638 37024 80680 37064
rect 80720 37024 80729 37064
rect 84343 37024 84352 37064
rect 84392 37024 84434 37064
rect 84474 37024 84516 37064
rect 84556 37024 84598 37064
rect 84638 37024 84680 37064
rect 84720 37024 84729 37064
rect 88343 37024 88352 37064
rect 88392 37024 88434 37064
rect 88474 37024 88516 37064
rect 88556 37024 88598 37064
rect 88638 37024 88680 37064
rect 88720 37024 88729 37064
rect 92343 37024 92352 37064
rect 92392 37024 92434 37064
rect 92474 37024 92516 37064
rect 92556 37024 92598 37064
rect 92638 37024 92680 37064
rect 92720 37024 92729 37064
rect 96343 37024 96352 37064
rect 96392 37024 96434 37064
rect 96474 37024 96516 37064
rect 96556 37024 96598 37064
rect 96638 37024 96680 37064
rect 96720 37024 96729 37064
rect 0 36668 80 36748
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 7103 36268 7112 36308
rect 7152 36268 7194 36308
rect 7234 36268 7276 36308
rect 7316 36268 7358 36308
rect 7398 36268 7440 36308
rect 7480 36268 7489 36308
rect 11103 36268 11112 36308
rect 11152 36268 11194 36308
rect 11234 36268 11276 36308
rect 11316 36268 11358 36308
rect 11398 36268 11440 36308
rect 11480 36268 11489 36308
rect 15103 36268 15112 36308
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15480 36268 15489 36308
rect 19103 36268 19112 36308
rect 19152 36268 19194 36308
rect 19234 36268 19276 36308
rect 19316 36268 19358 36308
rect 19398 36268 19440 36308
rect 19480 36268 19489 36308
rect 23103 36268 23112 36308
rect 23152 36268 23194 36308
rect 23234 36268 23276 36308
rect 23316 36268 23358 36308
rect 23398 36268 23440 36308
rect 23480 36268 23489 36308
rect 27103 36268 27112 36308
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27480 36268 27489 36308
rect 31103 36268 31112 36308
rect 31152 36268 31194 36308
rect 31234 36268 31276 36308
rect 31316 36268 31358 36308
rect 31398 36268 31440 36308
rect 31480 36268 31489 36308
rect 35103 36268 35112 36308
rect 35152 36268 35194 36308
rect 35234 36268 35276 36308
rect 35316 36268 35358 36308
rect 35398 36268 35440 36308
rect 35480 36268 35489 36308
rect 39103 36268 39112 36308
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39480 36268 39489 36308
rect 43103 36268 43112 36308
rect 43152 36268 43194 36308
rect 43234 36268 43276 36308
rect 43316 36268 43358 36308
rect 43398 36268 43440 36308
rect 43480 36268 43489 36308
rect 47103 36268 47112 36308
rect 47152 36268 47194 36308
rect 47234 36268 47276 36308
rect 47316 36268 47358 36308
rect 47398 36268 47440 36308
rect 47480 36268 47489 36308
rect 51103 36268 51112 36308
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51480 36268 51489 36308
rect 55103 36268 55112 36308
rect 55152 36268 55194 36308
rect 55234 36268 55276 36308
rect 55316 36268 55358 36308
rect 55398 36268 55440 36308
rect 55480 36268 55489 36308
rect 59103 36268 59112 36308
rect 59152 36268 59194 36308
rect 59234 36268 59276 36308
rect 59316 36268 59358 36308
rect 59398 36268 59440 36308
rect 59480 36268 59489 36308
rect 63103 36268 63112 36308
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63480 36268 63489 36308
rect 67103 36268 67112 36308
rect 67152 36268 67194 36308
rect 67234 36268 67276 36308
rect 67316 36268 67358 36308
rect 67398 36268 67440 36308
rect 67480 36268 67489 36308
rect 71103 36268 71112 36308
rect 71152 36268 71194 36308
rect 71234 36268 71276 36308
rect 71316 36268 71358 36308
rect 71398 36268 71440 36308
rect 71480 36268 71489 36308
rect 75103 36268 75112 36308
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75480 36268 75489 36308
rect 79103 36268 79112 36308
rect 79152 36268 79194 36308
rect 79234 36268 79276 36308
rect 79316 36268 79358 36308
rect 79398 36268 79440 36308
rect 79480 36268 79489 36308
rect 83103 36268 83112 36308
rect 83152 36268 83194 36308
rect 83234 36268 83276 36308
rect 83316 36268 83358 36308
rect 83398 36268 83440 36308
rect 83480 36268 83489 36308
rect 87103 36268 87112 36308
rect 87152 36268 87194 36308
rect 87234 36268 87276 36308
rect 87316 36268 87358 36308
rect 87398 36268 87440 36308
rect 87480 36268 87489 36308
rect 91103 36268 91112 36308
rect 91152 36268 91194 36308
rect 91234 36268 91276 36308
rect 91316 36268 91358 36308
rect 91398 36268 91440 36308
rect 91480 36268 91489 36308
rect 95103 36268 95112 36308
rect 95152 36268 95194 36308
rect 95234 36268 95276 36308
rect 95316 36268 95358 36308
rect 95398 36268 95440 36308
rect 95480 36268 95489 36308
rect 99103 36268 99112 36308
rect 99152 36268 99194 36308
rect 99234 36268 99276 36308
rect 99316 36268 99358 36308
rect 99398 36268 99440 36308
rect 99480 36268 99489 36308
rect 0 35828 80 35908
rect 76771 35720 76829 35721
rect 85219 35720 85277 35721
rect 76686 35680 76780 35720
rect 76820 35680 76829 35720
rect 85134 35680 85228 35720
rect 85268 35680 85277 35720
rect 76771 35679 76829 35680
rect 85219 35679 85277 35680
rect 92227 35720 92285 35721
rect 92227 35680 92236 35720
rect 92276 35680 92428 35720
rect 92468 35680 92477 35720
rect 92227 35679 92285 35680
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 8343 35512 8352 35552
rect 8392 35512 8434 35552
rect 8474 35512 8516 35552
rect 8556 35512 8598 35552
rect 8638 35512 8680 35552
rect 8720 35512 8729 35552
rect 12343 35512 12352 35552
rect 12392 35512 12434 35552
rect 12474 35512 12516 35552
rect 12556 35512 12598 35552
rect 12638 35512 12680 35552
rect 12720 35512 12729 35552
rect 16343 35512 16352 35552
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16720 35512 16729 35552
rect 20343 35512 20352 35552
rect 20392 35512 20434 35552
rect 20474 35512 20516 35552
rect 20556 35512 20598 35552
rect 20638 35512 20680 35552
rect 20720 35512 20729 35552
rect 24343 35512 24352 35552
rect 24392 35512 24434 35552
rect 24474 35512 24516 35552
rect 24556 35512 24598 35552
rect 24638 35512 24680 35552
rect 24720 35512 24729 35552
rect 28343 35512 28352 35552
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28720 35512 28729 35552
rect 32343 35512 32352 35552
rect 32392 35512 32434 35552
rect 32474 35512 32516 35552
rect 32556 35512 32598 35552
rect 32638 35512 32680 35552
rect 32720 35512 32729 35552
rect 36343 35512 36352 35552
rect 36392 35512 36434 35552
rect 36474 35512 36516 35552
rect 36556 35512 36598 35552
rect 36638 35512 36680 35552
rect 36720 35512 36729 35552
rect 40343 35512 40352 35552
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40720 35512 40729 35552
rect 44343 35512 44352 35552
rect 44392 35512 44434 35552
rect 44474 35512 44516 35552
rect 44556 35512 44598 35552
rect 44638 35512 44680 35552
rect 44720 35512 44729 35552
rect 48343 35512 48352 35552
rect 48392 35512 48434 35552
rect 48474 35512 48516 35552
rect 48556 35512 48598 35552
rect 48638 35512 48680 35552
rect 48720 35512 48729 35552
rect 52343 35512 52352 35552
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52720 35512 52729 35552
rect 56343 35512 56352 35552
rect 56392 35512 56434 35552
rect 56474 35512 56516 35552
rect 56556 35512 56598 35552
rect 56638 35512 56680 35552
rect 56720 35512 56729 35552
rect 60343 35512 60352 35552
rect 60392 35512 60434 35552
rect 60474 35512 60516 35552
rect 60556 35512 60598 35552
rect 60638 35512 60680 35552
rect 60720 35512 60729 35552
rect 64343 35512 64352 35552
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64720 35512 64729 35552
rect 68343 35512 68352 35552
rect 68392 35512 68434 35552
rect 68474 35512 68516 35552
rect 68556 35512 68598 35552
rect 68638 35512 68680 35552
rect 68720 35512 68729 35552
rect 72343 35512 72352 35552
rect 72392 35512 72434 35552
rect 72474 35512 72516 35552
rect 72556 35512 72598 35552
rect 72638 35512 72680 35552
rect 72720 35512 72729 35552
rect 76343 35512 76352 35552
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76720 35512 76729 35552
rect 80343 35512 80352 35552
rect 80392 35512 80434 35552
rect 80474 35512 80516 35552
rect 80556 35512 80598 35552
rect 80638 35512 80680 35552
rect 80720 35512 80729 35552
rect 84343 35512 84352 35552
rect 84392 35512 84434 35552
rect 84474 35512 84516 35552
rect 84556 35512 84598 35552
rect 84638 35512 84680 35552
rect 84720 35512 84729 35552
rect 88343 35512 88352 35552
rect 88392 35512 88434 35552
rect 88474 35512 88516 35552
rect 88556 35512 88598 35552
rect 88638 35512 88680 35552
rect 88720 35512 88729 35552
rect 92343 35512 92352 35552
rect 92392 35512 92434 35552
rect 92474 35512 92516 35552
rect 92556 35512 92598 35552
rect 92638 35512 92680 35552
rect 92720 35512 92729 35552
rect 96343 35512 96352 35552
rect 96392 35512 96434 35552
rect 96474 35512 96516 35552
rect 96556 35512 96598 35552
rect 96638 35512 96680 35552
rect 96720 35512 96729 35552
rect 89923 35300 89981 35301
rect 89838 35260 89932 35300
rect 89972 35260 89981 35300
rect 89923 35259 89981 35260
rect 76195 35176 76204 35216
rect 76244 35176 76684 35216
rect 76724 35176 76733 35216
rect 77251 35176 77260 35216
rect 77300 35176 77548 35216
rect 77588 35176 77836 35216
rect 77876 35176 77885 35216
rect 83875 35176 83884 35216
rect 83924 35176 84268 35216
rect 84308 35176 84652 35216
rect 84692 35176 84701 35216
rect 87619 35176 87628 35216
rect 87668 35176 88108 35216
rect 88148 35176 88492 35216
rect 88532 35176 88541 35216
rect 83884 35132 83924 35176
rect 73891 35092 73900 35132
rect 73940 35092 74092 35132
rect 74132 35092 74860 35132
rect 74900 35092 74909 35132
rect 75619 35092 75628 35132
rect 75668 35092 76108 35132
rect 76148 35092 76588 35132
rect 76628 35092 77068 35132
rect 77108 35092 78988 35132
rect 79028 35092 79037 35132
rect 81571 35092 81580 35132
rect 81620 35092 81772 35132
rect 81812 35092 82348 35132
rect 82388 35092 82397 35132
rect 82627 35092 82636 35132
rect 82676 35092 82685 35132
rect 83299 35092 83308 35132
rect 83348 35092 83500 35132
rect 83540 35092 83924 35132
rect 86083 35092 86092 35132
rect 86132 35092 86380 35132
rect 86420 35092 86572 35132
rect 86612 35092 87052 35132
rect 87092 35092 87436 35132
rect 87476 35092 88684 35132
rect 88724 35092 88733 35132
rect 89923 35092 89932 35132
rect 89972 35092 90220 35132
rect 90260 35092 90269 35132
rect 90673 35092 90682 35132
rect 90722 35092 91084 35132
rect 91124 35092 91468 35132
rect 91508 35092 91756 35132
rect 91796 35092 91805 35132
rect 92227 35092 92236 35132
rect 92276 35092 92428 35132
rect 92468 35092 92620 35132
rect 92660 35092 93100 35132
rect 93140 35092 93149 35132
rect 95203 35092 95212 35132
rect 95252 35092 95404 35132
rect 95444 35092 95884 35132
rect 95924 35092 96172 35132
rect 96212 35092 97804 35132
rect 97844 35092 97853 35132
rect 0 34988 80 35068
rect 75628 35048 75668 35092
rect 82636 35048 82676 35092
rect 73699 35008 73708 35048
rect 73748 35008 74476 35048
rect 74516 35008 75668 35048
rect 80131 35008 80140 35048
rect 80180 35008 80428 35048
rect 80468 35008 80620 35048
rect 80660 35008 80908 35048
rect 80948 35008 81388 35048
rect 81428 35008 82676 35048
rect 86467 35008 86476 35048
rect 86516 35008 87916 35048
rect 87956 35008 89356 35048
rect 89396 35008 89405 35048
rect 86659 34964 86717 34965
rect 86574 34924 86668 34964
rect 86708 34924 86717 34964
rect 86659 34923 86717 34924
rect 86947 34964 87005 34965
rect 86947 34924 86956 34964
rect 86996 34924 87244 34964
rect 87284 34924 87293 34964
rect 87715 34924 87724 34964
rect 87764 34924 88300 34964
rect 88340 34924 88349 34964
rect 95107 34924 95116 34964
rect 95156 34924 95788 34964
rect 95828 34924 95837 34964
rect 96163 34924 96172 34964
rect 96212 34924 96940 34964
rect 96980 34924 96989 34964
rect 86947 34923 87005 34924
rect 86668 34880 86708 34923
rect 86668 34840 90220 34880
rect 90260 34840 90269 34880
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 7103 34756 7112 34796
rect 7152 34756 7194 34796
rect 7234 34756 7276 34796
rect 7316 34756 7358 34796
rect 7398 34756 7440 34796
rect 7480 34756 7489 34796
rect 11103 34756 11112 34796
rect 11152 34756 11194 34796
rect 11234 34756 11276 34796
rect 11316 34756 11358 34796
rect 11398 34756 11440 34796
rect 11480 34756 11489 34796
rect 15103 34756 15112 34796
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15480 34756 15489 34796
rect 19103 34756 19112 34796
rect 19152 34756 19194 34796
rect 19234 34756 19276 34796
rect 19316 34756 19358 34796
rect 19398 34756 19440 34796
rect 19480 34756 19489 34796
rect 23103 34756 23112 34796
rect 23152 34756 23194 34796
rect 23234 34756 23276 34796
rect 23316 34756 23358 34796
rect 23398 34756 23440 34796
rect 23480 34756 23489 34796
rect 27103 34756 27112 34796
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27480 34756 27489 34796
rect 31103 34756 31112 34796
rect 31152 34756 31194 34796
rect 31234 34756 31276 34796
rect 31316 34756 31358 34796
rect 31398 34756 31440 34796
rect 31480 34756 31489 34796
rect 35103 34756 35112 34796
rect 35152 34756 35194 34796
rect 35234 34756 35276 34796
rect 35316 34756 35358 34796
rect 35398 34756 35440 34796
rect 35480 34756 35489 34796
rect 39103 34756 39112 34796
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39480 34756 39489 34796
rect 43103 34756 43112 34796
rect 43152 34756 43194 34796
rect 43234 34756 43276 34796
rect 43316 34756 43358 34796
rect 43398 34756 43440 34796
rect 43480 34756 43489 34796
rect 47103 34756 47112 34796
rect 47152 34756 47194 34796
rect 47234 34756 47276 34796
rect 47316 34756 47358 34796
rect 47398 34756 47440 34796
rect 47480 34756 47489 34796
rect 51103 34756 51112 34796
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51480 34756 51489 34796
rect 55103 34756 55112 34796
rect 55152 34756 55194 34796
rect 55234 34756 55276 34796
rect 55316 34756 55358 34796
rect 55398 34756 55440 34796
rect 55480 34756 55489 34796
rect 59103 34756 59112 34796
rect 59152 34756 59194 34796
rect 59234 34756 59276 34796
rect 59316 34756 59358 34796
rect 59398 34756 59440 34796
rect 59480 34756 59489 34796
rect 63103 34756 63112 34796
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63480 34756 63489 34796
rect 67103 34756 67112 34796
rect 67152 34756 67194 34796
rect 67234 34756 67276 34796
rect 67316 34756 67358 34796
rect 67398 34756 67440 34796
rect 67480 34756 67489 34796
rect 71103 34756 71112 34796
rect 71152 34756 71194 34796
rect 71234 34756 71276 34796
rect 71316 34756 71358 34796
rect 71398 34756 71440 34796
rect 71480 34756 71489 34796
rect 75103 34756 75112 34796
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75480 34756 75489 34796
rect 79103 34756 79112 34796
rect 79152 34756 79194 34796
rect 79234 34756 79276 34796
rect 79316 34756 79358 34796
rect 79398 34756 79440 34796
rect 79480 34756 79489 34796
rect 83103 34756 83112 34796
rect 83152 34756 83194 34796
rect 83234 34756 83276 34796
rect 83316 34756 83358 34796
rect 83398 34756 83440 34796
rect 83480 34756 83489 34796
rect 87103 34756 87112 34796
rect 87152 34756 87194 34796
rect 87234 34756 87276 34796
rect 87316 34756 87358 34796
rect 87398 34756 87440 34796
rect 87480 34756 87489 34796
rect 91103 34756 91112 34796
rect 91152 34756 91194 34796
rect 91234 34756 91276 34796
rect 91316 34756 91358 34796
rect 91398 34756 91440 34796
rect 91480 34756 91489 34796
rect 95103 34756 95112 34796
rect 95152 34756 95194 34796
rect 95234 34756 95276 34796
rect 95316 34756 95358 34796
rect 95398 34756 95440 34796
rect 95480 34756 95489 34796
rect 99103 34756 99112 34796
rect 99152 34756 99194 34796
rect 99234 34756 99276 34796
rect 99316 34756 99358 34796
rect 99398 34756 99440 34796
rect 99480 34756 99489 34796
rect 80227 34712 80285 34713
rect 80142 34672 80236 34712
rect 80276 34672 80285 34712
rect 80707 34672 80716 34712
rect 80756 34672 80765 34712
rect 80227 34671 80285 34672
rect 74659 34588 74668 34628
rect 74708 34588 80564 34628
rect 74851 34504 74860 34544
rect 74900 34504 74909 34544
rect 74860 34460 74900 34504
rect 69763 34420 69772 34460
rect 69812 34420 73420 34460
rect 73460 34420 73469 34460
rect 74860 34420 75148 34460
rect 75188 34420 75668 34460
rect 75628 34376 75668 34420
rect 75619 34336 75628 34376
rect 75668 34336 76204 34376
rect 76244 34336 76253 34376
rect 76963 34336 76972 34376
rect 77012 34336 77836 34376
rect 77876 34336 78220 34376
rect 78260 34336 78700 34376
rect 78740 34336 79756 34376
rect 79796 34336 79805 34376
rect 74467 34252 74476 34292
rect 74516 34252 74860 34292
rect 74900 34252 75916 34292
rect 75956 34252 77548 34292
rect 77588 34252 79276 34292
rect 79316 34252 79325 34292
rect 0 34148 80 34228
rect 80524 34208 80564 34588
rect 80716 34292 80756 34672
rect 86851 34628 86909 34629
rect 83299 34588 83308 34628
rect 83348 34588 83596 34628
rect 83636 34588 83884 34628
rect 83924 34588 84172 34628
rect 84212 34588 84221 34628
rect 85027 34588 85036 34628
rect 85076 34588 85116 34628
rect 86766 34588 86860 34628
rect 86900 34588 86909 34628
rect 85036 34544 85076 34588
rect 86851 34587 86909 34588
rect 82243 34504 82252 34544
rect 82292 34504 82636 34544
rect 82676 34504 82685 34544
rect 84643 34504 84652 34544
rect 84692 34504 85228 34544
rect 85268 34504 85420 34544
rect 85460 34504 85804 34544
rect 85844 34504 85853 34544
rect 90211 34504 90220 34544
rect 90260 34504 92620 34544
rect 92660 34504 92669 34544
rect 96835 34504 96844 34544
rect 96884 34504 97132 34544
rect 97172 34504 97181 34544
rect 80995 34420 81004 34460
rect 81044 34420 81196 34460
rect 81236 34420 81484 34460
rect 81524 34420 81868 34460
rect 81908 34420 83116 34460
rect 83156 34420 85036 34460
rect 85076 34420 85085 34460
rect 87811 34420 87820 34460
rect 87860 34420 88108 34460
rect 88148 34420 88300 34460
rect 88340 34420 88684 34460
rect 88724 34420 88733 34460
rect 90595 34420 90604 34460
rect 90644 34420 91180 34460
rect 91220 34420 91468 34460
rect 91508 34420 91756 34460
rect 91796 34420 91805 34460
rect 93091 34420 93100 34460
rect 93140 34420 93580 34460
rect 93620 34420 93629 34460
rect 93859 34420 93868 34460
rect 93908 34420 94060 34460
rect 94100 34420 94636 34460
rect 94676 34420 94685 34460
rect 96067 34420 96076 34460
rect 96116 34420 96460 34460
rect 96500 34420 97076 34460
rect 97507 34420 97516 34460
rect 97556 34420 97804 34460
rect 97844 34420 98324 34460
rect 97036 34376 97076 34420
rect 98284 34376 98324 34420
rect 81667 34336 81676 34376
rect 81716 34336 82156 34376
rect 82196 34336 82205 34376
rect 84739 34336 84748 34376
rect 84788 34336 84797 34376
rect 89155 34336 89164 34376
rect 89204 34336 89452 34376
rect 89492 34336 89644 34376
rect 89684 34336 89932 34376
rect 89972 34336 89981 34376
rect 92035 34336 92044 34376
rect 92084 34336 92236 34376
rect 92276 34336 92812 34376
rect 92852 34336 94252 34376
rect 94292 34336 95596 34376
rect 95636 34336 96268 34376
rect 96308 34336 96748 34376
rect 96788 34336 96797 34376
rect 97027 34336 97036 34376
rect 97076 34336 97900 34376
rect 97940 34336 97949 34376
rect 98275 34336 98284 34376
rect 98324 34336 98860 34376
rect 98900 34336 98909 34376
rect 84748 34292 84788 34336
rect 80716 34252 81004 34292
rect 81044 34252 81053 34292
rect 84172 34252 84788 34292
rect 89347 34252 89356 34292
rect 89396 34252 90988 34292
rect 91028 34252 91037 34292
rect 93571 34252 93580 34292
rect 93620 34252 95020 34292
rect 95060 34252 95069 34292
rect 76771 34168 76780 34208
rect 76820 34168 76829 34208
rect 78307 34168 78316 34208
rect 78356 34168 78604 34208
rect 78644 34168 78653 34208
rect 80323 34168 80332 34208
rect 80372 34168 80381 34208
rect 80524 34168 81920 34208
rect 83875 34168 83884 34208
rect 83924 34168 84076 34208
rect 84116 34168 84125 34208
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 8343 34000 8352 34040
rect 8392 34000 8434 34040
rect 8474 34000 8516 34040
rect 8556 34000 8598 34040
rect 8638 34000 8680 34040
rect 8720 34000 8729 34040
rect 12343 34000 12352 34040
rect 12392 34000 12434 34040
rect 12474 34000 12516 34040
rect 12556 34000 12598 34040
rect 12638 34000 12680 34040
rect 12720 34000 12729 34040
rect 16343 34000 16352 34040
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16720 34000 16729 34040
rect 20343 34000 20352 34040
rect 20392 34000 20434 34040
rect 20474 34000 20516 34040
rect 20556 34000 20598 34040
rect 20638 34000 20680 34040
rect 20720 34000 20729 34040
rect 24343 34000 24352 34040
rect 24392 34000 24434 34040
rect 24474 34000 24516 34040
rect 24556 34000 24598 34040
rect 24638 34000 24680 34040
rect 24720 34000 24729 34040
rect 28343 34000 28352 34040
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28720 34000 28729 34040
rect 32343 34000 32352 34040
rect 32392 34000 32434 34040
rect 32474 34000 32516 34040
rect 32556 34000 32598 34040
rect 32638 34000 32680 34040
rect 32720 34000 32729 34040
rect 36343 34000 36352 34040
rect 36392 34000 36434 34040
rect 36474 34000 36516 34040
rect 36556 34000 36598 34040
rect 36638 34000 36680 34040
rect 36720 34000 36729 34040
rect 40343 34000 40352 34040
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40720 34000 40729 34040
rect 44343 34000 44352 34040
rect 44392 34000 44434 34040
rect 44474 34000 44516 34040
rect 44556 34000 44598 34040
rect 44638 34000 44680 34040
rect 44720 34000 44729 34040
rect 48343 34000 48352 34040
rect 48392 34000 48434 34040
rect 48474 34000 48516 34040
rect 48556 34000 48598 34040
rect 48638 34000 48680 34040
rect 48720 34000 48729 34040
rect 52343 34000 52352 34040
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52720 34000 52729 34040
rect 56343 34000 56352 34040
rect 56392 34000 56434 34040
rect 56474 34000 56516 34040
rect 56556 34000 56598 34040
rect 56638 34000 56680 34040
rect 56720 34000 56729 34040
rect 60343 34000 60352 34040
rect 60392 34000 60434 34040
rect 60474 34000 60516 34040
rect 60556 34000 60598 34040
rect 60638 34000 60680 34040
rect 60720 34000 60729 34040
rect 64343 34000 64352 34040
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64720 34000 64729 34040
rect 68343 34000 68352 34040
rect 68392 34000 68434 34040
rect 68474 34000 68516 34040
rect 68556 34000 68598 34040
rect 68638 34000 68680 34040
rect 68720 34000 68729 34040
rect 72343 34000 72352 34040
rect 72392 34000 72434 34040
rect 72474 34000 72516 34040
rect 72556 34000 72598 34040
rect 72638 34000 72680 34040
rect 72720 34000 72729 34040
rect 76343 34000 76352 34040
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76720 34000 76729 34040
rect 76780 33872 76820 34168
rect 80332 34124 80372 34168
rect 76675 33832 76684 33872
rect 76724 33832 76820 33872
rect 80236 34084 80372 34124
rect 81880 34124 81920 34168
rect 84172 34124 84212 34252
rect 84355 34168 84364 34208
rect 84404 34168 84940 34208
rect 84980 34168 84989 34208
rect 86179 34168 86188 34208
rect 86228 34168 86764 34208
rect 86804 34168 86813 34208
rect 89059 34168 89068 34208
rect 89108 34168 89548 34208
rect 89588 34168 89597 34208
rect 90307 34168 90316 34208
rect 90356 34168 90604 34208
rect 90644 34168 90653 34208
rect 91939 34168 91948 34208
rect 91988 34168 92812 34208
rect 92852 34168 92861 34208
rect 93091 34168 93100 34208
rect 93140 34168 93484 34208
rect 93524 34168 93533 34208
rect 96643 34168 96652 34208
rect 96692 34168 96701 34208
rect 97891 34168 97900 34208
rect 97940 34168 98956 34208
rect 98996 34168 99005 34208
rect 96652 34124 96692 34168
rect 81880 34084 82060 34124
rect 82100 34084 82109 34124
rect 84163 34084 84172 34124
rect 84212 34084 84221 34124
rect 96652 34084 96940 34124
rect 96980 34084 96989 34124
rect 80236 33872 80276 34084
rect 80343 34000 80352 34040
rect 80392 34000 80434 34040
rect 80474 34000 80516 34040
rect 80556 34000 80598 34040
rect 80638 34000 80680 34040
rect 80720 34000 80729 34040
rect 83116 34000 83500 34040
rect 83540 34000 83549 34040
rect 84343 34000 84352 34040
rect 84392 34000 84434 34040
rect 84474 34000 84516 34040
rect 84556 34000 84598 34040
rect 84638 34000 84680 34040
rect 84720 34000 84729 34040
rect 87619 34000 87628 34040
rect 87668 34000 88244 34040
rect 88343 34000 88352 34040
rect 88392 34000 88434 34040
rect 88474 34000 88516 34040
rect 88556 34000 88598 34040
rect 88638 34000 88680 34040
rect 88720 34000 88729 34040
rect 92343 34000 92352 34040
rect 92392 34000 92434 34040
rect 92474 34000 92516 34040
rect 92556 34000 92598 34040
rect 92638 34000 92680 34040
rect 92720 34000 92729 34040
rect 96343 34000 96352 34040
rect 96392 34000 96434 34040
rect 96474 34000 96516 34040
rect 96556 34000 96598 34040
rect 96638 34000 96680 34040
rect 96720 34000 96729 34040
rect 96835 34000 96844 34040
rect 96884 34000 97996 34040
rect 98036 34000 98045 34040
rect 83116 33872 83156 34000
rect 88204 33872 88244 34000
rect 80236 33832 80428 33872
rect 80468 33832 80477 33872
rect 83107 33832 83116 33872
rect 83156 33832 83165 33872
rect 88204 33832 88300 33872
rect 88340 33832 88349 33872
rect 80227 33788 80285 33789
rect 80227 33748 80236 33788
rect 80276 33748 80332 33788
rect 80372 33748 80381 33788
rect 80227 33747 80285 33748
rect 0 33308 80 33388
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 7103 33244 7112 33284
rect 7152 33244 7194 33284
rect 7234 33244 7276 33284
rect 7316 33244 7358 33284
rect 7398 33244 7440 33284
rect 7480 33244 7489 33284
rect 11103 33244 11112 33284
rect 11152 33244 11194 33284
rect 11234 33244 11276 33284
rect 11316 33244 11358 33284
rect 11398 33244 11440 33284
rect 11480 33244 11489 33284
rect 15103 33244 15112 33284
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15480 33244 15489 33284
rect 19103 33244 19112 33284
rect 19152 33244 19194 33284
rect 19234 33244 19276 33284
rect 19316 33244 19358 33284
rect 19398 33244 19440 33284
rect 19480 33244 19489 33284
rect 23103 33244 23112 33284
rect 23152 33244 23194 33284
rect 23234 33244 23276 33284
rect 23316 33244 23358 33284
rect 23398 33244 23440 33284
rect 23480 33244 23489 33284
rect 27103 33244 27112 33284
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27480 33244 27489 33284
rect 31103 33244 31112 33284
rect 31152 33244 31194 33284
rect 31234 33244 31276 33284
rect 31316 33244 31358 33284
rect 31398 33244 31440 33284
rect 31480 33244 31489 33284
rect 35103 33244 35112 33284
rect 35152 33244 35194 33284
rect 35234 33244 35276 33284
rect 35316 33244 35358 33284
rect 35398 33244 35440 33284
rect 35480 33244 35489 33284
rect 39103 33244 39112 33284
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39480 33244 39489 33284
rect 43103 33244 43112 33284
rect 43152 33244 43194 33284
rect 43234 33244 43276 33284
rect 43316 33244 43358 33284
rect 43398 33244 43440 33284
rect 43480 33244 43489 33284
rect 47103 33244 47112 33284
rect 47152 33244 47194 33284
rect 47234 33244 47276 33284
rect 47316 33244 47358 33284
rect 47398 33244 47440 33284
rect 47480 33244 47489 33284
rect 51103 33244 51112 33284
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51480 33244 51489 33284
rect 55103 33244 55112 33284
rect 55152 33244 55194 33284
rect 55234 33244 55276 33284
rect 55316 33244 55358 33284
rect 55398 33244 55440 33284
rect 55480 33244 55489 33284
rect 59103 33244 59112 33284
rect 59152 33244 59194 33284
rect 59234 33244 59276 33284
rect 59316 33244 59358 33284
rect 59398 33244 59440 33284
rect 59480 33244 59489 33284
rect 63103 33244 63112 33284
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63480 33244 63489 33284
rect 67103 33244 67112 33284
rect 67152 33244 67194 33284
rect 67234 33244 67276 33284
rect 67316 33244 67358 33284
rect 67398 33244 67440 33284
rect 67480 33244 67489 33284
rect 74275 32908 74284 32948
rect 74324 32908 74764 32948
rect 74804 32908 74813 32948
rect 71788 32824 73100 32864
rect 71788 32780 71828 32824
rect 73060 32780 73100 32824
rect 71748 32740 71788 32780
rect 71828 32740 71837 32780
rect 73060 32740 74668 32780
rect 74708 32740 74717 32780
rect 75331 32740 75340 32780
rect 75380 32740 75628 32780
rect 75668 32740 75677 32780
rect 80227 32740 80236 32780
rect 80276 32740 80716 32780
rect 80756 32740 80765 32780
rect 81283 32740 81292 32780
rect 81332 32740 81868 32780
rect 81908 32740 81917 32780
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 8343 32488 8352 32528
rect 8392 32488 8434 32528
rect 8474 32488 8516 32528
rect 8556 32488 8598 32528
rect 8638 32488 8680 32528
rect 8720 32488 8729 32528
rect 12343 32488 12352 32528
rect 12392 32488 12434 32528
rect 12474 32488 12516 32528
rect 12556 32488 12598 32528
rect 12638 32488 12680 32528
rect 12720 32488 12729 32528
rect 16343 32488 16352 32528
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16720 32488 16729 32528
rect 20343 32488 20352 32528
rect 20392 32488 20434 32528
rect 20474 32488 20516 32528
rect 20556 32488 20598 32528
rect 20638 32488 20680 32528
rect 20720 32488 20729 32528
rect 24343 32488 24352 32528
rect 24392 32488 24434 32528
rect 24474 32488 24516 32528
rect 24556 32488 24598 32528
rect 24638 32488 24680 32528
rect 24720 32488 24729 32528
rect 28343 32488 28352 32528
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28720 32488 28729 32528
rect 32343 32488 32352 32528
rect 32392 32488 32434 32528
rect 32474 32488 32516 32528
rect 32556 32488 32598 32528
rect 32638 32488 32680 32528
rect 32720 32488 32729 32528
rect 36343 32488 36352 32528
rect 36392 32488 36434 32528
rect 36474 32488 36516 32528
rect 36556 32488 36598 32528
rect 36638 32488 36680 32528
rect 36720 32488 36729 32528
rect 40343 32488 40352 32528
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40720 32488 40729 32528
rect 44343 32488 44352 32528
rect 44392 32488 44434 32528
rect 44474 32488 44516 32528
rect 44556 32488 44598 32528
rect 44638 32488 44680 32528
rect 44720 32488 44729 32528
rect 48343 32488 48352 32528
rect 48392 32488 48434 32528
rect 48474 32488 48516 32528
rect 48556 32488 48598 32528
rect 48638 32488 48680 32528
rect 48720 32488 48729 32528
rect 52343 32488 52352 32528
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52720 32488 52729 32528
rect 56343 32488 56352 32528
rect 56392 32488 56434 32528
rect 56474 32488 56516 32528
rect 56556 32488 56598 32528
rect 56638 32488 56680 32528
rect 56720 32488 56729 32528
rect 60343 32488 60352 32528
rect 60392 32488 60434 32528
rect 60474 32488 60516 32528
rect 60556 32488 60598 32528
rect 60638 32488 60680 32528
rect 60720 32488 60729 32528
rect 64343 32488 64352 32528
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64720 32488 64729 32528
rect 68343 32488 68352 32528
rect 68392 32488 68434 32528
rect 68474 32488 68516 32528
rect 68556 32488 68598 32528
rect 68638 32488 68680 32528
rect 68720 32488 68729 32528
rect 76675 32488 76684 32528
rect 76724 32488 77356 32528
rect 77396 32488 77405 32528
rect 67555 32068 67564 32108
rect 67604 32068 73900 32108
rect 73940 32068 73949 32108
rect 68716 31984 73612 32024
rect 73652 31984 73661 32024
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 7103 31732 7112 31772
rect 7152 31732 7194 31772
rect 7234 31732 7276 31772
rect 7316 31732 7358 31772
rect 7398 31732 7440 31772
rect 7480 31732 7489 31772
rect 11103 31732 11112 31772
rect 11152 31732 11194 31772
rect 11234 31732 11276 31772
rect 11316 31732 11358 31772
rect 11398 31732 11440 31772
rect 11480 31732 11489 31772
rect 15103 31732 15112 31772
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15480 31732 15489 31772
rect 19103 31732 19112 31772
rect 19152 31732 19194 31772
rect 19234 31732 19276 31772
rect 19316 31732 19358 31772
rect 19398 31732 19440 31772
rect 19480 31732 19489 31772
rect 23103 31732 23112 31772
rect 23152 31732 23194 31772
rect 23234 31732 23276 31772
rect 23316 31732 23358 31772
rect 23398 31732 23440 31772
rect 23480 31732 23489 31772
rect 27103 31732 27112 31772
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27480 31732 27489 31772
rect 31103 31732 31112 31772
rect 31152 31732 31194 31772
rect 31234 31732 31276 31772
rect 31316 31732 31358 31772
rect 31398 31732 31440 31772
rect 31480 31732 31489 31772
rect 35103 31732 35112 31772
rect 35152 31732 35194 31772
rect 35234 31732 35276 31772
rect 35316 31732 35358 31772
rect 35398 31732 35440 31772
rect 35480 31732 35489 31772
rect 39103 31732 39112 31772
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39480 31732 39489 31772
rect 43103 31732 43112 31772
rect 43152 31732 43194 31772
rect 43234 31732 43276 31772
rect 43316 31732 43358 31772
rect 43398 31732 43440 31772
rect 43480 31732 43489 31772
rect 47103 31732 47112 31772
rect 47152 31732 47194 31772
rect 47234 31732 47276 31772
rect 47316 31732 47358 31772
rect 47398 31732 47440 31772
rect 47480 31732 47489 31772
rect 51103 31732 51112 31772
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51480 31732 51489 31772
rect 55103 31732 55112 31772
rect 55152 31732 55194 31772
rect 55234 31732 55276 31772
rect 55316 31732 55358 31772
rect 55398 31732 55440 31772
rect 55480 31732 55489 31772
rect 59103 31732 59112 31772
rect 59152 31732 59194 31772
rect 59234 31732 59276 31772
rect 59316 31732 59358 31772
rect 59398 31732 59440 31772
rect 59480 31732 59489 31772
rect 63103 31732 63112 31772
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63480 31732 63489 31772
rect 67103 31732 67112 31772
rect 67152 31732 67194 31772
rect 67234 31732 67276 31772
rect 67316 31732 67358 31772
rect 67398 31732 67440 31772
rect 67480 31732 67489 31772
rect 0 31628 80 31708
rect 67171 31564 67180 31604
rect 67220 31564 67564 31604
rect 67604 31564 67613 31604
rect 68716 31520 68756 31984
rect 69859 31900 69868 31940
rect 69908 31900 74668 31940
rect 74708 31900 74717 31940
rect 68899 31816 68908 31856
rect 68948 31816 74284 31856
rect 74324 31816 74333 31856
rect 69475 31732 69484 31772
rect 69524 31732 73228 31772
rect 73268 31732 73277 31772
rect 82723 31732 82732 31772
rect 82772 31732 82781 31772
rect 68812 31648 73268 31688
rect 68812 31604 68852 31648
rect 73228 31604 73268 31648
rect 82732 31604 82772 31732
rect 86947 31604 87005 31605
rect 68803 31564 68812 31604
rect 68852 31564 68861 31604
rect 69859 31564 69868 31604
rect 69908 31564 73100 31604
rect 73206 31564 73215 31604
rect 73255 31564 73268 31604
rect 82296 31564 82305 31604
rect 82345 31564 82772 31604
rect 83496 31564 83505 31604
rect 83545 31564 83788 31604
rect 83828 31564 83837 31604
rect 84696 31564 84705 31604
rect 84745 31564 84940 31604
rect 84980 31564 84989 31604
rect 86947 31564 86956 31604
rect 86996 31564 87215 31604
rect 87255 31564 87264 31604
rect 88195 31564 88204 31604
rect 88244 31564 88415 31604
rect 88455 31564 88464 31604
rect 97496 31564 97505 31604
rect 97545 31564 98188 31604
rect 98228 31564 98237 31604
rect 98296 31564 98305 31604
rect 98345 31564 99244 31604
rect 99284 31564 99293 31604
rect 73060 31520 73100 31564
rect 86947 31563 87005 31564
rect 76771 31520 76829 31521
rect 85219 31520 85277 31521
rect 86851 31520 86909 31521
rect 89923 31520 89981 31521
rect 92227 31520 92285 31521
rect 67651 31480 67660 31520
rect 67700 31480 68756 31520
rect 69187 31480 69196 31520
rect 69236 31480 69245 31520
rect 69571 31480 69580 31520
rect 69620 31480 72415 31520
rect 72455 31480 72464 31520
rect 73060 31480 73505 31520
rect 73545 31480 73554 31520
rect 76771 31480 76780 31520
rect 76855 31480 76915 31520
rect 85133 31480 85215 31520
rect 85268 31480 85277 31520
rect 86765 31480 86815 31520
rect 86855 31480 86860 31520
rect 86900 31480 86909 31520
rect 89837 31480 89905 31520
rect 89972 31480 89981 31520
rect 91096 31480 91105 31520
rect 91145 31480 91372 31520
rect 91412 31480 91421 31520
rect 92227 31480 92236 31520
rect 92276 31480 92415 31520
rect 92455 31480 92464 31520
rect 69196 31436 69236 31480
rect 76771 31479 76829 31480
rect 85219 31479 85277 31480
rect 86851 31479 86909 31480
rect 89923 31479 89981 31480
rect 92227 31479 92285 31480
rect 69196 31396 72815 31436
rect 72855 31396 72864 31436
rect 89496 31396 89505 31436
rect 89545 31396 89740 31436
rect 89780 31396 89789 31436
rect 90979 31396 90988 31436
rect 91028 31396 91615 31436
rect 91655 31396 91664 31436
rect 69667 31312 69676 31352
rect 69716 31312 72305 31352
rect 72345 31312 72354 31352
rect 75715 31312 75724 31352
rect 75764 31312 76015 31352
rect 76055 31312 76064 31352
rect 67267 31228 67276 31268
rect 67316 31228 67564 31268
rect 67604 31228 68620 31268
rect 68660 31228 69292 31268
rect 69332 31228 69772 31268
rect 69812 31228 69821 31268
rect 69379 31144 69388 31184
rect 69428 31144 69580 31184
rect 69620 31144 69629 31184
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 8343 30976 8352 31016
rect 8392 30976 8434 31016
rect 8474 30976 8516 31016
rect 8556 30976 8598 31016
rect 8638 30976 8680 31016
rect 8720 30976 8729 31016
rect 12343 30976 12352 31016
rect 12392 30976 12434 31016
rect 12474 30976 12516 31016
rect 12556 30976 12598 31016
rect 12638 30976 12680 31016
rect 12720 30976 12729 31016
rect 16343 30976 16352 31016
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16720 30976 16729 31016
rect 20343 30976 20352 31016
rect 20392 30976 20434 31016
rect 20474 30976 20516 31016
rect 20556 30976 20598 31016
rect 20638 30976 20680 31016
rect 20720 30976 20729 31016
rect 24343 30976 24352 31016
rect 24392 30976 24434 31016
rect 24474 30976 24516 31016
rect 24556 30976 24598 31016
rect 24638 30976 24680 31016
rect 24720 30976 24729 31016
rect 28343 30976 28352 31016
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28720 30976 28729 31016
rect 32343 30976 32352 31016
rect 32392 30976 32434 31016
rect 32474 30976 32516 31016
rect 32556 30976 32598 31016
rect 32638 30976 32680 31016
rect 32720 30976 32729 31016
rect 36343 30976 36352 31016
rect 36392 30976 36434 31016
rect 36474 30976 36516 31016
rect 36556 30976 36598 31016
rect 36638 30976 36680 31016
rect 36720 30976 36729 31016
rect 40343 30976 40352 31016
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40720 30976 40729 31016
rect 44343 30976 44352 31016
rect 44392 30976 44434 31016
rect 44474 30976 44516 31016
rect 44556 30976 44598 31016
rect 44638 30976 44680 31016
rect 44720 30976 44729 31016
rect 48343 30976 48352 31016
rect 48392 30976 48434 31016
rect 48474 30976 48516 31016
rect 48556 30976 48598 31016
rect 48638 30976 48680 31016
rect 48720 30976 48729 31016
rect 52343 30976 52352 31016
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52720 30976 52729 31016
rect 56343 30976 56352 31016
rect 56392 30976 56434 31016
rect 56474 30976 56516 31016
rect 56556 30976 56598 31016
rect 56638 30976 56680 31016
rect 56720 30976 56729 31016
rect 60343 30976 60352 31016
rect 60392 30976 60434 31016
rect 60474 30976 60516 31016
rect 60556 30976 60598 31016
rect 60638 30976 60680 31016
rect 60720 30976 60729 31016
rect 64343 30976 64352 31016
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64720 30976 64729 31016
rect 68343 30976 68352 31016
rect 68392 30976 68434 31016
rect 68474 30976 68516 31016
rect 68556 30976 68598 31016
rect 68638 30976 68680 31016
rect 68720 30976 68729 31016
rect 0 30788 80 30868
rect 69091 30808 69100 30848
rect 69140 30808 71884 30848
rect 71924 30808 71933 30848
rect 68515 30724 68524 30764
rect 68564 30724 69292 30764
rect 69332 30724 69341 30764
rect 67747 30640 67756 30680
rect 67796 30640 68044 30680
rect 68084 30640 69004 30680
rect 69044 30640 69053 30680
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 7103 30220 7112 30260
rect 7152 30220 7194 30260
rect 7234 30220 7276 30260
rect 7316 30220 7358 30260
rect 7398 30220 7440 30260
rect 7480 30220 7489 30260
rect 11103 30220 11112 30260
rect 11152 30220 11194 30260
rect 11234 30220 11276 30260
rect 11316 30220 11358 30260
rect 11398 30220 11440 30260
rect 11480 30220 11489 30260
rect 15103 30220 15112 30260
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15480 30220 15489 30260
rect 19103 30220 19112 30260
rect 19152 30220 19194 30260
rect 19234 30220 19276 30260
rect 19316 30220 19358 30260
rect 19398 30220 19440 30260
rect 19480 30220 19489 30260
rect 23103 30220 23112 30260
rect 23152 30220 23194 30260
rect 23234 30220 23276 30260
rect 23316 30220 23358 30260
rect 23398 30220 23440 30260
rect 23480 30220 23489 30260
rect 27103 30220 27112 30260
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27480 30220 27489 30260
rect 31103 30220 31112 30260
rect 31152 30220 31194 30260
rect 31234 30220 31276 30260
rect 31316 30220 31358 30260
rect 31398 30220 31440 30260
rect 31480 30220 31489 30260
rect 35103 30220 35112 30260
rect 35152 30220 35194 30260
rect 35234 30220 35276 30260
rect 35316 30220 35358 30260
rect 35398 30220 35440 30260
rect 35480 30220 35489 30260
rect 39103 30220 39112 30260
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39480 30220 39489 30260
rect 43103 30220 43112 30260
rect 43152 30220 43194 30260
rect 43234 30220 43276 30260
rect 43316 30220 43358 30260
rect 43398 30220 43440 30260
rect 43480 30220 43489 30260
rect 47103 30220 47112 30260
rect 47152 30220 47194 30260
rect 47234 30220 47276 30260
rect 47316 30220 47358 30260
rect 47398 30220 47440 30260
rect 47480 30220 47489 30260
rect 51103 30220 51112 30260
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51480 30220 51489 30260
rect 55103 30220 55112 30260
rect 55152 30220 55194 30260
rect 55234 30220 55276 30260
rect 55316 30220 55358 30260
rect 55398 30220 55440 30260
rect 55480 30220 55489 30260
rect 59103 30220 59112 30260
rect 59152 30220 59194 30260
rect 59234 30220 59276 30260
rect 59316 30220 59358 30260
rect 59398 30220 59440 30260
rect 59480 30220 59489 30260
rect 63103 30220 63112 30260
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63480 30220 63489 30260
rect 67103 30220 67112 30260
rect 67152 30220 67194 30260
rect 67234 30220 67276 30260
rect 67316 30220 67358 30260
rect 67398 30220 67440 30260
rect 67480 30220 67489 30260
rect 0 29948 80 30028
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 8343 29464 8352 29504
rect 8392 29464 8434 29504
rect 8474 29464 8516 29504
rect 8556 29464 8598 29504
rect 8638 29464 8680 29504
rect 8720 29464 8729 29504
rect 12343 29464 12352 29504
rect 12392 29464 12434 29504
rect 12474 29464 12516 29504
rect 12556 29464 12598 29504
rect 12638 29464 12680 29504
rect 12720 29464 12729 29504
rect 16343 29464 16352 29504
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16720 29464 16729 29504
rect 20343 29464 20352 29504
rect 20392 29464 20434 29504
rect 20474 29464 20516 29504
rect 20556 29464 20598 29504
rect 20638 29464 20680 29504
rect 20720 29464 20729 29504
rect 24343 29464 24352 29504
rect 24392 29464 24434 29504
rect 24474 29464 24516 29504
rect 24556 29464 24598 29504
rect 24638 29464 24680 29504
rect 24720 29464 24729 29504
rect 28343 29464 28352 29504
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28720 29464 28729 29504
rect 32343 29464 32352 29504
rect 32392 29464 32434 29504
rect 32474 29464 32516 29504
rect 32556 29464 32598 29504
rect 32638 29464 32680 29504
rect 32720 29464 32729 29504
rect 36343 29464 36352 29504
rect 36392 29464 36434 29504
rect 36474 29464 36516 29504
rect 36556 29464 36598 29504
rect 36638 29464 36680 29504
rect 36720 29464 36729 29504
rect 40343 29464 40352 29504
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40720 29464 40729 29504
rect 44343 29464 44352 29504
rect 44392 29464 44434 29504
rect 44474 29464 44516 29504
rect 44556 29464 44598 29504
rect 44638 29464 44680 29504
rect 44720 29464 44729 29504
rect 48343 29464 48352 29504
rect 48392 29464 48434 29504
rect 48474 29464 48516 29504
rect 48556 29464 48598 29504
rect 48638 29464 48680 29504
rect 48720 29464 48729 29504
rect 52343 29464 52352 29504
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52720 29464 52729 29504
rect 56343 29464 56352 29504
rect 56392 29464 56434 29504
rect 56474 29464 56516 29504
rect 56556 29464 56598 29504
rect 56638 29464 56680 29504
rect 56720 29464 56729 29504
rect 60343 29464 60352 29504
rect 60392 29464 60434 29504
rect 60474 29464 60516 29504
rect 60556 29464 60598 29504
rect 60638 29464 60680 29504
rect 60720 29464 60729 29504
rect 64343 29464 64352 29504
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64720 29464 64729 29504
rect 68343 29464 68352 29504
rect 68392 29464 68434 29504
rect 68474 29464 68516 29504
rect 68556 29464 68598 29504
rect 68638 29464 68680 29504
rect 68720 29464 68729 29504
rect 0 29108 80 29188
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 7103 28708 7112 28748
rect 7152 28708 7194 28748
rect 7234 28708 7276 28748
rect 7316 28708 7358 28748
rect 7398 28708 7440 28748
rect 7480 28708 7489 28748
rect 11103 28708 11112 28748
rect 11152 28708 11194 28748
rect 11234 28708 11276 28748
rect 11316 28708 11358 28748
rect 11398 28708 11440 28748
rect 11480 28708 11489 28748
rect 15103 28708 15112 28748
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15480 28708 15489 28748
rect 19103 28708 19112 28748
rect 19152 28708 19194 28748
rect 19234 28708 19276 28748
rect 19316 28708 19358 28748
rect 19398 28708 19440 28748
rect 19480 28708 19489 28748
rect 23103 28708 23112 28748
rect 23152 28708 23194 28748
rect 23234 28708 23276 28748
rect 23316 28708 23358 28748
rect 23398 28708 23440 28748
rect 23480 28708 23489 28748
rect 27103 28708 27112 28748
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27480 28708 27489 28748
rect 31103 28708 31112 28748
rect 31152 28708 31194 28748
rect 31234 28708 31276 28748
rect 31316 28708 31358 28748
rect 31398 28708 31440 28748
rect 31480 28708 31489 28748
rect 35103 28708 35112 28748
rect 35152 28708 35194 28748
rect 35234 28708 35276 28748
rect 35316 28708 35358 28748
rect 35398 28708 35440 28748
rect 35480 28708 35489 28748
rect 39103 28708 39112 28748
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39480 28708 39489 28748
rect 43103 28708 43112 28748
rect 43152 28708 43194 28748
rect 43234 28708 43276 28748
rect 43316 28708 43358 28748
rect 43398 28708 43440 28748
rect 43480 28708 43489 28748
rect 47103 28708 47112 28748
rect 47152 28708 47194 28748
rect 47234 28708 47276 28748
rect 47316 28708 47358 28748
rect 47398 28708 47440 28748
rect 47480 28708 47489 28748
rect 51103 28708 51112 28748
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51480 28708 51489 28748
rect 55103 28708 55112 28748
rect 55152 28708 55194 28748
rect 55234 28708 55276 28748
rect 55316 28708 55358 28748
rect 55398 28708 55440 28748
rect 55480 28708 55489 28748
rect 59103 28708 59112 28748
rect 59152 28708 59194 28748
rect 59234 28708 59276 28748
rect 59316 28708 59358 28748
rect 59398 28708 59440 28748
rect 59480 28708 59489 28748
rect 63103 28708 63112 28748
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63480 28708 63489 28748
rect 67103 28708 67112 28748
rect 67152 28708 67194 28748
rect 67234 28708 67276 28748
rect 67316 28708 67358 28748
rect 67398 28708 67440 28748
rect 67480 28708 67489 28748
rect 0 28268 80 28348
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 8343 27952 8352 27992
rect 8392 27952 8434 27992
rect 8474 27952 8516 27992
rect 8556 27952 8598 27992
rect 8638 27952 8680 27992
rect 8720 27952 8729 27992
rect 12343 27952 12352 27992
rect 12392 27952 12434 27992
rect 12474 27952 12516 27992
rect 12556 27952 12598 27992
rect 12638 27952 12680 27992
rect 12720 27952 12729 27992
rect 16343 27952 16352 27992
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16720 27952 16729 27992
rect 20343 27952 20352 27992
rect 20392 27952 20434 27992
rect 20474 27952 20516 27992
rect 20556 27952 20598 27992
rect 20638 27952 20680 27992
rect 20720 27952 20729 27992
rect 24343 27952 24352 27992
rect 24392 27952 24434 27992
rect 24474 27952 24516 27992
rect 24556 27952 24598 27992
rect 24638 27952 24680 27992
rect 24720 27952 24729 27992
rect 28343 27952 28352 27992
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28720 27952 28729 27992
rect 32343 27952 32352 27992
rect 32392 27952 32434 27992
rect 32474 27952 32516 27992
rect 32556 27952 32598 27992
rect 32638 27952 32680 27992
rect 32720 27952 32729 27992
rect 36343 27952 36352 27992
rect 36392 27952 36434 27992
rect 36474 27952 36516 27992
rect 36556 27952 36598 27992
rect 36638 27952 36680 27992
rect 36720 27952 36729 27992
rect 40343 27952 40352 27992
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40720 27952 40729 27992
rect 44343 27952 44352 27992
rect 44392 27952 44434 27992
rect 44474 27952 44516 27992
rect 44556 27952 44598 27992
rect 44638 27952 44680 27992
rect 44720 27952 44729 27992
rect 48343 27952 48352 27992
rect 48392 27952 48434 27992
rect 48474 27952 48516 27992
rect 48556 27952 48598 27992
rect 48638 27952 48680 27992
rect 48720 27952 48729 27992
rect 52343 27952 52352 27992
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52720 27952 52729 27992
rect 56343 27952 56352 27992
rect 56392 27952 56434 27992
rect 56474 27952 56516 27992
rect 56556 27952 56598 27992
rect 56638 27952 56680 27992
rect 56720 27952 56729 27992
rect 60343 27952 60352 27992
rect 60392 27952 60434 27992
rect 60474 27952 60516 27992
rect 60556 27952 60598 27992
rect 60638 27952 60680 27992
rect 60720 27952 60729 27992
rect 64343 27952 64352 27992
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64720 27952 64729 27992
rect 68343 27952 68352 27992
rect 68392 27952 68434 27992
rect 68474 27952 68516 27992
rect 68556 27952 68598 27992
rect 68638 27952 68680 27992
rect 68720 27952 68729 27992
rect 0 27428 80 27508
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 7103 27196 7112 27236
rect 7152 27196 7194 27236
rect 7234 27196 7276 27236
rect 7316 27196 7358 27236
rect 7398 27196 7440 27236
rect 7480 27196 7489 27236
rect 11103 27196 11112 27236
rect 11152 27196 11194 27236
rect 11234 27196 11276 27236
rect 11316 27196 11358 27236
rect 11398 27196 11440 27236
rect 11480 27196 11489 27236
rect 15103 27196 15112 27236
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15480 27196 15489 27236
rect 19103 27196 19112 27236
rect 19152 27196 19194 27236
rect 19234 27196 19276 27236
rect 19316 27196 19358 27236
rect 19398 27196 19440 27236
rect 19480 27196 19489 27236
rect 23103 27196 23112 27236
rect 23152 27196 23194 27236
rect 23234 27196 23276 27236
rect 23316 27196 23358 27236
rect 23398 27196 23440 27236
rect 23480 27196 23489 27236
rect 27103 27196 27112 27236
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27480 27196 27489 27236
rect 31103 27196 31112 27236
rect 31152 27196 31194 27236
rect 31234 27196 31276 27236
rect 31316 27196 31358 27236
rect 31398 27196 31440 27236
rect 31480 27196 31489 27236
rect 35103 27196 35112 27236
rect 35152 27196 35194 27236
rect 35234 27196 35276 27236
rect 35316 27196 35358 27236
rect 35398 27196 35440 27236
rect 35480 27196 35489 27236
rect 39103 27196 39112 27236
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39480 27196 39489 27236
rect 43103 27196 43112 27236
rect 43152 27196 43194 27236
rect 43234 27196 43276 27236
rect 43316 27196 43358 27236
rect 43398 27196 43440 27236
rect 43480 27196 43489 27236
rect 47103 27196 47112 27236
rect 47152 27196 47194 27236
rect 47234 27196 47276 27236
rect 47316 27196 47358 27236
rect 47398 27196 47440 27236
rect 47480 27196 47489 27236
rect 51103 27196 51112 27236
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51480 27196 51489 27236
rect 55103 27196 55112 27236
rect 55152 27196 55194 27236
rect 55234 27196 55276 27236
rect 55316 27196 55358 27236
rect 55398 27196 55440 27236
rect 55480 27196 55489 27236
rect 59103 27196 59112 27236
rect 59152 27196 59194 27236
rect 59234 27196 59276 27236
rect 59316 27196 59358 27236
rect 59398 27196 59440 27236
rect 59480 27196 59489 27236
rect 63103 27196 63112 27236
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63480 27196 63489 27236
rect 67103 27196 67112 27236
rect 67152 27196 67194 27236
rect 67234 27196 67276 27236
rect 67316 27196 67358 27236
rect 67398 27196 67440 27236
rect 67480 27196 67489 27236
rect 0 26588 80 26668
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 8343 26440 8352 26480
rect 8392 26440 8434 26480
rect 8474 26440 8516 26480
rect 8556 26440 8598 26480
rect 8638 26440 8680 26480
rect 8720 26440 8729 26480
rect 12343 26440 12352 26480
rect 12392 26440 12434 26480
rect 12474 26440 12516 26480
rect 12556 26440 12598 26480
rect 12638 26440 12680 26480
rect 12720 26440 12729 26480
rect 16343 26440 16352 26480
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16720 26440 16729 26480
rect 20343 26440 20352 26480
rect 20392 26440 20434 26480
rect 20474 26440 20516 26480
rect 20556 26440 20598 26480
rect 20638 26440 20680 26480
rect 20720 26440 20729 26480
rect 24343 26440 24352 26480
rect 24392 26440 24434 26480
rect 24474 26440 24516 26480
rect 24556 26440 24598 26480
rect 24638 26440 24680 26480
rect 24720 26440 24729 26480
rect 28343 26440 28352 26480
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28720 26440 28729 26480
rect 32343 26440 32352 26480
rect 32392 26440 32434 26480
rect 32474 26440 32516 26480
rect 32556 26440 32598 26480
rect 32638 26440 32680 26480
rect 32720 26440 32729 26480
rect 36343 26440 36352 26480
rect 36392 26440 36434 26480
rect 36474 26440 36516 26480
rect 36556 26440 36598 26480
rect 36638 26440 36680 26480
rect 36720 26440 36729 26480
rect 40343 26440 40352 26480
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40720 26440 40729 26480
rect 44343 26440 44352 26480
rect 44392 26440 44434 26480
rect 44474 26440 44516 26480
rect 44556 26440 44598 26480
rect 44638 26440 44680 26480
rect 44720 26440 44729 26480
rect 48343 26440 48352 26480
rect 48392 26440 48434 26480
rect 48474 26440 48516 26480
rect 48556 26440 48598 26480
rect 48638 26440 48680 26480
rect 48720 26440 48729 26480
rect 52343 26440 52352 26480
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52720 26440 52729 26480
rect 56343 26440 56352 26480
rect 56392 26440 56434 26480
rect 56474 26440 56516 26480
rect 56556 26440 56598 26480
rect 56638 26440 56680 26480
rect 56720 26440 56729 26480
rect 60343 26440 60352 26480
rect 60392 26440 60434 26480
rect 60474 26440 60516 26480
rect 60556 26440 60598 26480
rect 60638 26440 60680 26480
rect 60720 26440 60729 26480
rect 64343 26440 64352 26480
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64720 26440 64729 26480
rect 68343 26440 68352 26480
rect 68392 26440 68434 26480
rect 68474 26440 68516 26480
rect 68556 26440 68598 26480
rect 68638 26440 68680 26480
rect 68720 26440 68729 26480
rect 68611 26104 68620 26144
rect 68660 26104 68812 26144
rect 68852 26104 69292 26144
rect 69332 26104 69484 26144
rect 69524 26104 69772 26144
rect 69812 26104 69821 26144
rect 71779 26060 71837 26061
rect 68323 26020 68332 26060
rect 68372 26020 69100 26060
rect 69140 26020 69388 26060
rect 69428 26020 69580 26060
rect 69620 26020 71788 26060
rect 71828 26020 71837 26060
rect 71779 26019 71837 26020
rect 71875 25976 71933 25977
rect 68803 25936 68812 25976
rect 68852 25936 71884 25976
rect 71924 25936 71933 25976
rect 71875 25935 71933 25936
rect 72451 25892 72509 25893
rect 69571 25852 69580 25892
rect 69620 25852 72305 25892
rect 72345 25852 72354 25892
rect 72451 25852 72460 25892
rect 72500 25852 74305 25892
rect 74345 25852 74354 25892
rect 91896 25852 91905 25892
rect 91945 25852 92140 25892
rect 92180 25852 92189 25892
rect 72451 25851 72509 25852
rect 0 25748 80 25828
rect 94915 25808 94973 25809
rect 69187 25768 69196 25808
rect 69236 25768 72415 25808
rect 72455 25768 72464 25808
rect 72652 25768 72705 25808
rect 72745 25768 72754 25808
rect 76579 25768 76588 25808
rect 76628 25768 76815 25808
rect 76855 25768 76864 25808
rect 94915 25768 94924 25808
rect 94964 25768 95105 25808
rect 95145 25768 95154 25808
rect 72652 25724 72692 25768
rect 94915 25767 94973 25768
rect 95011 25724 95069 25725
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 7103 25684 7112 25724
rect 7152 25684 7194 25724
rect 7234 25684 7276 25724
rect 7316 25684 7358 25724
rect 7398 25684 7440 25724
rect 7480 25684 7489 25724
rect 11103 25684 11112 25724
rect 11152 25684 11194 25724
rect 11234 25684 11276 25724
rect 11316 25684 11358 25724
rect 11398 25684 11440 25724
rect 11480 25684 11489 25724
rect 15103 25684 15112 25724
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15480 25684 15489 25724
rect 19103 25684 19112 25724
rect 19152 25684 19194 25724
rect 19234 25684 19276 25724
rect 19316 25684 19358 25724
rect 19398 25684 19440 25724
rect 19480 25684 19489 25724
rect 23103 25684 23112 25724
rect 23152 25684 23194 25724
rect 23234 25684 23276 25724
rect 23316 25684 23358 25724
rect 23398 25684 23440 25724
rect 23480 25684 23489 25724
rect 27103 25684 27112 25724
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27480 25684 27489 25724
rect 31103 25684 31112 25724
rect 31152 25684 31194 25724
rect 31234 25684 31276 25724
rect 31316 25684 31358 25724
rect 31398 25684 31440 25724
rect 31480 25684 31489 25724
rect 35103 25684 35112 25724
rect 35152 25684 35194 25724
rect 35234 25684 35276 25724
rect 35316 25684 35358 25724
rect 35398 25684 35440 25724
rect 35480 25684 35489 25724
rect 39103 25684 39112 25724
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39480 25684 39489 25724
rect 43103 25684 43112 25724
rect 43152 25684 43194 25724
rect 43234 25684 43276 25724
rect 43316 25684 43358 25724
rect 43398 25684 43440 25724
rect 43480 25684 43489 25724
rect 47103 25684 47112 25724
rect 47152 25684 47194 25724
rect 47234 25684 47276 25724
rect 47316 25684 47358 25724
rect 47398 25684 47440 25724
rect 47480 25684 47489 25724
rect 51103 25684 51112 25724
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51480 25684 51489 25724
rect 55103 25684 55112 25724
rect 55152 25684 55194 25724
rect 55234 25684 55276 25724
rect 55316 25684 55358 25724
rect 55398 25684 55440 25724
rect 55480 25684 55489 25724
rect 59103 25684 59112 25724
rect 59152 25684 59194 25724
rect 59234 25684 59276 25724
rect 59316 25684 59358 25724
rect 59398 25684 59440 25724
rect 59480 25684 59489 25724
rect 63103 25684 63112 25724
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63480 25684 63489 25724
rect 67103 25684 67112 25724
rect 67152 25684 67194 25724
rect 67234 25684 67276 25724
rect 67316 25684 67358 25724
rect 67398 25684 67440 25724
rect 67480 25684 67489 25724
rect 68995 25684 69004 25724
rect 69044 25684 72692 25724
rect 72835 25684 72844 25724
rect 72884 25684 72893 25724
rect 73891 25684 73900 25724
rect 73940 25684 74415 25724
rect 74455 25684 74464 25724
rect 75811 25684 75820 25724
rect 75860 25684 76415 25724
rect 76455 25684 76464 25724
rect 84696 25684 84705 25724
rect 84745 25684 84940 25724
rect 84980 25684 84989 25724
rect 87206 25684 87215 25724
rect 87255 25684 87724 25724
rect 87764 25684 87773 25724
rect 90006 25684 90015 25724
rect 90055 25684 90508 25724
rect 90548 25684 90557 25724
rect 95011 25684 95020 25724
rect 95060 25684 95215 25724
rect 95255 25684 95264 25724
rect 72844 25640 72884 25684
rect 95011 25683 95069 25684
rect 67939 25600 67948 25640
rect 67988 25600 68468 25640
rect 68515 25600 68524 25640
rect 68564 25600 72884 25640
rect 72931 25640 72989 25641
rect 72931 25600 72940 25640
rect 72980 25600 81920 25640
rect 68428 25388 68468 25600
rect 72931 25599 72989 25600
rect 69859 25516 69868 25556
rect 69908 25516 73228 25556
rect 73268 25516 73277 25556
rect 81880 25472 81920 25600
rect 69955 25432 69964 25472
rect 70004 25432 73996 25472
rect 74036 25432 74045 25472
rect 81880 25432 99148 25472
rect 99188 25432 99197 25472
rect 59200 25348 68332 25388
rect 68372 25348 68381 25388
rect 68428 25348 73804 25388
rect 73844 25348 73853 25388
rect 59200 25304 59240 25348
rect 835 25264 844 25304
rect 884 25264 59240 25304
rect 67747 25264 67756 25304
rect 67796 25264 68620 25304
rect 68660 25264 69484 25304
rect 69524 25264 73036 25304
rect 73076 25264 73085 25304
rect 73228 25264 73460 25304
rect 73228 25220 73268 25264
rect 73420 25220 73460 25264
rect 69763 25180 69772 25220
rect 69812 25180 73268 25220
rect 73315 25180 73324 25220
rect 73364 25180 73373 25220
rect 73420 25180 73516 25220
rect 73556 25180 73565 25220
rect 74083 25180 74092 25220
rect 74132 25180 75628 25220
rect 75668 25180 75677 25220
rect 91363 25180 91372 25220
rect 91412 25180 92044 25220
rect 92084 25180 92093 25220
rect 73324 25136 73364 25180
rect 68899 25096 68908 25136
rect 68948 25096 73364 25136
rect 69283 25012 69292 25052
rect 69332 25012 69676 25052
rect 69716 25012 73324 25052
rect 73364 25012 73373 25052
rect 0 24968 80 24988
rect 0 24928 652 24968
rect 692 24928 701 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 8343 24928 8352 24968
rect 8392 24928 8434 24968
rect 8474 24928 8516 24968
rect 8556 24928 8598 24968
rect 8638 24928 8680 24968
rect 8720 24928 8729 24968
rect 12343 24928 12352 24968
rect 12392 24928 12434 24968
rect 12474 24928 12516 24968
rect 12556 24928 12598 24968
rect 12638 24928 12680 24968
rect 12720 24928 12729 24968
rect 16343 24928 16352 24968
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16720 24928 16729 24968
rect 20343 24928 20352 24968
rect 20392 24928 20434 24968
rect 20474 24928 20516 24968
rect 20556 24928 20598 24968
rect 20638 24928 20680 24968
rect 20720 24928 20729 24968
rect 24343 24928 24352 24968
rect 24392 24928 24434 24968
rect 24474 24928 24516 24968
rect 24556 24928 24598 24968
rect 24638 24928 24680 24968
rect 24720 24928 24729 24968
rect 28343 24928 28352 24968
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28720 24928 28729 24968
rect 32343 24928 32352 24968
rect 32392 24928 32434 24968
rect 32474 24928 32516 24968
rect 32556 24928 32598 24968
rect 32638 24928 32680 24968
rect 32720 24928 32729 24968
rect 36343 24928 36352 24968
rect 36392 24928 36434 24968
rect 36474 24928 36516 24968
rect 36556 24928 36598 24968
rect 36638 24928 36680 24968
rect 36720 24928 36729 24968
rect 40343 24928 40352 24968
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40720 24928 40729 24968
rect 44343 24928 44352 24968
rect 44392 24928 44434 24968
rect 44474 24928 44516 24968
rect 44556 24928 44598 24968
rect 44638 24928 44680 24968
rect 44720 24928 44729 24968
rect 48343 24928 48352 24968
rect 48392 24928 48434 24968
rect 48474 24928 48516 24968
rect 48556 24928 48598 24968
rect 48638 24928 48680 24968
rect 48720 24928 48729 24968
rect 52343 24928 52352 24968
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52720 24928 52729 24968
rect 56343 24928 56352 24968
rect 56392 24928 56434 24968
rect 56474 24928 56516 24968
rect 56556 24928 56598 24968
rect 56638 24928 56680 24968
rect 56720 24928 56729 24968
rect 60343 24928 60352 24968
rect 60392 24928 60434 24968
rect 60474 24928 60516 24968
rect 60556 24928 60598 24968
rect 60638 24928 60680 24968
rect 60720 24928 60729 24968
rect 64343 24928 64352 24968
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64720 24928 64729 24968
rect 68343 24928 68352 24968
rect 68392 24928 68434 24968
rect 68474 24928 68516 24968
rect 68556 24928 68598 24968
rect 68638 24928 68680 24968
rect 68720 24928 68729 24968
rect 0 24908 80 24928
rect 67555 24844 67564 24884
rect 67604 24844 75244 24884
rect 75284 24844 75293 24884
rect 95395 24676 95404 24716
rect 95444 24676 95692 24716
rect 95732 24676 95741 24716
rect 80035 24424 80044 24464
rect 80084 24424 80908 24464
rect 80948 24424 80957 24464
rect 80419 24340 80428 24380
rect 80468 24340 81196 24380
rect 81236 24340 81245 24380
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 7103 24172 7112 24212
rect 7152 24172 7194 24212
rect 7234 24172 7276 24212
rect 7316 24172 7358 24212
rect 7398 24172 7440 24212
rect 7480 24172 7489 24212
rect 11103 24172 11112 24212
rect 11152 24172 11194 24212
rect 11234 24172 11276 24212
rect 11316 24172 11358 24212
rect 11398 24172 11440 24212
rect 11480 24172 11489 24212
rect 15103 24172 15112 24212
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15480 24172 15489 24212
rect 19103 24172 19112 24212
rect 19152 24172 19194 24212
rect 19234 24172 19276 24212
rect 19316 24172 19358 24212
rect 19398 24172 19440 24212
rect 19480 24172 19489 24212
rect 23103 24172 23112 24212
rect 23152 24172 23194 24212
rect 23234 24172 23276 24212
rect 23316 24172 23358 24212
rect 23398 24172 23440 24212
rect 23480 24172 23489 24212
rect 27103 24172 27112 24212
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27480 24172 27489 24212
rect 31103 24172 31112 24212
rect 31152 24172 31194 24212
rect 31234 24172 31276 24212
rect 31316 24172 31358 24212
rect 31398 24172 31440 24212
rect 31480 24172 31489 24212
rect 35103 24172 35112 24212
rect 35152 24172 35194 24212
rect 35234 24172 35276 24212
rect 35316 24172 35358 24212
rect 35398 24172 35440 24212
rect 35480 24172 35489 24212
rect 39103 24172 39112 24212
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39480 24172 39489 24212
rect 43103 24172 43112 24212
rect 43152 24172 43194 24212
rect 43234 24172 43276 24212
rect 43316 24172 43358 24212
rect 43398 24172 43440 24212
rect 43480 24172 43489 24212
rect 47103 24172 47112 24212
rect 47152 24172 47194 24212
rect 47234 24172 47276 24212
rect 47316 24172 47358 24212
rect 47398 24172 47440 24212
rect 47480 24172 47489 24212
rect 51103 24172 51112 24212
rect 51152 24172 51194 24212
rect 51234 24172 51276 24212
rect 51316 24172 51358 24212
rect 51398 24172 51440 24212
rect 51480 24172 51489 24212
rect 55103 24172 55112 24212
rect 55152 24172 55194 24212
rect 55234 24172 55276 24212
rect 55316 24172 55358 24212
rect 55398 24172 55440 24212
rect 55480 24172 55489 24212
rect 59103 24172 59112 24212
rect 59152 24172 59194 24212
rect 59234 24172 59276 24212
rect 59316 24172 59358 24212
rect 59398 24172 59440 24212
rect 59480 24172 59489 24212
rect 63103 24172 63112 24212
rect 63152 24172 63194 24212
rect 63234 24172 63276 24212
rect 63316 24172 63358 24212
rect 63398 24172 63440 24212
rect 63480 24172 63489 24212
rect 67103 24172 67112 24212
rect 67152 24172 67194 24212
rect 67234 24172 67276 24212
rect 67316 24172 67358 24212
rect 67398 24172 67440 24212
rect 67480 24172 67489 24212
rect 0 24128 80 24148
rect 0 24088 652 24128
rect 692 24088 701 24128
rect 73123 24088 73132 24128
rect 73172 24088 74860 24128
rect 74900 24088 74909 24128
rect 0 24068 80 24088
rect 92419 24004 92428 24044
rect 92468 24004 93332 24044
rect 85411 23960 85469 23961
rect 85326 23920 85420 23960
rect 85460 23920 85469 23960
rect 90403 23920 90412 23960
rect 90452 23920 90740 23960
rect 85411 23919 85469 23920
rect 90700 23876 90740 23920
rect 93292 23876 93332 24004
rect 90700 23836 90796 23876
rect 90836 23836 90845 23876
rect 93292 23836 93580 23876
rect 93620 23836 93629 23876
rect 84259 23792 84317 23793
rect 835 23752 844 23792
rect 884 23752 2092 23792
rect 2132 23752 2141 23792
rect 84174 23752 84268 23792
rect 84308 23752 84317 23792
rect 84259 23751 84317 23752
rect 76579 23584 76588 23624
rect 76628 23584 76637 23624
rect 80707 23584 80716 23624
rect 80756 23584 80765 23624
rect 88387 23584 88396 23624
rect 88436 23584 88445 23624
rect 76588 23540 76628 23584
rect 80716 23540 80756 23584
rect 88396 23540 88436 23584
rect 76588 23500 76820 23540
rect 80716 23500 80852 23540
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 8343 23416 8352 23456
rect 8392 23416 8434 23456
rect 8474 23416 8516 23456
rect 8556 23416 8598 23456
rect 8638 23416 8680 23456
rect 8720 23416 8729 23456
rect 12343 23416 12352 23456
rect 12392 23416 12434 23456
rect 12474 23416 12516 23456
rect 12556 23416 12598 23456
rect 12638 23416 12680 23456
rect 12720 23416 12729 23456
rect 16343 23416 16352 23456
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16720 23416 16729 23456
rect 20343 23416 20352 23456
rect 20392 23416 20434 23456
rect 20474 23416 20516 23456
rect 20556 23416 20598 23456
rect 20638 23416 20680 23456
rect 20720 23416 20729 23456
rect 24343 23416 24352 23456
rect 24392 23416 24434 23456
rect 24474 23416 24516 23456
rect 24556 23416 24598 23456
rect 24638 23416 24680 23456
rect 24720 23416 24729 23456
rect 28343 23416 28352 23456
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28720 23416 28729 23456
rect 32343 23416 32352 23456
rect 32392 23416 32434 23456
rect 32474 23416 32516 23456
rect 32556 23416 32598 23456
rect 32638 23416 32680 23456
rect 32720 23416 32729 23456
rect 36343 23416 36352 23456
rect 36392 23416 36434 23456
rect 36474 23416 36516 23456
rect 36556 23416 36598 23456
rect 36638 23416 36680 23456
rect 36720 23416 36729 23456
rect 40343 23416 40352 23456
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40720 23416 40729 23456
rect 44343 23416 44352 23456
rect 44392 23416 44434 23456
rect 44474 23416 44516 23456
rect 44556 23416 44598 23456
rect 44638 23416 44680 23456
rect 44720 23416 44729 23456
rect 48343 23416 48352 23456
rect 48392 23416 48434 23456
rect 48474 23416 48516 23456
rect 48556 23416 48598 23456
rect 48638 23416 48680 23456
rect 48720 23416 48729 23456
rect 52343 23416 52352 23456
rect 52392 23416 52434 23456
rect 52474 23416 52516 23456
rect 52556 23416 52598 23456
rect 52638 23416 52680 23456
rect 52720 23416 52729 23456
rect 56343 23416 56352 23456
rect 56392 23416 56434 23456
rect 56474 23416 56516 23456
rect 56556 23416 56598 23456
rect 56638 23416 56680 23456
rect 56720 23416 56729 23456
rect 60343 23416 60352 23456
rect 60392 23416 60434 23456
rect 60474 23416 60516 23456
rect 60556 23416 60598 23456
rect 60638 23416 60680 23456
rect 60720 23416 60729 23456
rect 64343 23416 64352 23456
rect 64392 23416 64434 23456
rect 64474 23416 64516 23456
rect 64556 23416 64598 23456
rect 64638 23416 64680 23456
rect 64720 23416 64729 23456
rect 68343 23416 68352 23456
rect 68392 23416 68434 23456
rect 68474 23416 68516 23456
rect 68556 23416 68598 23456
rect 68638 23416 68680 23456
rect 68720 23416 68729 23456
rect 72343 23416 72352 23456
rect 72392 23416 72434 23456
rect 72474 23416 72516 23456
rect 72556 23416 72598 23456
rect 72638 23416 72680 23456
rect 72720 23416 72729 23456
rect 76343 23416 76352 23456
rect 76392 23416 76434 23456
rect 76474 23416 76516 23456
rect 76556 23416 76598 23456
rect 76638 23416 76680 23456
rect 76720 23416 76729 23456
rect 71779 23332 71788 23372
rect 71828 23332 75628 23372
rect 75668 23332 75677 23372
rect 0 23288 80 23308
rect 76780 23288 76820 23500
rect 80343 23416 80352 23456
rect 80392 23416 80434 23456
rect 80474 23416 80516 23456
rect 80556 23416 80598 23456
rect 80638 23416 80680 23456
rect 80720 23416 80729 23456
rect 80812 23288 80852 23500
rect 88204 23500 88436 23540
rect 84343 23416 84352 23456
rect 84392 23416 84434 23456
rect 84474 23416 84516 23456
rect 84556 23416 84598 23456
rect 84638 23416 84680 23456
rect 84720 23416 84729 23456
rect 83587 23288 83645 23289
rect 0 23248 652 23288
rect 692 23248 701 23288
rect 2083 23248 2092 23288
rect 2132 23248 68236 23288
rect 68276 23248 76300 23288
rect 76340 23248 76349 23288
rect 76675 23248 76684 23288
rect 76724 23248 76820 23288
rect 78403 23248 78412 23288
rect 78452 23248 79180 23288
rect 79220 23248 79229 23288
rect 80611 23248 80620 23288
rect 80660 23248 80852 23288
rect 83491 23248 83500 23288
rect 83540 23248 83596 23288
rect 83636 23248 83645 23288
rect 88204 23288 88244 23500
rect 88343 23416 88352 23456
rect 88392 23416 88434 23456
rect 88474 23416 88516 23456
rect 88556 23416 88598 23456
rect 88638 23416 88680 23456
rect 88720 23416 88729 23456
rect 92343 23416 92352 23456
rect 92392 23416 92434 23456
rect 92474 23416 92516 23456
rect 92556 23416 92598 23456
rect 92638 23416 92680 23456
rect 92720 23416 92729 23456
rect 96343 23416 96352 23456
rect 96392 23416 96434 23456
rect 96474 23416 96516 23456
rect 96556 23416 96598 23456
rect 96638 23416 96680 23456
rect 96720 23416 96729 23456
rect 88204 23248 88396 23288
rect 88436 23248 88445 23288
rect 89347 23248 89356 23288
rect 89396 23248 89644 23288
rect 89684 23248 89693 23288
rect 91171 23248 91180 23288
rect 91220 23248 91756 23288
rect 91796 23248 91805 23288
rect 93667 23248 93676 23288
rect 93716 23248 93964 23288
rect 94004 23248 94013 23288
rect 96067 23248 96076 23288
rect 96116 23248 96460 23288
rect 96500 23248 96509 23288
rect 0 23228 80 23248
rect 83587 23247 83645 23248
rect 80707 23164 80716 23204
rect 80756 23164 83788 23204
rect 83828 23164 85804 23204
rect 85844 23164 85853 23204
rect 88396 23164 91660 23204
rect 91700 23164 91709 23204
rect 86659 23120 86717 23121
rect 88396 23120 88436 23164
rect 835 23080 844 23120
rect 884 23080 1996 23120
rect 2036 23080 2045 23120
rect 80227 23080 80236 23120
rect 80276 23080 81004 23120
rect 81044 23080 81292 23120
rect 81332 23080 81580 23120
rect 81620 23080 81868 23120
rect 81908 23080 82156 23120
rect 82196 23080 82444 23120
rect 82484 23080 82493 23120
rect 82915 23080 82924 23120
rect 82964 23080 83212 23120
rect 83252 23080 84076 23120
rect 84116 23080 84364 23120
rect 84404 23080 84748 23120
rect 84788 23080 85132 23120
rect 85172 23080 85420 23120
rect 85460 23080 85469 23120
rect 86574 23080 86668 23120
rect 86708 23080 88436 23120
rect 89443 23080 89452 23120
rect 89492 23080 89836 23120
rect 89876 23080 90508 23120
rect 90548 23080 90892 23120
rect 90932 23080 91180 23120
rect 91220 23080 91229 23120
rect 95299 23080 95308 23120
rect 95348 23080 95692 23120
rect 95732 23080 95741 23120
rect 97795 23080 97804 23120
rect 97844 23080 98188 23120
rect 98228 23080 98237 23120
rect 86659 23079 86717 23080
rect 74755 22996 74764 23036
rect 74804 22996 75148 23036
rect 75188 22996 75724 23036
rect 75764 22996 76876 23036
rect 76916 22996 76925 23036
rect 78403 22996 78412 23036
rect 78452 22996 78988 23036
rect 79028 22996 79564 23036
rect 79604 22996 79756 23036
rect 79796 22996 79805 23036
rect 83971 22996 83980 23036
rect 84020 22996 84268 23036
rect 84308 22996 84317 23036
rect 85699 22996 85708 23036
rect 85748 22996 86284 23036
rect 86324 22996 86333 23036
rect 87523 22996 87532 23036
rect 87572 22996 87724 23036
rect 87764 22996 90316 23036
rect 90356 22996 90365 23036
rect 91843 22996 91852 23036
rect 91892 22996 92044 23036
rect 92084 22996 93484 23036
rect 93524 22996 93533 23036
rect 75619 22912 75628 22952
rect 75668 22912 76492 22952
rect 76532 22912 86476 22952
rect 86516 22912 86525 22952
rect 95683 22912 95692 22952
rect 95732 22912 96556 22952
rect 96596 22912 96844 22952
rect 96884 22912 97132 22952
rect 97172 22912 97420 22952
rect 97460 22912 97804 22952
rect 97844 22912 97853 22952
rect 87523 22868 87581 22869
rect 74563 22828 74572 22868
rect 74612 22828 75340 22868
rect 75380 22828 76108 22868
rect 76148 22828 77836 22868
rect 77876 22828 78796 22868
rect 78836 22828 78845 22868
rect 78988 22828 79276 22868
rect 79316 22828 79325 22868
rect 83299 22828 83308 22868
rect 83348 22828 83980 22868
rect 84020 22828 84029 22868
rect 87331 22828 87340 22868
rect 87380 22828 87532 22868
rect 87572 22828 87820 22868
rect 87860 22828 88108 22868
rect 88148 22828 88492 22868
rect 88532 22828 88780 22868
rect 88820 22828 88829 22868
rect 90307 22828 90316 22868
rect 90356 22828 90892 22868
rect 90932 22828 90941 22868
rect 91363 22828 91372 22868
rect 91412 22828 91421 22868
rect 78988 22700 79028 22828
rect 87523 22827 87581 22828
rect 91372 22784 91412 22828
rect 91372 22744 91604 22784
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 7103 22660 7112 22700
rect 7152 22660 7194 22700
rect 7234 22660 7276 22700
rect 7316 22660 7358 22700
rect 7398 22660 7440 22700
rect 7480 22660 7489 22700
rect 11103 22660 11112 22700
rect 11152 22660 11194 22700
rect 11234 22660 11276 22700
rect 11316 22660 11358 22700
rect 11398 22660 11440 22700
rect 11480 22660 11489 22700
rect 15103 22660 15112 22700
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15480 22660 15489 22700
rect 19103 22660 19112 22700
rect 19152 22660 19194 22700
rect 19234 22660 19276 22700
rect 19316 22660 19358 22700
rect 19398 22660 19440 22700
rect 19480 22660 19489 22700
rect 23103 22660 23112 22700
rect 23152 22660 23194 22700
rect 23234 22660 23276 22700
rect 23316 22660 23358 22700
rect 23398 22660 23440 22700
rect 23480 22660 23489 22700
rect 27103 22660 27112 22700
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27480 22660 27489 22700
rect 31103 22660 31112 22700
rect 31152 22660 31194 22700
rect 31234 22660 31276 22700
rect 31316 22660 31358 22700
rect 31398 22660 31440 22700
rect 31480 22660 31489 22700
rect 35103 22660 35112 22700
rect 35152 22660 35194 22700
rect 35234 22660 35276 22700
rect 35316 22660 35358 22700
rect 35398 22660 35440 22700
rect 35480 22660 35489 22700
rect 39103 22660 39112 22700
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39480 22660 39489 22700
rect 43103 22660 43112 22700
rect 43152 22660 43194 22700
rect 43234 22660 43276 22700
rect 43316 22660 43358 22700
rect 43398 22660 43440 22700
rect 43480 22660 43489 22700
rect 47103 22660 47112 22700
rect 47152 22660 47194 22700
rect 47234 22660 47276 22700
rect 47316 22660 47358 22700
rect 47398 22660 47440 22700
rect 47480 22660 47489 22700
rect 51103 22660 51112 22700
rect 51152 22660 51194 22700
rect 51234 22660 51276 22700
rect 51316 22660 51358 22700
rect 51398 22660 51440 22700
rect 51480 22660 51489 22700
rect 55103 22660 55112 22700
rect 55152 22660 55194 22700
rect 55234 22660 55276 22700
rect 55316 22660 55358 22700
rect 55398 22660 55440 22700
rect 55480 22660 55489 22700
rect 59103 22660 59112 22700
rect 59152 22660 59194 22700
rect 59234 22660 59276 22700
rect 59316 22660 59358 22700
rect 59398 22660 59440 22700
rect 59480 22660 59489 22700
rect 63103 22660 63112 22700
rect 63152 22660 63194 22700
rect 63234 22660 63276 22700
rect 63316 22660 63358 22700
rect 63398 22660 63440 22700
rect 63480 22660 63489 22700
rect 67103 22660 67112 22700
rect 67152 22660 67194 22700
rect 67234 22660 67276 22700
rect 67316 22660 67358 22700
rect 67398 22660 67440 22700
rect 67480 22660 67489 22700
rect 71103 22660 71112 22700
rect 71152 22660 71194 22700
rect 71234 22660 71276 22700
rect 71316 22660 71358 22700
rect 71398 22660 71440 22700
rect 71480 22660 71489 22700
rect 75103 22660 75112 22700
rect 75152 22660 75194 22700
rect 75234 22660 75276 22700
rect 75316 22660 75358 22700
rect 75398 22660 75440 22700
rect 75480 22660 75489 22700
rect 77251 22660 77260 22700
rect 77300 22660 77740 22700
rect 77780 22660 77789 22700
rect 78115 22660 78124 22700
rect 78164 22660 79028 22700
rect 79103 22660 79112 22700
rect 79152 22660 79194 22700
rect 79234 22660 79276 22700
rect 79316 22660 79358 22700
rect 79398 22660 79440 22700
rect 79480 22660 79489 22700
rect 83103 22660 83112 22700
rect 83152 22660 83194 22700
rect 83234 22660 83276 22700
rect 83316 22660 83358 22700
rect 83398 22660 83440 22700
rect 83480 22660 83489 22700
rect 83587 22660 83596 22700
rect 83636 22660 83788 22700
rect 83828 22660 83837 22700
rect 85891 22660 85900 22700
rect 85940 22660 86092 22700
rect 86132 22660 86572 22700
rect 86612 22660 86956 22700
rect 86996 22660 87005 22700
rect 87103 22660 87112 22700
rect 87152 22660 87194 22700
rect 87234 22660 87276 22700
rect 87316 22660 87358 22700
rect 87398 22660 87440 22700
rect 87480 22660 87489 22700
rect 91103 22660 91112 22700
rect 91152 22660 91194 22700
rect 91234 22660 91276 22700
rect 91316 22660 91358 22700
rect 91398 22660 91440 22700
rect 91480 22660 91489 22700
rect 85411 22532 85469 22533
rect 91564 22532 91604 22744
rect 92611 22660 92620 22700
rect 92660 22660 92908 22700
rect 92948 22660 93100 22700
rect 93140 22660 93292 22700
rect 93332 22660 93772 22700
rect 93812 22660 94060 22700
rect 94100 22660 94444 22700
rect 94484 22660 94493 22700
rect 95103 22660 95112 22700
rect 95152 22660 95194 22700
rect 95234 22660 95276 22700
rect 95316 22660 95358 22700
rect 95398 22660 95440 22700
rect 95480 22660 95489 22700
rect 95875 22660 95884 22700
rect 95924 22660 96364 22700
rect 96404 22660 96413 22700
rect 99103 22660 99112 22700
rect 99152 22660 99194 22700
rect 99234 22660 99276 22700
rect 99316 22660 99358 22700
rect 99398 22660 99440 22700
rect 99480 22660 99489 22700
rect 92227 22576 92236 22616
rect 92276 22576 92524 22616
rect 92564 22576 92573 22616
rect 75235 22492 75244 22532
rect 75284 22492 75436 22532
rect 75476 22492 80716 22532
rect 80756 22492 80765 22532
rect 85326 22492 85420 22532
rect 85460 22492 85469 22532
rect 87043 22492 87052 22532
rect 87092 22492 87628 22532
rect 87668 22492 87677 22532
rect 89347 22492 89356 22532
rect 89396 22492 89740 22532
rect 89780 22492 90124 22532
rect 90164 22492 90604 22532
rect 90644 22492 91276 22532
rect 91316 22492 91604 22532
rect 93475 22492 93484 22532
rect 93524 22492 95404 22532
rect 95444 22492 96076 22532
rect 96116 22492 96125 22532
rect 85411 22491 85469 22492
rect 0 22448 80 22468
rect 94915 22448 94973 22449
rect 0 22408 556 22448
rect 596 22408 605 22448
rect 86380 22408 86668 22448
rect 86708 22408 86717 22448
rect 90988 22408 91852 22448
rect 91892 22408 92276 22448
rect 0 22388 80 22408
rect 83587 22364 83645 22365
rect 86380 22364 86420 22408
rect 90988 22364 91028 22408
rect 92236 22364 92276 22408
rect 94915 22408 94924 22448
rect 94964 22408 95116 22448
rect 95156 22408 95165 22448
rect 95299 22408 95308 22448
rect 95348 22408 95788 22448
rect 95828 22408 95837 22448
rect 94915 22407 94973 22408
rect 77731 22324 77740 22364
rect 77780 22324 78124 22364
rect 78164 22324 78173 22364
rect 79939 22324 79948 22364
rect 79988 22324 80428 22364
rect 80468 22324 81676 22364
rect 81716 22324 82636 22364
rect 82676 22324 82685 22364
rect 83502 22324 83596 22364
rect 83636 22324 83645 22364
rect 83779 22324 83788 22364
rect 83828 22324 84556 22364
rect 84596 22324 84940 22364
rect 84980 22324 85612 22364
rect 85652 22324 85804 22364
rect 85844 22324 85853 22364
rect 86371 22324 86380 22364
rect 86420 22324 86429 22364
rect 86563 22324 86572 22364
rect 86612 22324 87628 22364
rect 87668 22324 88396 22364
rect 88436 22324 88876 22364
rect 88916 22324 88925 22364
rect 90499 22324 90508 22364
rect 90548 22324 90988 22364
rect 91028 22324 91037 22364
rect 92227 22324 92236 22364
rect 92276 22324 92285 22364
rect 93763 22324 93772 22364
rect 93812 22324 94924 22364
rect 94964 22324 94973 22364
rect 95683 22324 95692 22364
rect 95732 22324 96076 22364
rect 96116 22324 96364 22364
rect 96404 22324 97228 22364
rect 97268 22324 98188 22364
rect 98228 22324 98237 22364
rect 83587 22323 83645 22324
rect 74371 22240 74380 22280
rect 74420 22240 75052 22280
rect 75092 22240 75820 22280
rect 75860 22240 77164 22280
rect 77204 22240 78796 22280
rect 78836 22240 78845 22280
rect 86275 22240 86284 22280
rect 86324 22240 86956 22280
rect 86996 22240 87724 22280
rect 87764 22240 87773 22280
rect 91075 22240 91084 22280
rect 91124 22240 91948 22280
rect 91988 22240 91997 22280
rect 87523 22196 87581 22197
rect 87235 22156 87244 22196
rect 87284 22156 87532 22196
rect 87572 22156 88012 22196
rect 88052 22156 88061 22196
rect 87523 22155 87581 22156
rect 93772 22112 93812 22324
rect 75715 22072 75724 22112
rect 75764 22072 76108 22112
rect 76148 22072 76588 22112
rect 76628 22072 76820 22112
rect 92611 22072 92620 22112
rect 92660 22072 93484 22112
rect 93524 22072 93812 22112
rect 931 21988 940 22028
rect 980 21988 9388 22028
rect 9428 21988 9437 22028
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 8343 21904 8352 21944
rect 8392 21904 8434 21944
rect 8474 21904 8516 21944
rect 8556 21904 8598 21944
rect 8638 21904 8680 21944
rect 8720 21904 8729 21944
rect 12343 21904 12352 21944
rect 12392 21904 12434 21944
rect 12474 21904 12516 21944
rect 12556 21904 12598 21944
rect 12638 21904 12680 21944
rect 12720 21904 12729 21944
rect 16343 21904 16352 21944
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16720 21904 16729 21944
rect 20343 21904 20352 21944
rect 20392 21904 20434 21944
rect 20474 21904 20516 21944
rect 20556 21904 20598 21944
rect 20638 21904 20680 21944
rect 20720 21904 20729 21944
rect 24343 21904 24352 21944
rect 24392 21904 24434 21944
rect 24474 21904 24516 21944
rect 24556 21904 24598 21944
rect 24638 21904 24680 21944
rect 24720 21904 24729 21944
rect 28343 21904 28352 21944
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28720 21904 28729 21944
rect 32343 21904 32352 21944
rect 32392 21904 32434 21944
rect 32474 21904 32516 21944
rect 32556 21904 32598 21944
rect 32638 21904 32680 21944
rect 32720 21904 32729 21944
rect 36343 21904 36352 21944
rect 36392 21904 36434 21944
rect 36474 21904 36516 21944
rect 36556 21904 36598 21944
rect 36638 21904 36680 21944
rect 36720 21904 36729 21944
rect 40343 21904 40352 21944
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40720 21904 40729 21944
rect 44343 21904 44352 21944
rect 44392 21904 44434 21944
rect 44474 21904 44516 21944
rect 44556 21904 44598 21944
rect 44638 21904 44680 21944
rect 44720 21904 44729 21944
rect 48343 21904 48352 21944
rect 48392 21904 48434 21944
rect 48474 21904 48516 21944
rect 48556 21904 48598 21944
rect 48638 21904 48680 21944
rect 48720 21904 48729 21944
rect 52343 21904 52352 21944
rect 52392 21904 52434 21944
rect 52474 21904 52516 21944
rect 52556 21904 52598 21944
rect 52638 21904 52680 21944
rect 52720 21904 52729 21944
rect 56343 21904 56352 21944
rect 56392 21904 56434 21944
rect 56474 21904 56516 21944
rect 56556 21904 56598 21944
rect 56638 21904 56680 21944
rect 56720 21904 56729 21944
rect 60343 21904 60352 21944
rect 60392 21904 60434 21944
rect 60474 21904 60516 21944
rect 60556 21904 60598 21944
rect 60638 21904 60680 21944
rect 60720 21904 60729 21944
rect 64343 21904 64352 21944
rect 64392 21904 64434 21944
rect 64474 21904 64516 21944
rect 64556 21904 64598 21944
rect 64638 21904 64680 21944
rect 64720 21904 64729 21944
rect 68343 21904 68352 21944
rect 68392 21904 68434 21944
rect 68474 21904 68516 21944
rect 68556 21904 68598 21944
rect 68638 21904 68680 21944
rect 68720 21904 68729 21944
rect 72343 21904 72352 21944
rect 72392 21904 72434 21944
rect 72474 21904 72516 21944
rect 72556 21904 72598 21944
rect 72638 21904 72680 21944
rect 72720 21904 72729 21944
rect 76343 21904 76352 21944
rect 76392 21904 76434 21944
rect 76474 21904 76516 21944
rect 76556 21904 76598 21944
rect 76638 21904 76680 21944
rect 76720 21904 76729 21944
rect 76780 21860 76820 22072
rect 80343 21904 80352 21944
rect 80392 21904 80434 21944
rect 80474 21904 80516 21944
rect 80556 21904 80598 21944
rect 80638 21904 80680 21944
rect 80720 21904 80729 21944
rect 84343 21904 84352 21944
rect 84392 21904 84434 21944
rect 84474 21904 84516 21944
rect 84556 21904 84598 21944
rect 84638 21904 84680 21944
rect 84720 21904 84729 21944
rect 88343 21904 88352 21944
rect 88392 21904 88434 21944
rect 88474 21904 88516 21944
rect 88556 21904 88598 21944
rect 88638 21904 88680 21944
rect 88720 21904 88729 21944
rect 92343 21904 92352 21944
rect 92392 21904 92434 21944
rect 92474 21904 92516 21944
rect 92556 21904 92598 21944
rect 92638 21904 92680 21944
rect 92720 21904 92729 21944
rect 96343 21904 96352 21944
rect 96392 21904 96434 21944
rect 96474 21904 96516 21944
rect 96556 21904 96598 21944
rect 96638 21904 96680 21944
rect 96720 21904 96729 21944
rect 76588 21820 76820 21860
rect 76588 21776 76628 21820
rect 84259 21776 84317 21777
rect 95011 21776 95069 21777
rect 76579 21736 76588 21776
rect 76628 21736 76637 21776
rect 84259 21736 84268 21776
rect 84308 21736 84364 21776
rect 84404 21736 84413 21776
rect 95011 21736 95020 21776
rect 95060 21736 95212 21776
rect 95252 21736 95261 21776
rect 84259 21735 84317 21736
rect 95011 21735 95069 21736
rect 0 21608 80 21628
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 92707 21568 92716 21608
rect 92756 21568 93388 21608
rect 93428 21568 93437 21608
rect 0 21548 80 21568
rect 77539 21484 77548 21524
rect 77588 21484 77740 21524
rect 77780 21484 78892 21524
rect 78932 21484 79276 21524
rect 79316 21484 79325 21524
rect 80803 21484 80812 21524
rect 80852 21484 82156 21524
rect 82196 21484 82636 21524
rect 82676 21484 82685 21524
rect 83395 21484 83404 21524
rect 83444 21484 83788 21524
rect 83828 21484 84172 21524
rect 84212 21484 84221 21524
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 7103 21148 7112 21188
rect 7152 21148 7194 21188
rect 7234 21148 7276 21188
rect 7316 21148 7358 21188
rect 7398 21148 7440 21188
rect 7480 21148 7489 21188
rect 11103 21148 11112 21188
rect 11152 21148 11194 21188
rect 11234 21148 11276 21188
rect 11316 21148 11358 21188
rect 11398 21148 11440 21188
rect 11480 21148 11489 21188
rect 15103 21148 15112 21188
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15480 21148 15489 21188
rect 19103 21148 19112 21188
rect 19152 21148 19194 21188
rect 19234 21148 19276 21188
rect 19316 21148 19358 21188
rect 19398 21148 19440 21188
rect 19480 21148 19489 21188
rect 23103 21148 23112 21188
rect 23152 21148 23194 21188
rect 23234 21148 23276 21188
rect 23316 21148 23358 21188
rect 23398 21148 23440 21188
rect 23480 21148 23489 21188
rect 27103 21148 27112 21188
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27480 21148 27489 21188
rect 31103 21148 31112 21188
rect 31152 21148 31194 21188
rect 31234 21148 31276 21188
rect 31316 21148 31358 21188
rect 31398 21148 31440 21188
rect 31480 21148 31489 21188
rect 35103 21148 35112 21188
rect 35152 21148 35194 21188
rect 35234 21148 35276 21188
rect 35316 21148 35358 21188
rect 35398 21148 35440 21188
rect 35480 21148 35489 21188
rect 39103 21148 39112 21188
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39480 21148 39489 21188
rect 43103 21148 43112 21188
rect 43152 21148 43194 21188
rect 43234 21148 43276 21188
rect 43316 21148 43358 21188
rect 43398 21148 43440 21188
rect 43480 21148 43489 21188
rect 47103 21148 47112 21188
rect 47152 21148 47194 21188
rect 47234 21148 47276 21188
rect 47316 21148 47358 21188
rect 47398 21148 47440 21188
rect 47480 21148 47489 21188
rect 51103 21148 51112 21188
rect 51152 21148 51194 21188
rect 51234 21148 51276 21188
rect 51316 21148 51358 21188
rect 51398 21148 51440 21188
rect 51480 21148 51489 21188
rect 55103 21148 55112 21188
rect 55152 21148 55194 21188
rect 55234 21148 55276 21188
rect 55316 21148 55358 21188
rect 55398 21148 55440 21188
rect 55480 21148 55489 21188
rect 59103 21148 59112 21188
rect 59152 21148 59194 21188
rect 59234 21148 59276 21188
rect 59316 21148 59358 21188
rect 59398 21148 59440 21188
rect 59480 21148 59489 21188
rect 63103 21148 63112 21188
rect 63152 21148 63194 21188
rect 63234 21148 63276 21188
rect 63316 21148 63358 21188
rect 63398 21148 63440 21188
rect 63480 21148 63489 21188
rect 67103 21148 67112 21188
rect 67152 21148 67194 21188
rect 67234 21148 67276 21188
rect 67316 21148 67358 21188
rect 67398 21148 67440 21188
rect 67480 21148 67489 21188
rect 71103 21148 71112 21188
rect 71152 21148 71194 21188
rect 71234 21148 71276 21188
rect 71316 21148 71358 21188
rect 71398 21148 71440 21188
rect 71480 21148 71489 21188
rect 75103 21148 75112 21188
rect 75152 21148 75194 21188
rect 75234 21148 75276 21188
rect 75316 21148 75358 21188
rect 75398 21148 75440 21188
rect 75480 21148 75489 21188
rect 79103 21148 79112 21188
rect 79152 21148 79194 21188
rect 79234 21148 79276 21188
rect 79316 21148 79358 21188
rect 79398 21148 79440 21188
rect 79480 21148 79489 21188
rect 83103 21148 83112 21188
rect 83152 21148 83194 21188
rect 83234 21148 83276 21188
rect 83316 21148 83358 21188
rect 83398 21148 83440 21188
rect 83480 21148 83489 21188
rect 87103 21148 87112 21188
rect 87152 21148 87194 21188
rect 87234 21148 87276 21188
rect 87316 21148 87358 21188
rect 87398 21148 87440 21188
rect 87480 21148 87489 21188
rect 91103 21148 91112 21188
rect 91152 21148 91194 21188
rect 91234 21148 91276 21188
rect 91316 21148 91358 21188
rect 91398 21148 91440 21188
rect 91480 21148 91489 21188
rect 95103 21148 95112 21188
rect 95152 21148 95194 21188
rect 95234 21148 95276 21188
rect 95316 21148 95358 21188
rect 95398 21148 95440 21188
rect 95480 21148 95489 21188
rect 99103 21148 99112 21188
rect 99152 21148 99194 21188
rect 99234 21148 99276 21188
rect 99316 21148 99358 21188
rect 99398 21148 99440 21188
rect 99480 21148 99489 21188
rect 0 20768 80 20788
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 0 20708 80 20728
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 8343 20392 8352 20432
rect 8392 20392 8434 20432
rect 8474 20392 8516 20432
rect 8556 20392 8598 20432
rect 8638 20392 8680 20432
rect 8720 20392 8729 20432
rect 12343 20392 12352 20432
rect 12392 20392 12434 20432
rect 12474 20392 12516 20432
rect 12556 20392 12598 20432
rect 12638 20392 12680 20432
rect 12720 20392 12729 20432
rect 16343 20392 16352 20432
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16720 20392 16729 20432
rect 20343 20392 20352 20432
rect 20392 20392 20434 20432
rect 20474 20392 20516 20432
rect 20556 20392 20598 20432
rect 20638 20392 20680 20432
rect 20720 20392 20729 20432
rect 24343 20392 24352 20432
rect 24392 20392 24434 20432
rect 24474 20392 24516 20432
rect 24556 20392 24598 20432
rect 24638 20392 24680 20432
rect 24720 20392 24729 20432
rect 28343 20392 28352 20432
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28720 20392 28729 20432
rect 32343 20392 32352 20432
rect 32392 20392 32434 20432
rect 32474 20392 32516 20432
rect 32556 20392 32598 20432
rect 32638 20392 32680 20432
rect 32720 20392 32729 20432
rect 36343 20392 36352 20432
rect 36392 20392 36434 20432
rect 36474 20392 36516 20432
rect 36556 20392 36598 20432
rect 36638 20392 36680 20432
rect 36720 20392 36729 20432
rect 40343 20392 40352 20432
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40720 20392 40729 20432
rect 44343 20392 44352 20432
rect 44392 20392 44434 20432
rect 44474 20392 44516 20432
rect 44556 20392 44598 20432
rect 44638 20392 44680 20432
rect 44720 20392 44729 20432
rect 48343 20392 48352 20432
rect 48392 20392 48434 20432
rect 48474 20392 48516 20432
rect 48556 20392 48598 20432
rect 48638 20392 48680 20432
rect 48720 20392 48729 20432
rect 52343 20392 52352 20432
rect 52392 20392 52434 20432
rect 52474 20392 52516 20432
rect 52556 20392 52598 20432
rect 52638 20392 52680 20432
rect 52720 20392 52729 20432
rect 56343 20392 56352 20432
rect 56392 20392 56434 20432
rect 56474 20392 56516 20432
rect 56556 20392 56598 20432
rect 56638 20392 56680 20432
rect 56720 20392 56729 20432
rect 60343 20392 60352 20432
rect 60392 20392 60434 20432
rect 60474 20392 60516 20432
rect 60556 20392 60598 20432
rect 60638 20392 60680 20432
rect 60720 20392 60729 20432
rect 64343 20392 64352 20432
rect 64392 20392 64434 20432
rect 64474 20392 64516 20432
rect 64556 20392 64598 20432
rect 64638 20392 64680 20432
rect 64720 20392 64729 20432
rect 68343 20392 68352 20432
rect 68392 20392 68434 20432
rect 68474 20392 68516 20432
rect 68556 20392 68598 20432
rect 68638 20392 68680 20432
rect 68720 20392 68729 20432
rect 72343 20392 72352 20432
rect 72392 20392 72434 20432
rect 72474 20392 72516 20432
rect 72556 20392 72598 20432
rect 72638 20392 72680 20432
rect 72720 20392 72729 20432
rect 76343 20392 76352 20432
rect 76392 20392 76434 20432
rect 76474 20392 76516 20432
rect 76556 20392 76598 20432
rect 76638 20392 76680 20432
rect 76720 20392 76729 20432
rect 80343 20392 80352 20432
rect 80392 20392 80434 20432
rect 80474 20392 80516 20432
rect 80556 20392 80598 20432
rect 80638 20392 80680 20432
rect 80720 20392 80729 20432
rect 84343 20392 84352 20432
rect 84392 20392 84434 20432
rect 84474 20392 84516 20432
rect 84556 20392 84598 20432
rect 84638 20392 84680 20432
rect 84720 20392 84729 20432
rect 88343 20392 88352 20432
rect 88392 20392 88434 20432
rect 88474 20392 88516 20432
rect 88556 20392 88598 20432
rect 88638 20392 88680 20432
rect 88720 20392 88729 20432
rect 92343 20392 92352 20432
rect 92392 20392 92434 20432
rect 92474 20392 92516 20432
rect 92556 20392 92598 20432
rect 92638 20392 92680 20432
rect 92720 20392 92729 20432
rect 96343 20392 96352 20432
rect 96392 20392 96434 20432
rect 96474 20392 96516 20432
rect 96556 20392 96598 20432
rect 96638 20392 96680 20432
rect 96720 20392 96729 20432
rect 75724 19972 80620 20012
rect 80660 19972 86860 20012
rect 86900 19972 86909 20012
rect 0 19928 80 19948
rect 75724 19928 75764 19972
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 75715 19888 75724 19928
rect 75764 19888 75773 19928
rect 0 19868 80 19888
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 7103 19636 7112 19676
rect 7152 19636 7194 19676
rect 7234 19636 7276 19676
rect 7316 19636 7358 19676
rect 7398 19636 7440 19676
rect 7480 19636 7489 19676
rect 11103 19636 11112 19676
rect 11152 19636 11194 19676
rect 11234 19636 11276 19676
rect 11316 19636 11358 19676
rect 11398 19636 11440 19676
rect 11480 19636 11489 19676
rect 15103 19636 15112 19676
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15480 19636 15489 19676
rect 19103 19636 19112 19676
rect 19152 19636 19194 19676
rect 19234 19636 19276 19676
rect 19316 19636 19358 19676
rect 19398 19636 19440 19676
rect 19480 19636 19489 19676
rect 23103 19636 23112 19676
rect 23152 19636 23194 19676
rect 23234 19636 23276 19676
rect 23316 19636 23358 19676
rect 23398 19636 23440 19676
rect 23480 19636 23489 19676
rect 27103 19636 27112 19676
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27480 19636 27489 19676
rect 31103 19636 31112 19676
rect 31152 19636 31194 19676
rect 31234 19636 31276 19676
rect 31316 19636 31358 19676
rect 31398 19636 31440 19676
rect 31480 19636 31489 19676
rect 35103 19636 35112 19676
rect 35152 19636 35194 19676
rect 35234 19636 35276 19676
rect 35316 19636 35358 19676
rect 35398 19636 35440 19676
rect 35480 19636 35489 19676
rect 39103 19636 39112 19676
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39480 19636 39489 19676
rect 43103 19636 43112 19676
rect 43152 19636 43194 19676
rect 43234 19636 43276 19676
rect 43316 19636 43358 19676
rect 43398 19636 43440 19676
rect 43480 19636 43489 19676
rect 47103 19636 47112 19676
rect 47152 19636 47194 19676
rect 47234 19636 47276 19676
rect 47316 19636 47358 19676
rect 47398 19636 47440 19676
rect 47480 19636 47489 19676
rect 51103 19636 51112 19676
rect 51152 19636 51194 19676
rect 51234 19636 51276 19676
rect 51316 19636 51358 19676
rect 51398 19636 51440 19676
rect 51480 19636 51489 19676
rect 55103 19636 55112 19676
rect 55152 19636 55194 19676
rect 55234 19636 55276 19676
rect 55316 19636 55358 19676
rect 55398 19636 55440 19676
rect 55480 19636 55489 19676
rect 59103 19636 59112 19676
rect 59152 19636 59194 19676
rect 59234 19636 59276 19676
rect 59316 19636 59358 19676
rect 59398 19636 59440 19676
rect 59480 19636 59489 19676
rect 63103 19636 63112 19676
rect 63152 19636 63194 19676
rect 63234 19636 63276 19676
rect 63316 19636 63358 19676
rect 63398 19636 63440 19676
rect 63480 19636 63489 19676
rect 67103 19636 67112 19676
rect 67152 19636 67194 19676
rect 67234 19636 67276 19676
rect 67316 19636 67358 19676
rect 67398 19636 67440 19676
rect 67480 19636 67489 19676
rect 71103 19636 71112 19676
rect 71152 19636 71194 19676
rect 71234 19636 71276 19676
rect 71316 19636 71358 19676
rect 71398 19636 71440 19676
rect 71480 19636 71489 19676
rect 75103 19636 75112 19676
rect 75152 19636 75194 19676
rect 75234 19636 75276 19676
rect 75316 19636 75358 19676
rect 75398 19636 75440 19676
rect 75480 19636 75489 19676
rect 79103 19636 79112 19676
rect 79152 19636 79194 19676
rect 79234 19636 79276 19676
rect 79316 19636 79358 19676
rect 79398 19636 79440 19676
rect 79480 19636 79489 19676
rect 83103 19636 83112 19676
rect 83152 19636 83194 19676
rect 83234 19636 83276 19676
rect 83316 19636 83358 19676
rect 83398 19636 83440 19676
rect 83480 19636 83489 19676
rect 87103 19636 87112 19676
rect 87152 19636 87194 19676
rect 87234 19636 87276 19676
rect 87316 19636 87358 19676
rect 87398 19636 87440 19676
rect 87480 19636 87489 19676
rect 91103 19636 91112 19676
rect 91152 19636 91194 19676
rect 91234 19636 91276 19676
rect 91316 19636 91358 19676
rect 91398 19636 91440 19676
rect 91480 19636 91489 19676
rect 95103 19636 95112 19676
rect 95152 19636 95194 19676
rect 95234 19636 95276 19676
rect 95316 19636 95358 19676
rect 95398 19636 95440 19676
rect 95480 19636 95489 19676
rect 99103 19636 99112 19676
rect 99152 19636 99194 19676
rect 99234 19636 99276 19676
rect 99316 19636 99358 19676
rect 99398 19636 99440 19676
rect 99480 19636 99489 19676
rect 86755 19340 86813 19341
rect 80515 19300 80524 19340
rect 80564 19300 82060 19340
rect 82100 19300 82348 19340
rect 82388 19300 84076 19340
rect 84116 19300 85612 19340
rect 85652 19300 85661 19340
rect 86670 19300 86764 19340
rect 86804 19300 86956 19340
rect 86996 19300 87005 19340
rect 88195 19300 88204 19340
rect 88244 19300 88253 19340
rect 93091 19300 93100 19340
rect 93140 19300 94156 19340
rect 94196 19300 95788 19340
rect 95828 19300 97132 19340
rect 97172 19300 97181 19340
rect 86755 19299 86813 19300
rect 88204 19256 88244 19300
rect 71779 19216 71788 19256
rect 71828 19216 75436 19256
rect 75476 19216 75724 19256
rect 75764 19216 75773 19256
rect 75820 19216 76588 19256
rect 76628 19216 76637 19256
rect 86563 19216 86572 19256
rect 86612 19216 89932 19256
rect 89972 19216 93196 19256
rect 93236 19216 93245 19256
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 0 19028 80 19048
rect 75820 18920 75860 19216
rect 86956 19172 86996 19216
rect 81859 19132 81868 19172
rect 81908 19132 82636 19172
rect 82676 19132 83020 19172
rect 83060 19132 83069 19172
rect 86947 19132 86956 19172
rect 86996 19132 87005 19172
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 8343 18880 8352 18920
rect 8392 18880 8434 18920
rect 8474 18880 8516 18920
rect 8556 18880 8598 18920
rect 8638 18880 8680 18920
rect 8720 18880 8729 18920
rect 12343 18880 12352 18920
rect 12392 18880 12434 18920
rect 12474 18880 12516 18920
rect 12556 18880 12598 18920
rect 12638 18880 12680 18920
rect 12720 18880 12729 18920
rect 16343 18880 16352 18920
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16720 18880 16729 18920
rect 20343 18880 20352 18920
rect 20392 18880 20434 18920
rect 20474 18880 20516 18920
rect 20556 18880 20598 18920
rect 20638 18880 20680 18920
rect 20720 18880 20729 18920
rect 24343 18880 24352 18920
rect 24392 18880 24434 18920
rect 24474 18880 24516 18920
rect 24556 18880 24598 18920
rect 24638 18880 24680 18920
rect 24720 18880 24729 18920
rect 28343 18880 28352 18920
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28720 18880 28729 18920
rect 32343 18880 32352 18920
rect 32392 18880 32434 18920
rect 32474 18880 32516 18920
rect 32556 18880 32598 18920
rect 32638 18880 32680 18920
rect 32720 18880 32729 18920
rect 36343 18880 36352 18920
rect 36392 18880 36434 18920
rect 36474 18880 36516 18920
rect 36556 18880 36598 18920
rect 36638 18880 36680 18920
rect 36720 18880 36729 18920
rect 40343 18880 40352 18920
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40720 18880 40729 18920
rect 44343 18880 44352 18920
rect 44392 18880 44434 18920
rect 44474 18880 44516 18920
rect 44556 18880 44598 18920
rect 44638 18880 44680 18920
rect 44720 18880 44729 18920
rect 48343 18880 48352 18920
rect 48392 18880 48434 18920
rect 48474 18880 48516 18920
rect 48556 18880 48598 18920
rect 48638 18880 48680 18920
rect 48720 18880 48729 18920
rect 52343 18880 52352 18920
rect 52392 18880 52434 18920
rect 52474 18880 52516 18920
rect 52556 18880 52598 18920
rect 52638 18880 52680 18920
rect 52720 18880 52729 18920
rect 56343 18880 56352 18920
rect 56392 18880 56434 18920
rect 56474 18880 56516 18920
rect 56556 18880 56598 18920
rect 56638 18880 56680 18920
rect 56720 18880 56729 18920
rect 60343 18880 60352 18920
rect 60392 18880 60434 18920
rect 60474 18880 60516 18920
rect 60556 18880 60598 18920
rect 60638 18880 60680 18920
rect 60720 18880 60729 18920
rect 64343 18880 64352 18920
rect 64392 18880 64434 18920
rect 64474 18880 64516 18920
rect 64556 18880 64598 18920
rect 64638 18880 64680 18920
rect 64720 18880 64729 18920
rect 68343 18880 68352 18920
rect 68392 18880 68434 18920
rect 68474 18880 68516 18920
rect 68556 18880 68598 18920
rect 68638 18880 68680 18920
rect 68720 18880 68729 18920
rect 72343 18880 72352 18920
rect 72392 18880 72434 18920
rect 72474 18880 72516 18920
rect 72556 18880 72598 18920
rect 72638 18880 72680 18920
rect 72720 18880 72729 18920
rect 75139 18880 75148 18920
rect 75188 18880 75820 18920
rect 75860 18880 76204 18920
rect 76244 18880 76253 18920
rect 76343 18880 76352 18920
rect 76392 18880 76434 18920
rect 76474 18880 76516 18920
rect 76556 18880 76598 18920
rect 76638 18880 76680 18920
rect 76720 18880 76729 18920
rect 78115 18880 78124 18920
rect 78164 18880 78604 18920
rect 78644 18880 79372 18920
rect 79412 18880 79421 18920
rect 80343 18880 80352 18920
rect 80392 18880 80434 18920
rect 80474 18880 80516 18920
rect 80556 18880 80598 18920
rect 80638 18880 80680 18920
rect 80720 18880 80729 18920
rect 84343 18880 84352 18920
rect 84392 18880 84434 18920
rect 84474 18880 84516 18920
rect 84556 18880 84598 18920
rect 84638 18880 84680 18920
rect 84720 18880 84729 18920
rect 88343 18880 88352 18920
rect 88392 18880 88434 18920
rect 88474 18880 88516 18920
rect 88556 18880 88598 18920
rect 88638 18880 88680 18920
rect 88720 18880 88729 18920
rect 90115 18880 90124 18920
rect 90164 18880 90508 18920
rect 90548 18880 91372 18920
rect 91412 18880 91421 18920
rect 92343 18880 92352 18920
rect 92392 18880 92434 18920
rect 92474 18880 92516 18920
rect 92556 18880 92598 18920
rect 92638 18880 92680 18920
rect 92720 18880 92729 18920
rect 96343 18880 96352 18920
rect 96392 18880 96434 18920
rect 96474 18880 96516 18920
rect 96556 18880 96598 18920
rect 96638 18880 96680 18920
rect 96720 18880 96729 18920
rect 74563 18796 74572 18836
rect 74612 18796 74956 18836
rect 74996 18796 75628 18836
rect 75668 18796 76972 18836
rect 77012 18796 77021 18836
rect 77443 18796 77452 18836
rect 77492 18796 78220 18836
rect 78260 18796 78988 18836
rect 79028 18796 79037 18836
rect 68227 18544 68236 18584
rect 68276 18544 72940 18584
rect 72980 18544 73708 18584
rect 73748 18544 73757 18584
rect 74275 18544 74284 18584
rect 74324 18544 75244 18584
rect 75284 18544 76492 18584
rect 76532 18544 77452 18584
rect 77492 18544 77501 18584
rect 86563 18544 86572 18584
rect 86612 18544 87052 18584
rect 87092 18544 87436 18584
rect 87476 18544 89012 18584
rect 91459 18544 91468 18584
rect 91508 18544 91852 18584
rect 91892 18544 92236 18584
rect 92276 18544 92285 18584
rect 93187 18544 93196 18584
rect 93236 18544 95116 18584
rect 95156 18544 95165 18584
rect 88972 18500 89012 18544
rect 78403 18460 78412 18500
rect 78452 18460 78796 18500
rect 78836 18460 78845 18500
rect 79363 18460 79372 18500
rect 79412 18460 79852 18500
rect 79892 18460 79901 18500
rect 80035 18460 80044 18500
rect 80084 18460 80524 18500
rect 80564 18460 81004 18500
rect 81044 18460 81388 18500
rect 81428 18460 81437 18500
rect 83395 18460 83404 18500
rect 83444 18460 83788 18500
rect 83828 18460 84268 18500
rect 84308 18460 84652 18500
rect 84692 18460 85036 18500
rect 85076 18460 85085 18500
rect 85507 18460 85516 18500
rect 85556 18460 85900 18500
rect 85940 18460 86284 18500
rect 86324 18460 86333 18500
rect 87715 18460 87724 18500
rect 87764 18460 88012 18500
rect 88052 18460 88204 18500
rect 88244 18460 88588 18500
rect 88628 18460 88637 18500
rect 88963 18460 88972 18500
rect 89012 18460 89021 18500
rect 89539 18460 89548 18500
rect 89588 18460 89740 18500
rect 89780 18460 90124 18500
rect 90164 18460 90604 18500
rect 90644 18460 92620 18500
rect 92660 18460 92669 18500
rect 92899 18460 92908 18500
rect 92948 18460 93100 18500
rect 93140 18460 93149 18500
rect 94531 18292 94540 18332
rect 94580 18292 95212 18332
rect 95252 18292 95261 18332
rect 95491 18292 95500 18332
rect 95540 18292 95636 18332
rect 0 18248 80 18268
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 78979 18208 78988 18248
rect 79028 18208 79852 18248
rect 79892 18208 79901 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 7103 18124 7112 18164
rect 7152 18124 7194 18164
rect 7234 18124 7276 18164
rect 7316 18124 7358 18164
rect 7398 18124 7440 18164
rect 7480 18124 7489 18164
rect 11103 18124 11112 18164
rect 11152 18124 11194 18164
rect 11234 18124 11276 18164
rect 11316 18124 11358 18164
rect 11398 18124 11440 18164
rect 11480 18124 11489 18164
rect 15103 18124 15112 18164
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15480 18124 15489 18164
rect 19103 18124 19112 18164
rect 19152 18124 19194 18164
rect 19234 18124 19276 18164
rect 19316 18124 19358 18164
rect 19398 18124 19440 18164
rect 19480 18124 19489 18164
rect 23103 18124 23112 18164
rect 23152 18124 23194 18164
rect 23234 18124 23276 18164
rect 23316 18124 23358 18164
rect 23398 18124 23440 18164
rect 23480 18124 23489 18164
rect 27103 18124 27112 18164
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27480 18124 27489 18164
rect 31103 18124 31112 18164
rect 31152 18124 31194 18164
rect 31234 18124 31276 18164
rect 31316 18124 31358 18164
rect 31398 18124 31440 18164
rect 31480 18124 31489 18164
rect 35103 18124 35112 18164
rect 35152 18124 35194 18164
rect 35234 18124 35276 18164
rect 35316 18124 35358 18164
rect 35398 18124 35440 18164
rect 35480 18124 35489 18164
rect 39103 18124 39112 18164
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39480 18124 39489 18164
rect 43103 18124 43112 18164
rect 43152 18124 43194 18164
rect 43234 18124 43276 18164
rect 43316 18124 43358 18164
rect 43398 18124 43440 18164
rect 43480 18124 43489 18164
rect 47103 18124 47112 18164
rect 47152 18124 47194 18164
rect 47234 18124 47276 18164
rect 47316 18124 47358 18164
rect 47398 18124 47440 18164
rect 47480 18124 47489 18164
rect 51103 18124 51112 18164
rect 51152 18124 51194 18164
rect 51234 18124 51276 18164
rect 51316 18124 51358 18164
rect 51398 18124 51440 18164
rect 51480 18124 51489 18164
rect 55103 18124 55112 18164
rect 55152 18124 55194 18164
rect 55234 18124 55276 18164
rect 55316 18124 55358 18164
rect 55398 18124 55440 18164
rect 55480 18124 55489 18164
rect 59103 18124 59112 18164
rect 59152 18124 59194 18164
rect 59234 18124 59276 18164
rect 59316 18124 59358 18164
rect 59398 18124 59440 18164
rect 59480 18124 59489 18164
rect 63103 18124 63112 18164
rect 63152 18124 63194 18164
rect 63234 18124 63276 18164
rect 63316 18124 63358 18164
rect 63398 18124 63440 18164
rect 63480 18124 63489 18164
rect 67103 18124 67112 18164
rect 67152 18124 67194 18164
rect 67234 18124 67276 18164
rect 67316 18124 67358 18164
rect 67398 18124 67440 18164
rect 67480 18124 67489 18164
rect 71103 18124 71112 18164
rect 71152 18124 71194 18164
rect 71234 18124 71276 18164
rect 71316 18124 71358 18164
rect 71398 18124 71440 18164
rect 71480 18124 71489 18164
rect 75103 18124 75112 18164
rect 75152 18124 75194 18164
rect 75234 18124 75276 18164
rect 75316 18124 75358 18164
rect 75398 18124 75440 18164
rect 75480 18124 75489 18164
rect 79103 18124 79112 18164
rect 79152 18124 79194 18164
rect 79234 18124 79276 18164
rect 79316 18124 79358 18164
rect 79398 18124 79440 18164
rect 79480 18124 79489 18164
rect 83103 18124 83112 18164
rect 83152 18124 83194 18164
rect 83234 18124 83276 18164
rect 83316 18124 83358 18164
rect 83398 18124 83440 18164
rect 83480 18124 83489 18164
rect 87103 18124 87112 18164
rect 87152 18124 87194 18164
rect 87234 18124 87276 18164
rect 87316 18124 87358 18164
rect 87398 18124 87440 18164
rect 87480 18124 87489 18164
rect 91103 18124 91112 18164
rect 91152 18124 91194 18164
rect 91234 18124 91276 18164
rect 91316 18124 91358 18164
rect 91398 18124 91440 18164
rect 91480 18124 91489 18164
rect 95103 18124 95112 18164
rect 95152 18124 95194 18164
rect 95234 18124 95276 18164
rect 95316 18124 95358 18164
rect 95398 18124 95440 18164
rect 95480 18124 95489 18164
rect 95596 17996 95636 18292
rect 99103 18124 99112 18164
rect 99152 18124 99194 18164
rect 99234 18124 99276 18164
rect 99316 18124 99358 18164
rect 99398 18124 99440 18164
rect 99480 18124 99489 18164
rect 92803 17956 92812 17996
rect 92852 17956 93196 17996
rect 93236 17956 93245 17996
rect 95395 17956 95404 17996
rect 95444 17956 95884 17996
rect 95924 17956 96076 17996
rect 96116 17956 96364 17996
rect 96404 17956 96652 17996
rect 96692 17956 98476 17996
rect 98516 17956 98525 17996
rect 78787 17872 78796 17912
rect 78836 17872 79180 17912
rect 79220 17872 79468 17912
rect 79508 17872 79517 17912
rect 97315 17872 97324 17912
rect 97364 17872 97404 17912
rect 97324 17828 97364 17872
rect 73699 17788 73708 17828
rect 73748 17788 74092 17828
rect 74132 17788 74141 17828
rect 76579 17788 76588 17828
rect 76628 17788 76972 17828
rect 77012 17788 77021 17828
rect 77347 17788 77356 17828
rect 77396 17788 77740 17828
rect 77780 17788 78220 17828
rect 78260 17788 78269 17828
rect 84739 17788 84748 17828
rect 84788 17788 84940 17828
rect 84980 17788 85420 17828
rect 85460 17788 85469 17828
rect 93187 17788 93196 17828
rect 93236 17788 93772 17828
rect 93812 17788 94732 17828
rect 94772 17788 94924 17828
rect 94964 17788 94973 17828
rect 97027 17788 97036 17828
rect 97076 17788 97900 17828
rect 97940 17788 98708 17828
rect 98668 17744 98708 17788
rect 75811 17704 75820 17744
rect 75860 17704 76492 17744
rect 76532 17704 76541 17744
rect 81283 17704 81292 17744
rect 81332 17704 81484 17744
rect 81524 17704 81533 17744
rect 81955 17704 81964 17744
rect 82004 17704 82348 17744
rect 82388 17704 82397 17744
rect 83395 17704 83404 17744
rect 83444 17704 83788 17744
rect 83828 17704 84172 17744
rect 84212 17704 84221 17744
rect 86179 17704 86188 17744
rect 86228 17704 86572 17744
rect 86612 17704 87052 17744
rect 87092 17704 87436 17744
rect 87476 17704 87485 17744
rect 88579 17704 88588 17744
rect 88628 17704 89068 17744
rect 89108 17704 89117 17744
rect 89443 17704 89452 17744
rect 89492 17704 89932 17744
rect 89972 17704 90220 17744
rect 90260 17704 90269 17744
rect 90595 17704 90604 17744
rect 90644 17704 90988 17744
rect 91028 17704 91037 17744
rect 91363 17704 91372 17744
rect 91412 17704 91852 17744
rect 91892 17704 92236 17744
rect 92276 17704 92285 17744
rect 98659 17704 98668 17744
rect 98708 17704 98717 17744
rect 84643 17620 84652 17660
rect 84692 17620 84701 17660
rect 87907 17620 87916 17660
rect 87956 17620 88108 17660
rect 88148 17620 88157 17660
rect 92899 17620 92908 17660
rect 92948 17620 93484 17660
rect 93524 17620 93533 17660
rect 97891 17620 97900 17660
rect 97940 17620 98764 17660
rect 98804 17620 98813 17660
rect 84259 17576 84317 17577
rect 76675 17536 76684 17576
rect 76724 17536 76733 17576
rect 80707 17536 80716 17576
rect 80756 17536 81004 17576
rect 81044 17536 81053 17576
rect 84259 17536 84268 17576
rect 84308 17536 84460 17576
rect 84500 17536 84509 17576
rect 76684 17492 76724 17536
rect 84259 17535 84317 17536
rect 84652 17492 84692 17620
rect 88204 17536 88396 17576
rect 88436 17536 88445 17576
rect 76684 17452 76820 17492
rect 84652 17452 85036 17492
rect 85076 17452 85085 17492
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 8343 17368 8352 17408
rect 8392 17368 8434 17408
rect 8474 17368 8516 17408
rect 8556 17368 8598 17408
rect 8638 17368 8680 17408
rect 8720 17368 8729 17408
rect 12343 17368 12352 17408
rect 12392 17368 12434 17408
rect 12474 17368 12516 17408
rect 12556 17368 12598 17408
rect 12638 17368 12680 17408
rect 12720 17368 12729 17408
rect 16343 17368 16352 17408
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16720 17368 16729 17408
rect 20343 17368 20352 17408
rect 20392 17368 20434 17408
rect 20474 17368 20516 17408
rect 20556 17368 20598 17408
rect 20638 17368 20680 17408
rect 20720 17368 20729 17408
rect 24343 17368 24352 17408
rect 24392 17368 24434 17408
rect 24474 17368 24516 17408
rect 24556 17368 24598 17408
rect 24638 17368 24680 17408
rect 24720 17368 24729 17408
rect 28343 17368 28352 17408
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28720 17368 28729 17408
rect 32343 17368 32352 17408
rect 32392 17368 32434 17408
rect 32474 17368 32516 17408
rect 32556 17368 32598 17408
rect 32638 17368 32680 17408
rect 32720 17368 32729 17408
rect 36343 17368 36352 17408
rect 36392 17368 36434 17408
rect 36474 17368 36516 17408
rect 36556 17368 36598 17408
rect 36638 17368 36680 17408
rect 36720 17368 36729 17408
rect 40343 17368 40352 17408
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40720 17368 40729 17408
rect 44343 17368 44352 17408
rect 44392 17368 44434 17408
rect 44474 17368 44516 17408
rect 44556 17368 44598 17408
rect 44638 17368 44680 17408
rect 44720 17368 44729 17408
rect 48343 17368 48352 17408
rect 48392 17368 48434 17408
rect 48474 17368 48516 17408
rect 48556 17368 48598 17408
rect 48638 17368 48680 17408
rect 48720 17368 48729 17408
rect 52343 17368 52352 17408
rect 52392 17368 52434 17408
rect 52474 17368 52516 17408
rect 52556 17368 52598 17408
rect 52638 17368 52680 17408
rect 52720 17368 52729 17408
rect 56343 17368 56352 17408
rect 56392 17368 56434 17408
rect 56474 17368 56516 17408
rect 56556 17368 56598 17408
rect 56638 17368 56680 17408
rect 56720 17368 56729 17408
rect 60343 17368 60352 17408
rect 60392 17368 60434 17408
rect 60474 17368 60516 17408
rect 60556 17368 60598 17408
rect 60638 17368 60680 17408
rect 60720 17368 60729 17408
rect 64343 17368 64352 17408
rect 64392 17368 64434 17408
rect 64474 17368 64516 17408
rect 64556 17368 64598 17408
rect 64638 17368 64680 17408
rect 64720 17368 64729 17408
rect 68343 17368 68352 17408
rect 68392 17368 68434 17408
rect 68474 17368 68516 17408
rect 68556 17368 68598 17408
rect 68638 17368 68680 17408
rect 68720 17368 68729 17408
rect 72343 17368 72352 17408
rect 72392 17368 72434 17408
rect 72474 17368 72516 17408
rect 72556 17368 72598 17408
rect 72638 17368 72680 17408
rect 72720 17368 72729 17408
rect 76343 17368 76352 17408
rect 76392 17368 76434 17408
rect 76474 17368 76516 17408
rect 76556 17368 76598 17408
rect 76638 17368 76680 17408
rect 76720 17368 76729 17408
rect 0 17348 80 17368
rect 76780 17240 76820 17452
rect 80343 17368 80352 17408
rect 80392 17368 80434 17408
rect 80474 17368 80516 17408
rect 80556 17368 80598 17408
rect 80638 17368 80680 17408
rect 80720 17368 80729 17408
rect 84343 17368 84352 17408
rect 84392 17368 84434 17408
rect 84474 17368 84516 17408
rect 84556 17368 84598 17408
rect 84638 17368 84680 17408
rect 84720 17368 84729 17408
rect 76675 17200 76684 17240
rect 76724 17200 76820 17240
rect 88204 17240 88244 17536
rect 88343 17368 88352 17408
rect 88392 17368 88434 17408
rect 88474 17368 88516 17408
rect 88556 17368 88598 17408
rect 88638 17368 88680 17408
rect 88720 17368 88729 17408
rect 92343 17368 92352 17408
rect 92392 17368 92434 17408
rect 92474 17368 92516 17408
rect 92556 17368 92598 17408
rect 92638 17368 92680 17408
rect 92720 17368 92729 17408
rect 96343 17368 96352 17408
rect 96392 17368 96434 17408
rect 96474 17368 96516 17408
rect 96556 17368 96598 17408
rect 96638 17368 96680 17408
rect 96720 17368 96729 17408
rect 88204 17200 88396 17240
rect 88436 17200 88445 17240
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 7103 16612 7112 16652
rect 7152 16612 7194 16652
rect 7234 16612 7276 16652
rect 7316 16612 7358 16652
rect 7398 16612 7440 16652
rect 7480 16612 7489 16652
rect 11103 16612 11112 16652
rect 11152 16612 11194 16652
rect 11234 16612 11276 16652
rect 11316 16612 11358 16652
rect 11398 16612 11440 16652
rect 11480 16612 11489 16652
rect 15103 16612 15112 16652
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15480 16612 15489 16652
rect 19103 16612 19112 16652
rect 19152 16612 19194 16652
rect 19234 16612 19276 16652
rect 19316 16612 19358 16652
rect 19398 16612 19440 16652
rect 19480 16612 19489 16652
rect 23103 16612 23112 16652
rect 23152 16612 23194 16652
rect 23234 16612 23276 16652
rect 23316 16612 23358 16652
rect 23398 16612 23440 16652
rect 23480 16612 23489 16652
rect 27103 16612 27112 16652
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27480 16612 27489 16652
rect 31103 16612 31112 16652
rect 31152 16612 31194 16652
rect 31234 16612 31276 16652
rect 31316 16612 31358 16652
rect 31398 16612 31440 16652
rect 31480 16612 31489 16652
rect 35103 16612 35112 16652
rect 35152 16612 35194 16652
rect 35234 16612 35276 16652
rect 35316 16612 35358 16652
rect 35398 16612 35440 16652
rect 35480 16612 35489 16652
rect 39103 16612 39112 16652
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39480 16612 39489 16652
rect 43103 16612 43112 16652
rect 43152 16612 43194 16652
rect 43234 16612 43276 16652
rect 43316 16612 43358 16652
rect 43398 16612 43440 16652
rect 43480 16612 43489 16652
rect 47103 16612 47112 16652
rect 47152 16612 47194 16652
rect 47234 16612 47276 16652
rect 47316 16612 47358 16652
rect 47398 16612 47440 16652
rect 47480 16612 47489 16652
rect 51103 16612 51112 16652
rect 51152 16612 51194 16652
rect 51234 16612 51276 16652
rect 51316 16612 51358 16652
rect 51398 16612 51440 16652
rect 51480 16612 51489 16652
rect 55103 16612 55112 16652
rect 55152 16612 55194 16652
rect 55234 16612 55276 16652
rect 55316 16612 55358 16652
rect 55398 16612 55440 16652
rect 55480 16612 55489 16652
rect 59103 16612 59112 16652
rect 59152 16612 59194 16652
rect 59234 16612 59276 16652
rect 59316 16612 59358 16652
rect 59398 16612 59440 16652
rect 59480 16612 59489 16652
rect 63103 16612 63112 16652
rect 63152 16612 63194 16652
rect 63234 16612 63276 16652
rect 63316 16612 63358 16652
rect 63398 16612 63440 16652
rect 63480 16612 63489 16652
rect 67103 16612 67112 16652
rect 67152 16612 67194 16652
rect 67234 16612 67276 16652
rect 67316 16612 67358 16652
rect 67398 16612 67440 16652
rect 67480 16612 67489 16652
rect 0 16568 80 16588
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 74179 16528 74188 16568
rect 74228 16528 74668 16568
rect 74708 16528 74717 16568
rect 91171 16528 91180 16568
rect 91220 16528 91660 16568
rect 91700 16528 91709 16568
rect 0 16508 80 16528
rect 96739 16360 96748 16400
rect 96788 16360 97516 16400
rect 97556 16360 97565 16400
rect 71683 16024 71692 16064
rect 71732 16024 75340 16064
rect 75380 16024 75389 16064
rect 67363 15940 67372 15980
rect 67412 15940 73228 15980
rect 73268 15940 73277 15980
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 8343 15856 8352 15896
rect 8392 15856 8434 15896
rect 8474 15856 8516 15896
rect 8556 15856 8598 15896
rect 8638 15856 8680 15896
rect 8720 15856 8729 15896
rect 12343 15856 12352 15896
rect 12392 15856 12434 15896
rect 12474 15856 12516 15896
rect 12556 15856 12598 15896
rect 12638 15856 12680 15896
rect 12720 15856 12729 15896
rect 16343 15856 16352 15896
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16720 15856 16729 15896
rect 20343 15856 20352 15896
rect 20392 15856 20434 15896
rect 20474 15856 20516 15896
rect 20556 15856 20598 15896
rect 20638 15856 20680 15896
rect 20720 15856 20729 15896
rect 24343 15856 24352 15896
rect 24392 15856 24434 15896
rect 24474 15856 24516 15896
rect 24556 15856 24598 15896
rect 24638 15856 24680 15896
rect 24720 15856 24729 15896
rect 28343 15856 28352 15896
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28720 15856 28729 15896
rect 32343 15856 32352 15896
rect 32392 15856 32434 15896
rect 32474 15856 32516 15896
rect 32556 15856 32598 15896
rect 32638 15856 32680 15896
rect 32720 15856 32729 15896
rect 36343 15856 36352 15896
rect 36392 15856 36434 15896
rect 36474 15856 36516 15896
rect 36556 15856 36598 15896
rect 36638 15856 36680 15896
rect 36720 15856 36729 15896
rect 40343 15856 40352 15896
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40720 15856 40729 15896
rect 44343 15856 44352 15896
rect 44392 15856 44434 15896
rect 44474 15856 44516 15896
rect 44556 15856 44598 15896
rect 44638 15856 44680 15896
rect 44720 15856 44729 15896
rect 48343 15856 48352 15896
rect 48392 15856 48434 15896
rect 48474 15856 48516 15896
rect 48556 15856 48598 15896
rect 48638 15856 48680 15896
rect 48720 15856 48729 15896
rect 52343 15856 52352 15896
rect 52392 15856 52434 15896
rect 52474 15856 52516 15896
rect 52556 15856 52598 15896
rect 52638 15856 52680 15896
rect 52720 15856 52729 15896
rect 56343 15856 56352 15896
rect 56392 15856 56434 15896
rect 56474 15856 56516 15896
rect 56556 15856 56598 15896
rect 56638 15856 56680 15896
rect 56720 15856 56729 15896
rect 60343 15856 60352 15896
rect 60392 15856 60434 15896
rect 60474 15856 60516 15896
rect 60556 15856 60598 15896
rect 60638 15856 60680 15896
rect 60720 15856 60729 15896
rect 64343 15856 64352 15896
rect 64392 15856 64434 15896
rect 64474 15856 64516 15896
rect 64556 15856 64598 15896
rect 64638 15856 64680 15896
rect 64720 15856 64729 15896
rect 68343 15856 68352 15896
rect 68392 15856 68434 15896
rect 68474 15856 68516 15896
rect 68556 15856 68598 15896
rect 68638 15856 68680 15896
rect 68720 15856 68729 15896
rect 68803 15856 68812 15896
rect 68852 15856 73900 15896
rect 73940 15856 73949 15896
rect 69955 15772 69964 15812
rect 70004 15772 74284 15812
rect 74324 15772 74333 15812
rect 0 15728 80 15748
rect 0 15688 652 15728
rect 692 15688 701 15728
rect 69859 15688 69868 15728
rect 69908 15688 73652 15728
rect 89827 15688 89836 15728
rect 89876 15688 89885 15728
rect 0 15668 80 15688
rect 73612 15644 73652 15688
rect 69475 15604 69484 15644
rect 69524 15604 73132 15644
rect 73172 15604 73181 15644
rect 73603 15604 73612 15644
rect 73652 15604 73661 15644
rect 71779 15560 71837 15561
rect 84259 15560 84317 15561
rect 67171 15520 67180 15560
rect 67220 15520 67564 15560
rect 67604 15520 68428 15560
rect 68468 15520 69100 15560
rect 69140 15520 69149 15560
rect 71779 15520 71788 15560
rect 71828 15520 72815 15560
rect 72855 15520 72864 15560
rect 73027 15520 73036 15560
rect 73076 15520 73505 15560
rect 73545 15520 73554 15560
rect 77827 15520 77836 15560
rect 77876 15520 77885 15560
rect 78499 15520 78508 15560
rect 78548 15520 79215 15560
rect 79255 15520 79264 15560
rect 84259 15520 84268 15560
rect 84308 15520 84415 15560
rect 84455 15520 84464 15560
rect 84696 15520 84705 15560
rect 84745 15520 84940 15560
rect 84980 15520 84989 15560
rect 71779 15519 71837 15520
rect 1987 15436 1996 15476
rect 2036 15436 67756 15476
rect 67796 15436 71692 15476
rect 71732 15436 71741 15476
rect 71788 15436 72705 15476
rect 72745 15436 72754 15476
rect 71788 15224 71828 15436
rect 71875 15392 71933 15393
rect 77836 15392 77876 15520
rect 84259 15519 84317 15520
rect 89836 15476 89876 15688
rect 96067 15604 96076 15644
rect 96116 15604 96125 15644
rect 92131 15520 92140 15560
rect 92180 15520 92415 15560
rect 92455 15520 92464 15560
rect 89496 15436 89505 15476
rect 89545 15436 89876 15476
rect 96076 15392 96116 15604
rect 96163 15520 96172 15560
rect 96212 15520 96415 15560
rect 96455 15520 96464 15560
rect 98851 15476 98909 15477
rect 98406 15436 98415 15476
rect 98455 15436 98860 15476
rect 98900 15436 98909 15476
rect 98851 15435 98909 15436
rect 71875 15352 71884 15392
rect 71924 15352 72415 15392
rect 72455 15352 72464 15392
rect 75096 15352 75105 15392
rect 75145 15352 75724 15392
rect 75764 15352 75773 15392
rect 77836 15352 77905 15392
rect 77945 15352 77954 15392
rect 78806 15352 78815 15392
rect 78855 15352 78988 15392
rect 79028 15352 79037 15392
rect 96006 15352 96015 15392
rect 96055 15352 96116 15392
rect 98296 15352 98305 15392
rect 98345 15352 98956 15392
rect 98996 15352 99005 15392
rect 71875 15351 71933 15352
rect 71788 15184 71924 15224
rect 71884 15140 71924 15184
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 7103 15100 7112 15140
rect 7152 15100 7194 15140
rect 7234 15100 7276 15140
rect 7316 15100 7358 15140
rect 7398 15100 7440 15140
rect 7480 15100 7489 15140
rect 11103 15100 11112 15140
rect 11152 15100 11194 15140
rect 11234 15100 11276 15140
rect 11316 15100 11358 15140
rect 11398 15100 11440 15140
rect 11480 15100 11489 15140
rect 15103 15100 15112 15140
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15480 15100 15489 15140
rect 19103 15100 19112 15140
rect 19152 15100 19194 15140
rect 19234 15100 19276 15140
rect 19316 15100 19358 15140
rect 19398 15100 19440 15140
rect 19480 15100 19489 15140
rect 23103 15100 23112 15140
rect 23152 15100 23194 15140
rect 23234 15100 23276 15140
rect 23316 15100 23358 15140
rect 23398 15100 23440 15140
rect 23480 15100 23489 15140
rect 27103 15100 27112 15140
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27480 15100 27489 15140
rect 31103 15100 31112 15140
rect 31152 15100 31194 15140
rect 31234 15100 31276 15140
rect 31316 15100 31358 15140
rect 31398 15100 31440 15140
rect 31480 15100 31489 15140
rect 35103 15100 35112 15140
rect 35152 15100 35194 15140
rect 35234 15100 35276 15140
rect 35316 15100 35358 15140
rect 35398 15100 35440 15140
rect 35480 15100 35489 15140
rect 39103 15100 39112 15140
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39480 15100 39489 15140
rect 43103 15100 43112 15140
rect 43152 15100 43194 15140
rect 43234 15100 43276 15140
rect 43316 15100 43358 15140
rect 43398 15100 43440 15140
rect 43480 15100 43489 15140
rect 47103 15100 47112 15140
rect 47152 15100 47194 15140
rect 47234 15100 47276 15140
rect 47316 15100 47358 15140
rect 47398 15100 47440 15140
rect 47480 15100 47489 15140
rect 51103 15100 51112 15140
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51480 15100 51489 15140
rect 55103 15100 55112 15140
rect 55152 15100 55194 15140
rect 55234 15100 55276 15140
rect 55316 15100 55358 15140
rect 55398 15100 55440 15140
rect 55480 15100 55489 15140
rect 59103 15100 59112 15140
rect 59152 15100 59194 15140
rect 59234 15100 59276 15140
rect 59316 15100 59358 15140
rect 59398 15100 59440 15140
rect 59480 15100 59489 15140
rect 63103 15100 63112 15140
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63480 15100 63489 15140
rect 67103 15100 67112 15140
rect 67152 15100 67194 15140
rect 67234 15100 67276 15140
rect 67316 15100 67358 15140
rect 67398 15100 67440 15140
rect 67480 15100 67489 15140
rect 71683 15100 71692 15140
rect 71732 15100 71924 15140
rect 71779 15056 71837 15057
rect 69283 15016 69292 15056
rect 69332 15016 71788 15056
rect 71828 15016 71837 15056
rect 71779 15015 71837 15016
rect 835 14932 844 14972
rect 884 14932 1708 14972
rect 1748 14932 1757 14972
rect 69091 14932 69100 14972
rect 69140 14932 71884 14972
rect 71924 14932 71933 14972
rect 0 14888 80 14908
rect 71875 14888 71933 14889
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 69283 14848 69292 14888
rect 69332 14848 71884 14888
rect 71924 14848 71933 14888
rect 0 14828 80 14848
rect 71875 14847 71933 14848
rect 68035 14764 68044 14804
rect 68084 14764 71692 14804
rect 71732 14764 71741 14804
rect 68131 14680 68140 14720
rect 68180 14680 68620 14720
rect 68660 14680 69388 14720
rect 69428 14680 69437 14720
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 8343 14344 8352 14384
rect 8392 14344 8434 14384
rect 8474 14344 8516 14384
rect 8556 14344 8598 14384
rect 8638 14344 8680 14384
rect 8720 14344 8729 14384
rect 12343 14344 12352 14384
rect 12392 14344 12434 14384
rect 12474 14344 12516 14384
rect 12556 14344 12598 14384
rect 12638 14344 12680 14384
rect 12720 14344 12729 14384
rect 16343 14344 16352 14384
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16720 14344 16729 14384
rect 20343 14344 20352 14384
rect 20392 14344 20434 14384
rect 20474 14344 20516 14384
rect 20556 14344 20598 14384
rect 20638 14344 20680 14384
rect 20720 14344 20729 14384
rect 24343 14344 24352 14384
rect 24392 14344 24434 14384
rect 24474 14344 24516 14384
rect 24556 14344 24598 14384
rect 24638 14344 24680 14384
rect 24720 14344 24729 14384
rect 28343 14344 28352 14384
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28720 14344 28729 14384
rect 32343 14344 32352 14384
rect 32392 14344 32434 14384
rect 32474 14344 32516 14384
rect 32556 14344 32598 14384
rect 32638 14344 32680 14384
rect 32720 14344 32729 14384
rect 36343 14344 36352 14384
rect 36392 14344 36434 14384
rect 36474 14344 36516 14384
rect 36556 14344 36598 14384
rect 36638 14344 36680 14384
rect 36720 14344 36729 14384
rect 40343 14344 40352 14384
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40720 14344 40729 14384
rect 44343 14344 44352 14384
rect 44392 14344 44434 14384
rect 44474 14344 44516 14384
rect 44556 14344 44598 14384
rect 44638 14344 44680 14384
rect 44720 14344 44729 14384
rect 48343 14344 48352 14384
rect 48392 14344 48434 14384
rect 48474 14344 48516 14384
rect 48556 14344 48598 14384
rect 48638 14344 48680 14384
rect 48720 14344 48729 14384
rect 52343 14344 52352 14384
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52720 14344 52729 14384
rect 56343 14344 56352 14384
rect 56392 14344 56434 14384
rect 56474 14344 56516 14384
rect 56556 14344 56598 14384
rect 56638 14344 56680 14384
rect 56720 14344 56729 14384
rect 60343 14344 60352 14384
rect 60392 14344 60434 14384
rect 60474 14344 60516 14384
rect 60556 14344 60598 14384
rect 60638 14344 60680 14384
rect 60720 14344 60729 14384
rect 64343 14344 64352 14384
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64720 14344 64729 14384
rect 68343 14344 68352 14384
rect 68392 14344 68434 14384
rect 68474 14344 68516 14384
rect 68556 14344 68598 14384
rect 68638 14344 68680 14384
rect 68720 14344 68729 14384
rect 835 14176 844 14216
rect 884 14176 1324 14216
rect 1364 14176 1373 14216
rect 0 14048 80 14068
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 0 13988 80 14008
rect 9379 13924 9388 13964
rect 9428 13924 69004 13964
rect 69044 13924 69196 13964
rect 69236 13924 70060 13964
rect 70100 13924 70109 13964
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 7103 13588 7112 13628
rect 7152 13588 7194 13628
rect 7234 13588 7276 13628
rect 7316 13588 7358 13628
rect 7398 13588 7440 13628
rect 7480 13588 7489 13628
rect 11103 13588 11112 13628
rect 11152 13588 11194 13628
rect 11234 13588 11276 13628
rect 11316 13588 11358 13628
rect 11398 13588 11440 13628
rect 11480 13588 11489 13628
rect 15103 13588 15112 13628
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15480 13588 15489 13628
rect 19103 13588 19112 13628
rect 19152 13588 19194 13628
rect 19234 13588 19276 13628
rect 19316 13588 19358 13628
rect 19398 13588 19440 13628
rect 19480 13588 19489 13628
rect 23103 13588 23112 13628
rect 23152 13588 23194 13628
rect 23234 13588 23276 13628
rect 23316 13588 23358 13628
rect 23398 13588 23440 13628
rect 23480 13588 23489 13628
rect 27103 13588 27112 13628
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27480 13588 27489 13628
rect 31103 13588 31112 13628
rect 31152 13588 31194 13628
rect 31234 13588 31276 13628
rect 31316 13588 31358 13628
rect 31398 13588 31440 13628
rect 31480 13588 31489 13628
rect 35103 13588 35112 13628
rect 35152 13588 35194 13628
rect 35234 13588 35276 13628
rect 35316 13588 35358 13628
rect 35398 13588 35440 13628
rect 35480 13588 35489 13628
rect 39103 13588 39112 13628
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39480 13588 39489 13628
rect 43103 13588 43112 13628
rect 43152 13588 43194 13628
rect 43234 13588 43276 13628
rect 43316 13588 43358 13628
rect 43398 13588 43440 13628
rect 43480 13588 43489 13628
rect 47103 13588 47112 13628
rect 47152 13588 47194 13628
rect 47234 13588 47276 13628
rect 47316 13588 47358 13628
rect 47398 13588 47440 13628
rect 47480 13588 47489 13628
rect 51103 13588 51112 13628
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51480 13588 51489 13628
rect 55103 13588 55112 13628
rect 55152 13588 55194 13628
rect 55234 13588 55276 13628
rect 55316 13588 55358 13628
rect 55398 13588 55440 13628
rect 55480 13588 55489 13628
rect 59103 13588 59112 13628
rect 59152 13588 59194 13628
rect 59234 13588 59276 13628
rect 59316 13588 59358 13628
rect 59398 13588 59440 13628
rect 59480 13588 59489 13628
rect 63103 13588 63112 13628
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63480 13588 63489 13628
rect 67103 13588 67112 13628
rect 67152 13588 67194 13628
rect 67234 13588 67276 13628
rect 67316 13588 67358 13628
rect 67398 13588 67440 13628
rect 67480 13588 67489 13628
rect 835 13336 844 13376
rect 884 13336 1708 13376
rect 1748 13336 1757 13376
rect 0 13208 80 13228
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 0 13148 80 13168
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 8343 12832 8352 12872
rect 8392 12832 8434 12872
rect 8474 12832 8516 12872
rect 8556 12832 8598 12872
rect 8638 12832 8680 12872
rect 8720 12832 8729 12872
rect 12343 12832 12352 12872
rect 12392 12832 12434 12872
rect 12474 12832 12516 12872
rect 12556 12832 12598 12872
rect 12638 12832 12680 12872
rect 12720 12832 12729 12872
rect 16343 12832 16352 12872
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16720 12832 16729 12872
rect 20343 12832 20352 12872
rect 20392 12832 20434 12872
rect 20474 12832 20516 12872
rect 20556 12832 20598 12872
rect 20638 12832 20680 12872
rect 20720 12832 20729 12872
rect 24343 12832 24352 12872
rect 24392 12832 24434 12872
rect 24474 12832 24516 12872
rect 24556 12832 24598 12872
rect 24638 12832 24680 12872
rect 24720 12832 24729 12872
rect 28343 12832 28352 12872
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28720 12832 28729 12872
rect 32343 12832 32352 12872
rect 32392 12832 32434 12872
rect 32474 12832 32516 12872
rect 32556 12832 32598 12872
rect 32638 12832 32680 12872
rect 32720 12832 32729 12872
rect 36343 12832 36352 12872
rect 36392 12832 36434 12872
rect 36474 12832 36516 12872
rect 36556 12832 36598 12872
rect 36638 12832 36680 12872
rect 36720 12832 36729 12872
rect 40343 12832 40352 12872
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40720 12832 40729 12872
rect 44343 12832 44352 12872
rect 44392 12832 44434 12872
rect 44474 12832 44516 12872
rect 44556 12832 44598 12872
rect 44638 12832 44680 12872
rect 44720 12832 44729 12872
rect 48343 12832 48352 12872
rect 48392 12832 48434 12872
rect 48474 12832 48516 12872
rect 48556 12832 48598 12872
rect 48638 12832 48680 12872
rect 48720 12832 48729 12872
rect 52343 12832 52352 12872
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52720 12832 52729 12872
rect 56343 12832 56352 12872
rect 56392 12832 56434 12872
rect 56474 12832 56516 12872
rect 56556 12832 56598 12872
rect 56638 12832 56680 12872
rect 56720 12832 56729 12872
rect 60343 12832 60352 12872
rect 60392 12832 60434 12872
rect 60474 12832 60516 12872
rect 60556 12832 60598 12872
rect 60638 12832 60680 12872
rect 60720 12832 60729 12872
rect 64343 12832 64352 12872
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64720 12832 64729 12872
rect 68343 12832 68352 12872
rect 68392 12832 68434 12872
rect 68474 12832 68516 12872
rect 68556 12832 68598 12872
rect 68638 12832 68680 12872
rect 68720 12832 68729 12872
rect 0 12368 80 12388
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 0 12308 80 12328
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 7103 12076 7112 12116
rect 7152 12076 7194 12116
rect 7234 12076 7276 12116
rect 7316 12076 7358 12116
rect 7398 12076 7440 12116
rect 7480 12076 7489 12116
rect 11103 12076 11112 12116
rect 11152 12076 11194 12116
rect 11234 12076 11276 12116
rect 11316 12076 11358 12116
rect 11398 12076 11440 12116
rect 11480 12076 11489 12116
rect 15103 12076 15112 12116
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15480 12076 15489 12116
rect 19103 12076 19112 12116
rect 19152 12076 19194 12116
rect 19234 12076 19276 12116
rect 19316 12076 19358 12116
rect 19398 12076 19440 12116
rect 19480 12076 19489 12116
rect 23103 12076 23112 12116
rect 23152 12076 23194 12116
rect 23234 12076 23276 12116
rect 23316 12076 23358 12116
rect 23398 12076 23440 12116
rect 23480 12076 23489 12116
rect 27103 12076 27112 12116
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27480 12076 27489 12116
rect 31103 12076 31112 12116
rect 31152 12076 31194 12116
rect 31234 12076 31276 12116
rect 31316 12076 31358 12116
rect 31398 12076 31440 12116
rect 31480 12076 31489 12116
rect 35103 12076 35112 12116
rect 35152 12076 35194 12116
rect 35234 12076 35276 12116
rect 35316 12076 35358 12116
rect 35398 12076 35440 12116
rect 35480 12076 35489 12116
rect 39103 12076 39112 12116
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39480 12076 39489 12116
rect 43103 12076 43112 12116
rect 43152 12076 43194 12116
rect 43234 12076 43276 12116
rect 43316 12076 43358 12116
rect 43398 12076 43440 12116
rect 43480 12076 43489 12116
rect 47103 12076 47112 12116
rect 47152 12076 47194 12116
rect 47234 12076 47276 12116
rect 47316 12076 47358 12116
rect 47398 12076 47440 12116
rect 47480 12076 47489 12116
rect 51103 12076 51112 12116
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51480 12076 51489 12116
rect 55103 12076 55112 12116
rect 55152 12076 55194 12116
rect 55234 12076 55276 12116
rect 55316 12076 55358 12116
rect 55398 12076 55440 12116
rect 55480 12076 55489 12116
rect 59103 12076 59112 12116
rect 59152 12076 59194 12116
rect 59234 12076 59276 12116
rect 59316 12076 59358 12116
rect 59398 12076 59440 12116
rect 59480 12076 59489 12116
rect 63103 12076 63112 12116
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63480 12076 63489 12116
rect 67103 12076 67112 12116
rect 67152 12076 67194 12116
rect 67234 12076 67276 12116
rect 67316 12076 67358 12116
rect 67398 12076 67440 12116
rect 67480 12076 67489 12116
rect 835 11908 844 11948
rect 884 11908 1996 11948
rect 2036 11908 2045 11948
rect 835 11740 844 11780
rect 884 11740 1612 11780
rect 1652 11740 1661 11780
rect 0 11528 80 11548
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 0 11468 80 11488
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 8343 11320 8352 11360
rect 8392 11320 8434 11360
rect 8474 11320 8516 11360
rect 8556 11320 8598 11360
rect 8638 11320 8680 11360
rect 8720 11320 8729 11360
rect 12343 11320 12352 11360
rect 12392 11320 12434 11360
rect 12474 11320 12516 11360
rect 12556 11320 12598 11360
rect 12638 11320 12680 11360
rect 12720 11320 12729 11360
rect 16343 11320 16352 11360
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16720 11320 16729 11360
rect 20343 11320 20352 11360
rect 20392 11320 20434 11360
rect 20474 11320 20516 11360
rect 20556 11320 20598 11360
rect 20638 11320 20680 11360
rect 20720 11320 20729 11360
rect 24343 11320 24352 11360
rect 24392 11320 24434 11360
rect 24474 11320 24516 11360
rect 24556 11320 24598 11360
rect 24638 11320 24680 11360
rect 24720 11320 24729 11360
rect 28343 11320 28352 11360
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28720 11320 28729 11360
rect 32343 11320 32352 11360
rect 32392 11320 32434 11360
rect 32474 11320 32516 11360
rect 32556 11320 32598 11360
rect 32638 11320 32680 11360
rect 32720 11320 32729 11360
rect 36343 11320 36352 11360
rect 36392 11320 36434 11360
rect 36474 11320 36516 11360
rect 36556 11320 36598 11360
rect 36638 11320 36680 11360
rect 36720 11320 36729 11360
rect 40343 11320 40352 11360
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40720 11320 40729 11360
rect 44343 11320 44352 11360
rect 44392 11320 44434 11360
rect 44474 11320 44516 11360
rect 44556 11320 44598 11360
rect 44638 11320 44680 11360
rect 44720 11320 44729 11360
rect 48343 11320 48352 11360
rect 48392 11320 48434 11360
rect 48474 11320 48516 11360
rect 48556 11320 48598 11360
rect 48638 11320 48680 11360
rect 48720 11320 48729 11360
rect 52343 11320 52352 11360
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52720 11320 52729 11360
rect 56343 11320 56352 11360
rect 56392 11320 56434 11360
rect 56474 11320 56516 11360
rect 56556 11320 56598 11360
rect 56638 11320 56680 11360
rect 56720 11320 56729 11360
rect 60343 11320 60352 11360
rect 60392 11320 60434 11360
rect 60474 11320 60516 11360
rect 60556 11320 60598 11360
rect 60638 11320 60680 11360
rect 60720 11320 60729 11360
rect 64343 11320 64352 11360
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64720 11320 64729 11360
rect 68343 11320 68352 11360
rect 68392 11320 68434 11360
rect 68474 11320 68516 11360
rect 68556 11320 68598 11360
rect 68638 11320 68680 11360
rect 68720 11320 68729 11360
rect 68515 10984 68524 11024
rect 68564 10984 69772 11024
rect 69812 10984 69821 11024
rect 1603 10900 1612 10940
rect 1652 10900 1804 10940
rect 1844 10900 2188 10940
rect 2228 10900 2237 10940
rect 835 10816 844 10856
rect 884 10816 1420 10856
rect 1460 10816 1469 10856
rect 643 10732 652 10772
rect 692 10732 701 10772
rect 0 10688 80 10708
rect 652 10688 692 10732
rect 0 10648 692 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 7103 10564 7112 10604
rect 7152 10564 7194 10604
rect 7234 10564 7276 10604
rect 7316 10564 7358 10604
rect 7398 10564 7440 10604
rect 7480 10564 7489 10604
rect 11103 10564 11112 10604
rect 11152 10564 11194 10604
rect 11234 10564 11276 10604
rect 11316 10564 11358 10604
rect 11398 10564 11440 10604
rect 11480 10564 11489 10604
rect 15103 10564 15112 10604
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15480 10564 15489 10604
rect 19103 10564 19112 10604
rect 19152 10564 19194 10604
rect 19234 10564 19276 10604
rect 19316 10564 19358 10604
rect 19398 10564 19440 10604
rect 19480 10564 19489 10604
rect 23103 10564 23112 10604
rect 23152 10564 23194 10604
rect 23234 10564 23276 10604
rect 23316 10564 23358 10604
rect 23398 10564 23440 10604
rect 23480 10564 23489 10604
rect 27103 10564 27112 10604
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27480 10564 27489 10604
rect 31103 10564 31112 10604
rect 31152 10564 31194 10604
rect 31234 10564 31276 10604
rect 31316 10564 31358 10604
rect 31398 10564 31440 10604
rect 31480 10564 31489 10604
rect 35103 10564 35112 10604
rect 35152 10564 35194 10604
rect 35234 10564 35276 10604
rect 35316 10564 35358 10604
rect 35398 10564 35440 10604
rect 35480 10564 35489 10604
rect 39103 10564 39112 10604
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39480 10564 39489 10604
rect 43103 10564 43112 10604
rect 43152 10564 43194 10604
rect 43234 10564 43276 10604
rect 43316 10564 43358 10604
rect 43398 10564 43440 10604
rect 43480 10564 43489 10604
rect 47103 10564 47112 10604
rect 47152 10564 47194 10604
rect 47234 10564 47276 10604
rect 47316 10564 47358 10604
rect 47398 10564 47440 10604
rect 47480 10564 47489 10604
rect 51103 10564 51112 10604
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51480 10564 51489 10604
rect 55103 10564 55112 10604
rect 55152 10564 55194 10604
rect 55234 10564 55276 10604
rect 55316 10564 55358 10604
rect 55398 10564 55440 10604
rect 55480 10564 55489 10604
rect 59103 10564 59112 10604
rect 59152 10564 59194 10604
rect 59234 10564 59276 10604
rect 59316 10564 59358 10604
rect 59398 10564 59440 10604
rect 59480 10564 59489 10604
rect 63103 10564 63112 10604
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63480 10564 63489 10604
rect 67103 10564 67112 10604
rect 67152 10564 67194 10604
rect 67234 10564 67276 10604
rect 67316 10564 67358 10604
rect 67398 10564 67440 10604
rect 67480 10564 67489 10604
rect 835 10312 844 10352
rect 884 10312 1324 10352
rect 1364 10312 1373 10352
rect 67459 10144 67468 10184
rect 67508 10144 68524 10184
rect 68564 10144 68573 10184
rect 69379 10144 69388 10184
rect 69428 10144 69676 10184
rect 69716 10144 69725 10184
rect 67651 10060 67660 10100
rect 67700 10060 70732 10100
rect 70772 10060 70781 10100
rect 68323 9976 68332 10016
rect 68372 9976 68716 10016
rect 68756 9976 69004 10016
rect 69044 9976 69388 10016
rect 69428 9976 69437 10016
rect 69763 9892 69772 9932
rect 69812 9892 73215 9932
rect 73255 9892 73264 9932
rect 73896 9892 73905 9932
rect 73945 9892 73954 9932
rect 0 9848 80 9868
rect 73900 9848 73940 9892
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 8343 9808 8352 9848
rect 8392 9808 8434 9848
rect 8474 9808 8516 9848
rect 8556 9808 8598 9848
rect 8638 9808 8680 9848
rect 8720 9808 8729 9848
rect 12343 9808 12352 9848
rect 12392 9808 12434 9848
rect 12474 9808 12516 9848
rect 12556 9808 12598 9848
rect 12638 9808 12680 9848
rect 12720 9808 12729 9848
rect 16343 9808 16352 9848
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16720 9808 16729 9848
rect 20343 9808 20352 9848
rect 20392 9808 20434 9848
rect 20474 9808 20516 9848
rect 20556 9808 20598 9848
rect 20638 9808 20680 9848
rect 20720 9808 20729 9848
rect 24343 9808 24352 9848
rect 24392 9808 24434 9848
rect 24474 9808 24516 9848
rect 24556 9808 24598 9848
rect 24638 9808 24680 9848
rect 24720 9808 24729 9848
rect 28343 9808 28352 9848
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28720 9808 28729 9848
rect 32343 9808 32352 9848
rect 32392 9808 32434 9848
rect 32474 9808 32516 9848
rect 32556 9808 32598 9848
rect 32638 9808 32680 9848
rect 32720 9808 32729 9848
rect 36343 9808 36352 9848
rect 36392 9808 36434 9848
rect 36474 9808 36516 9848
rect 36556 9808 36598 9848
rect 36638 9808 36680 9848
rect 36720 9808 36729 9848
rect 40343 9808 40352 9848
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40720 9808 40729 9848
rect 44343 9808 44352 9848
rect 44392 9808 44434 9848
rect 44474 9808 44516 9848
rect 44556 9808 44598 9848
rect 44638 9808 44680 9848
rect 44720 9808 44729 9848
rect 48343 9808 48352 9848
rect 48392 9808 48434 9848
rect 48474 9808 48516 9848
rect 48556 9808 48598 9848
rect 48638 9808 48680 9848
rect 48720 9808 48729 9848
rect 52343 9808 52352 9848
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52720 9808 52729 9848
rect 56343 9808 56352 9848
rect 56392 9808 56434 9848
rect 56474 9808 56516 9848
rect 56556 9808 56598 9848
rect 56638 9808 56680 9848
rect 56720 9808 56729 9848
rect 60343 9808 60352 9848
rect 60392 9808 60434 9848
rect 60474 9808 60516 9848
rect 60556 9808 60598 9848
rect 60638 9808 60680 9848
rect 60720 9808 60729 9848
rect 64343 9808 64352 9848
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64720 9808 64729 9848
rect 68343 9808 68352 9848
rect 68392 9808 68434 9848
rect 68474 9808 68516 9848
rect 68556 9808 68598 9848
rect 68638 9808 68680 9848
rect 68720 9808 68729 9848
rect 69571 9808 69580 9848
rect 69620 9808 72305 9848
rect 72345 9808 72354 9848
rect 73228 9808 73940 9848
rect 74947 9808 74956 9848
rect 74996 9808 75215 9848
rect 75255 9808 75264 9848
rect 79496 9808 79505 9848
rect 79545 9808 79756 9848
rect 79796 9808 79805 9848
rect 82296 9808 82305 9848
rect 82345 9808 82540 9848
rect 82580 9808 82589 9848
rect 91496 9808 91505 9848
rect 91545 9808 91756 9848
rect 91796 9808 91805 9848
rect 92995 9808 93004 9848
rect 93044 9808 93215 9848
rect 93255 9808 93264 9848
rect 0 9788 80 9808
rect 73228 9764 73268 9808
rect 80131 9764 80189 9765
rect 83587 9764 83645 9765
rect 89059 9764 89117 9765
rect 69859 9724 69868 9764
rect 69908 9724 72415 9764
rect 72455 9724 72464 9764
rect 73219 9724 73228 9764
rect 73268 9724 73277 9764
rect 74563 9724 74572 9764
rect 74612 9724 75505 9764
rect 75545 9724 75554 9764
rect 80131 9724 80140 9764
rect 80180 9724 80305 9764
rect 80345 9724 80354 9764
rect 83520 9724 83596 9764
rect 83655 9724 83664 9764
rect 87206 9724 87215 9764
rect 87255 9724 87724 9764
rect 87764 9724 87773 9764
rect 89010 9724 89068 9764
rect 89145 9724 89154 9764
rect 92696 9724 92705 9764
rect 92745 9724 92908 9764
rect 92948 9724 92957 9764
rect 95875 9724 95884 9764
rect 95924 9724 96305 9764
rect 96345 9724 96354 9764
rect 80131 9723 80189 9724
rect 83587 9723 83645 9724
rect 89059 9723 89117 9724
rect 70723 9640 70732 9680
rect 70772 9640 73324 9680
rect 73364 9640 73373 9680
rect 68227 9556 68236 9596
rect 68276 9556 72844 9596
rect 72884 9556 72893 9596
rect 98851 9512 98909 9513
rect 69187 9472 69196 9512
rect 69236 9472 73132 9512
rect 73172 9472 73181 9512
rect 97507 9472 97516 9512
rect 97556 9472 98860 9512
rect 98900 9472 98909 9512
rect 98851 9471 98909 9472
rect 69475 9388 69484 9428
rect 69524 9388 73612 9428
rect 73652 9388 73661 9428
rect 835 9304 844 9344
rect 884 9304 1324 9344
rect 1364 9304 1373 9344
rect 69187 9304 69196 9344
rect 69236 9304 72652 9344
rect 72692 9304 72701 9344
rect 69667 9220 69676 9260
rect 69716 9220 73228 9260
rect 73268 9220 73277 9260
rect 69955 9136 69964 9176
rect 70004 9136 74380 9176
rect 74420 9136 74429 9176
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 7103 9052 7112 9092
rect 7152 9052 7194 9092
rect 7234 9052 7276 9092
rect 7316 9052 7358 9092
rect 7398 9052 7440 9092
rect 7480 9052 7489 9092
rect 11103 9052 11112 9092
rect 11152 9052 11194 9092
rect 11234 9052 11276 9092
rect 11316 9052 11358 9092
rect 11398 9052 11440 9092
rect 11480 9052 11489 9092
rect 15103 9052 15112 9092
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15480 9052 15489 9092
rect 19103 9052 19112 9092
rect 19152 9052 19194 9092
rect 19234 9052 19276 9092
rect 19316 9052 19358 9092
rect 19398 9052 19440 9092
rect 19480 9052 19489 9092
rect 23103 9052 23112 9092
rect 23152 9052 23194 9092
rect 23234 9052 23276 9092
rect 23316 9052 23358 9092
rect 23398 9052 23440 9092
rect 23480 9052 23489 9092
rect 27103 9052 27112 9092
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27480 9052 27489 9092
rect 31103 9052 31112 9092
rect 31152 9052 31194 9092
rect 31234 9052 31276 9092
rect 31316 9052 31358 9092
rect 31398 9052 31440 9092
rect 31480 9052 31489 9092
rect 35103 9052 35112 9092
rect 35152 9052 35194 9092
rect 35234 9052 35276 9092
rect 35316 9052 35358 9092
rect 35398 9052 35440 9092
rect 35480 9052 35489 9092
rect 39103 9052 39112 9092
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39480 9052 39489 9092
rect 43103 9052 43112 9092
rect 43152 9052 43194 9092
rect 43234 9052 43276 9092
rect 43316 9052 43358 9092
rect 43398 9052 43440 9092
rect 43480 9052 43489 9092
rect 47103 9052 47112 9092
rect 47152 9052 47194 9092
rect 47234 9052 47276 9092
rect 47316 9052 47358 9092
rect 47398 9052 47440 9092
rect 47480 9052 47489 9092
rect 51103 9052 51112 9092
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51480 9052 51489 9092
rect 55103 9052 55112 9092
rect 55152 9052 55194 9092
rect 55234 9052 55276 9092
rect 55316 9052 55358 9092
rect 55398 9052 55440 9092
rect 55480 9052 55489 9092
rect 59103 9052 59112 9092
rect 59152 9052 59194 9092
rect 59234 9052 59276 9092
rect 59316 9052 59358 9092
rect 59398 9052 59440 9092
rect 59480 9052 59489 9092
rect 63103 9052 63112 9092
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63480 9052 63489 9092
rect 67103 9052 67112 9092
rect 67152 9052 67194 9092
rect 67234 9052 67276 9092
rect 67316 9052 67358 9092
rect 67398 9052 67440 9092
rect 67480 9052 67489 9092
rect 0 9008 80 9028
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 0 8948 80 8968
rect 85603 8840 85661 8841
rect 835 8800 844 8840
rect 884 8800 1420 8840
rect 1460 8800 1469 8840
rect 68995 8800 69004 8840
rect 69044 8800 73324 8840
rect 73364 8800 73373 8840
rect 85518 8800 85612 8840
rect 85652 8800 85661 8840
rect 85603 8799 85661 8800
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 8343 8296 8352 8336
rect 8392 8296 8434 8336
rect 8474 8296 8516 8336
rect 8556 8296 8598 8336
rect 8638 8296 8680 8336
rect 8720 8296 8729 8336
rect 12343 8296 12352 8336
rect 12392 8296 12434 8336
rect 12474 8296 12516 8336
rect 12556 8296 12598 8336
rect 12638 8296 12680 8336
rect 12720 8296 12729 8336
rect 16343 8296 16352 8336
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16720 8296 16729 8336
rect 20343 8296 20352 8336
rect 20392 8296 20434 8336
rect 20474 8296 20516 8336
rect 20556 8296 20598 8336
rect 20638 8296 20680 8336
rect 20720 8296 20729 8336
rect 24343 8296 24352 8336
rect 24392 8296 24434 8336
rect 24474 8296 24516 8336
rect 24556 8296 24598 8336
rect 24638 8296 24680 8336
rect 24720 8296 24729 8336
rect 28343 8296 28352 8336
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28720 8296 28729 8336
rect 32343 8296 32352 8336
rect 32392 8296 32434 8336
rect 32474 8296 32516 8336
rect 32556 8296 32598 8336
rect 32638 8296 32680 8336
rect 32720 8296 32729 8336
rect 36343 8296 36352 8336
rect 36392 8296 36434 8336
rect 36474 8296 36516 8336
rect 36556 8296 36598 8336
rect 36638 8296 36680 8336
rect 36720 8296 36729 8336
rect 40343 8296 40352 8336
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40720 8296 40729 8336
rect 44343 8296 44352 8336
rect 44392 8296 44434 8336
rect 44474 8296 44516 8336
rect 44556 8296 44598 8336
rect 44638 8296 44680 8336
rect 44720 8296 44729 8336
rect 48343 8296 48352 8336
rect 48392 8296 48434 8336
rect 48474 8296 48516 8336
rect 48556 8296 48598 8336
rect 48638 8296 48680 8336
rect 48720 8296 48729 8336
rect 52343 8296 52352 8336
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52720 8296 52729 8336
rect 56343 8296 56352 8336
rect 56392 8296 56434 8336
rect 56474 8296 56516 8336
rect 56556 8296 56598 8336
rect 56638 8296 56680 8336
rect 56720 8296 56729 8336
rect 60343 8296 60352 8336
rect 60392 8296 60434 8336
rect 60474 8296 60516 8336
rect 60556 8296 60598 8336
rect 60638 8296 60680 8336
rect 60720 8296 60729 8336
rect 64343 8296 64352 8336
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64720 8296 64729 8336
rect 68343 8296 68352 8336
rect 68392 8296 68434 8336
rect 68474 8296 68516 8336
rect 68556 8296 68598 8336
rect 68638 8296 68680 8336
rect 68720 8296 68729 8336
rect 81571 8212 81580 8252
rect 81620 8212 82252 8252
rect 82292 8212 82301 8252
rect 0 8168 80 8188
rect 0 8128 652 8168
rect 692 8128 701 8168
rect 69763 8128 69772 8168
rect 69812 8128 86188 8168
rect 86228 8128 86237 8168
rect 0 8108 80 8128
rect 82915 7916 82973 7917
rect 82915 7876 82924 7916
rect 82964 7876 83116 7916
rect 83156 7876 83165 7916
rect 82915 7875 82973 7876
rect 95587 7832 95645 7833
rect 835 7792 844 7832
rect 884 7792 1516 7832
rect 1556 7792 1565 7832
rect 95395 7792 95404 7832
rect 95444 7792 95596 7832
rect 95636 7792 95645 7832
rect 95587 7791 95645 7792
rect 74755 7708 74764 7748
rect 74804 7708 75052 7748
rect 75092 7708 75101 7748
rect 95203 7708 95212 7748
rect 95252 7708 96172 7748
rect 96212 7708 96221 7748
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 7103 7540 7112 7580
rect 7152 7540 7194 7580
rect 7234 7540 7276 7580
rect 7316 7540 7358 7580
rect 7398 7540 7440 7580
rect 7480 7540 7489 7580
rect 11103 7540 11112 7580
rect 11152 7540 11194 7580
rect 11234 7540 11276 7580
rect 11316 7540 11358 7580
rect 11398 7540 11440 7580
rect 11480 7540 11489 7580
rect 15103 7540 15112 7580
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15480 7540 15489 7580
rect 19103 7540 19112 7580
rect 19152 7540 19194 7580
rect 19234 7540 19276 7580
rect 19316 7540 19358 7580
rect 19398 7540 19440 7580
rect 19480 7540 19489 7580
rect 23103 7540 23112 7580
rect 23152 7540 23194 7580
rect 23234 7540 23276 7580
rect 23316 7540 23358 7580
rect 23398 7540 23440 7580
rect 23480 7540 23489 7580
rect 27103 7540 27112 7580
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27480 7540 27489 7580
rect 31103 7540 31112 7580
rect 31152 7540 31194 7580
rect 31234 7540 31276 7580
rect 31316 7540 31358 7580
rect 31398 7540 31440 7580
rect 31480 7540 31489 7580
rect 35103 7540 35112 7580
rect 35152 7540 35194 7580
rect 35234 7540 35276 7580
rect 35316 7540 35358 7580
rect 35398 7540 35440 7580
rect 35480 7540 35489 7580
rect 39103 7540 39112 7580
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39480 7540 39489 7580
rect 43103 7540 43112 7580
rect 43152 7540 43194 7580
rect 43234 7540 43276 7580
rect 43316 7540 43358 7580
rect 43398 7540 43440 7580
rect 43480 7540 43489 7580
rect 47103 7540 47112 7580
rect 47152 7540 47194 7580
rect 47234 7540 47276 7580
rect 47316 7540 47358 7580
rect 47398 7540 47440 7580
rect 47480 7540 47489 7580
rect 51103 7540 51112 7580
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51480 7540 51489 7580
rect 55103 7540 55112 7580
rect 55152 7540 55194 7580
rect 55234 7540 55276 7580
rect 55316 7540 55358 7580
rect 55398 7540 55440 7580
rect 55480 7540 55489 7580
rect 59103 7540 59112 7580
rect 59152 7540 59194 7580
rect 59234 7540 59276 7580
rect 59316 7540 59358 7580
rect 59398 7540 59440 7580
rect 59480 7540 59489 7580
rect 63103 7540 63112 7580
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63480 7540 63489 7580
rect 67103 7540 67112 7580
rect 67152 7540 67194 7580
rect 67234 7540 67276 7580
rect 67316 7540 67358 7580
rect 67398 7540 67440 7580
rect 67480 7540 67489 7580
rect 71103 7540 71112 7580
rect 71152 7540 71194 7580
rect 71234 7540 71276 7580
rect 71316 7540 71358 7580
rect 71398 7540 71440 7580
rect 71480 7540 71489 7580
rect 74179 7540 74188 7580
rect 74228 7540 74860 7580
rect 74900 7540 74909 7580
rect 75103 7540 75112 7580
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75480 7540 75489 7580
rect 78019 7540 78028 7580
rect 78068 7540 78316 7580
rect 78356 7540 78365 7580
rect 79103 7540 79112 7580
rect 79152 7540 79194 7580
rect 79234 7540 79276 7580
rect 79316 7540 79358 7580
rect 79398 7540 79440 7580
rect 79480 7540 79489 7580
rect 81667 7540 81676 7580
rect 81716 7540 81964 7580
rect 82004 7540 82013 7580
rect 83103 7540 83112 7580
rect 83152 7540 83194 7580
rect 83234 7540 83276 7580
rect 83316 7540 83358 7580
rect 83398 7540 83440 7580
rect 83480 7540 83489 7580
rect 84451 7540 84460 7580
rect 84500 7540 85708 7580
rect 85748 7540 85757 7580
rect 86467 7540 86476 7580
rect 86516 7540 86996 7580
rect 87103 7540 87112 7580
rect 87152 7540 87194 7580
rect 87234 7540 87276 7580
rect 87316 7540 87358 7580
rect 87398 7540 87440 7580
rect 87480 7540 87489 7580
rect 88003 7540 88012 7580
rect 88052 7540 88972 7580
rect 89012 7540 89021 7580
rect 91103 7540 91112 7580
rect 91152 7540 91194 7580
rect 91234 7540 91276 7580
rect 91316 7540 91358 7580
rect 91398 7540 91440 7580
rect 91480 7540 91489 7580
rect 92419 7540 92428 7580
rect 92468 7540 93292 7580
rect 93332 7540 93341 7580
rect 95103 7540 95112 7580
rect 95152 7540 95194 7580
rect 95234 7540 95276 7580
rect 95316 7540 95358 7580
rect 95398 7540 95440 7580
rect 95480 7540 95489 7580
rect 96835 7540 96844 7580
rect 96884 7540 97132 7580
rect 97172 7540 97181 7580
rect 99103 7540 99112 7580
rect 99152 7540 99194 7580
rect 99234 7540 99276 7580
rect 99316 7540 99358 7580
rect 99398 7540 99440 7580
rect 99480 7540 99489 7580
rect 74659 7456 74668 7496
rect 74708 7456 74717 7496
rect 74668 7412 74708 7456
rect 76771 7412 76829 7413
rect 86659 7412 86717 7413
rect 74668 7372 75244 7412
rect 75284 7372 75293 7412
rect 76579 7372 76588 7412
rect 76628 7372 76780 7412
rect 76820 7372 76829 7412
rect 77059 7372 77068 7412
rect 77108 7372 77452 7412
rect 77492 7372 77501 7412
rect 77635 7372 77644 7412
rect 77684 7372 78028 7412
rect 78068 7372 78077 7412
rect 80899 7372 80908 7412
rect 80948 7372 81676 7412
rect 81716 7372 81725 7412
rect 83875 7372 83884 7412
rect 83924 7372 84076 7412
rect 84116 7372 84125 7412
rect 84643 7372 84652 7412
rect 84692 7372 84844 7412
rect 84884 7372 84893 7412
rect 86574 7372 86668 7412
rect 86708 7372 86717 7412
rect 86956 7412 86996 7540
rect 86956 7372 87148 7412
rect 87188 7372 87197 7412
rect 89635 7372 89644 7412
rect 89684 7372 89836 7412
rect 89876 7372 89885 7412
rect 90019 7372 90028 7412
rect 90068 7372 90604 7412
rect 90644 7372 90653 7412
rect 90883 7372 90892 7412
rect 90932 7372 91852 7412
rect 91892 7372 91901 7412
rect 93475 7372 93484 7412
rect 93524 7372 93676 7412
rect 93716 7372 93725 7412
rect 96451 7372 96460 7412
rect 96500 7372 96844 7412
rect 96884 7372 96893 7412
rect 76771 7371 76829 7372
rect 86659 7371 86717 7372
rect 0 7328 80 7348
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 74275 7288 74284 7328
rect 74324 7288 74476 7328
rect 74516 7288 75148 7328
rect 75188 7288 75197 7328
rect 76588 7288 77260 7328
rect 77300 7288 77309 7328
rect 79651 7288 79660 7328
rect 79700 7288 80044 7328
rect 80084 7288 80093 7328
rect 86275 7288 86284 7328
rect 86324 7288 87244 7328
rect 87284 7288 87293 7328
rect 91171 7288 91180 7328
rect 91220 7288 91756 7328
rect 91796 7288 91805 7328
rect 92323 7288 92332 7328
rect 92372 7288 93100 7328
rect 93140 7288 93388 7328
rect 93428 7288 93437 7328
rect 93955 7288 93964 7328
rect 94004 7288 94924 7328
rect 94964 7288 95308 7328
rect 95348 7288 95357 7328
rect 0 7268 80 7288
rect 71779 7204 71788 7244
rect 71828 7204 74668 7244
rect 74708 7204 74717 7244
rect 75427 7204 75436 7244
rect 75476 7204 75724 7244
rect 75764 7204 75773 7244
rect 76588 7076 76628 7288
rect 76867 7204 76876 7244
rect 76916 7204 77644 7244
rect 77684 7204 77693 7244
rect 77827 7204 77836 7244
rect 77876 7204 79084 7244
rect 79124 7204 80236 7244
rect 80276 7204 80285 7244
rect 80707 7204 80716 7244
rect 80756 7204 81100 7244
rect 81140 7204 82252 7244
rect 82292 7204 82828 7244
rect 82868 7204 84268 7244
rect 84308 7204 85228 7244
rect 85268 7204 85277 7244
rect 86083 7204 86092 7244
rect 86132 7204 86476 7244
rect 86516 7204 88012 7244
rect 88052 7204 88061 7244
rect 88291 7204 88300 7244
rect 88340 7204 88588 7244
rect 88628 7204 89068 7244
rect 89108 7204 89117 7244
rect 90979 7204 90988 7244
rect 91028 7204 91564 7244
rect 91604 7204 91613 7244
rect 92131 7204 92140 7244
rect 92180 7204 92524 7244
rect 92564 7204 94156 7244
rect 94196 7204 94292 7244
rect 95683 7204 95692 7244
rect 95732 7204 96076 7244
rect 96116 7204 96125 7244
rect 96259 7204 96268 7244
rect 96308 7204 96652 7244
rect 96692 7204 97612 7244
rect 97652 7204 97804 7244
rect 97844 7204 98188 7244
rect 98228 7204 98237 7244
rect 77836 7160 77876 7204
rect 94252 7160 94292 7204
rect 76675 7120 76684 7160
rect 76724 7120 77260 7160
rect 77300 7120 77876 7160
rect 80899 7120 80908 7160
rect 80948 7120 81292 7160
rect 81332 7120 81920 7160
rect 82627 7120 82636 7160
rect 82676 7120 83116 7160
rect 83156 7120 83308 7160
rect 83348 7120 83357 7160
rect 83779 7120 83788 7160
rect 83828 7120 84076 7160
rect 84116 7120 84844 7160
rect 84884 7120 85612 7160
rect 85652 7120 85661 7160
rect 86947 7120 86956 7160
rect 86996 7120 87436 7160
rect 87476 7120 87485 7160
rect 89443 7120 89452 7160
rect 89492 7120 89836 7160
rect 89876 7120 90713 7160
rect 90753 7120 90892 7160
rect 90932 7120 91756 7160
rect 91796 7120 91805 7160
rect 93763 7120 93772 7160
rect 93812 7120 94196 7160
rect 94252 7120 94732 7160
rect 94772 7120 96500 7160
rect 96931 7120 96940 7160
rect 96980 7120 97228 7160
rect 97268 7120 97277 7160
rect 81880 7076 81920 7120
rect 82915 7076 82973 7077
rect 94156 7076 94196 7120
rect 96460 7076 96500 7120
rect 74083 7036 74092 7076
rect 74132 7036 75052 7076
rect 75092 7036 75764 7076
rect 76579 7036 76588 7076
rect 76628 7036 76637 7076
rect 77635 7036 77644 7076
rect 77684 7036 78412 7076
rect 78452 7036 78700 7076
rect 78740 7036 78749 7076
rect 81880 7036 81961 7076
rect 82001 7036 82010 7076
rect 82830 7036 82924 7076
rect 82964 7036 82973 7076
rect 87235 7036 87244 7076
rect 87284 7036 87532 7076
rect 87572 7036 87820 7076
rect 87860 7036 87869 7076
rect 88003 7036 88012 7076
rect 88052 7036 90028 7076
rect 90068 7036 91372 7076
rect 91412 7036 91421 7076
rect 92707 7036 92716 7076
rect 92756 7036 93676 7076
rect 93716 7036 93725 7076
rect 94147 7036 94156 7076
rect 94196 7036 94205 7076
rect 96451 7036 96460 7076
rect 96500 7036 96509 7076
rect 75724 6992 75764 7036
rect 82915 7035 82973 7036
rect 88195 6992 88253 6993
rect 74380 6952 74860 6992
rect 74900 6952 75436 6992
rect 75476 6952 75485 6992
rect 75715 6952 75724 6992
rect 75764 6952 77452 6992
rect 77492 6952 78124 6992
rect 78164 6952 79372 6992
rect 79412 6952 79421 6992
rect 80515 6952 80524 6992
rect 80564 6952 81772 6992
rect 81812 6952 84556 6992
rect 84596 6952 84605 6992
rect 85987 6952 85996 6992
rect 86036 6952 86956 6992
rect 86996 6952 87005 6992
rect 88195 6952 88204 6992
rect 88244 6952 88396 6992
rect 88436 6952 88445 6992
rect 93763 6952 93772 6992
rect 93812 6952 94444 6992
rect 94484 6952 94493 6992
rect 74380 6824 74420 6952
rect 80524 6908 80564 6952
rect 88195 6951 88253 6952
rect 75139 6868 75148 6908
rect 75188 6868 80564 6908
rect 86659 6868 86668 6908
rect 86708 6868 90316 6908
rect 90356 6868 94348 6908
rect 94388 6868 94397 6908
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 8343 6784 8352 6824
rect 8392 6784 8434 6824
rect 8474 6784 8516 6824
rect 8556 6784 8598 6824
rect 8638 6784 8680 6824
rect 8720 6784 8729 6824
rect 12343 6784 12352 6824
rect 12392 6784 12434 6824
rect 12474 6784 12516 6824
rect 12556 6784 12598 6824
rect 12638 6784 12680 6824
rect 12720 6784 12729 6824
rect 16343 6784 16352 6824
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16720 6784 16729 6824
rect 20343 6784 20352 6824
rect 20392 6784 20434 6824
rect 20474 6784 20516 6824
rect 20556 6784 20598 6824
rect 20638 6784 20680 6824
rect 20720 6784 20729 6824
rect 24343 6784 24352 6824
rect 24392 6784 24434 6824
rect 24474 6784 24516 6824
rect 24556 6784 24598 6824
rect 24638 6784 24680 6824
rect 24720 6784 24729 6824
rect 28343 6784 28352 6824
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28720 6784 28729 6824
rect 32343 6784 32352 6824
rect 32392 6784 32434 6824
rect 32474 6784 32516 6824
rect 32556 6784 32598 6824
rect 32638 6784 32680 6824
rect 32720 6784 32729 6824
rect 36343 6784 36352 6824
rect 36392 6784 36434 6824
rect 36474 6784 36516 6824
rect 36556 6784 36598 6824
rect 36638 6784 36680 6824
rect 36720 6784 36729 6824
rect 40343 6784 40352 6824
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40720 6784 40729 6824
rect 44343 6784 44352 6824
rect 44392 6784 44434 6824
rect 44474 6784 44516 6824
rect 44556 6784 44598 6824
rect 44638 6784 44680 6824
rect 44720 6784 44729 6824
rect 48343 6784 48352 6824
rect 48392 6784 48434 6824
rect 48474 6784 48516 6824
rect 48556 6784 48598 6824
rect 48638 6784 48680 6824
rect 48720 6784 48729 6824
rect 52343 6784 52352 6824
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52720 6784 52729 6824
rect 56343 6784 56352 6824
rect 56392 6784 56434 6824
rect 56474 6784 56516 6824
rect 56556 6784 56598 6824
rect 56638 6784 56680 6824
rect 56720 6784 56729 6824
rect 60343 6784 60352 6824
rect 60392 6784 60434 6824
rect 60474 6784 60516 6824
rect 60556 6784 60598 6824
rect 60638 6784 60680 6824
rect 60720 6784 60729 6824
rect 64343 6784 64352 6824
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64720 6784 64729 6824
rect 68343 6784 68352 6824
rect 68392 6784 68434 6824
rect 68474 6784 68516 6824
rect 68556 6784 68598 6824
rect 68638 6784 68680 6824
rect 68720 6784 68729 6824
rect 72343 6784 72352 6824
rect 72392 6784 72434 6824
rect 72474 6784 72516 6824
rect 72556 6784 72598 6824
rect 72638 6784 72680 6824
rect 72720 6784 72729 6824
rect 74371 6784 74380 6824
rect 74420 6784 74429 6824
rect 76343 6784 76352 6824
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76720 6784 76729 6824
rect 80343 6784 80352 6824
rect 80392 6784 80434 6824
rect 80474 6784 80516 6824
rect 80556 6784 80598 6824
rect 80638 6784 80680 6824
rect 80720 6784 80729 6824
rect 84343 6784 84352 6824
rect 84392 6784 84434 6824
rect 84474 6784 84516 6824
rect 84556 6784 84598 6824
rect 84638 6784 84680 6824
rect 84720 6784 84729 6824
rect 88343 6784 88352 6824
rect 88392 6784 88434 6824
rect 88474 6784 88516 6824
rect 88556 6784 88598 6824
rect 88638 6784 88680 6824
rect 88720 6784 88729 6824
rect 92343 6784 92352 6824
rect 92392 6784 92434 6824
rect 92474 6784 92516 6824
rect 92556 6784 92598 6824
rect 92638 6784 92680 6824
rect 92720 6784 92729 6824
rect 96343 6784 96352 6824
rect 96392 6784 96434 6824
rect 96474 6784 96516 6824
rect 96556 6784 96598 6824
rect 96638 6784 96680 6824
rect 96720 6784 96729 6824
rect 95587 6740 95645 6741
rect 95299 6700 95308 6740
rect 95348 6700 95596 6740
rect 95636 6700 95645 6740
rect 95587 6699 95645 6700
rect 88195 6656 88253 6657
rect 835 6616 844 6656
rect 884 6616 1324 6656
rect 1364 6616 1373 6656
rect 75148 6616 75340 6656
rect 75380 6616 76588 6656
rect 76628 6616 76637 6656
rect 88195 6616 88204 6656
rect 88244 6616 88492 6656
rect 88532 6616 88541 6656
rect 93667 6616 93676 6656
rect 93716 6616 94540 6656
rect 94580 6616 95692 6656
rect 95732 6616 97996 6656
rect 98036 6616 98045 6656
rect 0 6488 80 6508
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 0 6428 80 6448
rect 75148 6404 75188 6616
rect 88195 6615 88253 6616
rect 86083 6532 86092 6572
rect 86132 6532 86860 6572
rect 86900 6532 86909 6572
rect 96067 6532 96076 6572
rect 96116 6532 96125 6572
rect 75427 6448 75436 6488
rect 75476 6448 76108 6488
rect 76148 6448 76300 6488
rect 76340 6448 76349 6488
rect 88099 6448 88108 6488
rect 88148 6448 88588 6488
rect 88628 6448 88876 6488
rect 88916 6448 88925 6488
rect 95116 6448 95884 6488
rect 95924 6448 95933 6488
rect 95116 6404 95156 6448
rect 74563 6364 74572 6404
rect 74612 6364 74764 6404
rect 74804 6364 75148 6404
rect 75188 6364 75197 6404
rect 77731 6364 77740 6404
rect 77780 6364 78124 6404
rect 78164 6364 78604 6404
rect 78644 6364 78892 6404
rect 78932 6364 78941 6404
rect 82051 6364 82060 6404
rect 82100 6364 82540 6404
rect 82580 6364 82732 6404
rect 82772 6364 82781 6404
rect 83203 6364 83212 6404
rect 83252 6364 83692 6404
rect 83732 6364 84172 6404
rect 84212 6364 84556 6404
rect 84596 6364 84605 6404
rect 85027 6364 85036 6404
rect 85076 6364 85228 6404
rect 85268 6364 85612 6404
rect 85652 6364 86092 6404
rect 86132 6364 86141 6404
rect 89635 6364 89644 6404
rect 89684 6364 90412 6404
rect 90452 6364 90892 6404
rect 90932 6364 90941 6404
rect 91363 6364 91372 6404
rect 91412 6364 91660 6404
rect 91700 6364 92140 6404
rect 92180 6364 92524 6404
rect 92564 6364 92573 6404
rect 94051 6364 94060 6404
rect 94100 6364 94444 6404
rect 94484 6364 94924 6404
rect 94964 6364 95116 6404
rect 95156 6364 95165 6404
rect 96076 6320 96116 6532
rect 92995 6280 93004 6320
rect 93044 6280 93388 6320
rect 93428 6280 93868 6320
rect 93908 6280 93917 6320
rect 95875 6280 95884 6320
rect 95924 6280 96364 6320
rect 96404 6280 96940 6320
rect 96980 6280 97324 6320
rect 97364 6280 97373 6320
rect 95971 6196 95980 6236
rect 96020 6196 96172 6236
rect 96212 6196 96221 6236
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 7103 6028 7112 6068
rect 7152 6028 7194 6068
rect 7234 6028 7276 6068
rect 7316 6028 7358 6068
rect 7398 6028 7440 6068
rect 7480 6028 7489 6068
rect 11103 6028 11112 6068
rect 11152 6028 11194 6068
rect 11234 6028 11276 6068
rect 11316 6028 11358 6068
rect 11398 6028 11440 6068
rect 11480 6028 11489 6068
rect 15103 6028 15112 6068
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15480 6028 15489 6068
rect 19103 6028 19112 6068
rect 19152 6028 19194 6068
rect 19234 6028 19276 6068
rect 19316 6028 19358 6068
rect 19398 6028 19440 6068
rect 19480 6028 19489 6068
rect 23103 6028 23112 6068
rect 23152 6028 23194 6068
rect 23234 6028 23276 6068
rect 23316 6028 23358 6068
rect 23398 6028 23440 6068
rect 23480 6028 23489 6068
rect 27103 6028 27112 6068
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27480 6028 27489 6068
rect 31103 6028 31112 6068
rect 31152 6028 31194 6068
rect 31234 6028 31276 6068
rect 31316 6028 31358 6068
rect 31398 6028 31440 6068
rect 31480 6028 31489 6068
rect 35103 6028 35112 6068
rect 35152 6028 35194 6068
rect 35234 6028 35276 6068
rect 35316 6028 35358 6068
rect 35398 6028 35440 6068
rect 35480 6028 35489 6068
rect 39103 6028 39112 6068
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39480 6028 39489 6068
rect 43103 6028 43112 6068
rect 43152 6028 43194 6068
rect 43234 6028 43276 6068
rect 43316 6028 43358 6068
rect 43398 6028 43440 6068
rect 43480 6028 43489 6068
rect 47103 6028 47112 6068
rect 47152 6028 47194 6068
rect 47234 6028 47276 6068
rect 47316 6028 47358 6068
rect 47398 6028 47440 6068
rect 47480 6028 47489 6068
rect 51103 6028 51112 6068
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51480 6028 51489 6068
rect 55103 6028 55112 6068
rect 55152 6028 55194 6068
rect 55234 6028 55276 6068
rect 55316 6028 55358 6068
rect 55398 6028 55440 6068
rect 55480 6028 55489 6068
rect 59103 6028 59112 6068
rect 59152 6028 59194 6068
rect 59234 6028 59276 6068
rect 59316 6028 59358 6068
rect 59398 6028 59440 6068
rect 59480 6028 59489 6068
rect 63103 6028 63112 6068
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63480 6028 63489 6068
rect 67103 6028 67112 6068
rect 67152 6028 67194 6068
rect 67234 6028 67276 6068
rect 67316 6028 67358 6068
rect 67398 6028 67440 6068
rect 67480 6028 67489 6068
rect 71103 6028 71112 6068
rect 71152 6028 71194 6068
rect 71234 6028 71276 6068
rect 71316 6028 71358 6068
rect 71398 6028 71440 6068
rect 71480 6028 71489 6068
rect 75103 6028 75112 6068
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75480 6028 75489 6068
rect 79103 6028 79112 6068
rect 79152 6028 79194 6068
rect 79234 6028 79276 6068
rect 79316 6028 79358 6068
rect 79398 6028 79440 6068
rect 79480 6028 79489 6068
rect 83103 6028 83112 6068
rect 83152 6028 83194 6068
rect 83234 6028 83276 6068
rect 83316 6028 83358 6068
rect 83398 6028 83440 6068
rect 83480 6028 83489 6068
rect 87103 6028 87112 6068
rect 87152 6028 87194 6068
rect 87234 6028 87276 6068
rect 87316 6028 87358 6068
rect 87398 6028 87440 6068
rect 87480 6028 87489 6068
rect 91103 6028 91112 6068
rect 91152 6028 91194 6068
rect 91234 6028 91276 6068
rect 91316 6028 91358 6068
rect 91398 6028 91440 6068
rect 91480 6028 91489 6068
rect 95103 6028 95112 6068
rect 95152 6028 95194 6068
rect 95234 6028 95276 6068
rect 95316 6028 95358 6068
rect 95398 6028 95440 6068
rect 95480 6028 95489 6068
rect 99103 6028 99112 6068
rect 99152 6028 99194 6068
rect 99234 6028 99276 6068
rect 99316 6028 99358 6068
rect 99398 6028 99440 6068
rect 99480 6028 99489 6068
rect 76771 5900 76829 5901
rect 80131 5900 80189 5901
rect 83587 5900 83645 5901
rect 85603 5900 85661 5901
rect 89059 5900 89117 5901
rect 76675 5860 76684 5900
rect 76724 5860 76780 5900
rect 76820 5860 76829 5900
rect 80046 5860 80140 5900
rect 80180 5860 80189 5900
rect 83502 5860 83596 5900
rect 83636 5860 83645 5900
rect 85507 5860 85516 5900
rect 85556 5860 85612 5900
rect 85652 5860 85661 5900
rect 88974 5860 89068 5900
rect 89108 5860 89117 5900
rect 76771 5859 76829 5860
rect 80131 5859 80189 5860
rect 83587 5859 83645 5860
rect 85603 5859 85661 5860
rect 89059 5859 89117 5860
rect 835 5776 844 5816
rect 884 5776 1804 5816
rect 1844 5776 1853 5816
rect 86179 5776 86188 5816
rect 86228 5776 96940 5816
rect 96980 5776 98380 5816
rect 98420 5776 98668 5816
rect 98708 5776 98717 5816
rect 0 5648 80 5668
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 93283 5608 93292 5648
rect 93332 5608 93676 5648
rect 93716 5608 93725 5648
rect 0 5588 80 5608
rect 835 5440 844 5480
rect 884 5440 1420 5480
rect 1460 5440 1469 5480
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 8343 5272 8352 5312
rect 8392 5272 8434 5312
rect 8474 5272 8516 5312
rect 8556 5272 8598 5312
rect 8638 5272 8680 5312
rect 8720 5272 8729 5312
rect 12343 5272 12352 5312
rect 12392 5272 12434 5312
rect 12474 5272 12516 5312
rect 12556 5272 12598 5312
rect 12638 5272 12680 5312
rect 12720 5272 12729 5312
rect 16343 5272 16352 5312
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16720 5272 16729 5312
rect 20343 5272 20352 5312
rect 20392 5272 20434 5312
rect 20474 5272 20516 5312
rect 20556 5272 20598 5312
rect 20638 5272 20680 5312
rect 20720 5272 20729 5312
rect 24343 5272 24352 5312
rect 24392 5272 24434 5312
rect 24474 5272 24516 5312
rect 24556 5272 24598 5312
rect 24638 5272 24680 5312
rect 24720 5272 24729 5312
rect 28343 5272 28352 5312
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28720 5272 28729 5312
rect 32343 5272 32352 5312
rect 32392 5272 32434 5312
rect 32474 5272 32516 5312
rect 32556 5272 32598 5312
rect 32638 5272 32680 5312
rect 32720 5272 32729 5312
rect 36343 5272 36352 5312
rect 36392 5272 36434 5312
rect 36474 5272 36516 5312
rect 36556 5272 36598 5312
rect 36638 5272 36680 5312
rect 36720 5272 36729 5312
rect 40343 5272 40352 5312
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40720 5272 40729 5312
rect 44343 5272 44352 5312
rect 44392 5272 44434 5312
rect 44474 5272 44516 5312
rect 44556 5272 44598 5312
rect 44638 5272 44680 5312
rect 44720 5272 44729 5312
rect 48343 5272 48352 5312
rect 48392 5272 48434 5312
rect 48474 5272 48516 5312
rect 48556 5272 48598 5312
rect 48638 5272 48680 5312
rect 48720 5272 48729 5312
rect 52343 5272 52352 5312
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52720 5272 52729 5312
rect 56343 5272 56352 5312
rect 56392 5272 56434 5312
rect 56474 5272 56516 5312
rect 56556 5272 56598 5312
rect 56638 5272 56680 5312
rect 56720 5272 56729 5312
rect 60343 5272 60352 5312
rect 60392 5272 60434 5312
rect 60474 5272 60516 5312
rect 60556 5272 60598 5312
rect 60638 5272 60680 5312
rect 60720 5272 60729 5312
rect 64343 5272 64352 5312
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64720 5272 64729 5312
rect 68343 5272 68352 5312
rect 68392 5272 68434 5312
rect 68474 5272 68516 5312
rect 68556 5272 68598 5312
rect 68638 5272 68680 5312
rect 68720 5272 68729 5312
rect 72343 5272 72352 5312
rect 72392 5272 72434 5312
rect 72474 5272 72516 5312
rect 72556 5272 72598 5312
rect 72638 5272 72680 5312
rect 72720 5272 72729 5312
rect 76343 5272 76352 5312
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76720 5272 76729 5312
rect 80343 5272 80352 5312
rect 80392 5272 80434 5312
rect 80474 5272 80516 5312
rect 80556 5272 80598 5312
rect 80638 5272 80680 5312
rect 80720 5272 80729 5312
rect 84343 5272 84352 5312
rect 84392 5272 84434 5312
rect 84474 5272 84516 5312
rect 84556 5272 84598 5312
rect 84638 5272 84680 5312
rect 84720 5272 84729 5312
rect 88343 5272 88352 5312
rect 88392 5272 88434 5312
rect 88474 5272 88516 5312
rect 88556 5272 88598 5312
rect 88638 5272 88680 5312
rect 88720 5272 88729 5312
rect 92343 5272 92352 5312
rect 92392 5272 92434 5312
rect 92474 5272 92516 5312
rect 92556 5272 92598 5312
rect 92638 5272 92680 5312
rect 92720 5272 92729 5312
rect 96343 5272 96352 5312
rect 96392 5272 96434 5312
rect 96474 5272 96516 5312
rect 96556 5272 96598 5312
rect 96638 5272 96680 5312
rect 96720 5272 96729 5312
rect 0 4808 80 4828
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 0 4748 80 4768
rect 739 4684 748 4724
rect 788 4684 1996 4724
rect 2036 4684 2045 4724
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 7103 4516 7112 4556
rect 7152 4516 7194 4556
rect 7234 4516 7276 4556
rect 7316 4516 7358 4556
rect 7398 4516 7440 4556
rect 7480 4516 7489 4556
rect 11103 4516 11112 4556
rect 11152 4516 11194 4556
rect 11234 4516 11276 4556
rect 11316 4516 11358 4556
rect 11398 4516 11440 4556
rect 11480 4516 11489 4556
rect 15103 4516 15112 4556
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15480 4516 15489 4556
rect 19103 4516 19112 4556
rect 19152 4516 19194 4556
rect 19234 4516 19276 4556
rect 19316 4516 19358 4556
rect 19398 4516 19440 4556
rect 19480 4516 19489 4556
rect 23103 4516 23112 4556
rect 23152 4516 23194 4556
rect 23234 4516 23276 4556
rect 23316 4516 23358 4556
rect 23398 4516 23440 4556
rect 23480 4516 23489 4556
rect 27103 4516 27112 4556
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27480 4516 27489 4556
rect 31103 4516 31112 4556
rect 31152 4516 31194 4556
rect 31234 4516 31276 4556
rect 31316 4516 31358 4556
rect 31398 4516 31440 4556
rect 31480 4516 31489 4556
rect 35103 4516 35112 4556
rect 35152 4516 35194 4556
rect 35234 4516 35276 4556
rect 35316 4516 35358 4556
rect 35398 4516 35440 4556
rect 35480 4516 35489 4556
rect 39103 4516 39112 4556
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39480 4516 39489 4556
rect 43103 4516 43112 4556
rect 43152 4516 43194 4556
rect 43234 4516 43276 4556
rect 43316 4516 43358 4556
rect 43398 4516 43440 4556
rect 43480 4516 43489 4556
rect 47103 4516 47112 4556
rect 47152 4516 47194 4556
rect 47234 4516 47276 4556
rect 47316 4516 47358 4556
rect 47398 4516 47440 4556
rect 47480 4516 47489 4556
rect 51103 4516 51112 4556
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51480 4516 51489 4556
rect 55103 4516 55112 4556
rect 55152 4516 55194 4556
rect 55234 4516 55276 4556
rect 55316 4516 55358 4556
rect 55398 4516 55440 4556
rect 55480 4516 55489 4556
rect 59103 4516 59112 4556
rect 59152 4516 59194 4556
rect 59234 4516 59276 4556
rect 59316 4516 59358 4556
rect 59398 4516 59440 4556
rect 59480 4516 59489 4556
rect 63103 4516 63112 4556
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63480 4516 63489 4556
rect 67103 4516 67112 4556
rect 67152 4516 67194 4556
rect 67234 4516 67276 4556
rect 67316 4516 67358 4556
rect 67398 4516 67440 4556
rect 67480 4516 67489 4556
rect 71103 4516 71112 4556
rect 71152 4516 71194 4556
rect 71234 4516 71276 4556
rect 71316 4516 71358 4556
rect 71398 4516 71440 4556
rect 71480 4516 71489 4556
rect 75103 4516 75112 4556
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75480 4516 75489 4556
rect 79103 4516 79112 4556
rect 79152 4516 79194 4556
rect 79234 4516 79276 4556
rect 79316 4516 79358 4556
rect 79398 4516 79440 4556
rect 79480 4516 79489 4556
rect 83103 4516 83112 4556
rect 83152 4516 83194 4556
rect 83234 4516 83276 4556
rect 83316 4516 83358 4556
rect 83398 4516 83440 4556
rect 83480 4516 83489 4556
rect 87103 4516 87112 4556
rect 87152 4516 87194 4556
rect 87234 4516 87276 4556
rect 87316 4516 87358 4556
rect 87398 4516 87440 4556
rect 87480 4516 87489 4556
rect 91103 4516 91112 4556
rect 91152 4516 91194 4556
rect 91234 4516 91276 4556
rect 91316 4516 91358 4556
rect 91398 4516 91440 4556
rect 91480 4516 91489 4556
rect 95103 4516 95112 4556
rect 95152 4516 95194 4556
rect 95234 4516 95276 4556
rect 95316 4516 95358 4556
rect 95398 4516 95440 4556
rect 95480 4516 95489 4556
rect 99103 4516 99112 4556
rect 99152 4516 99194 4556
rect 99234 4516 99276 4556
rect 99316 4516 99358 4556
rect 99398 4516 99440 4556
rect 99480 4516 99489 4556
rect 835 4180 844 4220
rect 884 4180 1612 4220
rect 1652 4180 1661 4220
rect 0 3968 80 3988
rect 0 3928 652 3968
rect 692 3928 701 3968
rect 0 3908 80 3928
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 8343 3760 8352 3800
rect 8392 3760 8434 3800
rect 8474 3760 8516 3800
rect 8556 3760 8598 3800
rect 8638 3760 8680 3800
rect 8720 3760 8729 3800
rect 12343 3760 12352 3800
rect 12392 3760 12434 3800
rect 12474 3760 12516 3800
rect 12556 3760 12598 3800
rect 12638 3760 12680 3800
rect 12720 3760 12729 3800
rect 16343 3760 16352 3800
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16720 3760 16729 3800
rect 20343 3760 20352 3800
rect 20392 3760 20434 3800
rect 20474 3760 20516 3800
rect 20556 3760 20598 3800
rect 20638 3760 20680 3800
rect 20720 3760 20729 3800
rect 24343 3760 24352 3800
rect 24392 3760 24434 3800
rect 24474 3760 24516 3800
rect 24556 3760 24598 3800
rect 24638 3760 24680 3800
rect 24720 3760 24729 3800
rect 28343 3760 28352 3800
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28720 3760 28729 3800
rect 32343 3760 32352 3800
rect 32392 3760 32434 3800
rect 32474 3760 32516 3800
rect 32556 3760 32598 3800
rect 32638 3760 32680 3800
rect 32720 3760 32729 3800
rect 36343 3760 36352 3800
rect 36392 3760 36434 3800
rect 36474 3760 36516 3800
rect 36556 3760 36598 3800
rect 36638 3760 36680 3800
rect 36720 3760 36729 3800
rect 40343 3760 40352 3800
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40720 3760 40729 3800
rect 44343 3760 44352 3800
rect 44392 3760 44434 3800
rect 44474 3760 44516 3800
rect 44556 3760 44598 3800
rect 44638 3760 44680 3800
rect 44720 3760 44729 3800
rect 48343 3760 48352 3800
rect 48392 3760 48434 3800
rect 48474 3760 48516 3800
rect 48556 3760 48598 3800
rect 48638 3760 48680 3800
rect 48720 3760 48729 3800
rect 52343 3760 52352 3800
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52720 3760 52729 3800
rect 56343 3760 56352 3800
rect 56392 3760 56434 3800
rect 56474 3760 56516 3800
rect 56556 3760 56598 3800
rect 56638 3760 56680 3800
rect 56720 3760 56729 3800
rect 60343 3760 60352 3800
rect 60392 3760 60434 3800
rect 60474 3760 60516 3800
rect 60556 3760 60598 3800
rect 60638 3760 60680 3800
rect 60720 3760 60729 3800
rect 64343 3760 64352 3800
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64720 3760 64729 3800
rect 68343 3760 68352 3800
rect 68392 3760 68434 3800
rect 68474 3760 68516 3800
rect 68556 3760 68598 3800
rect 68638 3760 68680 3800
rect 68720 3760 68729 3800
rect 72343 3760 72352 3800
rect 72392 3760 72434 3800
rect 72474 3760 72516 3800
rect 72556 3760 72598 3800
rect 72638 3760 72680 3800
rect 72720 3760 72729 3800
rect 76343 3760 76352 3800
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76720 3760 76729 3800
rect 80343 3760 80352 3800
rect 80392 3760 80434 3800
rect 80474 3760 80516 3800
rect 80556 3760 80598 3800
rect 80638 3760 80680 3800
rect 80720 3760 80729 3800
rect 84343 3760 84352 3800
rect 84392 3760 84434 3800
rect 84474 3760 84516 3800
rect 84556 3760 84598 3800
rect 84638 3760 84680 3800
rect 84720 3760 84729 3800
rect 88343 3760 88352 3800
rect 88392 3760 88434 3800
rect 88474 3760 88516 3800
rect 88556 3760 88598 3800
rect 88638 3760 88680 3800
rect 88720 3760 88729 3800
rect 92343 3760 92352 3800
rect 92392 3760 92434 3800
rect 92474 3760 92516 3800
rect 92556 3760 92598 3800
rect 92638 3760 92680 3800
rect 92720 3760 92729 3800
rect 96343 3760 96352 3800
rect 96392 3760 96434 3800
rect 96474 3760 96516 3800
rect 96556 3760 96598 3800
rect 96638 3760 96680 3800
rect 96720 3760 96729 3800
rect 643 3172 652 3212
rect 692 3172 701 3212
rect 0 3128 80 3148
rect 652 3128 692 3172
rect 0 3088 692 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 7103 3004 7112 3044
rect 7152 3004 7194 3044
rect 7234 3004 7276 3044
rect 7316 3004 7358 3044
rect 7398 3004 7440 3044
rect 7480 3004 7489 3044
rect 11103 3004 11112 3044
rect 11152 3004 11194 3044
rect 11234 3004 11276 3044
rect 11316 3004 11358 3044
rect 11398 3004 11440 3044
rect 11480 3004 11489 3044
rect 15103 3004 15112 3044
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15480 3004 15489 3044
rect 19103 3004 19112 3044
rect 19152 3004 19194 3044
rect 19234 3004 19276 3044
rect 19316 3004 19358 3044
rect 19398 3004 19440 3044
rect 19480 3004 19489 3044
rect 23103 3004 23112 3044
rect 23152 3004 23194 3044
rect 23234 3004 23276 3044
rect 23316 3004 23358 3044
rect 23398 3004 23440 3044
rect 23480 3004 23489 3044
rect 27103 3004 27112 3044
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27480 3004 27489 3044
rect 31103 3004 31112 3044
rect 31152 3004 31194 3044
rect 31234 3004 31276 3044
rect 31316 3004 31358 3044
rect 31398 3004 31440 3044
rect 31480 3004 31489 3044
rect 35103 3004 35112 3044
rect 35152 3004 35194 3044
rect 35234 3004 35276 3044
rect 35316 3004 35358 3044
rect 35398 3004 35440 3044
rect 35480 3004 35489 3044
rect 39103 3004 39112 3044
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39480 3004 39489 3044
rect 43103 3004 43112 3044
rect 43152 3004 43194 3044
rect 43234 3004 43276 3044
rect 43316 3004 43358 3044
rect 43398 3004 43440 3044
rect 43480 3004 43489 3044
rect 47103 3004 47112 3044
rect 47152 3004 47194 3044
rect 47234 3004 47276 3044
rect 47316 3004 47358 3044
rect 47398 3004 47440 3044
rect 47480 3004 47489 3044
rect 51103 3004 51112 3044
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51480 3004 51489 3044
rect 55103 3004 55112 3044
rect 55152 3004 55194 3044
rect 55234 3004 55276 3044
rect 55316 3004 55358 3044
rect 55398 3004 55440 3044
rect 55480 3004 55489 3044
rect 59103 3004 59112 3044
rect 59152 3004 59194 3044
rect 59234 3004 59276 3044
rect 59316 3004 59358 3044
rect 59398 3004 59440 3044
rect 59480 3004 59489 3044
rect 63103 3004 63112 3044
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63480 3004 63489 3044
rect 67103 3004 67112 3044
rect 67152 3004 67194 3044
rect 67234 3004 67276 3044
rect 67316 3004 67358 3044
rect 67398 3004 67440 3044
rect 67480 3004 67489 3044
rect 71103 3004 71112 3044
rect 71152 3004 71194 3044
rect 71234 3004 71276 3044
rect 71316 3004 71358 3044
rect 71398 3004 71440 3044
rect 71480 3004 71489 3044
rect 75103 3004 75112 3044
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75480 3004 75489 3044
rect 79103 3004 79112 3044
rect 79152 3004 79194 3044
rect 79234 3004 79276 3044
rect 79316 3004 79358 3044
rect 79398 3004 79440 3044
rect 79480 3004 79489 3044
rect 83103 3004 83112 3044
rect 83152 3004 83194 3044
rect 83234 3004 83276 3044
rect 83316 3004 83358 3044
rect 83398 3004 83440 3044
rect 83480 3004 83489 3044
rect 87103 3004 87112 3044
rect 87152 3004 87194 3044
rect 87234 3004 87276 3044
rect 87316 3004 87358 3044
rect 87398 3004 87440 3044
rect 87480 3004 87489 3044
rect 91103 3004 91112 3044
rect 91152 3004 91194 3044
rect 91234 3004 91276 3044
rect 91316 3004 91358 3044
rect 91398 3004 91440 3044
rect 91480 3004 91489 3044
rect 95103 3004 95112 3044
rect 95152 3004 95194 3044
rect 95234 3004 95276 3044
rect 95316 3004 95358 3044
rect 95398 3004 95440 3044
rect 95480 3004 95489 3044
rect 99103 3004 99112 3044
rect 99152 3004 99194 3044
rect 99234 3004 99276 3044
rect 99316 3004 99358 3044
rect 99398 3004 99440 3044
rect 99480 3004 99489 3044
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 8343 2248 8352 2288
rect 8392 2248 8434 2288
rect 8474 2248 8516 2288
rect 8556 2248 8598 2288
rect 8638 2248 8680 2288
rect 8720 2248 8729 2288
rect 12343 2248 12352 2288
rect 12392 2248 12434 2288
rect 12474 2248 12516 2288
rect 12556 2248 12598 2288
rect 12638 2248 12680 2288
rect 12720 2248 12729 2288
rect 16343 2248 16352 2288
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16720 2248 16729 2288
rect 20343 2248 20352 2288
rect 20392 2248 20434 2288
rect 20474 2248 20516 2288
rect 20556 2248 20598 2288
rect 20638 2248 20680 2288
rect 20720 2248 20729 2288
rect 24343 2248 24352 2288
rect 24392 2248 24434 2288
rect 24474 2248 24516 2288
rect 24556 2248 24598 2288
rect 24638 2248 24680 2288
rect 24720 2248 24729 2288
rect 28343 2248 28352 2288
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28720 2248 28729 2288
rect 32343 2248 32352 2288
rect 32392 2248 32434 2288
rect 32474 2248 32516 2288
rect 32556 2248 32598 2288
rect 32638 2248 32680 2288
rect 32720 2248 32729 2288
rect 36343 2248 36352 2288
rect 36392 2248 36434 2288
rect 36474 2248 36516 2288
rect 36556 2248 36598 2288
rect 36638 2248 36680 2288
rect 36720 2248 36729 2288
rect 40343 2248 40352 2288
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40720 2248 40729 2288
rect 44343 2248 44352 2288
rect 44392 2248 44434 2288
rect 44474 2248 44516 2288
rect 44556 2248 44598 2288
rect 44638 2248 44680 2288
rect 44720 2248 44729 2288
rect 48343 2248 48352 2288
rect 48392 2248 48434 2288
rect 48474 2248 48516 2288
rect 48556 2248 48598 2288
rect 48638 2248 48680 2288
rect 48720 2248 48729 2288
rect 52343 2248 52352 2288
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52720 2248 52729 2288
rect 56343 2248 56352 2288
rect 56392 2248 56434 2288
rect 56474 2248 56516 2288
rect 56556 2248 56598 2288
rect 56638 2248 56680 2288
rect 56720 2248 56729 2288
rect 60343 2248 60352 2288
rect 60392 2248 60434 2288
rect 60474 2248 60516 2288
rect 60556 2248 60598 2288
rect 60638 2248 60680 2288
rect 60720 2248 60729 2288
rect 64343 2248 64352 2288
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64720 2248 64729 2288
rect 68343 2248 68352 2288
rect 68392 2248 68434 2288
rect 68474 2248 68516 2288
rect 68556 2248 68598 2288
rect 68638 2248 68680 2288
rect 68720 2248 68729 2288
rect 72343 2248 72352 2288
rect 72392 2248 72434 2288
rect 72474 2248 72516 2288
rect 72556 2248 72598 2288
rect 72638 2248 72680 2288
rect 72720 2248 72729 2288
rect 76343 2248 76352 2288
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76720 2248 76729 2288
rect 80343 2248 80352 2288
rect 80392 2248 80434 2288
rect 80474 2248 80516 2288
rect 80556 2248 80598 2288
rect 80638 2248 80680 2288
rect 80720 2248 80729 2288
rect 84343 2248 84352 2288
rect 84392 2248 84434 2288
rect 84474 2248 84516 2288
rect 84556 2248 84598 2288
rect 84638 2248 84680 2288
rect 84720 2248 84729 2288
rect 88343 2248 88352 2288
rect 88392 2248 88434 2288
rect 88474 2248 88516 2288
rect 88556 2248 88598 2288
rect 88638 2248 88680 2288
rect 88720 2248 88729 2288
rect 92343 2248 92352 2288
rect 92392 2248 92434 2288
rect 92474 2248 92516 2288
rect 92556 2248 92598 2288
rect 92638 2248 92680 2288
rect 92720 2248 92729 2288
rect 96343 2248 96352 2288
rect 96392 2248 96434 2288
rect 96474 2248 96516 2288
rect 96556 2248 96598 2288
rect 96638 2248 96680 2288
rect 96720 2248 96729 2288
rect 0 2228 80 2248
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 7103 1492 7112 1532
rect 7152 1492 7194 1532
rect 7234 1492 7276 1532
rect 7316 1492 7358 1532
rect 7398 1492 7440 1532
rect 7480 1492 7489 1532
rect 11103 1492 11112 1532
rect 11152 1492 11194 1532
rect 11234 1492 11276 1532
rect 11316 1492 11358 1532
rect 11398 1492 11440 1532
rect 11480 1492 11489 1532
rect 15103 1492 15112 1532
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15480 1492 15489 1532
rect 19103 1492 19112 1532
rect 19152 1492 19194 1532
rect 19234 1492 19276 1532
rect 19316 1492 19358 1532
rect 19398 1492 19440 1532
rect 19480 1492 19489 1532
rect 23103 1492 23112 1532
rect 23152 1492 23194 1532
rect 23234 1492 23276 1532
rect 23316 1492 23358 1532
rect 23398 1492 23440 1532
rect 23480 1492 23489 1532
rect 27103 1492 27112 1532
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27480 1492 27489 1532
rect 31103 1492 31112 1532
rect 31152 1492 31194 1532
rect 31234 1492 31276 1532
rect 31316 1492 31358 1532
rect 31398 1492 31440 1532
rect 31480 1492 31489 1532
rect 35103 1492 35112 1532
rect 35152 1492 35194 1532
rect 35234 1492 35276 1532
rect 35316 1492 35358 1532
rect 35398 1492 35440 1532
rect 35480 1492 35489 1532
rect 39103 1492 39112 1532
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39480 1492 39489 1532
rect 43103 1492 43112 1532
rect 43152 1492 43194 1532
rect 43234 1492 43276 1532
rect 43316 1492 43358 1532
rect 43398 1492 43440 1532
rect 43480 1492 43489 1532
rect 47103 1492 47112 1532
rect 47152 1492 47194 1532
rect 47234 1492 47276 1532
rect 47316 1492 47358 1532
rect 47398 1492 47440 1532
rect 47480 1492 47489 1532
rect 51103 1492 51112 1532
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51480 1492 51489 1532
rect 55103 1492 55112 1532
rect 55152 1492 55194 1532
rect 55234 1492 55276 1532
rect 55316 1492 55358 1532
rect 55398 1492 55440 1532
rect 55480 1492 55489 1532
rect 59103 1492 59112 1532
rect 59152 1492 59194 1532
rect 59234 1492 59276 1532
rect 59316 1492 59358 1532
rect 59398 1492 59440 1532
rect 59480 1492 59489 1532
rect 63103 1492 63112 1532
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63480 1492 63489 1532
rect 67103 1492 67112 1532
rect 67152 1492 67194 1532
rect 67234 1492 67276 1532
rect 67316 1492 67358 1532
rect 67398 1492 67440 1532
rect 67480 1492 67489 1532
rect 71103 1492 71112 1532
rect 71152 1492 71194 1532
rect 71234 1492 71276 1532
rect 71316 1492 71358 1532
rect 71398 1492 71440 1532
rect 71480 1492 71489 1532
rect 75103 1492 75112 1532
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75480 1492 75489 1532
rect 79103 1492 79112 1532
rect 79152 1492 79194 1532
rect 79234 1492 79276 1532
rect 79316 1492 79358 1532
rect 79398 1492 79440 1532
rect 79480 1492 79489 1532
rect 83103 1492 83112 1532
rect 83152 1492 83194 1532
rect 83234 1492 83276 1532
rect 83316 1492 83358 1532
rect 83398 1492 83440 1532
rect 83480 1492 83489 1532
rect 87103 1492 87112 1532
rect 87152 1492 87194 1532
rect 87234 1492 87276 1532
rect 87316 1492 87358 1532
rect 87398 1492 87440 1532
rect 87480 1492 87489 1532
rect 91103 1492 91112 1532
rect 91152 1492 91194 1532
rect 91234 1492 91276 1532
rect 91316 1492 91358 1532
rect 91398 1492 91440 1532
rect 91480 1492 91489 1532
rect 95103 1492 95112 1532
rect 95152 1492 95194 1532
rect 95234 1492 95276 1532
rect 95316 1492 95358 1532
rect 95398 1492 95440 1532
rect 95480 1492 95489 1532
rect 99103 1492 99112 1532
rect 99152 1492 99194 1532
rect 99234 1492 99276 1532
rect 99316 1492 99358 1532
rect 99398 1492 99440 1532
rect 99480 1492 99489 1532
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 8343 736 8352 776
rect 8392 736 8434 776
rect 8474 736 8516 776
rect 8556 736 8598 776
rect 8638 736 8680 776
rect 8720 736 8729 776
rect 12343 736 12352 776
rect 12392 736 12434 776
rect 12474 736 12516 776
rect 12556 736 12598 776
rect 12638 736 12680 776
rect 12720 736 12729 776
rect 16343 736 16352 776
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16720 736 16729 776
rect 20343 736 20352 776
rect 20392 736 20434 776
rect 20474 736 20516 776
rect 20556 736 20598 776
rect 20638 736 20680 776
rect 20720 736 20729 776
rect 24343 736 24352 776
rect 24392 736 24434 776
rect 24474 736 24516 776
rect 24556 736 24598 776
rect 24638 736 24680 776
rect 24720 736 24729 776
rect 28343 736 28352 776
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28720 736 28729 776
rect 32343 736 32352 776
rect 32392 736 32434 776
rect 32474 736 32516 776
rect 32556 736 32598 776
rect 32638 736 32680 776
rect 32720 736 32729 776
rect 36343 736 36352 776
rect 36392 736 36434 776
rect 36474 736 36516 776
rect 36556 736 36598 776
rect 36638 736 36680 776
rect 36720 736 36729 776
rect 40343 736 40352 776
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40720 736 40729 776
rect 44343 736 44352 776
rect 44392 736 44434 776
rect 44474 736 44516 776
rect 44556 736 44598 776
rect 44638 736 44680 776
rect 44720 736 44729 776
rect 48343 736 48352 776
rect 48392 736 48434 776
rect 48474 736 48516 776
rect 48556 736 48598 776
rect 48638 736 48680 776
rect 48720 736 48729 776
rect 52343 736 52352 776
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52720 736 52729 776
rect 56343 736 56352 776
rect 56392 736 56434 776
rect 56474 736 56516 776
rect 56556 736 56598 776
rect 56638 736 56680 776
rect 56720 736 56729 776
rect 60343 736 60352 776
rect 60392 736 60434 776
rect 60474 736 60516 776
rect 60556 736 60598 776
rect 60638 736 60680 776
rect 60720 736 60729 776
rect 64343 736 64352 776
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64720 736 64729 776
rect 68343 736 68352 776
rect 68392 736 68434 776
rect 68474 736 68516 776
rect 68556 736 68598 776
rect 68638 736 68680 776
rect 68720 736 68729 776
rect 72343 736 72352 776
rect 72392 736 72434 776
rect 72474 736 72516 776
rect 72556 736 72598 776
rect 72638 736 72680 776
rect 72720 736 72729 776
rect 76343 736 76352 776
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76720 736 76729 776
rect 80343 736 80352 776
rect 80392 736 80434 776
rect 80474 736 80516 776
rect 80556 736 80598 776
rect 80638 736 80680 776
rect 80720 736 80729 776
rect 84343 736 84352 776
rect 84392 736 84434 776
rect 84474 736 84516 776
rect 84556 736 84598 776
rect 84638 736 84680 776
rect 84720 736 84729 776
rect 88343 736 88352 776
rect 88392 736 88434 776
rect 88474 736 88516 776
rect 88556 736 88598 776
rect 88638 736 88680 776
rect 88720 736 88729 776
rect 92343 736 92352 776
rect 92392 736 92434 776
rect 92474 736 92516 776
rect 92556 736 92598 776
rect 92638 736 92680 776
rect 92720 736 92729 776
rect 96343 736 96352 776
rect 96392 736 96434 776
rect 96474 736 96516 776
rect 96556 736 96598 776
rect 96638 736 96680 776
rect 96720 736 96729 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 8352 38536 8392 38576
rect 8434 38536 8474 38576
rect 8516 38536 8556 38576
rect 8598 38536 8638 38576
rect 8680 38536 8720 38576
rect 12352 38536 12392 38576
rect 12434 38536 12474 38576
rect 12516 38536 12556 38576
rect 12598 38536 12638 38576
rect 12680 38536 12720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 20352 38536 20392 38576
rect 20434 38536 20474 38576
rect 20516 38536 20556 38576
rect 20598 38536 20638 38576
rect 20680 38536 20720 38576
rect 24352 38536 24392 38576
rect 24434 38536 24474 38576
rect 24516 38536 24556 38576
rect 24598 38536 24638 38576
rect 24680 38536 24720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 32352 38536 32392 38576
rect 32434 38536 32474 38576
rect 32516 38536 32556 38576
rect 32598 38536 32638 38576
rect 32680 38536 32720 38576
rect 36352 38536 36392 38576
rect 36434 38536 36474 38576
rect 36516 38536 36556 38576
rect 36598 38536 36638 38576
rect 36680 38536 36720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 44352 38536 44392 38576
rect 44434 38536 44474 38576
rect 44516 38536 44556 38576
rect 44598 38536 44638 38576
rect 44680 38536 44720 38576
rect 48352 38536 48392 38576
rect 48434 38536 48474 38576
rect 48516 38536 48556 38576
rect 48598 38536 48638 38576
rect 48680 38536 48720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 56352 38536 56392 38576
rect 56434 38536 56474 38576
rect 56516 38536 56556 38576
rect 56598 38536 56638 38576
rect 56680 38536 56720 38576
rect 60352 38536 60392 38576
rect 60434 38536 60474 38576
rect 60516 38536 60556 38576
rect 60598 38536 60638 38576
rect 60680 38536 60720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 68352 38536 68392 38576
rect 68434 38536 68474 38576
rect 68516 38536 68556 38576
rect 68598 38536 68638 38576
rect 68680 38536 68720 38576
rect 72352 38536 72392 38576
rect 72434 38536 72474 38576
rect 72516 38536 72556 38576
rect 72598 38536 72638 38576
rect 72680 38536 72720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 80352 38536 80392 38576
rect 80434 38536 80474 38576
rect 80516 38536 80556 38576
rect 80598 38536 80638 38576
rect 80680 38536 80720 38576
rect 84352 38536 84392 38576
rect 84434 38536 84474 38576
rect 84516 38536 84556 38576
rect 84598 38536 84638 38576
rect 84680 38536 84720 38576
rect 88352 38536 88392 38576
rect 88434 38536 88474 38576
rect 88516 38536 88556 38576
rect 88598 38536 88638 38576
rect 88680 38536 88720 38576
rect 92352 38536 92392 38576
rect 92434 38536 92474 38576
rect 92516 38536 92556 38576
rect 92598 38536 92638 38576
rect 92680 38536 92720 38576
rect 96352 38536 96392 38576
rect 96434 38536 96474 38576
rect 96516 38536 96556 38576
rect 96598 38536 96638 38576
rect 96680 38536 96720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 7112 37780 7152 37820
rect 7194 37780 7234 37820
rect 7276 37780 7316 37820
rect 7358 37780 7398 37820
rect 7440 37780 7480 37820
rect 11112 37780 11152 37820
rect 11194 37780 11234 37820
rect 11276 37780 11316 37820
rect 11358 37780 11398 37820
rect 11440 37780 11480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 19112 37780 19152 37820
rect 19194 37780 19234 37820
rect 19276 37780 19316 37820
rect 19358 37780 19398 37820
rect 19440 37780 19480 37820
rect 23112 37780 23152 37820
rect 23194 37780 23234 37820
rect 23276 37780 23316 37820
rect 23358 37780 23398 37820
rect 23440 37780 23480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 31112 37780 31152 37820
rect 31194 37780 31234 37820
rect 31276 37780 31316 37820
rect 31358 37780 31398 37820
rect 31440 37780 31480 37820
rect 35112 37780 35152 37820
rect 35194 37780 35234 37820
rect 35276 37780 35316 37820
rect 35358 37780 35398 37820
rect 35440 37780 35480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 43112 37780 43152 37820
rect 43194 37780 43234 37820
rect 43276 37780 43316 37820
rect 43358 37780 43398 37820
rect 43440 37780 43480 37820
rect 47112 37780 47152 37820
rect 47194 37780 47234 37820
rect 47276 37780 47316 37820
rect 47358 37780 47398 37820
rect 47440 37780 47480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 55112 37780 55152 37820
rect 55194 37780 55234 37820
rect 55276 37780 55316 37820
rect 55358 37780 55398 37820
rect 55440 37780 55480 37820
rect 59112 37780 59152 37820
rect 59194 37780 59234 37820
rect 59276 37780 59316 37820
rect 59358 37780 59398 37820
rect 59440 37780 59480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 67112 37780 67152 37820
rect 67194 37780 67234 37820
rect 67276 37780 67316 37820
rect 67358 37780 67398 37820
rect 67440 37780 67480 37820
rect 71112 37780 71152 37820
rect 71194 37780 71234 37820
rect 71276 37780 71316 37820
rect 71358 37780 71398 37820
rect 71440 37780 71480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 79112 37780 79152 37820
rect 79194 37780 79234 37820
rect 79276 37780 79316 37820
rect 79358 37780 79398 37820
rect 79440 37780 79480 37820
rect 83112 37780 83152 37820
rect 83194 37780 83234 37820
rect 83276 37780 83316 37820
rect 83358 37780 83398 37820
rect 83440 37780 83480 37820
rect 87112 37780 87152 37820
rect 87194 37780 87234 37820
rect 87276 37780 87316 37820
rect 87358 37780 87398 37820
rect 87440 37780 87480 37820
rect 91112 37780 91152 37820
rect 91194 37780 91234 37820
rect 91276 37780 91316 37820
rect 91358 37780 91398 37820
rect 91440 37780 91480 37820
rect 95112 37780 95152 37820
rect 95194 37780 95234 37820
rect 95276 37780 95316 37820
rect 95358 37780 95398 37820
rect 95440 37780 95480 37820
rect 99112 37780 99152 37820
rect 99194 37780 99234 37820
rect 99276 37780 99316 37820
rect 99358 37780 99398 37820
rect 99440 37780 99480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 8352 37024 8392 37064
rect 8434 37024 8474 37064
rect 8516 37024 8556 37064
rect 8598 37024 8638 37064
rect 8680 37024 8720 37064
rect 12352 37024 12392 37064
rect 12434 37024 12474 37064
rect 12516 37024 12556 37064
rect 12598 37024 12638 37064
rect 12680 37024 12720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 20352 37024 20392 37064
rect 20434 37024 20474 37064
rect 20516 37024 20556 37064
rect 20598 37024 20638 37064
rect 20680 37024 20720 37064
rect 24352 37024 24392 37064
rect 24434 37024 24474 37064
rect 24516 37024 24556 37064
rect 24598 37024 24638 37064
rect 24680 37024 24720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 32352 37024 32392 37064
rect 32434 37024 32474 37064
rect 32516 37024 32556 37064
rect 32598 37024 32638 37064
rect 32680 37024 32720 37064
rect 36352 37024 36392 37064
rect 36434 37024 36474 37064
rect 36516 37024 36556 37064
rect 36598 37024 36638 37064
rect 36680 37024 36720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 44352 37024 44392 37064
rect 44434 37024 44474 37064
rect 44516 37024 44556 37064
rect 44598 37024 44638 37064
rect 44680 37024 44720 37064
rect 48352 37024 48392 37064
rect 48434 37024 48474 37064
rect 48516 37024 48556 37064
rect 48598 37024 48638 37064
rect 48680 37024 48720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 56352 37024 56392 37064
rect 56434 37024 56474 37064
rect 56516 37024 56556 37064
rect 56598 37024 56638 37064
rect 56680 37024 56720 37064
rect 60352 37024 60392 37064
rect 60434 37024 60474 37064
rect 60516 37024 60556 37064
rect 60598 37024 60638 37064
rect 60680 37024 60720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 68352 37024 68392 37064
rect 68434 37024 68474 37064
rect 68516 37024 68556 37064
rect 68598 37024 68638 37064
rect 68680 37024 68720 37064
rect 72352 37024 72392 37064
rect 72434 37024 72474 37064
rect 72516 37024 72556 37064
rect 72598 37024 72638 37064
rect 72680 37024 72720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 80352 37024 80392 37064
rect 80434 37024 80474 37064
rect 80516 37024 80556 37064
rect 80598 37024 80638 37064
rect 80680 37024 80720 37064
rect 84352 37024 84392 37064
rect 84434 37024 84474 37064
rect 84516 37024 84556 37064
rect 84598 37024 84638 37064
rect 84680 37024 84720 37064
rect 88352 37024 88392 37064
rect 88434 37024 88474 37064
rect 88516 37024 88556 37064
rect 88598 37024 88638 37064
rect 88680 37024 88720 37064
rect 92352 37024 92392 37064
rect 92434 37024 92474 37064
rect 92516 37024 92556 37064
rect 92598 37024 92638 37064
rect 92680 37024 92720 37064
rect 96352 37024 96392 37064
rect 96434 37024 96474 37064
rect 96516 37024 96556 37064
rect 96598 37024 96638 37064
rect 96680 37024 96720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 7112 36268 7152 36308
rect 7194 36268 7234 36308
rect 7276 36268 7316 36308
rect 7358 36268 7398 36308
rect 7440 36268 7480 36308
rect 11112 36268 11152 36308
rect 11194 36268 11234 36308
rect 11276 36268 11316 36308
rect 11358 36268 11398 36308
rect 11440 36268 11480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 19112 36268 19152 36308
rect 19194 36268 19234 36308
rect 19276 36268 19316 36308
rect 19358 36268 19398 36308
rect 19440 36268 19480 36308
rect 23112 36268 23152 36308
rect 23194 36268 23234 36308
rect 23276 36268 23316 36308
rect 23358 36268 23398 36308
rect 23440 36268 23480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 31112 36268 31152 36308
rect 31194 36268 31234 36308
rect 31276 36268 31316 36308
rect 31358 36268 31398 36308
rect 31440 36268 31480 36308
rect 35112 36268 35152 36308
rect 35194 36268 35234 36308
rect 35276 36268 35316 36308
rect 35358 36268 35398 36308
rect 35440 36268 35480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 43112 36268 43152 36308
rect 43194 36268 43234 36308
rect 43276 36268 43316 36308
rect 43358 36268 43398 36308
rect 43440 36268 43480 36308
rect 47112 36268 47152 36308
rect 47194 36268 47234 36308
rect 47276 36268 47316 36308
rect 47358 36268 47398 36308
rect 47440 36268 47480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 55112 36268 55152 36308
rect 55194 36268 55234 36308
rect 55276 36268 55316 36308
rect 55358 36268 55398 36308
rect 55440 36268 55480 36308
rect 59112 36268 59152 36308
rect 59194 36268 59234 36308
rect 59276 36268 59316 36308
rect 59358 36268 59398 36308
rect 59440 36268 59480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 67112 36268 67152 36308
rect 67194 36268 67234 36308
rect 67276 36268 67316 36308
rect 67358 36268 67398 36308
rect 67440 36268 67480 36308
rect 71112 36268 71152 36308
rect 71194 36268 71234 36308
rect 71276 36268 71316 36308
rect 71358 36268 71398 36308
rect 71440 36268 71480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 79112 36268 79152 36308
rect 79194 36268 79234 36308
rect 79276 36268 79316 36308
rect 79358 36268 79398 36308
rect 79440 36268 79480 36308
rect 83112 36268 83152 36308
rect 83194 36268 83234 36308
rect 83276 36268 83316 36308
rect 83358 36268 83398 36308
rect 83440 36268 83480 36308
rect 87112 36268 87152 36308
rect 87194 36268 87234 36308
rect 87276 36268 87316 36308
rect 87358 36268 87398 36308
rect 87440 36268 87480 36308
rect 91112 36268 91152 36308
rect 91194 36268 91234 36308
rect 91276 36268 91316 36308
rect 91358 36268 91398 36308
rect 91440 36268 91480 36308
rect 95112 36268 95152 36308
rect 95194 36268 95234 36308
rect 95276 36268 95316 36308
rect 95358 36268 95398 36308
rect 95440 36268 95480 36308
rect 99112 36268 99152 36308
rect 99194 36268 99234 36308
rect 99276 36268 99316 36308
rect 99358 36268 99398 36308
rect 99440 36268 99480 36308
rect 76780 35680 76820 35720
rect 85228 35680 85268 35720
rect 92236 35680 92276 35720
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 8352 35512 8392 35552
rect 8434 35512 8474 35552
rect 8516 35512 8556 35552
rect 8598 35512 8638 35552
rect 8680 35512 8720 35552
rect 12352 35512 12392 35552
rect 12434 35512 12474 35552
rect 12516 35512 12556 35552
rect 12598 35512 12638 35552
rect 12680 35512 12720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 20352 35512 20392 35552
rect 20434 35512 20474 35552
rect 20516 35512 20556 35552
rect 20598 35512 20638 35552
rect 20680 35512 20720 35552
rect 24352 35512 24392 35552
rect 24434 35512 24474 35552
rect 24516 35512 24556 35552
rect 24598 35512 24638 35552
rect 24680 35512 24720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 32352 35512 32392 35552
rect 32434 35512 32474 35552
rect 32516 35512 32556 35552
rect 32598 35512 32638 35552
rect 32680 35512 32720 35552
rect 36352 35512 36392 35552
rect 36434 35512 36474 35552
rect 36516 35512 36556 35552
rect 36598 35512 36638 35552
rect 36680 35512 36720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 44352 35512 44392 35552
rect 44434 35512 44474 35552
rect 44516 35512 44556 35552
rect 44598 35512 44638 35552
rect 44680 35512 44720 35552
rect 48352 35512 48392 35552
rect 48434 35512 48474 35552
rect 48516 35512 48556 35552
rect 48598 35512 48638 35552
rect 48680 35512 48720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 56352 35512 56392 35552
rect 56434 35512 56474 35552
rect 56516 35512 56556 35552
rect 56598 35512 56638 35552
rect 56680 35512 56720 35552
rect 60352 35512 60392 35552
rect 60434 35512 60474 35552
rect 60516 35512 60556 35552
rect 60598 35512 60638 35552
rect 60680 35512 60720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 68352 35512 68392 35552
rect 68434 35512 68474 35552
rect 68516 35512 68556 35552
rect 68598 35512 68638 35552
rect 68680 35512 68720 35552
rect 72352 35512 72392 35552
rect 72434 35512 72474 35552
rect 72516 35512 72556 35552
rect 72598 35512 72638 35552
rect 72680 35512 72720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 80352 35512 80392 35552
rect 80434 35512 80474 35552
rect 80516 35512 80556 35552
rect 80598 35512 80638 35552
rect 80680 35512 80720 35552
rect 84352 35512 84392 35552
rect 84434 35512 84474 35552
rect 84516 35512 84556 35552
rect 84598 35512 84638 35552
rect 84680 35512 84720 35552
rect 88352 35512 88392 35552
rect 88434 35512 88474 35552
rect 88516 35512 88556 35552
rect 88598 35512 88638 35552
rect 88680 35512 88720 35552
rect 92352 35512 92392 35552
rect 92434 35512 92474 35552
rect 92516 35512 92556 35552
rect 92598 35512 92638 35552
rect 92680 35512 92720 35552
rect 96352 35512 96392 35552
rect 96434 35512 96474 35552
rect 96516 35512 96556 35552
rect 96598 35512 96638 35552
rect 96680 35512 96720 35552
rect 89932 35260 89972 35300
rect 86668 34924 86708 34964
rect 86956 34924 86996 34964
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 7112 34756 7152 34796
rect 7194 34756 7234 34796
rect 7276 34756 7316 34796
rect 7358 34756 7398 34796
rect 7440 34756 7480 34796
rect 11112 34756 11152 34796
rect 11194 34756 11234 34796
rect 11276 34756 11316 34796
rect 11358 34756 11398 34796
rect 11440 34756 11480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 19112 34756 19152 34796
rect 19194 34756 19234 34796
rect 19276 34756 19316 34796
rect 19358 34756 19398 34796
rect 19440 34756 19480 34796
rect 23112 34756 23152 34796
rect 23194 34756 23234 34796
rect 23276 34756 23316 34796
rect 23358 34756 23398 34796
rect 23440 34756 23480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 31112 34756 31152 34796
rect 31194 34756 31234 34796
rect 31276 34756 31316 34796
rect 31358 34756 31398 34796
rect 31440 34756 31480 34796
rect 35112 34756 35152 34796
rect 35194 34756 35234 34796
rect 35276 34756 35316 34796
rect 35358 34756 35398 34796
rect 35440 34756 35480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 43112 34756 43152 34796
rect 43194 34756 43234 34796
rect 43276 34756 43316 34796
rect 43358 34756 43398 34796
rect 43440 34756 43480 34796
rect 47112 34756 47152 34796
rect 47194 34756 47234 34796
rect 47276 34756 47316 34796
rect 47358 34756 47398 34796
rect 47440 34756 47480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 55112 34756 55152 34796
rect 55194 34756 55234 34796
rect 55276 34756 55316 34796
rect 55358 34756 55398 34796
rect 55440 34756 55480 34796
rect 59112 34756 59152 34796
rect 59194 34756 59234 34796
rect 59276 34756 59316 34796
rect 59358 34756 59398 34796
rect 59440 34756 59480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 67112 34756 67152 34796
rect 67194 34756 67234 34796
rect 67276 34756 67316 34796
rect 67358 34756 67398 34796
rect 67440 34756 67480 34796
rect 71112 34756 71152 34796
rect 71194 34756 71234 34796
rect 71276 34756 71316 34796
rect 71358 34756 71398 34796
rect 71440 34756 71480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 79112 34756 79152 34796
rect 79194 34756 79234 34796
rect 79276 34756 79316 34796
rect 79358 34756 79398 34796
rect 79440 34756 79480 34796
rect 83112 34756 83152 34796
rect 83194 34756 83234 34796
rect 83276 34756 83316 34796
rect 83358 34756 83398 34796
rect 83440 34756 83480 34796
rect 87112 34756 87152 34796
rect 87194 34756 87234 34796
rect 87276 34756 87316 34796
rect 87358 34756 87398 34796
rect 87440 34756 87480 34796
rect 91112 34756 91152 34796
rect 91194 34756 91234 34796
rect 91276 34756 91316 34796
rect 91358 34756 91398 34796
rect 91440 34756 91480 34796
rect 95112 34756 95152 34796
rect 95194 34756 95234 34796
rect 95276 34756 95316 34796
rect 95358 34756 95398 34796
rect 95440 34756 95480 34796
rect 99112 34756 99152 34796
rect 99194 34756 99234 34796
rect 99276 34756 99316 34796
rect 99358 34756 99398 34796
rect 99440 34756 99480 34796
rect 80236 34672 80276 34712
rect 86860 34588 86900 34628
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 8352 34000 8392 34040
rect 8434 34000 8474 34040
rect 8516 34000 8556 34040
rect 8598 34000 8638 34040
rect 8680 34000 8720 34040
rect 12352 34000 12392 34040
rect 12434 34000 12474 34040
rect 12516 34000 12556 34040
rect 12598 34000 12638 34040
rect 12680 34000 12720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 20352 34000 20392 34040
rect 20434 34000 20474 34040
rect 20516 34000 20556 34040
rect 20598 34000 20638 34040
rect 20680 34000 20720 34040
rect 24352 34000 24392 34040
rect 24434 34000 24474 34040
rect 24516 34000 24556 34040
rect 24598 34000 24638 34040
rect 24680 34000 24720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 32352 34000 32392 34040
rect 32434 34000 32474 34040
rect 32516 34000 32556 34040
rect 32598 34000 32638 34040
rect 32680 34000 32720 34040
rect 36352 34000 36392 34040
rect 36434 34000 36474 34040
rect 36516 34000 36556 34040
rect 36598 34000 36638 34040
rect 36680 34000 36720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 44352 34000 44392 34040
rect 44434 34000 44474 34040
rect 44516 34000 44556 34040
rect 44598 34000 44638 34040
rect 44680 34000 44720 34040
rect 48352 34000 48392 34040
rect 48434 34000 48474 34040
rect 48516 34000 48556 34040
rect 48598 34000 48638 34040
rect 48680 34000 48720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 56352 34000 56392 34040
rect 56434 34000 56474 34040
rect 56516 34000 56556 34040
rect 56598 34000 56638 34040
rect 56680 34000 56720 34040
rect 60352 34000 60392 34040
rect 60434 34000 60474 34040
rect 60516 34000 60556 34040
rect 60598 34000 60638 34040
rect 60680 34000 60720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 68352 34000 68392 34040
rect 68434 34000 68474 34040
rect 68516 34000 68556 34040
rect 68598 34000 68638 34040
rect 68680 34000 68720 34040
rect 72352 34000 72392 34040
rect 72434 34000 72474 34040
rect 72516 34000 72556 34040
rect 72598 34000 72638 34040
rect 72680 34000 72720 34040
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 80352 34000 80392 34040
rect 80434 34000 80474 34040
rect 80516 34000 80556 34040
rect 80598 34000 80638 34040
rect 80680 34000 80720 34040
rect 84352 34000 84392 34040
rect 84434 34000 84474 34040
rect 84516 34000 84556 34040
rect 84598 34000 84638 34040
rect 84680 34000 84720 34040
rect 88352 34000 88392 34040
rect 88434 34000 88474 34040
rect 88516 34000 88556 34040
rect 88598 34000 88638 34040
rect 88680 34000 88720 34040
rect 92352 34000 92392 34040
rect 92434 34000 92474 34040
rect 92516 34000 92556 34040
rect 92598 34000 92638 34040
rect 92680 34000 92720 34040
rect 96352 34000 96392 34040
rect 96434 34000 96474 34040
rect 96516 34000 96556 34040
rect 96598 34000 96638 34040
rect 96680 34000 96720 34040
rect 80236 33748 80276 33788
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 7112 33244 7152 33284
rect 7194 33244 7234 33284
rect 7276 33244 7316 33284
rect 7358 33244 7398 33284
rect 7440 33244 7480 33284
rect 11112 33244 11152 33284
rect 11194 33244 11234 33284
rect 11276 33244 11316 33284
rect 11358 33244 11398 33284
rect 11440 33244 11480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 19112 33244 19152 33284
rect 19194 33244 19234 33284
rect 19276 33244 19316 33284
rect 19358 33244 19398 33284
rect 19440 33244 19480 33284
rect 23112 33244 23152 33284
rect 23194 33244 23234 33284
rect 23276 33244 23316 33284
rect 23358 33244 23398 33284
rect 23440 33244 23480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 31112 33244 31152 33284
rect 31194 33244 31234 33284
rect 31276 33244 31316 33284
rect 31358 33244 31398 33284
rect 31440 33244 31480 33284
rect 35112 33244 35152 33284
rect 35194 33244 35234 33284
rect 35276 33244 35316 33284
rect 35358 33244 35398 33284
rect 35440 33244 35480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 43112 33244 43152 33284
rect 43194 33244 43234 33284
rect 43276 33244 43316 33284
rect 43358 33244 43398 33284
rect 43440 33244 43480 33284
rect 47112 33244 47152 33284
rect 47194 33244 47234 33284
rect 47276 33244 47316 33284
rect 47358 33244 47398 33284
rect 47440 33244 47480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 55112 33244 55152 33284
rect 55194 33244 55234 33284
rect 55276 33244 55316 33284
rect 55358 33244 55398 33284
rect 55440 33244 55480 33284
rect 59112 33244 59152 33284
rect 59194 33244 59234 33284
rect 59276 33244 59316 33284
rect 59358 33244 59398 33284
rect 59440 33244 59480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 67112 33244 67152 33284
rect 67194 33244 67234 33284
rect 67276 33244 67316 33284
rect 67358 33244 67398 33284
rect 67440 33244 67480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 8352 32488 8392 32528
rect 8434 32488 8474 32528
rect 8516 32488 8556 32528
rect 8598 32488 8638 32528
rect 8680 32488 8720 32528
rect 12352 32488 12392 32528
rect 12434 32488 12474 32528
rect 12516 32488 12556 32528
rect 12598 32488 12638 32528
rect 12680 32488 12720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 20352 32488 20392 32528
rect 20434 32488 20474 32528
rect 20516 32488 20556 32528
rect 20598 32488 20638 32528
rect 20680 32488 20720 32528
rect 24352 32488 24392 32528
rect 24434 32488 24474 32528
rect 24516 32488 24556 32528
rect 24598 32488 24638 32528
rect 24680 32488 24720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 32352 32488 32392 32528
rect 32434 32488 32474 32528
rect 32516 32488 32556 32528
rect 32598 32488 32638 32528
rect 32680 32488 32720 32528
rect 36352 32488 36392 32528
rect 36434 32488 36474 32528
rect 36516 32488 36556 32528
rect 36598 32488 36638 32528
rect 36680 32488 36720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 44352 32488 44392 32528
rect 44434 32488 44474 32528
rect 44516 32488 44556 32528
rect 44598 32488 44638 32528
rect 44680 32488 44720 32528
rect 48352 32488 48392 32528
rect 48434 32488 48474 32528
rect 48516 32488 48556 32528
rect 48598 32488 48638 32528
rect 48680 32488 48720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 56352 32488 56392 32528
rect 56434 32488 56474 32528
rect 56516 32488 56556 32528
rect 56598 32488 56638 32528
rect 56680 32488 56720 32528
rect 60352 32488 60392 32528
rect 60434 32488 60474 32528
rect 60516 32488 60556 32528
rect 60598 32488 60638 32528
rect 60680 32488 60720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 68352 32488 68392 32528
rect 68434 32488 68474 32528
rect 68516 32488 68556 32528
rect 68598 32488 68638 32528
rect 68680 32488 68720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 7112 31732 7152 31772
rect 7194 31732 7234 31772
rect 7276 31732 7316 31772
rect 7358 31732 7398 31772
rect 7440 31732 7480 31772
rect 11112 31732 11152 31772
rect 11194 31732 11234 31772
rect 11276 31732 11316 31772
rect 11358 31732 11398 31772
rect 11440 31732 11480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 19112 31732 19152 31772
rect 19194 31732 19234 31772
rect 19276 31732 19316 31772
rect 19358 31732 19398 31772
rect 19440 31732 19480 31772
rect 23112 31732 23152 31772
rect 23194 31732 23234 31772
rect 23276 31732 23316 31772
rect 23358 31732 23398 31772
rect 23440 31732 23480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 31112 31732 31152 31772
rect 31194 31732 31234 31772
rect 31276 31732 31316 31772
rect 31358 31732 31398 31772
rect 31440 31732 31480 31772
rect 35112 31732 35152 31772
rect 35194 31732 35234 31772
rect 35276 31732 35316 31772
rect 35358 31732 35398 31772
rect 35440 31732 35480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 43112 31732 43152 31772
rect 43194 31732 43234 31772
rect 43276 31732 43316 31772
rect 43358 31732 43398 31772
rect 43440 31732 43480 31772
rect 47112 31732 47152 31772
rect 47194 31732 47234 31772
rect 47276 31732 47316 31772
rect 47358 31732 47398 31772
rect 47440 31732 47480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 55112 31732 55152 31772
rect 55194 31732 55234 31772
rect 55276 31732 55316 31772
rect 55358 31732 55398 31772
rect 55440 31732 55480 31772
rect 59112 31732 59152 31772
rect 59194 31732 59234 31772
rect 59276 31732 59316 31772
rect 59358 31732 59398 31772
rect 59440 31732 59480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 67112 31732 67152 31772
rect 67194 31732 67234 31772
rect 67276 31732 67316 31772
rect 67358 31732 67398 31772
rect 67440 31732 67480 31772
rect 86956 31564 86996 31604
rect 76780 31480 76815 31520
rect 76815 31480 76820 31520
rect 85228 31480 85255 31520
rect 85255 31480 85268 31520
rect 86860 31480 86900 31520
rect 89932 31480 89945 31520
rect 89945 31480 89972 31520
rect 92236 31480 92276 31520
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 8352 30976 8392 31016
rect 8434 30976 8474 31016
rect 8516 30976 8556 31016
rect 8598 30976 8638 31016
rect 8680 30976 8720 31016
rect 12352 30976 12392 31016
rect 12434 30976 12474 31016
rect 12516 30976 12556 31016
rect 12598 30976 12638 31016
rect 12680 30976 12720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 20352 30976 20392 31016
rect 20434 30976 20474 31016
rect 20516 30976 20556 31016
rect 20598 30976 20638 31016
rect 20680 30976 20720 31016
rect 24352 30976 24392 31016
rect 24434 30976 24474 31016
rect 24516 30976 24556 31016
rect 24598 30976 24638 31016
rect 24680 30976 24720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 32352 30976 32392 31016
rect 32434 30976 32474 31016
rect 32516 30976 32556 31016
rect 32598 30976 32638 31016
rect 32680 30976 32720 31016
rect 36352 30976 36392 31016
rect 36434 30976 36474 31016
rect 36516 30976 36556 31016
rect 36598 30976 36638 31016
rect 36680 30976 36720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 44352 30976 44392 31016
rect 44434 30976 44474 31016
rect 44516 30976 44556 31016
rect 44598 30976 44638 31016
rect 44680 30976 44720 31016
rect 48352 30976 48392 31016
rect 48434 30976 48474 31016
rect 48516 30976 48556 31016
rect 48598 30976 48638 31016
rect 48680 30976 48720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 56352 30976 56392 31016
rect 56434 30976 56474 31016
rect 56516 30976 56556 31016
rect 56598 30976 56638 31016
rect 56680 30976 56720 31016
rect 60352 30976 60392 31016
rect 60434 30976 60474 31016
rect 60516 30976 60556 31016
rect 60598 30976 60638 31016
rect 60680 30976 60720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 68352 30976 68392 31016
rect 68434 30976 68474 31016
rect 68516 30976 68556 31016
rect 68598 30976 68638 31016
rect 68680 30976 68720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 7112 30220 7152 30260
rect 7194 30220 7234 30260
rect 7276 30220 7316 30260
rect 7358 30220 7398 30260
rect 7440 30220 7480 30260
rect 11112 30220 11152 30260
rect 11194 30220 11234 30260
rect 11276 30220 11316 30260
rect 11358 30220 11398 30260
rect 11440 30220 11480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 19112 30220 19152 30260
rect 19194 30220 19234 30260
rect 19276 30220 19316 30260
rect 19358 30220 19398 30260
rect 19440 30220 19480 30260
rect 23112 30220 23152 30260
rect 23194 30220 23234 30260
rect 23276 30220 23316 30260
rect 23358 30220 23398 30260
rect 23440 30220 23480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 31112 30220 31152 30260
rect 31194 30220 31234 30260
rect 31276 30220 31316 30260
rect 31358 30220 31398 30260
rect 31440 30220 31480 30260
rect 35112 30220 35152 30260
rect 35194 30220 35234 30260
rect 35276 30220 35316 30260
rect 35358 30220 35398 30260
rect 35440 30220 35480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 43112 30220 43152 30260
rect 43194 30220 43234 30260
rect 43276 30220 43316 30260
rect 43358 30220 43398 30260
rect 43440 30220 43480 30260
rect 47112 30220 47152 30260
rect 47194 30220 47234 30260
rect 47276 30220 47316 30260
rect 47358 30220 47398 30260
rect 47440 30220 47480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 55112 30220 55152 30260
rect 55194 30220 55234 30260
rect 55276 30220 55316 30260
rect 55358 30220 55398 30260
rect 55440 30220 55480 30260
rect 59112 30220 59152 30260
rect 59194 30220 59234 30260
rect 59276 30220 59316 30260
rect 59358 30220 59398 30260
rect 59440 30220 59480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 67112 30220 67152 30260
rect 67194 30220 67234 30260
rect 67276 30220 67316 30260
rect 67358 30220 67398 30260
rect 67440 30220 67480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 8352 29464 8392 29504
rect 8434 29464 8474 29504
rect 8516 29464 8556 29504
rect 8598 29464 8638 29504
rect 8680 29464 8720 29504
rect 12352 29464 12392 29504
rect 12434 29464 12474 29504
rect 12516 29464 12556 29504
rect 12598 29464 12638 29504
rect 12680 29464 12720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 20352 29464 20392 29504
rect 20434 29464 20474 29504
rect 20516 29464 20556 29504
rect 20598 29464 20638 29504
rect 20680 29464 20720 29504
rect 24352 29464 24392 29504
rect 24434 29464 24474 29504
rect 24516 29464 24556 29504
rect 24598 29464 24638 29504
rect 24680 29464 24720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 32352 29464 32392 29504
rect 32434 29464 32474 29504
rect 32516 29464 32556 29504
rect 32598 29464 32638 29504
rect 32680 29464 32720 29504
rect 36352 29464 36392 29504
rect 36434 29464 36474 29504
rect 36516 29464 36556 29504
rect 36598 29464 36638 29504
rect 36680 29464 36720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 44352 29464 44392 29504
rect 44434 29464 44474 29504
rect 44516 29464 44556 29504
rect 44598 29464 44638 29504
rect 44680 29464 44720 29504
rect 48352 29464 48392 29504
rect 48434 29464 48474 29504
rect 48516 29464 48556 29504
rect 48598 29464 48638 29504
rect 48680 29464 48720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 56352 29464 56392 29504
rect 56434 29464 56474 29504
rect 56516 29464 56556 29504
rect 56598 29464 56638 29504
rect 56680 29464 56720 29504
rect 60352 29464 60392 29504
rect 60434 29464 60474 29504
rect 60516 29464 60556 29504
rect 60598 29464 60638 29504
rect 60680 29464 60720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 68352 29464 68392 29504
rect 68434 29464 68474 29504
rect 68516 29464 68556 29504
rect 68598 29464 68638 29504
rect 68680 29464 68720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 7112 28708 7152 28748
rect 7194 28708 7234 28748
rect 7276 28708 7316 28748
rect 7358 28708 7398 28748
rect 7440 28708 7480 28748
rect 11112 28708 11152 28748
rect 11194 28708 11234 28748
rect 11276 28708 11316 28748
rect 11358 28708 11398 28748
rect 11440 28708 11480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 19112 28708 19152 28748
rect 19194 28708 19234 28748
rect 19276 28708 19316 28748
rect 19358 28708 19398 28748
rect 19440 28708 19480 28748
rect 23112 28708 23152 28748
rect 23194 28708 23234 28748
rect 23276 28708 23316 28748
rect 23358 28708 23398 28748
rect 23440 28708 23480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 31112 28708 31152 28748
rect 31194 28708 31234 28748
rect 31276 28708 31316 28748
rect 31358 28708 31398 28748
rect 31440 28708 31480 28748
rect 35112 28708 35152 28748
rect 35194 28708 35234 28748
rect 35276 28708 35316 28748
rect 35358 28708 35398 28748
rect 35440 28708 35480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 43112 28708 43152 28748
rect 43194 28708 43234 28748
rect 43276 28708 43316 28748
rect 43358 28708 43398 28748
rect 43440 28708 43480 28748
rect 47112 28708 47152 28748
rect 47194 28708 47234 28748
rect 47276 28708 47316 28748
rect 47358 28708 47398 28748
rect 47440 28708 47480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 55112 28708 55152 28748
rect 55194 28708 55234 28748
rect 55276 28708 55316 28748
rect 55358 28708 55398 28748
rect 55440 28708 55480 28748
rect 59112 28708 59152 28748
rect 59194 28708 59234 28748
rect 59276 28708 59316 28748
rect 59358 28708 59398 28748
rect 59440 28708 59480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 67112 28708 67152 28748
rect 67194 28708 67234 28748
rect 67276 28708 67316 28748
rect 67358 28708 67398 28748
rect 67440 28708 67480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 8352 27952 8392 27992
rect 8434 27952 8474 27992
rect 8516 27952 8556 27992
rect 8598 27952 8638 27992
rect 8680 27952 8720 27992
rect 12352 27952 12392 27992
rect 12434 27952 12474 27992
rect 12516 27952 12556 27992
rect 12598 27952 12638 27992
rect 12680 27952 12720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 20352 27952 20392 27992
rect 20434 27952 20474 27992
rect 20516 27952 20556 27992
rect 20598 27952 20638 27992
rect 20680 27952 20720 27992
rect 24352 27952 24392 27992
rect 24434 27952 24474 27992
rect 24516 27952 24556 27992
rect 24598 27952 24638 27992
rect 24680 27952 24720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 32352 27952 32392 27992
rect 32434 27952 32474 27992
rect 32516 27952 32556 27992
rect 32598 27952 32638 27992
rect 32680 27952 32720 27992
rect 36352 27952 36392 27992
rect 36434 27952 36474 27992
rect 36516 27952 36556 27992
rect 36598 27952 36638 27992
rect 36680 27952 36720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 44352 27952 44392 27992
rect 44434 27952 44474 27992
rect 44516 27952 44556 27992
rect 44598 27952 44638 27992
rect 44680 27952 44720 27992
rect 48352 27952 48392 27992
rect 48434 27952 48474 27992
rect 48516 27952 48556 27992
rect 48598 27952 48638 27992
rect 48680 27952 48720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 56352 27952 56392 27992
rect 56434 27952 56474 27992
rect 56516 27952 56556 27992
rect 56598 27952 56638 27992
rect 56680 27952 56720 27992
rect 60352 27952 60392 27992
rect 60434 27952 60474 27992
rect 60516 27952 60556 27992
rect 60598 27952 60638 27992
rect 60680 27952 60720 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 68352 27952 68392 27992
rect 68434 27952 68474 27992
rect 68516 27952 68556 27992
rect 68598 27952 68638 27992
rect 68680 27952 68720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 7112 27196 7152 27236
rect 7194 27196 7234 27236
rect 7276 27196 7316 27236
rect 7358 27196 7398 27236
rect 7440 27196 7480 27236
rect 11112 27196 11152 27236
rect 11194 27196 11234 27236
rect 11276 27196 11316 27236
rect 11358 27196 11398 27236
rect 11440 27196 11480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 19112 27196 19152 27236
rect 19194 27196 19234 27236
rect 19276 27196 19316 27236
rect 19358 27196 19398 27236
rect 19440 27196 19480 27236
rect 23112 27196 23152 27236
rect 23194 27196 23234 27236
rect 23276 27196 23316 27236
rect 23358 27196 23398 27236
rect 23440 27196 23480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 31112 27196 31152 27236
rect 31194 27196 31234 27236
rect 31276 27196 31316 27236
rect 31358 27196 31398 27236
rect 31440 27196 31480 27236
rect 35112 27196 35152 27236
rect 35194 27196 35234 27236
rect 35276 27196 35316 27236
rect 35358 27196 35398 27236
rect 35440 27196 35480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 43112 27196 43152 27236
rect 43194 27196 43234 27236
rect 43276 27196 43316 27236
rect 43358 27196 43398 27236
rect 43440 27196 43480 27236
rect 47112 27196 47152 27236
rect 47194 27196 47234 27236
rect 47276 27196 47316 27236
rect 47358 27196 47398 27236
rect 47440 27196 47480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 55112 27196 55152 27236
rect 55194 27196 55234 27236
rect 55276 27196 55316 27236
rect 55358 27196 55398 27236
rect 55440 27196 55480 27236
rect 59112 27196 59152 27236
rect 59194 27196 59234 27236
rect 59276 27196 59316 27236
rect 59358 27196 59398 27236
rect 59440 27196 59480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 67112 27196 67152 27236
rect 67194 27196 67234 27236
rect 67276 27196 67316 27236
rect 67358 27196 67398 27236
rect 67440 27196 67480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 8352 26440 8392 26480
rect 8434 26440 8474 26480
rect 8516 26440 8556 26480
rect 8598 26440 8638 26480
rect 8680 26440 8720 26480
rect 12352 26440 12392 26480
rect 12434 26440 12474 26480
rect 12516 26440 12556 26480
rect 12598 26440 12638 26480
rect 12680 26440 12720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 20352 26440 20392 26480
rect 20434 26440 20474 26480
rect 20516 26440 20556 26480
rect 20598 26440 20638 26480
rect 20680 26440 20720 26480
rect 24352 26440 24392 26480
rect 24434 26440 24474 26480
rect 24516 26440 24556 26480
rect 24598 26440 24638 26480
rect 24680 26440 24720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 32352 26440 32392 26480
rect 32434 26440 32474 26480
rect 32516 26440 32556 26480
rect 32598 26440 32638 26480
rect 32680 26440 32720 26480
rect 36352 26440 36392 26480
rect 36434 26440 36474 26480
rect 36516 26440 36556 26480
rect 36598 26440 36638 26480
rect 36680 26440 36720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 44352 26440 44392 26480
rect 44434 26440 44474 26480
rect 44516 26440 44556 26480
rect 44598 26440 44638 26480
rect 44680 26440 44720 26480
rect 48352 26440 48392 26480
rect 48434 26440 48474 26480
rect 48516 26440 48556 26480
rect 48598 26440 48638 26480
rect 48680 26440 48720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 56352 26440 56392 26480
rect 56434 26440 56474 26480
rect 56516 26440 56556 26480
rect 56598 26440 56638 26480
rect 56680 26440 56720 26480
rect 60352 26440 60392 26480
rect 60434 26440 60474 26480
rect 60516 26440 60556 26480
rect 60598 26440 60638 26480
rect 60680 26440 60720 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 68352 26440 68392 26480
rect 68434 26440 68474 26480
rect 68516 26440 68556 26480
rect 68598 26440 68638 26480
rect 68680 26440 68720 26480
rect 71788 26020 71828 26060
rect 71884 25936 71924 25976
rect 72460 25852 72500 25892
rect 94924 25768 94964 25808
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 7112 25684 7152 25724
rect 7194 25684 7234 25724
rect 7276 25684 7316 25724
rect 7358 25684 7398 25724
rect 7440 25684 7480 25724
rect 11112 25684 11152 25724
rect 11194 25684 11234 25724
rect 11276 25684 11316 25724
rect 11358 25684 11398 25724
rect 11440 25684 11480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 19112 25684 19152 25724
rect 19194 25684 19234 25724
rect 19276 25684 19316 25724
rect 19358 25684 19398 25724
rect 19440 25684 19480 25724
rect 23112 25684 23152 25724
rect 23194 25684 23234 25724
rect 23276 25684 23316 25724
rect 23358 25684 23398 25724
rect 23440 25684 23480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 31112 25684 31152 25724
rect 31194 25684 31234 25724
rect 31276 25684 31316 25724
rect 31358 25684 31398 25724
rect 31440 25684 31480 25724
rect 35112 25684 35152 25724
rect 35194 25684 35234 25724
rect 35276 25684 35316 25724
rect 35358 25684 35398 25724
rect 35440 25684 35480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 43112 25684 43152 25724
rect 43194 25684 43234 25724
rect 43276 25684 43316 25724
rect 43358 25684 43398 25724
rect 43440 25684 43480 25724
rect 47112 25684 47152 25724
rect 47194 25684 47234 25724
rect 47276 25684 47316 25724
rect 47358 25684 47398 25724
rect 47440 25684 47480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 55112 25684 55152 25724
rect 55194 25684 55234 25724
rect 55276 25684 55316 25724
rect 55358 25684 55398 25724
rect 55440 25684 55480 25724
rect 59112 25684 59152 25724
rect 59194 25684 59234 25724
rect 59276 25684 59316 25724
rect 59358 25684 59398 25724
rect 59440 25684 59480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 67112 25684 67152 25724
rect 67194 25684 67234 25724
rect 67276 25684 67316 25724
rect 67358 25684 67398 25724
rect 67440 25684 67480 25724
rect 95020 25684 95060 25724
rect 72940 25600 72980 25640
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 8352 24928 8392 24968
rect 8434 24928 8474 24968
rect 8516 24928 8556 24968
rect 8598 24928 8638 24968
rect 8680 24928 8720 24968
rect 12352 24928 12392 24968
rect 12434 24928 12474 24968
rect 12516 24928 12556 24968
rect 12598 24928 12638 24968
rect 12680 24928 12720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 20352 24928 20392 24968
rect 20434 24928 20474 24968
rect 20516 24928 20556 24968
rect 20598 24928 20638 24968
rect 20680 24928 20720 24968
rect 24352 24928 24392 24968
rect 24434 24928 24474 24968
rect 24516 24928 24556 24968
rect 24598 24928 24638 24968
rect 24680 24928 24720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 32352 24928 32392 24968
rect 32434 24928 32474 24968
rect 32516 24928 32556 24968
rect 32598 24928 32638 24968
rect 32680 24928 32720 24968
rect 36352 24928 36392 24968
rect 36434 24928 36474 24968
rect 36516 24928 36556 24968
rect 36598 24928 36638 24968
rect 36680 24928 36720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 44352 24928 44392 24968
rect 44434 24928 44474 24968
rect 44516 24928 44556 24968
rect 44598 24928 44638 24968
rect 44680 24928 44720 24968
rect 48352 24928 48392 24968
rect 48434 24928 48474 24968
rect 48516 24928 48556 24968
rect 48598 24928 48638 24968
rect 48680 24928 48720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 56352 24928 56392 24968
rect 56434 24928 56474 24968
rect 56516 24928 56556 24968
rect 56598 24928 56638 24968
rect 56680 24928 56720 24968
rect 60352 24928 60392 24968
rect 60434 24928 60474 24968
rect 60516 24928 60556 24968
rect 60598 24928 60638 24968
rect 60680 24928 60720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 68352 24928 68392 24968
rect 68434 24928 68474 24968
rect 68516 24928 68556 24968
rect 68598 24928 68638 24968
rect 68680 24928 68720 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 7112 24172 7152 24212
rect 7194 24172 7234 24212
rect 7276 24172 7316 24212
rect 7358 24172 7398 24212
rect 7440 24172 7480 24212
rect 11112 24172 11152 24212
rect 11194 24172 11234 24212
rect 11276 24172 11316 24212
rect 11358 24172 11398 24212
rect 11440 24172 11480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 19112 24172 19152 24212
rect 19194 24172 19234 24212
rect 19276 24172 19316 24212
rect 19358 24172 19398 24212
rect 19440 24172 19480 24212
rect 23112 24172 23152 24212
rect 23194 24172 23234 24212
rect 23276 24172 23316 24212
rect 23358 24172 23398 24212
rect 23440 24172 23480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 31112 24172 31152 24212
rect 31194 24172 31234 24212
rect 31276 24172 31316 24212
rect 31358 24172 31398 24212
rect 31440 24172 31480 24212
rect 35112 24172 35152 24212
rect 35194 24172 35234 24212
rect 35276 24172 35316 24212
rect 35358 24172 35398 24212
rect 35440 24172 35480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 43112 24172 43152 24212
rect 43194 24172 43234 24212
rect 43276 24172 43316 24212
rect 43358 24172 43398 24212
rect 43440 24172 43480 24212
rect 47112 24172 47152 24212
rect 47194 24172 47234 24212
rect 47276 24172 47316 24212
rect 47358 24172 47398 24212
rect 47440 24172 47480 24212
rect 51112 24172 51152 24212
rect 51194 24172 51234 24212
rect 51276 24172 51316 24212
rect 51358 24172 51398 24212
rect 51440 24172 51480 24212
rect 55112 24172 55152 24212
rect 55194 24172 55234 24212
rect 55276 24172 55316 24212
rect 55358 24172 55398 24212
rect 55440 24172 55480 24212
rect 59112 24172 59152 24212
rect 59194 24172 59234 24212
rect 59276 24172 59316 24212
rect 59358 24172 59398 24212
rect 59440 24172 59480 24212
rect 63112 24172 63152 24212
rect 63194 24172 63234 24212
rect 63276 24172 63316 24212
rect 63358 24172 63398 24212
rect 63440 24172 63480 24212
rect 67112 24172 67152 24212
rect 67194 24172 67234 24212
rect 67276 24172 67316 24212
rect 67358 24172 67398 24212
rect 67440 24172 67480 24212
rect 85420 23920 85460 23960
rect 84268 23752 84308 23792
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 8352 23416 8392 23456
rect 8434 23416 8474 23456
rect 8516 23416 8556 23456
rect 8598 23416 8638 23456
rect 8680 23416 8720 23456
rect 12352 23416 12392 23456
rect 12434 23416 12474 23456
rect 12516 23416 12556 23456
rect 12598 23416 12638 23456
rect 12680 23416 12720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 20352 23416 20392 23456
rect 20434 23416 20474 23456
rect 20516 23416 20556 23456
rect 20598 23416 20638 23456
rect 20680 23416 20720 23456
rect 24352 23416 24392 23456
rect 24434 23416 24474 23456
rect 24516 23416 24556 23456
rect 24598 23416 24638 23456
rect 24680 23416 24720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 32352 23416 32392 23456
rect 32434 23416 32474 23456
rect 32516 23416 32556 23456
rect 32598 23416 32638 23456
rect 32680 23416 32720 23456
rect 36352 23416 36392 23456
rect 36434 23416 36474 23456
rect 36516 23416 36556 23456
rect 36598 23416 36638 23456
rect 36680 23416 36720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 44352 23416 44392 23456
rect 44434 23416 44474 23456
rect 44516 23416 44556 23456
rect 44598 23416 44638 23456
rect 44680 23416 44720 23456
rect 48352 23416 48392 23456
rect 48434 23416 48474 23456
rect 48516 23416 48556 23456
rect 48598 23416 48638 23456
rect 48680 23416 48720 23456
rect 52352 23416 52392 23456
rect 52434 23416 52474 23456
rect 52516 23416 52556 23456
rect 52598 23416 52638 23456
rect 52680 23416 52720 23456
rect 56352 23416 56392 23456
rect 56434 23416 56474 23456
rect 56516 23416 56556 23456
rect 56598 23416 56638 23456
rect 56680 23416 56720 23456
rect 60352 23416 60392 23456
rect 60434 23416 60474 23456
rect 60516 23416 60556 23456
rect 60598 23416 60638 23456
rect 60680 23416 60720 23456
rect 64352 23416 64392 23456
rect 64434 23416 64474 23456
rect 64516 23416 64556 23456
rect 64598 23416 64638 23456
rect 64680 23416 64720 23456
rect 68352 23416 68392 23456
rect 68434 23416 68474 23456
rect 68516 23416 68556 23456
rect 68598 23416 68638 23456
rect 68680 23416 68720 23456
rect 72352 23416 72392 23456
rect 72434 23416 72474 23456
rect 72516 23416 72556 23456
rect 72598 23416 72638 23456
rect 72680 23416 72720 23456
rect 76352 23416 76392 23456
rect 76434 23416 76474 23456
rect 76516 23416 76556 23456
rect 76598 23416 76638 23456
rect 76680 23416 76720 23456
rect 80352 23416 80392 23456
rect 80434 23416 80474 23456
rect 80516 23416 80556 23456
rect 80598 23416 80638 23456
rect 80680 23416 80720 23456
rect 84352 23416 84392 23456
rect 84434 23416 84474 23456
rect 84516 23416 84556 23456
rect 84598 23416 84638 23456
rect 84680 23416 84720 23456
rect 83596 23248 83636 23288
rect 88352 23416 88392 23456
rect 88434 23416 88474 23456
rect 88516 23416 88556 23456
rect 88598 23416 88638 23456
rect 88680 23416 88720 23456
rect 92352 23416 92392 23456
rect 92434 23416 92474 23456
rect 92516 23416 92556 23456
rect 92598 23416 92638 23456
rect 92680 23416 92720 23456
rect 96352 23416 96392 23456
rect 96434 23416 96474 23456
rect 96516 23416 96556 23456
rect 96598 23416 96638 23456
rect 96680 23416 96720 23456
rect 86668 23080 86708 23120
rect 87532 22828 87572 22868
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 7112 22660 7152 22700
rect 7194 22660 7234 22700
rect 7276 22660 7316 22700
rect 7358 22660 7398 22700
rect 7440 22660 7480 22700
rect 11112 22660 11152 22700
rect 11194 22660 11234 22700
rect 11276 22660 11316 22700
rect 11358 22660 11398 22700
rect 11440 22660 11480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 19112 22660 19152 22700
rect 19194 22660 19234 22700
rect 19276 22660 19316 22700
rect 19358 22660 19398 22700
rect 19440 22660 19480 22700
rect 23112 22660 23152 22700
rect 23194 22660 23234 22700
rect 23276 22660 23316 22700
rect 23358 22660 23398 22700
rect 23440 22660 23480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 31112 22660 31152 22700
rect 31194 22660 31234 22700
rect 31276 22660 31316 22700
rect 31358 22660 31398 22700
rect 31440 22660 31480 22700
rect 35112 22660 35152 22700
rect 35194 22660 35234 22700
rect 35276 22660 35316 22700
rect 35358 22660 35398 22700
rect 35440 22660 35480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 43112 22660 43152 22700
rect 43194 22660 43234 22700
rect 43276 22660 43316 22700
rect 43358 22660 43398 22700
rect 43440 22660 43480 22700
rect 47112 22660 47152 22700
rect 47194 22660 47234 22700
rect 47276 22660 47316 22700
rect 47358 22660 47398 22700
rect 47440 22660 47480 22700
rect 51112 22660 51152 22700
rect 51194 22660 51234 22700
rect 51276 22660 51316 22700
rect 51358 22660 51398 22700
rect 51440 22660 51480 22700
rect 55112 22660 55152 22700
rect 55194 22660 55234 22700
rect 55276 22660 55316 22700
rect 55358 22660 55398 22700
rect 55440 22660 55480 22700
rect 59112 22660 59152 22700
rect 59194 22660 59234 22700
rect 59276 22660 59316 22700
rect 59358 22660 59398 22700
rect 59440 22660 59480 22700
rect 63112 22660 63152 22700
rect 63194 22660 63234 22700
rect 63276 22660 63316 22700
rect 63358 22660 63398 22700
rect 63440 22660 63480 22700
rect 67112 22660 67152 22700
rect 67194 22660 67234 22700
rect 67276 22660 67316 22700
rect 67358 22660 67398 22700
rect 67440 22660 67480 22700
rect 71112 22660 71152 22700
rect 71194 22660 71234 22700
rect 71276 22660 71316 22700
rect 71358 22660 71398 22700
rect 71440 22660 71480 22700
rect 75112 22660 75152 22700
rect 75194 22660 75234 22700
rect 75276 22660 75316 22700
rect 75358 22660 75398 22700
rect 75440 22660 75480 22700
rect 79112 22660 79152 22700
rect 79194 22660 79234 22700
rect 79276 22660 79316 22700
rect 79358 22660 79398 22700
rect 79440 22660 79480 22700
rect 83112 22660 83152 22700
rect 83194 22660 83234 22700
rect 83276 22660 83316 22700
rect 83358 22660 83398 22700
rect 83440 22660 83480 22700
rect 87112 22660 87152 22700
rect 87194 22660 87234 22700
rect 87276 22660 87316 22700
rect 87358 22660 87398 22700
rect 87440 22660 87480 22700
rect 91112 22660 91152 22700
rect 91194 22660 91234 22700
rect 91276 22660 91316 22700
rect 91358 22660 91398 22700
rect 91440 22660 91480 22700
rect 95112 22660 95152 22700
rect 95194 22660 95234 22700
rect 95276 22660 95316 22700
rect 95358 22660 95398 22700
rect 95440 22660 95480 22700
rect 99112 22660 99152 22700
rect 99194 22660 99234 22700
rect 99276 22660 99316 22700
rect 99358 22660 99398 22700
rect 99440 22660 99480 22700
rect 85420 22492 85460 22532
rect 94924 22408 94964 22448
rect 83596 22324 83636 22364
rect 87532 22156 87572 22196
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 8352 21904 8392 21944
rect 8434 21904 8474 21944
rect 8516 21904 8556 21944
rect 8598 21904 8638 21944
rect 8680 21904 8720 21944
rect 12352 21904 12392 21944
rect 12434 21904 12474 21944
rect 12516 21904 12556 21944
rect 12598 21904 12638 21944
rect 12680 21904 12720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 20352 21904 20392 21944
rect 20434 21904 20474 21944
rect 20516 21904 20556 21944
rect 20598 21904 20638 21944
rect 20680 21904 20720 21944
rect 24352 21904 24392 21944
rect 24434 21904 24474 21944
rect 24516 21904 24556 21944
rect 24598 21904 24638 21944
rect 24680 21904 24720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 32352 21904 32392 21944
rect 32434 21904 32474 21944
rect 32516 21904 32556 21944
rect 32598 21904 32638 21944
rect 32680 21904 32720 21944
rect 36352 21904 36392 21944
rect 36434 21904 36474 21944
rect 36516 21904 36556 21944
rect 36598 21904 36638 21944
rect 36680 21904 36720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 44352 21904 44392 21944
rect 44434 21904 44474 21944
rect 44516 21904 44556 21944
rect 44598 21904 44638 21944
rect 44680 21904 44720 21944
rect 48352 21904 48392 21944
rect 48434 21904 48474 21944
rect 48516 21904 48556 21944
rect 48598 21904 48638 21944
rect 48680 21904 48720 21944
rect 52352 21904 52392 21944
rect 52434 21904 52474 21944
rect 52516 21904 52556 21944
rect 52598 21904 52638 21944
rect 52680 21904 52720 21944
rect 56352 21904 56392 21944
rect 56434 21904 56474 21944
rect 56516 21904 56556 21944
rect 56598 21904 56638 21944
rect 56680 21904 56720 21944
rect 60352 21904 60392 21944
rect 60434 21904 60474 21944
rect 60516 21904 60556 21944
rect 60598 21904 60638 21944
rect 60680 21904 60720 21944
rect 64352 21904 64392 21944
rect 64434 21904 64474 21944
rect 64516 21904 64556 21944
rect 64598 21904 64638 21944
rect 64680 21904 64720 21944
rect 68352 21904 68392 21944
rect 68434 21904 68474 21944
rect 68516 21904 68556 21944
rect 68598 21904 68638 21944
rect 68680 21904 68720 21944
rect 72352 21904 72392 21944
rect 72434 21904 72474 21944
rect 72516 21904 72556 21944
rect 72598 21904 72638 21944
rect 72680 21904 72720 21944
rect 76352 21904 76392 21944
rect 76434 21904 76474 21944
rect 76516 21904 76556 21944
rect 76598 21904 76638 21944
rect 76680 21904 76720 21944
rect 80352 21904 80392 21944
rect 80434 21904 80474 21944
rect 80516 21904 80556 21944
rect 80598 21904 80638 21944
rect 80680 21904 80720 21944
rect 84352 21904 84392 21944
rect 84434 21904 84474 21944
rect 84516 21904 84556 21944
rect 84598 21904 84638 21944
rect 84680 21904 84720 21944
rect 88352 21904 88392 21944
rect 88434 21904 88474 21944
rect 88516 21904 88556 21944
rect 88598 21904 88638 21944
rect 88680 21904 88720 21944
rect 92352 21904 92392 21944
rect 92434 21904 92474 21944
rect 92516 21904 92556 21944
rect 92598 21904 92638 21944
rect 92680 21904 92720 21944
rect 96352 21904 96392 21944
rect 96434 21904 96474 21944
rect 96516 21904 96556 21944
rect 96598 21904 96638 21944
rect 96680 21904 96720 21944
rect 84268 21736 84308 21776
rect 95020 21736 95060 21776
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 7112 21148 7152 21188
rect 7194 21148 7234 21188
rect 7276 21148 7316 21188
rect 7358 21148 7398 21188
rect 7440 21148 7480 21188
rect 11112 21148 11152 21188
rect 11194 21148 11234 21188
rect 11276 21148 11316 21188
rect 11358 21148 11398 21188
rect 11440 21148 11480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 19112 21148 19152 21188
rect 19194 21148 19234 21188
rect 19276 21148 19316 21188
rect 19358 21148 19398 21188
rect 19440 21148 19480 21188
rect 23112 21148 23152 21188
rect 23194 21148 23234 21188
rect 23276 21148 23316 21188
rect 23358 21148 23398 21188
rect 23440 21148 23480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 31112 21148 31152 21188
rect 31194 21148 31234 21188
rect 31276 21148 31316 21188
rect 31358 21148 31398 21188
rect 31440 21148 31480 21188
rect 35112 21148 35152 21188
rect 35194 21148 35234 21188
rect 35276 21148 35316 21188
rect 35358 21148 35398 21188
rect 35440 21148 35480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 43112 21148 43152 21188
rect 43194 21148 43234 21188
rect 43276 21148 43316 21188
rect 43358 21148 43398 21188
rect 43440 21148 43480 21188
rect 47112 21148 47152 21188
rect 47194 21148 47234 21188
rect 47276 21148 47316 21188
rect 47358 21148 47398 21188
rect 47440 21148 47480 21188
rect 51112 21148 51152 21188
rect 51194 21148 51234 21188
rect 51276 21148 51316 21188
rect 51358 21148 51398 21188
rect 51440 21148 51480 21188
rect 55112 21148 55152 21188
rect 55194 21148 55234 21188
rect 55276 21148 55316 21188
rect 55358 21148 55398 21188
rect 55440 21148 55480 21188
rect 59112 21148 59152 21188
rect 59194 21148 59234 21188
rect 59276 21148 59316 21188
rect 59358 21148 59398 21188
rect 59440 21148 59480 21188
rect 63112 21148 63152 21188
rect 63194 21148 63234 21188
rect 63276 21148 63316 21188
rect 63358 21148 63398 21188
rect 63440 21148 63480 21188
rect 67112 21148 67152 21188
rect 67194 21148 67234 21188
rect 67276 21148 67316 21188
rect 67358 21148 67398 21188
rect 67440 21148 67480 21188
rect 71112 21148 71152 21188
rect 71194 21148 71234 21188
rect 71276 21148 71316 21188
rect 71358 21148 71398 21188
rect 71440 21148 71480 21188
rect 75112 21148 75152 21188
rect 75194 21148 75234 21188
rect 75276 21148 75316 21188
rect 75358 21148 75398 21188
rect 75440 21148 75480 21188
rect 79112 21148 79152 21188
rect 79194 21148 79234 21188
rect 79276 21148 79316 21188
rect 79358 21148 79398 21188
rect 79440 21148 79480 21188
rect 83112 21148 83152 21188
rect 83194 21148 83234 21188
rect 83276 21148 83316 21188
rect 83358 21148 83398 21188
rect 83440 21148 83480 21188
rect 87112 21148 87152 21188
rect 87194 21148 87234 21188
rect 87276 21148 87316 21188
rect 87358 21148 87398 21188
rect 87440 21148 87480 21188
rect 91112 21148 91152 21188
rect 91194 21148 91234 21188
rect 91276 21148 91316 21188
rect 91358 21148 91398 21188
rect 91440 21148 91480 21188
rect 95112 21148 95152 21188
rect 95194 21148 95234 21188
rect 95276 21148 95316 21188
rect 95358 21148 95398 21188
rect 95440 21148 95480 21188
rect 99112 21148 99152 21188
rect 99194 21148 99234 21188
rect 99276 21148 99316 21188
rect 99358 21148 99398 21188
rect 99440 21148 99480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 8352 20392 8392 20432
rect 8434 20392 8474 20432
rect 8516 20392 8556 20432
rect 8598 20392 8638 20432
rect 8680 20392 8720 20432
rect 12352 20392 12392 20432
rect 12434 20392 12474 20432
rect 12516 20392 12556 20432
rect 12598 20392 12638 20432
rect 12680 20392 12720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 20352 20392 20392 20432
rect 20434 20392 20474 20432
rect 20516 20392 20556 20432
rect 20598 20392 20638 20432
rect 20680 20392 20720 20432
rect 24352 20392 24392 20432
rect 24434 20392 24474 20432
rect 24516 20392 24556 20432
rect 24598 20392 24638 20432
rect 24680 20392 24720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 32352 20392 32392 20432
rect 32434 20392 32474 20432
rect 32516 20392 32556 20432
rect 32598 20392 32638 20432
rect 32680 20392 32720 20432
rect 36352 20392 36392 20432
rect 36434 20392 36474 20432
rect 36516 20392 36556 20432
rect 36598 20392 36638 20432
rect 36680 20392 36720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 44352 20392 44392 20432
rect 44434 20392 44474 20432
rect 44516 20392 44556 20432
rect 44598 20392 44638 20432
rect 44680 20392 44720 20432
rect 48352 20392 48392 20432
rect 48434 20392 48474 20432
rect 48516 20392 48556 20432
rect 48598 20392 48638 20432
rect 48680 20392 48720 20432
rect 52352 20392 52392 20432
rect 52434 20392 52474 20432
rect 52516 20392 52556 20432
rect 52598 20392 52638 20432
rect 52680 20392 52720 20432
rect 56352 20392 56392 20432
rect 56434 20392 56474 20432
rect 56516 20392 56556 20432
rect 56598 20392 56638 20432
rect 56680 20392 56720 20432
rect 60352 20392 60392 20432
rect 60434 20392 60474 20432
rect 60516 20392 60556 20432
rect 60598 20392 60638 20432
rect 60680 20392 60720 20432
rect 64352 20392 64392 20432
rect 64434 20392 64474 20432
rect 64516 20392 64556 20432
rect 64598 20392 64638 20432
rect 64680 20392 64720 20432
rect 68352 20392 68392 20432
rect 68434 20392 68474 20432
rect 68516 20392 68556 20432
rect 68598 20392 68638 20432
rect 68680 20392 68720 20432
rect 72352 20392 72392 20432
rect 72434 20392 72474 20432
rect 72516 20392 72556 20432
rect 72598 20392 72638 20432
rect 72680 20392 72720 20432
rect 76352 20392 76392 20432
rect 76434 20392 76474 20432
rect 76516 20392 76556 20432
rect 76598 20392 76638 20432
rect 76680 20392 76720 20432
rect 80352 20392 80392 20432
rect 80434 20392 80474 20432
rect 80516 20392 80556 20432
rect 80598 20392 80638 20432
rect 80680 20392 80720 20432
rect 84352 20392 84392 20432
rect 84434 20392 84474 20432
rect 84516 20392 84556 20432
rect 84598 20392 84638 20432
rect 84680 20392 84720 20432
rect 88352 20392 88392 20432
rect 88434 20392 88474 20432
rect 88516 20392 88556 20432
rect 88598 20392 88638 20432
rect 88680 20392 88720 20432
rect 92352 20392 92392 20432
rect 92434 20392 92474 20432
rect 92516 20392 92556 20432
rect 92598 20392 92638 20432
rect 92680 20392 92720 20432
rect 96352 20392 96392 20432
rect 96434 20392 96474 20432
rect 96516 20392 96556 20432
rect 96598 20392 96638 20432
rect 96680 20392 96720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 7112 19636 7152 19676
rect 7194 19636 7234 19676
rect 7276 19636 7316 19676
rect 7358 19636 7398 19676
rect 7440 19636 7480 19676
rect 11112 19636 11152 19676
rect 11194 19636 11234 19676
rect 11276 19636 11316 19676
rect 11358 19636 11398 19676
rect 11440 19636 11480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 19112 19636 19152 19676
rect 19194 19636 19234 19676
rect 19276 19636 19316 19676
rect 19358 19636 19398 19676
rect 19440 19636 19480 19676
rect 23112 19636 23152 19676
rect 23194 19636 23234 19676
rect 23276 19636 23316 19676
rect 23358 19636 23398 19676
rect 23440 19636 23480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 31112 19636 31152 19676
rect 31194 19636 31234 19676
rect 31276 19636 31316 19676
rect 31358 19636 31398 19676
rect 31440 19636 31480 19676
rect 35112 19636 35152 19676
rect 35194 19636 35234 19676
rect 35276 19636 35316 19676
rect 35358 19636 35398 19676
rect 35440 19636 35480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 43112 19636 43152 19676
rect 43194 19636 43234 19676
rect 43276 19636 43316 19676
rect 43358 19636 43398 19676
rect 43440 19636 43480 19676
rect 47112 19636 47152 19676
rect 47194 19636 47234 19676
rect 47276 19636 47316 19676
rect 47358 19636 47398 19676
rect 47440 19636 47480 19676
rect 51112 19636 51152 19676
rect 51194 19636 51234 19676
rect 51276 19636 51316 19676
rect 51358 19636 51398 19676
rect 51440 19636 51480 19676
rect 55112 19636 55152 19676
rect 55194 19636 55234 19676
rect 55276 19636 55316 19676
rect 55358 19636 55398 19676
rect 55440 19636 55480 19676
rect 59112 19636 59152 19676
rect 59194 19636 59234 19676
rect 59276 19636 59316 19676
rect 59358 19636 59398 19676
rect 59440 19636 59480 19676
rect 63112 19636 63152 19676
rect 63194 19636 63234 19676
rect 63276 19636 63316 19676
rect 63358 19636 63398 19676
rect 63440 19636 63480 19676
rect 67112 19636 67152 19676
rect 67194 19636 67234 19676
rect 67276 19636 67316 19676
rect 67358 19636 67398 19676
rect 67440 19636 67480 19676
rect 71112 19636 71152 19676
rect 71194 19636 71234 19676
rect 71276 19636 71316 19676
rect 71358 19636 71398 19676
rect 71440 19636 71480 19676
rect 75112 19636 75152 19676
rect 75194 19636 75234 19676
rect 75276 19636 75316 19676
rect 75358 19636 75398 19676
rect 75440 19636 75480 19676
rect 79112 19636 79152 19676
rect 79194 19636 79234 19676
rect 79276 19636 79316 19676
rect 79358 19636 79398 19676
rect 79440 19636 79480 19676
rect 83112 19636 83152 19676
rect 83194 19636 83234 19676
rect 83276 19636 83316 19676
rect 83358 19636 83398 19676
rect 83440 19636 83480 19676
rect 87112 19636 87152 19676
rect 87194 19636 87234 19676
rect 87276 19636 87316 19676
rect 87358 19636 87398 19676
rect 87440 19636 87480 19676
rect 91112 19636 91152 19676
rect 91194 19636 91234 19676
rect 91276 19636 91316 19676
rect 91358 19636 91398 19676
rect 91440 19636 91480 19676
rect 95112 19636 95152 19676
rect 95194 19636 95234 19676
rect 95276 19636 95316 19676
rect 95358 19636 95398 19676
rect 95440 19636 95480 19676
rect 99112 19636 99152 19676
rect 99194 19636 99234 19676
rect 99276 19636 99316 19676
rect 99358 19636 99398 19676
rect 99440 19636 99480 19676
rect 86764 19300 86804 19340
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 8352 18880 8392 18920
rect 8434 18880 8474 18920
rect 8516 18880 8556 18920
rect 8598 18880 8638 18920
rect 8680 18880 8720 18920
rect 12352 18880 12392 18920
rect 12434 18880 12474 18920
rect 12516 18880 12556 18920
rect 12598 18880 12638 18920
rect 12680 18880 12720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 20352 18880 20392 18920
rect 20434 18880 20474 18920
rect 20516 18880 20556 18920
rect 20598 18880 20638 18920
rect 20680 18880 20720 18920
rect 24352 18880 24392 18920
rect 24434 18880 24474 18920
rect 24516 18880 24556 18920
rect 24598 18880 24638 18920
rect 24680 18880 24720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 32352 18880 32392 18920
rect 32434 18880 32474 18920
rect 32516 18880 32556 18920
rect 32598 18880 32638 18920
rect 32680 18880 32720 18920
rect 36352 18880 36392 18920
rect 36434 18880 36474 18920
rect 36516 18880 36556 18920
rect 36598 18880 36638 18920
rect 36680 18880 36720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 44352 18880 44392 18920
rect 44434 18880 44474 18920
rect 44516 18880 44556 18920
rect 44598 18880 44638 18920
rect 44680 18880 44720 18920
rect 48352 18880 48392 18920
rect 48434 18880 48474 18920
rect 48516 18880 48556 18920
rect 48598 18880 48638 18920
rect 48680 18880 48720 18920
rect 52352 18880 52392 18920
rect 52434 18880 52474 18920
rect 52516 18880 52556 18920
rect 52598 18880 52638 18920
rect 52680 18880 52720 18920
rect 56352 18880 56392 18920
rect 56434 18880 56474 18920
rect 56516 18880 56556 18920
rect 56598 18880 56638 18920
rect 56680 18880 56720 18920
rect 60352 18880 60392 18920
rect 60434 18880 60474 18920
rect 60516 18880 60556 18920
rect 60598 18880 60638 18920
rect 60680 18880 60720 18920
rect 64352 18880 64392 18920
rect 64434 18880 64474 18920
rect 64516 18880 64556 18920
rect 64598 18880 64638 18920
rect 64680 18880 64720 18920
rect 68352 18880 68392 18920
rect 68434 18880 68474 18920
rect 68516 18880 68556 18920
rect 68598 18880 68638 18920
rect 68680 18880 68720 18920
rect 72352 18880 72392 18920
rect 72434 18880 72474 18920
rect 72516 18880 72556 18920
rect 72598 18880 72638 18920
rect 72680 18880 72720 18920
rect 76352 18880 76392 18920
rect 76434 18880 76474 18920
rect 76516 18880 76556 18920
rect 76598 18880 76638 18920
rect 76680 18880 76720 18920
rect 80352 18880 80392 18920
rect 80434 18880 80474 18920
rect 80516 18880 80556 18920
rect 80598 18880 80638 18920
rect 80680 18880 80720 18920
rect 84352 18880 84392 18920
rect 84434 18880 84474 18920
rect 84516 18880 84556 18920
rect 84598 18880 84638 18920
rect 84680 18880 84720 18920
rect 88352 18880 88392 18920
rect 88434 18880 88474 18920
rect 88516 18880 88556 18920
rect 88598 18880 88638 18920
rect 88680 18880 88720 18920
rect 92352 18880 92392 18920
rect 92434 18880 92474 18920
rect 92516 18880 92556 18920
rect 92598 18880 92638 18920
rect 92680 18880 92720 18920
rect 96352 18880 96392 18920
rect 96434 18880 96474 18920
rect 96516 18880 96556 18920
rect 96598 18880 96638 18920
rect 96680 18880 96720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 7112 18124 7152 18164
rect 7194 18124 7234 18164
rect 7276 18124 7316 18164
rect 7358 18124 7398 18164
rect 7440 18124 7480 18164
rect 11112 18124 11152 18164
rect 11194 18124 11234 18164
rect 11276 18124 11316 18164
rect 11358 18124 11398 18164
rect 11440 18124 11480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 19112 18124 19152 18164
rect 19194 18124 19234 18164
rect 19276 18124 19316 18164
rect 19358 18124 19398 18164
rect 19440 18124 19480 18164
rect 23112 18124 23152 18164
rect 23194 18124 23234 18164
rect 23276 18124 23316 18164
rect 23358 18124 23398 18164
rect 23440 18124 23480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 31112 18124 31152 18164
rect 31194 18124 31234 18164
rect 31276 18124 31316 18164
rect 31358 18124 31398 18164
rect 31440 18124 31480 18164
rect 35112 18124 35152 18164
rect 35194 18124 35234 18164
rect 35276 18124 35316 18164
rect 35358 18124 35398 18164
rect 35440 18124 35480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 43112 18124 43152 18164
rect 43194 18124 43234 18164
rect 43276 18124 43316 18164
rect 43358 18124 43398 18164
rect 43440 18124 43480 18164
rect 47112 18124 47152 18164
rect 47194 18124 47234 18164
rect 47276 18124 47316 18164
rect 47358 18124 47398 18164
rect 47440 18124 47480 18164
rect 51112 18124 51152 18164
rect 51194 18124 51234 18164
rect 51276 18124 51316 18164
rect 51358 18124 51398 18164
rect 51440 18124 51480 18164
rect 55112 18124 55152 18164
rect 55194 18124 55234 18164
rect 55276 18124 55316 18164
rect 55358 18124 55398 18164
rect 55440 18124 55480 18164
rect 59112 18124 59152 18164
rect 59194 18124 59234 18164
rect 59276 18124 59316 18164
rect 59358 18124 59398 18164
rect 59440 18124 59480 18164
rect 63112 18124 63152 18164
rect 63194 18124 63234 18164
rect 63276 18124 63316 18164
rect 63358 18124 63398 18164
rect 63440 18124 63480 18164
rect 67112 18124 67152 18164
rect 67194 18124 67234 18164
rect 67276 18124 67316 18164
rect 67358 18124 67398 18164
rect 67440 18124 67480 18164
rect 71112 18124 71152 18164
rect 71194 18124 71234 18164
rect 71276 18124 71316 18164
rect 71358 18124 71398 18164
rect 71440 18124 71480 18164
rect 75112 18124 75152 18164
rect 75194 18124 75234 18164
rect 75276 18124 75316 18164
rect 75358 18124 75398 18164
rect 75440 18124 75480 18164
rect 79112 18124 79152 18164
rect 79194 18124 79234 18164
rect 79276 18124 79316 18164
rect 79358 18124 79398 18164
rect 79440 18124 79480 18164
rect 83112 18124 83152 18164
rect 83194 18124 83234 18164
rect 83276 18124 83316 18164
rect 83358 18124 83398 18164
rect 83440 18124 83480 18164
rect 87112 18124 87152 18164
rect 87194 18124 87234 18164
rect 87276 18124 87316 18164
rect 87358 18124 87398 18164
rect 87440 18124 87480 18164
rect 91112 18124 91152 18164
rect 91194 18124 91234 18164
rect 91276 18124 91316 18164
rect 91358 18124 91398 18164
rect 91440 18124 91480 18164
rect 95112 18124 95152 18164
rect 95194 18124 95234 18164
rect 95276 18124 95316 18164
rect 95358 18124 95398 18164
rect 95440 18124 95480 18164
rect 99112 18124 99152 18164
rect 99194 18124 99234 18164
rect 99276 18124 99316 18164
rect 99358 18124 99398 18164
rect 99440 18124 99480 18164
rect 84268 17536 84308 17576
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 8352 17368 8392 17408
rect 8434 17368 8474 17408
rect 8516 17368 8556 17408
rect 8598 17368 8638 17408
rect 8680 17368 8720 17408
rect 12352 17368 12392 17408
rect 12434 17368 12474 17408
rect 12516 17368 12556 17408
rect 12598 17368 12638 17408
rect 12680 17368 12720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 20352 17368 20392 17408
rect 20434 17368 20474 17408
rect 20516 17368 20556 17408
rect 20598 17368 20638 17408
rect 20680 17368 20720 17408
rect 24352 17368 24392 17408
rect 24434 17368 24474 17408
rect 24516 17368 24556 17408
rect 24598 17368 24638 17408
rect 24680 17368 24720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 32352 17368 32392 17408
rect 32434 17368 32474 17408
rect 32516 17368 32556 17408
rect 32598 17368 32638 17408
rect 32680 17368 32720 17408
rect 36352 17368 36392 17408
rect 36434 17368 36474 17408
rect 36516 17368 36556 17408
rect 36598 17368 36638 17408
rect 36680 17368 36720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 44352 17368 44392 17408
rect 44434 17368 44474 17408
rect 44516 17368 44556 17408
rect 44598 17368 44638 17408
rect 44680 17368 44720 17408
rect 48352 17368 48392 17408
rect 48434 17368 48474 17408
rect 48516 17368 48556 17408
rect 48598 17368 48638 17408
rect 48680 17368 48720 17408
rect 52352 17368 52392 17408
rect 52434 17368 52474 17408
rect 52516 17368 52556 17408
rect 52598 17368 52638 17408
rect 52680 17368 52720 17408
rect 56352 17368 56392 17408
rect 56434 17368 56474 17408
rect 56516 17368 56556 17408
rect 56598 17368 56638 17408
rect 56680 17368 56720 17408
rect 60352 17368 60392 17408
rect 60434 17368 60474 17408
rect 60516 17368 60556 17408
rect 60598 17368 60638 17408
rect 60680 17368 60720 17408
rect 64352 17368 64392 17408
rect 64434 17368 64474 17408
rect 64516 17368 64556 17408
rect 64598 17368 64638 17408
rect 64680 17368 64720 17408
rect 68352 17368 68392 17408
rect 68434 17368 68474 17408
rect 68516 17368 68556 17408
rect 68598 17368 68638 17408
rect 68680 17368 68720 17408
rect 72352 17368 72392 17408
rect 72434 17368 72474 17408
rect 72516 17368 72556 17408
rect 72598 17368 72638 17408
rect 72680 17368 72720 17408
rect 76352 17368 76392 17408
rect 76434 17368 76474 17408
rect 76516 17368 76556 17408
rect 76598 17368 76638 17408
rect 76680 17368 76720 17408
rect 80352 17368 80392 17408
rect 80434 17368 80474 17408
rect 80516 17368 80556 17408
rect 80598 17368 80638 17408
rect 80680 17368 80720 17408
rect 84352 17368 84392 17408
rect 84434 17368 84474 17408
rect 84516 17368 84556 17408
rect 84598 17368 84638 17408
rect 84680 17368 84720 17408
rect 88352 17368 88392 17408
rect 88434 17368 88474 17408
rect 88516 17368 88556 17408
rect 88598 17368 88638 17408
rect 88680 17368 88720 17408
rect 92352 17368 92392 17408
rect 92434 17368 92474 17408
rect 92516 17368 92556 17408
rect 92598 17368 92638 17408
rect 92680 17368 92720 17408
rect 96352 17368 96392 17408
rect 96434 17368 96474 17408
rect 96516 17368 96556 17408
rect 96598 17368 96638 17408
rect 96680 17368 96720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 7112 16612 7152 16652
rect 7194 16612 7234 16652
rect 7276 16612 7316 16652
rect 7358 16612 7398 16652
rect 7440 16612 7480 16652
rect 11112 16612 11152 16652
rect 11194 16612 11234 16652
rect 11276 16612 11316 16652
rect 11358 16612 11398 16652
rect 11440 16612 11480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 19112 16612 19152 16652
rect 19194 16612 19234 16652
rect 19276 16612 19316 16652
rect 19358 16612 19398 16652
rect 19440 16612 19480 16652
rect 23112 16612 23152 16652
rect 23194 16612 23234 16652
rect 23276 16612 23316 16652
rect 23358 16612 23398 16652
rect 23440 16612 23480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 31112 16612 31152 16652
rect 31194 16612 31234 16652
rect 31276 16612 31316 16652
rect 31358 16612 31398 16652
rect 31440 16612 31480 16652
rect 35112 16612 35152 16652
rect 35194 16612 35234 16652
rect 35276 16612 35316 16652
rect 35358 16612 35398 16652
rect 35440 16612 35480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 43112 16612 43152 16652
rect 43194 16612 43234 16652
rect 43276 16612 43316 16652
rect 43358 16612 43398 16652
rect 43440 16612 43480 16652
rect 47112 16612 47152 16652
rect 47194 16612 47234 16652
rect 47276 16612 47316 16652
rect 47358 16612 47398 16652
rect 47440 16612 47480 16652
rect 51112 16612 51152 16652
rect 51194 16612 51234 16652
rect 51276 16612 51316 16652
rect 51358 16612 51398 16652
rect 51440 16612 51480 16652
rect 55112 16612 55152 16652
rect 55194 16612 55234 16652
rect 55276 16612 55316 16652
rect 55358 16612 55398 16652
rect 55440 16612 55480 16652
rect 59112 16612 59152 16652
rect 59194 16612 59234 16652
rect 59276 16612 59316 16652
rect 59358 16612 59398 16652
rect 59440 16612 59480 16652
rect 63112 16612 63152 16652
rect 63194 16612 63234 16652
rect 63276 16612 63316 16652
rect 63358 16612 63398 16652
rect 63440 16612 63480 16652
rect 67112 16612 67152 16652
rect 67194 16612 67234 16652
rect 67276 16612 67316 16652
rect 67358 16612 67398 16652
rect 67440 16612 67480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 8352 15856 8392 15896
rect 8434 15856 8474 15896
rect 8516 15856 8556 15896
rect 8598 15856 8638 15896
rect 8680 15856 8720 15896
rect 12352 15856 12392 15896
rect 12434 15856 12474 15896
rect 12516 15856 12556 15896
rect 12598 15856 12638 15896
rect 12680 15856 12720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 20352 15856 20392 15896
rect 20434 15856 20474 15896
rect 20516 15856 20556 15896
rect 20598 15856 20638 15896
rect 20680 15856 20720 15896
rect 24352 15856 24392 15896
rect 24434 15856 24474 15896
rect 24516 15856 24556 15896
rect 24598 15856 24638 15896
rect 24680 15856 24720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 32352 15856 32392 15896
rect 32434 15856 32474 15896
rect 32516 15856 32556 15896
rect 32598 15856 32638 15896
rect 32680 15856 32720 15896
rect 36352 15856 36392 15896
rect 36434 15856 36474 15896
rect 36516 15856 36556 15896
rect 36598 15856 36638 15896
rect 36680 15856 36720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 44352 15856 44392 15896
rect 44434 15856 44474 15896
rect 44516 15856 44556 15896
rect 44598 15856 44638 15896
rect 44680 15856 44720 15896
rect 48352 15856 48392 15896
rect 48434 15856 48474 15896
rect 48516 15856 48556 15896
rect 48598 15856 48638 15896
rect 48680 15856 48720 15896
rect 52352 15856 52392 15896
rect 52434 15856 52474 15896
rect 52516 15856 52556 15896
rect 52598 15856 52638 15896
rect 52680 15856 52720 15896
rect 56352 15856 56392 15896
rect 56434 15856 56474 15896
rect 56516 15856 56556 15896
rect 56598 15856 56638 15896
rect 56680 15856 56720 15896
rect 60352 15856 60392 15896
rect 60434 15856 60474 15896
rect 60516 15856 60556 15896
rect 60598 15856 60638 15896
rect 60680 15856 60720 15896
rect 64352 15856 64392 15896
rect 64434 15856 64474 15896
rect 64516 15856 64556 15896
rect 64598 15856 64638 15896
rect 64680 15856 64720 15896
rect 68352 15856 68392 15896
rect 68434 15856 68474 15896
rect 68516 15856 68556 15896
rect 68598 15856 68638 15896
rect 68680 15856 68720 15896
rect 71788 15520 71828 15560
rect 84268 15520 84308 15560
rect 98860 15436 98900 15476
rect 71884 15352 71924 15392
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 7112 15100 7152 15140
rect 7194 15100 7234 15140
rect 7276 15100 7316 15140
rect 7358 15100 7398 15140
rect 7440 15100 7480 15140
rect 11112 15100 11152 15140
rect 11194 15100 11234 15140
rect 11276 15100 11316 15140
rect 11358 15100 11398 15140
rect 11440 15100 11480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 19112 15100 19152 15140
rect 19194 15100 19234 15140
rect 19276 15100 19316 15140
rect 19358 15100 19398 15140
rect 19440 15100 19480 15140
rect 23112 15100 23152 15140
rect 23194 15100 23234 15140
rect 23276 15100 23316 15140
rect 23358 15100 23398 15140
rect 23440 15100 23480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 31112 15100 31152 15140
rect 31194 15100 31234 15140
rect 31276 15100 31316 15140
rect 31358 15100 31398 15140
rect 31440 15100 31480 15140
rect 35112 15100 35152 15140
rect 35194 15100 35234 15140
rect 35276 15100 35316 15140
rect 35358 15100 35398 15140
rect 35440 15100 35480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 43112 15100 43152 15140
rect 43194 15100 43234 15140
rect 43276 15100 43316 15140
rect 43358 15100 43398 15140
rect 43440 15100 43480 15140
rect 47112 15100 47152 15140
rect 47194 15100 47234 15140
rect 47276 15100 47316 15140
rect 47358 15100 47398 15140
rect 47440 15100 47480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 55112 15100 55152 15140
rect 55194 15100 55234 15140
rect 55276 15100 55316 15140
rect 55358 15100 55398 15140
rect 55440 15100 55480 15140
rect 59112 15100 59152 15140
rect 59194 15100 59234 15140
rect 59276 15100 59316 15140
rect 59358 15100 59398 15140
rect 59440 15100 59480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 67112 15100 67152 15140
rect 67194 15100 67234 15140
rect 67276 15100 67316 15140
rect 67358 15100 67398 15140
rect 67440 15100 67480 15140
rect 71788 15016 71828 15056
rect 71884 14848 71924 14888
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 8352 14344 8392 14384
rect 8434 14344 8474 14384
rect 8516 14344 8556 14384
rect 8598 14344 8638 14384
rect 8680 14344 8720 14384
rect 12352 14344 12392 14384
rect 12434 14344 12474 14384
rect 12516 14344 12556 14384
rect 12598 14344 12638 14384
rect 12680 14344 12720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 20352 14344 20392 14384
rect 20434 14344 20474 14384
rect 20516 14344 20556 14384
rect 20598 14344 20638 14384
rect 20680 14344 20720 14384
rect 24352 14344 24392 14384
rect 24434 14344 24474 14384
rect 24516 14344 24556 14384
rect 24598 14344 24638 14384
rect 24680 14344 24720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 32352 14344 32392 14384
rect 32434 14344 32474 14384
rect 32516 14344 32556 14384
rect 32598 14344 32638 14384
rect 32680 14344 32720 14384
rect 36352 14344 36392 14384
rect 36434 14344 36474 14384
rect 36516 14344 36556 14384
rect 36598 14344 36638 14384
rect 36680 14344 36720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 44352 14344 44392 14384
rect 44434 14344 44474 14384
rect 44516 14344 44556 14384
rect 44598 14344 44638 14384
rect 44680 14344 44720 14384
rect 48352 14344 48392 14384
rect 48434 14344 48474 14384
rect 48516 14344 48556 14384
rect 48598 14344 48638 14384
rect 48680 14344 48720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 56352 14344 56392 14384
rect 56434 14344 56474 14384
rect 56516 14344 56556 14384
rect 56598 14344 56638 14384
rect 56680 14344 56720 14384
rect 60352 14344 60392 14384
rect 60434 14344 60474 14384
rect 60516 14344 60556 14384
rect 60598 14344 60638 14384
rect 60680 14344 60720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 68352 14344 68392 14384
rect 68434 14344 68474 14384
rect 68516 14344 68556 14384
rect 68598 14344 68638 14384
rect 68680 14344 68720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 7112 13588 7152 13628
rect 7194 13588 7234 13628
rect 7276 13588 7316 13628
rect 7358 13588 7398 13628
rect 7440 13588 7480 13628
rect 11112 13588 11152 13628
rect 11194 13588 11234 13628
rect 11276 13588 11316 13628
rect 11358 13588 11398 13628
rect 11440 13588 11480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 19112 13588 19152 13628
rect 19194 13588 19234 13628
rect 19276 13588 19316 13628
rect 19358 13588 19398 13628
rect 19440 13588 19480 13628
rect 23112 13588 23152 13628
rect 23194 13588 23234 13628
rect 23276 13588 23316 13628
rect 23358 13588 23398 13628
rect 23440 13588 23480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 31112 13588 31152 13628
rect 31194 13588 31234 13628
rect 31276 13588 31316 13628
rect 31358 13588 31398 13628
rect 31440 13588 31480 13628
rect 35112 13588 35152 13628
rect 35194 13588 35234 13628
rect 35276 13588 35316 13628
rect 35358 13588 35398 13628
rect 35440 13588 35480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 43112 13588 43152 13628
rect 43194 13588 43234 13628
rect 43276 13588 43316 13628
rect 43358 13588 43398 13628
rect 43440 13588 43480 13628
rect 47112 13588 47152 13628
rect 47194 13588 47234 13628
rect 47276 13588 47316 13628
rect 47358 13588 47398 13628
rect 47440 13588 47480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 55112 13588 55152 13628
rect 55194 13588 55234 13628
rect 55276 13588 55316 13628
rect 55358 13588 55398 13628
rect 55440 13588 55480 13628
rect 59112 13588 59152 13628
rect 59194 13588 59234 13628
rect 59276 13588 59316 13628
rect 59358 13588 59398 13628
rect 59440 13588 59480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 67112 13588 67152 13628
rect 67194 13588 67234 13628
rect 67276 13588 67316 13628
rect 67358 13588 67398 13628
rect 67440 13588 67480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 8352 12832 8392 12872
rect 8434 12832 8474 12872
rect 8516 12832 8556 12872
rect 8598 12832 8638 12872
rect 8680 12832 8720 12872
rect 12352 12832 12392 12872
rect 12434 12832 12474 12872
rect 12516 12832 12556 12872
rect 12598 12832 12638 12872
rect 12680 12832 12720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 20352 12832 20392 12872
rect 20434 12832 20474 12872
rect 20516 12832 20556 12872
rect 20598 12832 20638 12872
rect 20680 12832 20720 12872
rect 24352 12832 24392 12872
rect 24434 12832 24474 12872
rect 24516 12832 24556 12872
rect 24598 12832 24638 12872
rect 24680 12832 24720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 32352 12832 32392 12872
rect 32434 12832 32474 12872
rect 32516 12832 32556 12872
rect 32598 12832 32638 12872
rect 32680 12832 32720 12872
rect 36352 12832 36392 12872
rect 36434 12832 36474 12872
rect 36516 12832 36556 12872
rect 36598 12832 36638 12872
rect 36680 12832 36720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 44352 12832 44392 12872
rect 44434 12832 44474 12872
rect 44516 12832 44556 12872
rect 44598 12832 44638 12872
rect 44680 12832 44720 12872
rect 48352 12832 48392 12872
rect 48434 12832 48474 12872
rect 48516 12832 48556 12872
rect 48598 12832 48638 12872
rect 48680 12832 48720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 56352 12832 56392 12872
rect 56434 12832 56474 12872
rect 56516 12832 56556 12872
rect 56598 12832 56638 12872
rect 56680 12832 56720 12872
rect 60352 12832 60392 12872
rect 60434 12832 60474 12872
rect 60516 12832 60556 12872
rect 60598 12832 60638 12872
rect 60680 12832 60720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 68352 12832 68392 12872
rect 68434 12832 68474 12872
rect 68516 12832 68556 12872
rect 68598 12832 68638 12872
rect 68680 12832 68720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 7112 12076 7152 12116
rect 7194 12076 7234 12116
rect 7276 12076 7316 12116
rect 7358 12076 7398 12116
rect 7440 12076 7480 12116
rect 11112 12076 11152 12116
rect 11194 12076 11234 12116
rect 11276 12076 11316 12116
rect 11358 12076 11398 12116
rect 11440 12076 11480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 19112 12076 19152 12116
rect 19194 12076 19234 12116
rect 19276 12076 19316 12116
rect 19358 12076 19398 12116
rect 19440 12076 19480 12116
rect 23112 12076 23152 12116
rect 23194 12076 23234 12116
rect 23276 12076 23316 12116
rect 23358 12076 23398 12116
rect 23440 12076 23480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 31112 12076 31152 12116
rect 31194 12076 31234 12116
rect 31276 12076 31316 12116
rect 31358 12076 31398 12116
rect 31440 12076 31480 12116
rect 35112 12076 35152 12116
rect 35194 12076 35234 12116
rect 35276 12076 35316 12116
rect 35358 12076 35398 12116
rect 35440 12076 35480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 43112 12076 43152 12116
rect 43194 12076 43234 12116
rect 43276 12076 43316 12116
rect 43358 12076 43398 12116
rect 43440 12076 43480 12116
rect 47112 12076 47152 12116
rect 47194 12076 47234 12116
rect 47276 12076 47316 12116
rect 47358 12076 47398 12116
rect 47440 12076 47480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 55112 12076 55152 12116
rect 55194 12076 55234 12116
rect 55276 12076 55316 12116
rect 55358 12076 55398 12116
rect 55440 12076 55480 12116
rect 59112 12076 59152 12116
rect 59194 12076 59234 12116
rect 59276 12076 59316 12116
rect 59358 12076 59398 12116
rect 59440 12076 59480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 67112 12076 67152 12116
rect 67194 12076 67234 12116
rect 67276 12076 67316 12116
rect 67358 12076 67398 12116
rect 67440 12076 67480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 8352 11320 8392 11360
rect 8434 11320 8474 11360
rect 8516 11320 8556 11360
rect 8598 11320 8638 11360
rect 8680 11320 8720 11360
rect 12352 11320 12392 11360
rect 12434 11320 12474 11360
rect 12516 11320 12556 11360
rect 12598 11320 12638 11360
rect 12680 11320 12720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 20352 11320 20392 11360
rect 20434 11320 20474 11360
rect 20516 11320 20556 11360
rect 20598 11320 20638 11360
rect 20680 11320 20720 11360
rect 24352 11320 24392 11360
rect 24434 11320 24474 11360
rect 24516 11320 24556 11360
rect 24598 11320 24638 11360
rect 24680 11320 24720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 32352 11320 32392 11360
rect 32434 11320 32474 11360
rect 32516 11320 32556 11360
rect 32598 11320 32638 11360
rect 32680 11320 32720 11360
rect 36352 11320 36392 11360
rect 36434 11320 36474 11360
rect 36516 11320 36556 11360
rect 36598 11320 36638 11360
rect 36680 11320 36720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 44352 11320 44392 11360
rect 44434 11320 44474 11360
rect 44516 11320 44556 11360
rect 44598 11320 44638 11360
rect 44680 11320 44720 11360
rect 48352 11320 48392 11360
rect 48434 11320 48474 11360
rect 48516 11320 48556 11360
rect 48598 11320 48638 11360
rect 48680 11320 48720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 56352 11320 56392 11360
rect 56434 11320 56474 11360
rect 56516 11320 56556 11360
rect 56598 11320 56638 11360
rect 56680 11320 56720 11360
rect 60352 11320 60392 11360
rect 60434 11320 60474 11360
rect 60516 11320 60556 11360
rect 60598 11320 60638 11360
rect 60680 11320 60720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 68352 11320 68392 11360
rect 68434 11320 68474 11360
rect 68516 11320 68556 11360
rect 68598 11320 68638 11360
rect 68680 11320 68720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 7112 10564 7152 10604
rect 7194 10564 7234 10604
rect 7276 10564 7316 10604
rect 7358 10564 7398 10604
rect 7440 10564 7480 10604
rect 11112 10564 11152 10604
rect 11194 10564 11234 10604
rect 11276 10564 11316 10604
rect 11358 10564 11398 10604
rect 11440 10564 11480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 19112 10564 19152 10604
rect 19194 10564 19234 10604
rect 19276 10564 19316 10604
rect 19358 10564 19398 10604
rect 19440 10564 19480 10604
rect 23112 10564 23152 10604
rect 23194 10564 23234 10604
rect 23276 10564 23316 10604
rect 23358 10564 23398 10604
rect 23440 10564 23480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 31112 10564 31152 10604
rect 31194 10564 31234 10604
rect 31276 10564 31316 10604
rect 31358 10564 31398 10604
rect 31440 10564 31480 10604
rect 35112 10564 35152 10604
rect 35194 10564 35234 10604
rect 35276 10564 35316 10604
rect 35358 10564 35398 10604
rect 35440 10564 35480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 43112 10564 43152 10604
rect 43194 10564 43234 10604
rect 43276 10564 43316 10604
rect 43358 10564 43398 10604
rect 43440 10564 43480 10604
rect 47112 10564 47152 10604
rect 47194 10564 47234 10604
rect 47276 10564 47316 10604
rect 47358 10564 47398 10604
rect 47440 10564 47480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 55112 10564 55152 10604
rect 55194 10564 55234 10604
rect 55276 10564 55316 10604
rect 55358 10564 55398 10604
rect 55440 10564 55480 10604
rect 59112 10564 59152 10604
rect 59194 10564 59234 10604
rect 59276 10564 59316 10604
rect 59358 10564 59398 10604
rect 59440 10564 59480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 67112 10564 67152 10604
rect 67194 10564 67234 10604
rect 67276 10564 67316 10604
rect 67358 10564 67398 10604
rect 67440 10564 67480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 8352 9808 8392 9848
rect 8434 9808 8474 9848
rect 8516 9808 8556 9848
rect 8598 9808 8638 9848
rect 8680 9808 8720 9848
rect 12352 9808 12392 9848
rect 12434 9808 12474 9848
rect 12516 9808 12556 9848
rect 12598 9808 12638 9848
rect 12680 9808 12720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 20352 9808 20392 9848
rect 20434 9808 20474 9848
rect 20516 9808 20556 9848
rect 20598 9808 20638 9848
rect 20680 9808 20720 9848
rect 24352 9808 24392 9848
rect 24434 9808 24474 9848
rect 24516 9808 24556 9848
rect 24598 9808 24638 9848
rect 24680 9808 24720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 32352 9808 32392 9848
rect 32434 9808 32474 9848
rect 32516 9808 32556 9848
rect 32598 9808 32638 9848
rect 32680 9808 32720 9848
rect 36352 9808 36392 9848
rect 36434 9808 36474 9848
rect 36516 9808 36556 9848
rect 36598 9808 36638 9848
rect 36680 9808 36720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 44352 9808 44392 9848
rect 44434 9808 44474 9848
rect 44516 9808 44556 9848
rect 44598 9808 44638 9848
rect 44680 9808 44720 9848
rect 48352 9808 48392 9848
rect 48434 9808 48474 9848
rect 48516 9808 48556 9848
rect 48598 9808 48638 9848
rect 48680 9808 48720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 56352 9808 56392 9848
rect 56434 9808 56474 9848
rect 56516 9808 56556 9848
rect 56598 9808 56638 9848
rect 56680 9808 56720 9848
rect 60352 9808 60392 9848
rect 60434 9808 60474 9848
rect 60516 9808 60556 9848
rect 60598 9808 60638 9848
rect 60680 9808 60720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 68352 9808 68392 9848
rect 68434 9808 68474 9848
rect 68516 9808 68556 9848
rect 68598 9808 68638 9848
rect 68680 9808 68720 9848
rect 80140 9724 80180 9764
rect 83596 9724 83615 9764
rect 83615 9724 83636 9764
rect 89068 9724 89105 9764
rect 89105 9724 89108 9764
rect 98860 9472 98900 9512
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 7112 9052 7152 9092
rect 7194 9052 7234 9092
rect 7276 9052 7316 9092
rect 7358 9052 7398 9092
rect 7440 9052 7480 9092
rect 11112 9052 11152 9092
rect 11194 9052 11234 9092
rect 11276 9052 11316 9092
rect 11358 9052 11398 9092
rect 11440 9052 11480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 19112 9052 19152 9092
rect 19194 9052 19234 9092
rect 19276 9052 19316 9092
rect 19358 9052 19398 9092
rect 19440 9052 19480 9092
rect 23112 9052 23152 9092
rect 23194 9052 23234 9092
rect 23276 9052 23316 9092
rect 23358 9052 23398 9092
rect 23440 9052 23480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 31112 9052 31152 9092
rect 31194 9052 31234 9092
rect 31276 9052 31316 9092
rect 31358 9052 31398 9092
rect 31440 9052 31480 9092
rect 35112 9052 35152 9092
rect 35194 9052 35234 9092
rect 35276 9052 35316 9092
rect 35358 9052 35398 9092
rect 35440 9052 35480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 43112 9052 43152 9092
rect 43194 9052 43234 9092
rect 43276 9052 43316 9092
rect 43358 9052 43398 9092
rect 43440 9052 43480 9092
rect 47112 9052 47152 9092
rect 47194 9052 47234 9092
rect 47276 9052 47316 9092
rect 47358 9052 47398 9092
rect 47440 9052 47480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 55112 9052 55152 9092
rect 55194 9052 55234 9092
rect 55276 9052 55316 9092
rect 55358 9052 55398 9092
rect 55440 9052 55480 9092
rect 59112 9052 59152 9092
rect 59194 9052 59234 9092
rect 59276 9052 59316 9092
rect 59358 9052 59398 9092
rect 59440 9052 59480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 67112 9052 67152 9092
rect 67194 9052 67234 9092
rect 67276 9052 67316 9092
rect 67358 9052 67398 9092
rect 67440 9052 67480 9092
rect 85612 8800 85652 8840
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 8352 8296 8392 8336
rect 8434 8296 8474 8336
rect 8516 8296 8556 8336
rect 8598 8296 8638 8336
rect 8680 8296 8720 8336
rect 12352 8296 12392 8336
rect 12434 8296 12474 8336
rect 12516 8296 12556 8336
rect 12598 8296 12638 8336
rect 12680 8296 12720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 20352 8296 20392 8336
rect 20434 8296 20474 8336
rect 20516 8296 20556 8336
rect 20598 8296 20638 8336
rect 20680 8296 20720 8336
rect 24352 8296 24392 8336
rect 24434 8296 24474 8336
rect 24516 8296 24556 8336
rect 24598 8296 24638 8336
rect 24680 8296 24720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 32352 8296 32392 8336
rect 32434 8296 32474 8336
rect 32516 8296 32556 8336
rect 32598 8296 32638 8336
rect 32680 8296 32720 8336
rect 36352 8296 36392 8336
rect 36434 8296 36474 8336
rect 36516 8296 36556 8336
rect 36598 8296 36638 8336
rect 36680 8296 36720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 44352 8296 44392 8336
rect 44434 8296 44474 8336
rect 44516 8296 44556 8336
rect 44598 8296 44638 8336
rect 44680 8296 44720 8336
rect 48352 8296 48392 8336
rect 48434 8296 48474 8336
rect 48516 8296 48556 8336
rect 48598 8296 48638 8336
rect 48680 8296 48720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 56352 8296 56392 8336
rect 56434 8296 56474 8336
rect 56516 8296 56556 8336
rect 56598 8296 56638 8336
rect 56680 8296 56720 8336
rect 60352 8296 60392 8336
rect 60434 8296 60474 8336
rect 60516 8296 60556 8336
rect 60598 8296 60638 8336
rect 60680 8296 60720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 68352 8296 68392 8336
rect 68434 8296 68474 8336
rect 68516 8296 68556 8336
rect 68598 8296 68638 8336
rect 68680 8296 68720 8336
rect 82924 7876 82964 7916
rect 95596 7792 95636 7832
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 7112 7540 7152 7580
rect 7194 7540 7234 7580
rect 7276 7540 7316 7580
rect 7358 7540 7398 7580
rect 7440 7540 7480 7580
rect 11112 7540 11152 7580
rect 11194 7540 11234 7580
rect 11276 7540 11316 7580
rect 11358 7540 11398 7580
rect 11440 7540 11480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 19112 7540 19152 7580
rect 19194 7540 19234 7580
rect 19276 7540 19316 7580
rect 19358 7540 19398 7580
rect 19440 7540 19480 7580
rect 23112 7540 23152 7580
rect 23194 7540 23234 7580
rect 23276 7540 23316 7580
rect 23358 7540 23398 7580
rect 23440 7540 23480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 31112 7540 31152 7580
rect 31194 7540 31234 7580
rect 31276 7540 31316 7580
rect 31358 7540 31398 7580
rect 31440 7540 31480 7580
rect 35112 7540 35152 7580
rect 35194 7540 35234 7580
rect 35276 7540 35316 7580
rect 35358 7540 35398 7580
rect 35440 7540 35480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 43112 7540 43152 7580
rect 43194 7540 43234 7580
rect 43276 7540 43316 7580
rect 43358 7540 43398 7580
rect 43440 7540 43480 7580
rect 47112 7540 47152 7580
rect 47194 7540 47234 7580
rect 47276 7540 47316 7580
rect 47358 7540 47398 7580
rect 47440 7540 47480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 55112 7540 55152 7580
rect 55194 7540 55234 7580
rect 55276 7540 55316 7580
rect 55358 7540 55398 7580
rect 55440 7540 55480 7580
rect 59112 7540 59152 7580
rect 59194 7540 59234 7580
rect 59276 7540 59316 7580
rect 59358 7540 59398 7580
rect 59440 7540 59480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 67112 7540 67152 7580
rect 67194 7540 67234 7580
rect 67276 7540 67316 7580
rect 67358 7540 67398 7580
rect 67440 7540 67480 7580
rect 71112 7540 71152 7580
rect 71194 7540 71234 7580
rect 71276 7540 71316 7580
rect 71358 7540 71398 7580
rect 71440 7540 71480 7580
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 79112 7540 79152 7580
rect 79194 7540 79234 7580
rect 79276 7540 79316 7580
rect 79358 7540 79398 7580
rect 79440 7540 79480 7580
rect 83112 7540 83152 7580
rect 83194 7540 83234 7580
rect 83276 7540 83316 7580
rect 83358 7540 83398 7580
rect 83440 7540 83480 7580
rect 87112 7540 87152 7580
rect 87194 7540 87234 7580
rect 87276 7540 87316 7580
rect 87358 7540 87398 7580
rect 87440 7540 87480 7580
rect 91112 7540 91152 7580
rect 91194 7540 91234 7580
rect 91276 7540 91316 7580
rect 91358 7540 91398 7580
rect 91440 7540 91480 7580
rect 95112 7540 95152 7580
rect 95194 7540 95234 7580
rect 95276 7540 95316 7580
rect 95358 7540 95398 7580
rect 95440 7540 95480 7580
rect 99112 7540 99152 7580
rect 99194 7540 99234 7580
rect 99276 7540 99316 7580
rect 99358 7540 99398 7580
rect 99440 7540 99480 7580
rect 76780 7372 76820 7412
rect 86668 7372 86708 7412
rect 82924 7036 82964 7076
rect 88204 6952 88244 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 8352 6784 8392 6824
rect 8434 6784 8474 6824
rect 8516 6784 8556 6824
rect 8598 6784 8638 6824
rect 8680 6784 8720 6824
rect 12352 6784 12392 6824
rect 12434 6784 12474 6824
rect 12516 6784 12556 6824
rect 12598 6784 12638 6824
rect 12680 6784 12720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 20352 6784 20392 6824
rect 20434 6784 20474 6824
rect 20516 6784 20556 6824
rect 20598 6784 20638 6824
rect 20680 6784 20720 6824
rect 24352 6784 24392 6824
rect 24434 6784 24474 6824
rect 24516 6784 24556 6824
rect 24598 6784 24638 6824
rect 24680 6784 24720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 32352 6784 32392 6824
rect 32434 6784 32474 6824
rect 32516 6784 32556 6824
rect 32598 6784 32638 6824
rect 32680 6784 32720 6824
rect 36352 6784 36392 6824
rect 36434 6784 36474 6824
rect 36516 6784 36556 6824
rect 36598 6784 36638 6824
rect 36680 6784 36720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 44352 6784 44392 6824
rect 44434 6784 44474 6824
rect 44516 6784 44556 6824
rect 44598 6784 44638 6824
rect 44680 6784 44720 6824
rect 48352 6784 48392 6824
rect 48434 6784 48474 6824
rect 48516 6784 48556 6824
rect 48598 6784 48638 6824
rect 48680 6784 48720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 56352 6784 56392 6824
rect 56434 6784 56474 6824
rect 56516 6784 56556 6824
rect 56598 6784 56638 6824
rect 56680 6784 56720 6824
rect 60352 6784 60392 6824
rect 60434 6784 60474 6824
rect 60516 6784 60556 6824
rect 60598 6784 60638 6824
rect 60680 6784 60720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 68352 6784 68392 6824
rect 68434 6784 68474 6824
rect 68516 6784 68556 6824
rect 68598 6784 68638 6824
rect 68680 6784 68720 6824
rect 72352 6784 72392 6824
rect 72434 6784 72474 6824
rect 72516 6784 72556 6824
rect 72598 6784 72638 6824
rect 72680 6784 72720 6824
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 80352 6784 80392 6824
rect 80434 6784 80474 6824
rect 80516 6784 80556 6824
rect 80598 6784 80638 6824
rect 80680 6784 80720 6824
rect 84352 6784 84392 6824
rect 84434 6784 84474 6824
rect 84516 6784 84556 6824
rect 84598 6784 84638 6824
rect 84680 6784 84720 6824
rect 88352 6784 88392 6824
rect 88434 6784 88474 6824
rect 88516 6784 88556 6824
rect 88598 6784 88638 6824
rect 88680 6784 88720 6824
rect 92352 6784 92392 6824
rect 92434 6784 92474 6824
rect 92516 6784 92556 6824
rect 92598 6784 92638 6824
rect 92680 6784 92720 6824
rect 96352 6784 96392 6824
rect 96434 6784 96474 6824
rect 96516 6784 96556 6824
rect 96598 6784 96638 6824
rect 96680 6784 96720 6824
rect 95596 6700 95636 6740
rect 88204 6616 88244 6656
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 7112 6028 7152 6068
rect 7194 6028 7234 6068
rect 7276 6028 7316 6068
rect 7358 6028 7398 6068
rect 7440 6028 7480 6068
rect 11112 6028 11152 6068
rect 11194 6028 11234 6068
rect 11276 6028 11316 6068
rect 11358 6028 11398 6068
rect 11440 6028 11480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 19112 6028 19152 6068
rect 19194 6028 19234 6068
rect 19276 6028 19316 6068
rect 19358 6028 19398 6068
rect 19440 6028 19480 6068
rect 23112 6028 23152 6068
rect 23194 6028 23234 6068
rect 23276 6028 23316 6068
rect 23358 6028 23398 6068
rect 23440 6028 23480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 31112 6028 31152 6068
rect 31194 6028 31234 6068
rect 31276 6028 31316 6068
rect 31358 6028 31398 6068
rect 31440 6028 31480 6068
rect 35112 6028 35152 6068
rect 35194 6028 35234 6068
rect 35276 6028 35316 6068
rect 35358 6028 35398 6068
rect 35440 6028 35480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 43112 6028 43152 6068
rect 43194 6028 43234 6068
rect 43276 6028 43316 6068
rect 43358 6028 43398 6068
rect 43440 6028 43480 6068
rect 47112 6028 47152 6068
rect 47194 6028 47234 6068
rect 47276 6028 47316 6068
rect 47358 6028 47398 6068
rect 47440 6028 47480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 55112 6028 55152 6068
rect 55194 6028 55234 6068
rect 55276 6028 55316 6068
rect 55358 6028 55398 6068
rect 55440 6028 55480 6068
rect 59112 6028 59152 6068
rect 59194 6028 59234 6068
rect 59276 6028 59316 6068
rect 59358 6028 59398 6068
rect 59440 6028 59480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 67112 6028 67152 6068
rect 67194 6028 67234 6068
rect 67276 6028 67316 6068
rect 67358 6028 67398 6068
rect 67440 6028 67480 6068
rect 71112 6028 71152 6068
rect 71194 6028 71234 6068
rect 71276 6028 71316 6068
rect 71358 6028 71398 6068
rect 71440 6028 71480 6068
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 79112 6028 79152 6068
rect 79194 6028 79234 6068
rect 79276 6028 79316 6068
rect 79358 6028 79398 6068
rect 79440 6028 79480 6068
rect 83112 6028 83152 6068
rect 83194 6028 83234 6068
rect 83276 6028 83316 6068
rect 83358 6028 83398 6068
rect 83440 6028 83480 6068
rect 87112 6028 87152 6068
rect 87194 6028 87234 6068
rect 87276 6028 87316 6068
rect 87358 6028 87398 6068
rect 87440 6028 87480 6068
rect 91112 6028 91152 6068
rect 91194 6028 91234 6068
rect 91276 6028 91316 6068
rect 91358 6028 91398 6068
rect 91440 6028 91480 6068
rect 95112 6028 95152 6068
rect 95194 6028 95234 6068
rect 95276 6028 95316 6068
rect 95358 6028 95398 6068
rect 95440 6028 95480 6068
rect 99112 6028 99152 6068
rect 99194 6028 99234 6068
rect 99276 6028 99316 6068
rect 99358 6028 99398 6068
rect 99440 6028 99480 6068
rect 76780 5860 76820 5900
rect 80140 5860 80180 5900
rect 83596 5860 83636 5900
rect 85612 5860 85652 5900
rect 89068 5860 89108 5900
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 8352 5272 8392 5312
rect 8434 5272 8474 5312
rect 8516 5272 8556 5312
rect 8598 5272 8638 5312
rect 8680 5272 8720 5312
rect 12352 5272 12392 5312
rect 12434 5272 12474 5312
rect 12516 5272 12556 5312
rect 12598 5272 12638 5312
rect 12680 5272 12720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 20352 5272 20392 5312
rect 20434 5272 20474 5312
rect 20516 5272 20556 5312
rect 20598 5272 20638 5312
rect 20680 5272 20720 5312
rect 24352 5272 24392 5312
rect 24434 5272 24474 5312
rect 24516 5272 24556 5312
rect 24598 5272 24638 5312
rect 24680 5272 24720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 32352 5272 32392 5312
rect 32434 5272 32474 5312
rect 32516 5272 32556 5312
rect 32598 5272 32638 5312
rect 32680 5272 32720 5312
rect 36352 5272 36392 5312
rect 36434 5272 36474 5312
rect 36516 5272 36556 5312
rect 36598 5272 36638 5312
rect 36680 5272 36720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 44352 5272 44392 5312
rect 44434 5272 44474 5312
rect 44516 5272 44556 5312
rect 44598 5272 44638 5312
rect 44680 5272 44720 5312
rect 48352 5272 48392 5312
rect 48434 5272 48474 5312
rect 48516 5272 48556 5312
rect 48598 5272 48638 5312
rect 48680 5272 48720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 56352 5272 56392 5312
rect 56434 5272 56474 5312
rect 56516 5272 56556 5312
rect 56598 5272 56638 5312
rect 56680 5272 56720 5312
rect 60352 5272 60392 5312
rect 60434 5272 60474 5312
rect 60516 5272 60556 5312
rect 60598 5272 60638 5312
rect 60680 5272 60720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 68352 5272 68392 5312
rect 68434 5272 68474 5312
rect 68516 5272 68556 5312
rect 68598 5272 68638 5312
rect 68680 5272 68720 5312
rect 72352 5272 72392 5312
rect 72434 5272 72474 5312
rect 72516 5272 72556 5312
rect 72598 5272 72638 5312
rect 72680 5272 72720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 80352 5272 80392 5312
rect 80434 5272 80474 5312
rect 80516 5272 80556 5312
rect 80598 5272 80638 5312
rect 80680 5272 80720 5312
rect 84352 5272 84392 5312
rect 84434 5272 84474 5312
rect 84516 5272 84556 5312
rect 84598 5272 84638 5312
rect 84680 5272 84720 5312
rect 88352 5272 88392 5312
rect 88434 5272 88474 5312
rect 88516 5272 88556 5312
rect 88598 5272 88638 5312
rect 88680 5272 88720 5312
rect 92352 5272 92392 5312
rect 92434 5272 92474 5312
rect 92516 5272 92556 5312
rect 92598 5272 92638 5312
rect 92680 5272 92720 5312
rect 96352 5272 96392 5312
rect 96434 5272 96474 5312
rect 96516 5272 96556 5312
rect 96598 5272 96638 5312
rect 96680 5272 96720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 7112 4516 7152 4556
rect 7194 4516 7234 4556
rect 7276 4516 7316 4556
rect 7358 4516 7398 4556
rect 7440 4516 7480 4556
rect 11112 4516 11152 4556
rect 11194 4516 11234 4556
rect 11276 4516 11316 4556
rect 11358 4516 11398 4556
rect 11440 4516 11480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 19112 4516 19152 4556
rect 19194 4516 19234 4556
rect 19276 4516 19316 4556
rect 19358 4516 19398 4556
rect 19440 4516 19480 4556
rect 23112 4516 23152 4556
rect 23194 4516 23234 4556
rect 23276 4516 23316 4556
rect 23358 4516 23398 4556
rect 23440 4516 23480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 31112 4516 31152 4556
rect 31194 4516 31234 4556
rect 31276 4516 31316 4556
rect 31358 4516 31398 4556
rect 31440 4516 31480 4556
rect 35112 4516 35152 4556
rect 35194 4516 35234 4556
rect 35276 4516 35316 4556
rect 35358 4516 35398 4556
rect 35440 4516 35480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 43112 4516 43152 4556
rect 43194 4516 43234 4556
rect 43276 4516 43316 4556
rect 43358 4516 43398 4556
rect 43440 4516 43480 4556
rect 47112 4516 47152 4556
rect 47194 4516 47234 4556
rect 47276 4516 47316 4556
rect 47358 4516 47398 4556
rect 47440 4516 47480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 55112 4516 55152 4556
rect 55194 4516 55234 4556
rect 55276 4516 55316 4556
rect 55358 4516 55398 4556
rect 55440 4516 55480 4556
rect 59112 4516 59152 4556
rect 59194 4516 59234 4556
rect 59276 4516 59316 4556
rect 59358 4516 59398 4556
rect 59440 4516 59480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 67112 4516 67152 4556
rect 67194 4516 67234 4556
rect 67276 4516 67316 4556
rect 67358 4516 67398 4556
rect 67440 4516 67480 4556
rect 71112 4516 71152 4556
rect 71194 4516 71234 4556
rect 71276 4516 71316 4556
rect 71358 4516 71398 4556
rect 71440 4516 71480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 79112 4516 79152 4556
rect 79194 4516 79234 4556
rect 79276 4516 79316 4556
rect 79358 4516 79398 4556
rect 79440 4516 79480 4556
rect 83112 4516 83152 4556
rect 83194 4516 83234 4556
rect 83276 4516 83316 4556
rect 83358 4516 83398 4556
rect 83440 4516 83480 4556
rect 87112 4516 87152 4556
rect 87194 4516 87234 4556
rect 87276 4516 87316 4556
rect 87358 4516 87398 4556
rect 87440 4516 87480 4556
rect 91112 4516 91152 4556
rect 91194 4516 91234 4556
rect 91276 4516 91316 4556
rect 91358 4516 91398 4556
rect 91440 4516 91480 4556
rect 95112 4516 95152 4556
rect 95194 4516 95234 4556
rect 95276 4516 95316 4556
rect 95358 4516 95398 4556
rect 95440 4516 95480 4556
rect 99112 4516 99152 4556
rect 99194 4516 99234 4556
rect 99276 4516 99316 4556
rect 99358 4516 99398 4556
rect 99440 4516 99480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 8352 3760 8392 3800
rect 8434 3760 8474 3800
rect 8516 3760 8556 3800
rect 8598 3760 8638 3800
rect 8680 3760 8720 3800
rect 12352 3760 12392 3800
rect 12434 3760 12474 3800
rect 12516 3760 12556 3800
rect 12598 3760 12638 3800
rect 12680 3760 12720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 20352 3760 20392 3800
rect 20434 3760 20474 3800
rect 20516 3760 20556 3800
rect 20598 3760 20638 3800
rect 20680 3760 20720 3800
rect 24352 3760 24392 3800
rect 24434 3760 24474 3800
rect 24516 3760 24556 3800
rect 24598 3760 24638 3800
rect 24680 3760 24720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 32352 3760 32392 3800
rect 32434 3760 32474 3800
rect 32516 3760 32556 3800
rect 32598 3760 32638 3800
rect 32680 3760 32720 3800
rect 36352 3760 36392 3800
rect 36434 3760 36474 3800
rect 36516 3760 36556 3800
rect 36598 3760 36638 3800
rect 36680 3760 36720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 44352 3760 44392 3800
rect 44434 3760 44474 3800
rect 44516 3760 44556 3800
rect 44598 3760 44638 3800
rect 44680 3760 44720 3800
rect 48352 3760 48392 3800
rect 48434 3760 48474 3800
rect 48516 3760 48556 3800
rect 48598 3760 48638 3800
rect 48680 3760 48720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 56352 3760 56392 3800
rect 56434 3760 56474 3800
rect 56516 3760 56556 3800
rect 56598 3760 56638 3800
rect 56680 3760 56720 3800
rect 60352 3760 60392 3800
rect 60434 3760 60474 3800
rect 60516 3760 60556 3800
rect 60598 3760 60638 3800
rect 60680 3760 60720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 68352 3760 68392 3800
rect 68434 3760 68474 3800
rect 68516 3760 68556 3800
rect 68598 3760 68638 3800
rect 68680 3760 68720 3800
rect 72352 3760 72392 3800
rect 72434 3760 72474 3800
rect 72516 3760 72556 3800
rect 72598 3760 72638 3800
rect 72680 3760 72720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 80352 3760 80392 3800
rect 80434 3760 80474 3800
rect 80516 3760 80556 3800
rect 80598 3760 80638 3800
rect 80680 3760 80720 3800
rect 84352 3760 84392 3800
rect 84434 3760 84474 3800
rect 84516 3760 84556 3800
rect 84598 3760 84638 3800
rect 84680 3760 84720 3800
rect 88352 3760 88392 3800
rect 88434 3760 88474 3800
rect 88516 3760 88556 3800
rect 88598 3760 88638 3800
rect 88680 3760 88720 3800
rect 92352 3760 92392 3800
rect 92434 3760 92474 3800
rect 92516 3760 92556 3800
rect 92598 3760 92638 3800
rect 92680 3760 92720 3800
rect 96352 3760 96392 3800
rect 96434 3760 96474 3800
rect 96516 3760 96556 3800
rect 96598 3760 96638 3800
rect 96680 3760 96720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 7112 3004 7152 3044
rect 7194 3004 7234 3044
rect 7276 3004 7316 3044
rect 7358 3004 7398 3044
rect 7440 3004 7480 3044
rect 11112 3004 11152 3044
rect 11194 3004 11234 3044
rect 11276 3004 11316 3044
rect 11358 3004 11398 3044
rect 11440 3004 11480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 19112 3004 19152 3044
rect 19194 3004 19234 3044
rect 19276 3004 19316 3044
rect 19358 3004 19398 3044
rect 19440 3004 19480 3044
rect 23112 3004 23152 3044
rect 23194 3004 23234 3044
rect 23276 3004 23316 3044
rect 23358 3004 23398 3044
rect 23440 3004 23480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 31112 3004 31152 3044
rect 31194 3004 31234 3044
rect 31276 3004 31316 3044
rect 31358 3004 31398 3044
rect 31440 3004 31480 3044
rect 35112 3004 35152 3044
rect 35194 3004 35234 3044
rect 35276 3004 35316 3044
rect 35358 3004 35398 3044
rect 35440 3004 35480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 43112 3004 43152 3044
rect 43194 3004 43234 3044
rect 43276 3004 43316 3044
rect 43358 3004 43398 3044
rect 43440 3004 43480 3044
rect 47112 3004 47152 3044
rect 47194 3004 47234 3044
rect 47276 3004 47316 3044
rect 47358 3004 47398 3044
rect 47440 3004 47480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 55112 3004 55152 3044
rect 55194 3004 55234 3044
rect 55276 3004 55316 3044
rect 55358 3004 55398 3044
rect 55440 3004 55480 3044
rect 59112 3004 59152 3044
rect 59194 3004 59234 3044
rect 59276 3004 59316 3044
rect 59358 3004 59398 3044
rect 59440 3004 59480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 67112 3004 67152 3044
rect 67194 3004 67234 3044
rect 67276 3004 67316 3044
rect 67358 3004 67398 3044
rect 67440 3004 67480 3044
rect 71112 3004 71152 3044
rect 71194 3004 71234 3044
rect 71276 3004 71316 3044
rect 71358 3004 71398 3044
rect 71440 3004 71480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 79112 3004 79152 3044
rect 79194 3004 79234 3044
rect 79276 3004 79316 3044
rect 79358 3004 79398 3044
rect 79440 3004 79480 3044
rect 83112 3004 83152 3044
rect 83194 3004 83234 3044
rect 83276 3004 83316 3044
rect 83358 3004 83398 3044
rect 83440 3004 83480 3044
rect 87112 3004 87152 3044
rect 87194 3004 87234 3044
rect 87276 3004 87316 3044
rect 87358 3004 87398 3044
rect 87440 3004 87480 3044
rect 91112 3004 91152 3044
rect 91194 3004 91234 3044
rect 91276 3004 91316 3044
rect 91358 3004 91398 3044
rect 91440 3004 91480 3044
rect 95112 3004 95152 3044
rect 95194 3004 95234 3044
rect 95276 3004 95316 3044
rect 95358 3004 95398 3044
rect 95440 3004 95480 3044
rect 99112 3004 99152 3044
rect 99194 3004 99234 3044
rect 99276 3004 99316 3044
rect 99358 3004 99398 3044
rect 99440 3004 99480 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 8352 2248 8392 2288
rect 8434 2248 8474 2288
rect 8516 2248 8556 2288
rect 8598 2248 8638 2288
rect 8680 2248 8720 2288
rect 12352 2248 12392 2288
rect 12434 2248 12474 2288
rect 12516 2248 12556 2288
rect 12598 2248 12638 2288
rect 12680 2248 12720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 20352 2248 20392 2288
rect 20434 2248 20474 2288
rect 20516 2248 20556 2288
rect 20598 2248 20638 2288
rect 20680 2248 20720 2288
rect 24352 2248 24392 2288
rect 24434 2248 24474 2288
rect 24516 2248 24556 2288
rect 24598 2248 24638 2288
rect 24680 2248 24720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 32352 2248 32392 2288
rect 32434 2248 32474 2288
rect 32516 2248 32556 2288
rect 32598 2248 32638 2288
rect 32680 2248 32720 2288
rect 36352 2248 36392 2288
rect 36434 2248 36474 2288
rect 36516 2248 36556 2288
rect 36598 2248 36638 2288
rect 36680 2248 36720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 44352 2248 44392 2288
rect 44434 2248 44474 2288
rect 44516 2248 44556 2288
rect 44598 2248 44638 2288
rect 44680 2248 44720 2288
rect 48352 2248 48392 2288
rect 48434 2248 48474 2288
rect 48516 2248 48556 2288
rect 48598 2248 48638 2288
rect 48680 2248 48720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 56352 2248 56392 2288
rect 56434 2248 56474 2288
rect 56516 2248 56556 2288
rect 56598 2248 56638 2288
rect 56680 2248 56720 2288
rect 60352 2248 60392 2288
rect 60434 2248 60474 2288
rect 60516 2248 60556 2288
rect 60598 2248 60638 2288
rect 60680 2248 60720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 68352 2248 68392 2288
rect 68434 2248 68474 2288
rect 68516 2248 68556 2288
rect 68598 2248 68638 2288
rect 68680 2248 68720 2288
rect 72352 2248 72392 2288
rect 72434 2248 72474 2288
rect 72516 2248 72556 2288
rect 72598 2248 72638 2288
rect 72680 2248 72720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 80352 2248 80392 2288
rect 80434 2248 80474 2288
rect 80516 2248 80556 2288
rect 80598 2248 80638 2288
rect 80680 2248 80720 2288
rect 84352 2248 84392 2288
rect 84434 2248 84474 2288
rect 84516 2248 84556 2288
rect 84598 2248 84638 2288
rect 84680 2248 84720 2288
rect 88352 2248 88392 2288
rect 88434 2248 88474 2288
rect 88516 2248 88556 2288
rect 88598 2248 88638 2288
rect 88680 2248 88720 2288
rect 92352 2248 92392 2288
rect 92434 2248 92474 2288
rect 92516 2248 92556 2288
rect 92598 2248 92638 2288
rect 92680 2248 92720 2288
rect 96352 2248 96392 2288
rect 96434 2248 96474 2288
rect 96516 2248 96556 2288
rect 96598 2248 96638 2288
rect 96680 2248 96720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 7112 1492 7152 1532
rect 7194 1492 7234 1532
rect 7276 1492 7316 1532
rect 7358 1492 7398 1532
rect 7440 1492 7480 1532
rect 11112 1492 11152 1532
rect 11194 1492 11234 1532
rect 11276 1492 11316 1532
rect 11358 1492 11398 1532
rect 11440 1492 11480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 19112 1492 19152 1532
rect 19194 1492 19234 1532
rect 19276 1492 19316 1532
rect 19358 1492 19398 1532
rect 19440 1492 19480 1532
rect 23112 1492 23152 1532
rect 23194 1492 23234 1532
rect 23276 1492 23316 1532
rect 23358 1492 23398 1532
rect 23440 1492 23480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 31112 1492 31152 1532
rect 31194 1492 31234 1532
rect 31276 1492 31316 1532
rect 31358 1492 31398 1532
rect 31440 1492 31480 1532
rect 35112 1492 35152 1532
rect 35194 1492 35234 1532
rect 35276 1492 35316 1532
rect 35358 1492 35398 1532
rect 35440 1492 35480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 43112 1492 43152 1532
rect 43194 1492 43234 1532
rect 43276 1492 43316 1532
rect 43358 1492 43398 1532
rect 43440 1492 43480 1532
rect 47112 1492 47152 1532
rect 47194 1492 47234 1532
rect 47276 1492 47316 1532
rect 47358 1492 47398 1532
rect 47440 1492 47480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 55112 1492 55152 1532
rect 55194 1492 55234 1532
rect 55276 1492 55316 1532
rect 55358 1492 55398 1532
rect 55440 1492 55480 1532
rect 59112 1492 59152 1532
rect 59194 1492 59234 1532
rect 59276 1492 59316 1532
rect 59358 1492 59398 1532
rect 59440 1492 59480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 67112 1492 67152 1532
rect 67194 1492 67234 1532
rect 67276 1492 67316 1532
rect 67358 1492 67398 1532
rect 67440 1492 67480 1532
rect 71112 1492 71152 1532
rect 71194 1492 71234 1532
rect 71276 1492 71316 1532
rect 71358 1492 71398 1532
rect 71440 1492 71480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 79112 1492 79152 1532
rect 79194 1492 79234 1532
rect 79276 1492 79316 1532
rect 79358 1492 79398 1532
rect 79440 1492 79480 1532
rect 83112 1492 83152 1532
rect 83194 1492 83234 1532
rect 83276 1492 83316 1532
rect 83358 1492 83398 1532
rect 83440 1492 83480 1532
rect 87112 1492 87152 1532
rect 87194 1492 87234 1532
rect 87276 1492 87316 1532
rect 87358 1492 87398 1532
rect 87440 1492 87480 1532
rect 91112 1492 91152 1532
rect 91194 1492 91234 1532
rect 91276 1492 91316 1532
rect 91358 1492 91398 1532
rect 91440 1492 91480 1532
rect 95112 1492 95152 1532
rect 95194 1492 95234 1532
rect 95276 1492 95316 1532
rect 95358 1492 95398 1532
rect 95440 1492 95480 1532
rect 99112 1492 99152 1532
rect 99194 1492 99234 1532
rect 99276 1492 99316 1532
rect 99358 1492 99398 1532
rect 99440 1492 99480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 8352 736 8392 776
rect 8434 736 8474 776
rect 8516 736 8556 776
rect 8598 736 8638 776
rect 8680 736 8720 776
rect 12352 736 12392 776
rect 12434 736 12474 776
rect 12516 736 12556 776
rect 12598 736 12638 776
rect 12680 736 12720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 20352 736 20392 776
rect 20434 736 20474 776
rect 20516 736 20556 776
rect 20598 736 20638 776
rect 20680 736 20720 776
rect 24352 736 24392 776
rect 24434 736 24474 776
rect 24516 736 24556 776
rect 24598 736 24638 776
rect 24680 736 24720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 32352 736 32392 776
rect 32434 736 32474 776
rect 32516 736 32556 776
rect 32598 736 32638 776
rect 32680 736 32720 776
rect 36352 736 36392 776
rect 36434 736 36474 776
rect 36516 736 36556 776
rect 36598 736 36638 776
rect 36680 736 36720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 44352 736 44392 776
rect 44434 736 44474 776
rect 44516 736 44556 776
rect 44598 736 44638 776
rect 44680 736 44720 776
rect 48352 736 48392 776
rect 48434 736 48474 776
rect 48516 736 48556 776
rect 48598 736 48638 776
rect 48680 736 48720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 56352 736 56392 776
rect 56434 736 56474 776
rect 56516 736 56556 776
rect 56598 736 56638 776
rect 56680 736 56720 776
rect 60352 736 60392 776
rect 60434 736 60474 776
rect 60516 736 60556 776
rect 60598 736 60638 776
rect 60680 736 60720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 68352 736 68392 776
rect 68434 736 68474 776
rect 68516 736 68556 776
rect 68598 736 68638 776
rect 68680 736 68720 776
rect 72352 736 72392 776
rect 72434 736 72474 776
rect 72516 736 72556 776
rect 72598 736 72638 776
rect 72680 736 72720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
rect 80352 736 80392 776
rect 80434 736 80474 776
rect 80516 736 80556 776
rect 80598 736 80638 776
rect 80680 736 80720 776
rect 84352 736 84392 776
rect 84434 736 84474 776
rect 84516 736 84556 776
rect 84598 736 84638 776
rect 84680 736 84720 776
rect 88352 736 88392 776
rect 88434 736 88474 776
rect 88516 736 88556 776
rect 88598 736 88638 776
rect 88680 736 88720 776
rect 92352 736 92392 776
rect 92434 736 92474 776
rect 92516 736 92556 776
rect 92598 736 92638 776
rect 92680 736 92720 776
rect 96352 736 96392 776
rect 96434 736 96474 776
rect 96516 736 96556 776
rect 96598 736 96638 776
rect 96680 736 96720 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 8352 38576 8720 38585
rect 8392 38536 8434 38576
rect 8474 38536 8516 38576
rect 8556 38536 8598 38576
rect 8638 38536 8680 38576
rect 8352 38527 8720 38536
rect 12352 38576 12720 38585
rect 12392 38536 12434 38576
rect 12474 38536 12516 38576
rect 12556 38536 12598 38576
rect 12638 38536 12680 38576
rect 12352 38527 12720 38536
rect 16352 38576 16720 38585
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16352 38527 16720 38536
rect 20352 38576 20720 38585
rect 20392 38536 20434 38576
rect 20474 38536 20516 38576
rect 20556 38536 20598 38576
rect 20638 38536 20680 38576
rect 20352 38527 20720 38536
rect 24352 38576 24720 38585
rect 24392 38536 24434 38576
rect 24474 38536 24516 38576
rect 24556 38536 24598 38576
rect 24638 38536 24680 38576
rect 24352 38527 24720 38536
rect 28352 38576 28720 38585
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28352 38527 28720 38536
rect 32352 38576 32720 38585
rect 32392 38536 32434 38576
rect 32474 38536 32516 38576
rect 32556 38536 32598 38576
rect 32638 38536 32680 38576
rect 32352 38527 32720 38536
rect 36352 38576 36720 38585
rect 36392 38536 36434 38576
rect 36474 38536 36516 38576
rect 36556 38536 36598 38576
rect 36638 38536 36680 38576
rect 36352 38527 36720 38536
rect 40352 38576 40720 38585
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40352 38527 40720 38536
rect 44352 38576 44720 38585
rect 44392 38536 44434 38576
rect 44474 38536 44516 38576
rect 44556 38536 44598 38576
rect 44638 38536 44680 38576
rect 44352 38527 44720 38536
rect 48352 38576 48720 38585
rect 48392 38536 48434 38576
rect 48474 38536 48516 38576
rect 48556 38536 48598 38576
rect 48638 38536 48680 38576
rect 48352 38527 48720 38536
rect 52352 38576 52720 38585
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52352 38527 52720 38536
rect 56352 38576 56720 38585
rect 56392 38536 56434 38576
rect 56474 38536 56516 38576
rect 56556 38536 56598 38576
rect 56638 38536 56680 38576
rect 56352 38527 56720 38536
rect 60352 38576 60720 38585
rect 60392 38536 60434 38576
rect 60474 38536 60516 38576
rect 60556 38536 60598 38576
rect 60638 38536 60680 38576
rect 60352 38527 60720 38536
rect 64352 38576 64720 38585
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64352 38527 64720 38536
rect 68352 38576 68720 38585
rect 68392 38536 68434 38576
rect 68474 38536 68516 38576
rect 68556 38536 68598 38576
rect 68638 38536 68680 38576
rect 68352 38527 68720 38536
rect 72352 38576 72720 38585
rect 72392 38536 72434 38576
rect 72474 38536 72516 38576
rect 72556 38536 72598 38576
rect 72638 38536 72680 38576
rect 72352 38527 72720 38536
rect 76352 38576 76720 38585
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76352 38527 76720 38536
rect 80352 38576 80720 38585
rect 80392 38536 80434 38576
rect 80474 38536 80516 38576
rect 80556 38536 80598 38576
rect 80638 38536 80680 38576
rect 80352 38527 80720 38536
rect 84352 38576 84720 38585
rect 84392 38536 84434 38576
rect 84474 38536 84516 38576
rect 84556 38536 84598 38576
rect 84638 38536 84680 38576
rect 84352 38527 84720 38536
rect 88352 38576 88720 38585
rect 88392 38536 88434 38576
rect 88474 38536 88516 38576
rect 88556 38536 88598 38576
rect 88638 38536 88680 38576
rect 88352 38527 88720 38536
rect 92352 38576 92720 38585
rect 92392 38536 92434 38576
rect 92474 38536 92516 38576
rect 92556 38536 92598 38576
rect 92638 38536 92680 38576
rect 92352 38527 92720 38536
rect 96352 38576 96720 38585
rect 96392 38536 96434 38576
rect 96474 38536 96516 38576
rect 96556 38536 96598 38576
rect 96638 38536 96680 38576
rect 96352 38527 96720 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 7112 37820 7480 37829
rect 7152 37780 7194 37820
rect 7234 37780 7276 37820
rect 7316 37780 7358 37820
rect 7398 37780 7440 37820
rect 7112 37771 7480 37780
rect 11112 37820 11480 37829
rect 11152 37780 11194 37820
rect 11234 37780 11276 37820
rect 11316 37780 11358 37820
rect 11398 37780 11440 37820
rect 11112 37771 11480 37780
rect 15112 37820 15480 37829
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15112 37771 15480 37780
rect 19112 37820 19480 37829
rect 19152 37780 19194 37820
rect 19234 37780 19276 37820
rect 19316 37780 19358 37820
rect 19398 37780 19440 37820
rect 19112 37771 19480 37780
rect 23112 37820 23480 37829
rect 23152 37780 23194 37820
rect 23234 37780 23276 37820
rect 23316 37780 23358 37820
rect 23398 37780 23440 37820
rect 23112 37771 23480 37780
rect 27112 37820 27480 37829
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27112 37771 27480 37780
rect 31112 37820 31480 37829
rect 31152 37780 31194 37820
rect 31234 37780 31276 37820
rect 31316 37780 31358 37820
rect 31398 37780 31440 37820
rect 31112 37771 31480 37780
rect 35112 37820 35480 37829
rect 35152 37780 35194 37820
rect 35234 37780 35276 37820
rect 35316 37780 35358 37820
rect 35398 37780 35440 37820
rect 35112 37771 35480 37780
rect 39112 37820 39480 37829
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39112 37771 39480 37780
rect 43112 37820 43480 37829
rect 43152 37780 43194 37820
rect 43234 37780 43276 37820
rect 43316 37780 43358 37820
rect 43398 37780 43440 37820
rect 43112 37771 43480 37780
rect 47112 37820 47480 37829
rect 47152 37780 47194 37820
rect 47234 37780 47276 37820
rect 47316 37780 47358 37820
rect 47398 37780 47440 37820
rect 47112 37771 47480 37780
rect 51112 37820 51480 37829
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51112 37771 51480 37780
rect 55112 37820 55480 37829
rect 55152 37780 55194 37820
rect 55234 37780 55276 37820
rect 55316 37780 55358 37820
rect 55398 37780 55440 37820
rect 55112 37771 55480 37780
rect 59112 37820 59480 37829
rect 59152 37780 59194 37820
rect 59234 37780 59276 37820
rect 59316 37780 59358 37820
rect 59398 37780 59440 37820
rect 59112 37771 59480 37780
rect 63112 37820 63480 37829
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63112 37771 63480 37780
rect 67112 37820 67480 37829
rect 67152 37780 67194 37820
rect 67234 37780 67276 37820
rect 67316 37780 67358 37820
rect 67398 37780 67440 37820
rect 67112 37771 67480 37780
rect 71112 37820 71480 37829
rect 71152 37780 71194 37820
rect 71234 37780 71276 37820
rect 71316 37780 71358 37820
rect 71398 37780 71440 37820
rect 71112 37771 71480 37780
rect 75112 37820 75480 37829
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75112 37771 75480 37780
rect 79112 37820 79480 37829
rect 79152 37780 79194 37820
rect 79234 37780 79276 37820
rect 79316 37780 79358 37820
rect 79398 37780 79440 37820
rect 79112 37771 79480 37780
rect 83112 37820 83480 37829
rect 83152 37780 83194 37820
rect 83234 37780 83276 37820
rect 83316 37780 83358 37820
rect 83398 37780 83440 37820
rect 83112 37771 83480 37780
rect 87112 37820 87480 37829
rect 87152 37780 87194 37820
rect 87234 37780 87276 37820
rect 87316 37780 87358 37820
rect 87398 37780 87440 37820
rect 87112 37771 87480 37780
rect 91112 37820 91480 37829
rect 91152 37780 91194 37820
rect 91234 37780 91276 37820
rect 91316 37780 91358 37820
rect 91398 37780 91440 37820
rect 91112 37771 91480 37780
rect 95112 37820 95480 37829
rect 95152 37780 95194 37820
rect 95234 37780 95276 37820
rect 95316 37780 95358 37820
rect 95398 37780 95440 37820
rect 95112 37771 95480 37780
rect 99112 37820 99480 37829
rect 99152 37780 99194 37820
rect 99234 37780 99276 37820
rect 99316 37780 99358 37820
rect 99398 37780 99440 37820
rect 99112 37771 99480 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 8352 37064 8720 37073
rect 8392 37024 8434 37064
rect 8474 37024 8516 37064
rect 8556 37024 8598 37064
rect 8638 37024 8680 37064
rect 8352 37015 8720 37024
rect 12352 37064 12720 37073
rect 12392 37024 12434 37064
rect 12474 37024 12516 37064
rect 12556 37024 12598 37064
rect 12638 37024 12680 37064
rect 12352 37015 12720 37024
rect 16352 37064 16720 37073
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16352 37015 16720 37024
rect 20352 37064 20720 37073
rect 20392 37024 20434 37064
rect 20474 37024 20516 37064
rect 20556 37024 20598 37064
rect 20638 37024 20680 37064
rect 20352 37015 20720 37024
rect 24352 37064 24720 37073
rect 24392 37024 24434 37064
rect 24474 37024 24516 37064
rect 24556 37024 24598 37064
rect 24638 37024 24680 37064
rect 24352 37015 24720 37024
rect 28352 37064 28720 37073
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28352 37015 28720 37024
rect 32352 37064 32720 37073
rect 32392 37024 32434 37064
rect 32474 37024 32516 37064
rect 32556 37024 32598 37064
rect 32638 37024 32680 37064
rect 32352 37015 32720 37024
rect 36352 37064 36720 37073
rect 36392 37024 36434 37064
rect 36474 37024 36516 37064
rect 36556 37024 36598 37064
rect 36638 37024 36680 37064
rect 36352 37015 36720 37024
rect 40352 37064 40720 37073
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40352 37015 40720 37024
rect 44352 37064 44720 37073
rect 44392 37024 44434 37064
rect 44474 37024 44516 37064
rect 44556 37024 44598 37064
rect 44638 37024 44680 37064
rect 44352 37015 44720 37024
rect 48352 37064 48720 37073
rect 48392 37024 48434 37064
rect 48474 37024 48516 37064
rect 48556 37024 48598 37064
rect 48638 37024 48680 37064
rect 48352 37015 48720 37024
rect 52352 37064 52720 37073
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52352 37015 52720 37024
rect 56352 37064 56720 37073
rect 56392 37024 56434 37064
rect 56474 37024 56516 37064
rect 56556 37024 56598 37064
rect 56638 37024 56680 37064
rect 56352 37015 56720 37024
rect 60352 37064 60720 37073
rect 60392 37024 60434 37064
rect 60474 37024 60516 37064
rect 60556 37024 60598 37064
rect 60638 37024 60680 37064
rect 60352 37015 60720 37024
rect 64352 37064 64720 37073
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64352 37015 64720 37024
rect 68352 37064 68720 37073
rect 68392 37024 68434 37064
rect 68474 37024 68516 37064
rect 68556 37024 68598 37064
rect 68638 37024 68680 37064
rect 68352 37015 68720 37024
rect 72352 37064 72720 37073
rect 72392 37024 72434 37064
rect 72474 37024 72516 37064
rect 72556 37024 72598 37064
rect 72638 37024 72680 37064
rect 72352 37015 72720 37024
rect 76352 37064 76720 37073
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76352 37015 76720 37024
rect 80352 37064 80720 37073
rect 80392 37024 80434 37064
rect 80474 37024 80516 37064
rect 80556 37024 80598 37064
rect 80638 37024 80680 37064
rect 80352 37015 80720 37024
rect 84352 37064 84720 37073
rect 84392 37024 84434 37064
rect 84474 37024 84516 37064
rect 84556 37024 84598 37064
rect 84638 37024 84680 37064
rect 84352 37015 84720 37024
rect 88352 37064 88720 37073
rect 88392 37024 88434 37064
rect 88474 37024 88516 37064
rect 88556 37024 88598 37064
rect 88638 37024 88680 37064
rect 88352 37015 88720 37024
rect 92352 37064 92720 37073
rect 92392 37024 92434 37064
rect 92474 37024 92516 37064
rect 92556 37024 92598 37064
rect 92638 37024 92680 37064
rect 92352 37015 92720 37024
rect 96352 37064 96720 37073
rect 96392 37024 96434 37064
rect 96474 37024 96516 37064
rect 96556 37024 96598 37064
rect 96638 37024 96680 37064
rect 96352 37015 96720 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 7112 36308 7480 36317
rect 7152 36268 7194 36308
rect 7234 36268 7276 36308
rect 7316 36268 7358 36308
rect 7398 36268 7440 36308
rect 7112 36259 7480 36268
rect 11112 36308 11480 36317
rect 11152 36268 11194 36308
rect 11234 36268 11276 36308
rect 11316 36268 11358 36308
rect 11398 36268 11440 36308
rect 11112 36259 11480 36268
rect 15112 36308 15480 36317
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15112 36259 15480 36268
rect 19112 36308 19480 36317
rect 19152 36268 19194 36308
rect 19234 36268 19276 36308
rect 19316 36268 19358 36308
rect 19398 36268 19440 36308
rect 19112 36259 19480 36268
rect 23112 36308 23480 36317
rect 23152 36268 23194 36308
rect 23234 36268 23276 36308
rect 23316 36268 23358 36308
rect 23398 36268 23440 36308
rect 23112 36259 23480 36268
rect 27112 36308 27480 36317
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27112 36259 27480 36268
rect 31112 36308 31480 36317
rect 31152 36268 31194 36308
rect 31234 36268 31276 36308
rect 31316 36268 31358 36308
rect 31398 36268 31440 36308
rect 31112 36259 31480 36268
rect 35112 36308 35480 36317
rect 35152 36268 35194 36308
rect 35234 36268 35276 36308
rect 35316 36268 35358 36308
rect 35398 36268 35440 36308
rect 35112 36259 35480 36268
rect 39112 36308 39480 36317
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39112 36259 39480 36268
rect 43112 36308 43480 36317
rect 43152 36268 43194 36308
rect 43234 36268 43276 36308
rect 43316 36268 43358 36308
rect 43398 36268 43440 36308
rect 43112 36259 43480 36268
rect 47112 36308 47480 36317
rect 47152 36268 47194 36308
rect 47234 36268 47276 36308
rect 47316 36268 47358 36308
rect 47398 36268 47440 36308
rect 47112 36259 47480 36268
rect 51112 36308 51480 36317
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51112 36259 51480 36268
rect 55112 36308 55480 36317
rect 55152 36268 55194 36308
rect 55234 36268 55276 36308
rect 55316 36268 55358 36308
rect 55398 36268 55440 36308
rect 55112 36259 55480 36268
rect 59112 36308 59480 36317
rect 59152 36268 59194 36308
rect 59234 36268 59276 36308
rect 59316 36268 59358 36308
rect 59398 36268 59440 36308
rect 59112 36259 59480 36268
rect 63112 36308 63480 36317
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63112 36259 63480 36268
rect 67112 36308 67480 36317
rect 67152 36268 67194 36308
rect 67234 36268 67276 36308
rect 67316 36268 67358 36308
rect 67398 36268 67440 36308
rect 67112 36259 67480 36268
rect 71112 36308 71480 36317
rect 71152 36268 71194 36308
rect 71234 36268 71276 36308
rect 71316 36268 71358 36308
rect 71398 36268 71440 36308
rect 71112 36259 71480 36268
rect 75112 36308 75480 36317
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75112 36259 75480 36268
rect 79112 36308 79480 36317
rect 79152 36268 79194 36308
rect 79234 36268 79276 36308
rect 79316 36268 79358 36308
rect 79398 36268 79440 36308
rect 79112 36259 79480 36268
rect 83112 36308 83480 36317
rect 83152 36268 83194 36308
rect 83234 36268 83276 36308
rect 83316 36268 83358 36308
rect 83398 36268 83440 36308
rect 83112 36259 83480 36268
rect 87112 36308 87480 36317
rect 87152 36268 87194 36308
rect 87234 36268 87276 36308
rect 87316 36268 87358 36308
rect 87398 36268 87440 36308
rect 87112 36259 87480 36268
rect 91112 36308 91480 36317
rect 91152 36268 91194 36308
rect 91234 36268 91276 36308
rect 91316 36268 91358 36308
rect 91398 36268 91440 36308
rect 91112 36259 91480 36268
rect 95112 36308 95480 36317
rect 95152 36268 95194 36308
rect 95234 36268 95276 36308
rect 95316 36268 95358 36308
rect 95398 36268 95440 36308
rect 95112 36259 95480 36268
rect 99112 36308 99480 36317
rect 99152 36268 99194 36308
rect 99234 36268 99276 36308
rect 99316 36268 99358 36308
rect 99398 36268 99440 36308
rect 99112 36259 99480 36268
rect 76780 35720 76820 35729
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 8352 35552 8720 35561
rect 8392 35512 8434 35552
rect 8474 35512 8516 35552
rect 8556 35512 8598 35552
rect 8638 35512 8680 35552
rect 8352 35503 8720 35512
rect 12352 35552 12720 35561
rect 12392 35512 12434 35552
rect 12474 35512 12516 35552
rect 12556 35512 12598 35552
rect 12638 35512 12680 35552
rect 12352 35503 12720 35512
rect 16352 35552 16720 35561
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16352 35503 16720 35512
rect 20352 35552 20720 35561
rect 20392 35512 20434 35552
rect 20474 35512 20516 35552
rect 20556 35512 20598 35552
rect 20638 35512 20680 35552
rect 20352 35503 20720 35512
rect 24352 35552 24720 35561
rect 24392 35512 24434 35552
rect 24474 35512 24516 35552
rect 24556 35512 24598 35552
rect 24638 35512 24680 35552
rect 24352 35503 24720 35512
rect 28352 35552 28720 35561
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28352 35503 28720 35512
rect 32352 35552 32720 35561
rect 32392 35512 32434 35552
rect 32474 35512 32516 35552
rect 32556 35512 32598 35552
rect 32638 35512 32680 35552
rect 32352 35503 32720 35512
rect 36352 35552 36720 35561
rect 36392 35512 36434 35552
rect 36474 35512 36516 35552
rect 36556 35512 36598 35552
rect 36638 35512 36680 35552
rect 36352 35503 36720 35512
rect 40352 35552 40720 35561
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40352 35503 40720 35512
rect 44352 35552 44720 35561
rect 44392 35512 44434 35552
rect 44474 35512 44516 35552
rect 44556 35512 44598 35552
rect 44638 35512 44680 35552
rect 44352 35503 44720 35512
rect 48352 35552 48720 35561
rect 48392 35512 48434 35552
rect 48474 35512 48516 35552
rect 48556 35512 48598 35552
rect 48638 35512 48680 35552
rect 48352 35503 48720 35512
rect 52352 35552 52720 35561
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52352 35503 52720 35512
rect 56352 35552 56720 35561
rect 56392 35512 56434 35552
rect 56474 35512 56516 35552
rect 56556 35512 56598 35552
rect 56638 35512 56680 35552
rect 56352 35503 56720 35512
rect 60352 35552 60720 35561
rect 60392 35512 60434 35552
rect 60474 35512 60516 35552
rect 60556 35512 60598 35552
rect 60638 35512 60680 35552
rect 60352 35503 60720 35512
rect 64352 35552 64720 35561
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64352 35503 64720 35512
rect 68352 35552 68720 35561
rect 68392 35512 68434 35552
rect 68474 35512 68516 35552
rect 68556 35512 68598 35552
rect 68638 35512 68680 35552
rect 68352 35503 68720 35512
rect 72352 35552 72720 35561
rect 72392 35512 72434 35552
rect 72474 35512 72516 35552
rect 72556 35512 72598 35552
rect 72638 35512 72680 35552
rect 72352 35503 72720 35512
rect 76352 35552 76720 35561
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76352 35503 76720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 7112 34796 7480 34805
rect 7152 34756 7194 34796
rect 7234 34756 7276 34796
rect 7316 34756 7358 34796
rect 7398 34756 7440 34796
rect 7112 34747 7480 34756
rect 11112 34796 11480 34805
rect 11152 34756 11194 34796
rect 11234 34756 11276 34796
rect 11316 34756 11358 34796
rect 11398 34756 11440 34796
rect 11112 34747 11480 34756
rect 15112 34796 15480 34805
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15112 34747 15480 34756
rect 19112 34796 19480 34805
rect 19152 34756 19194 34796
rect 19234 34756 19276 34796
rect 19316 34756 19358 34796
rect 19398 34756 19440 34796
rect 19112 34747 19480 34756
rect 23112 34796 23480 34805
rect 23152 34756 23194 34796
rect 23234 34756 23276 34796
rect 23316 34756 23358 34796
rect 23398 34756 23440 34796
rect 23112 34747 23480 34756
rect 27112 34796 27480 34805
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27112 34747 27480 34756
rect 31112 34796 31480 34805
rect 31152 34756 31194 34796
rect 31234 34756 31276 34796
rect 31316 34756 31358 34796
rect 31398 34756 31440 34796
rect 31112 34747 31480 34756
rect 35112 34796 35480 34805
rect 35152 34756 35194 34796
rect 35234 34756 35276 34796
rect 35316 34756 35358 34796
rect 35398 34756 35440 34796
rect 35112 34747 35480 34756
rect 39112 34796 39480 34805
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39112 34747 39480 34756
rect 43112 34796 43480 34805
rect 43152 34756 43194 34796
rect 43234 34756 43276 34796
rect 43316 34756 43358 34796
rect 43398 34756 43440 34796
rect 43112 34747 43480 34756
rect 47112 34796 47480 34805
rect 47152 34756 47194 34796
rect 47234 34756 47276 34796
rect 47316 34756 47358 34796
rect 47398 34756 47440 34796
rect 47112 34747 47480 34756
rect 51112 34796 51480 34805
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51112 34747 51480 34756
rect 55112 34796 55480 34805
rect 55152 34756 55194 34796
rect 55234 34756 55276 34796
rect 55316 34756 55358 34796
rect 55398 34756 55440 34796
rect 55112 34747 55480 34756
rect 59112 34796 59480 34805
rect 59152 34756 59194 34796
rect 59234 34756 59276 34796
rect 59316 34756 59358 34796
rect 59398 34756 59440 34796
rect 59112 34747 59480 34756
rect 63112 34796 63480 34805
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63112 34747 63480 34756
rect 67112 34796 67480 34805
rect 67152 34756 67194 34796
rect 67234 34756 67276 34796
rect 67316 34756 67358 34796
rect 67398 34756 67440 34796
rect 67112 34747 67480 34756
rect 71112 34796 71480 34805
rect 71152 34756 71194 34796
rect 71234 34756 71276 34796
rect 71316 34756 71358 34796
rect 71398 34756 71440 34796
rect 71112 34747 71480 34756
rect 75112 34796 75480 34805
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75112 34747 75480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 8352 34040 8720 34049
rect 8392 34000 8434 34040
rect 8474 34000 8516 34040
rect 8556 34000 8598 34040
rect 8638 34000 8680 34040
rect 8352 33991 8720 34000
rect 12352 34040 12720 34049
rect 12392 34000 12434 34040
rect 12474 34000 12516 34040
rect 12556 34000 12598 34040
rect 12638 34000 12680 34040
rect 12352 33991 12720 34000
rect 16352 34040 16720 34049
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16352 33991 16720 34000
rect 20352 34040 20720 34049
rect 20392 34000 20434 34040
rect 20474 34000 20516 34040
rect 20556 34000 20598 34040
rect 20638 34000 20680 34040
rect 20352 33991 20720 34000
rect 24352 34040 24720 34049
rect 24392 34000 24434 34040
rect 24474 34000 24516 34040
rect 24556 34000 24598 34040
rect 24638 34000 24680 34040
rect 24352 33991 24720 34000
rect 28352 34040 28720 34049
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28352 33991 28720 34000
rect 32352 34040 32720 34049
rect 32392 34000 32434 34040
rect 32474 34000 32516 34040
rect 32556 34000 32598 34040
rect 32638 34000 32680 34040
rect 32352 33991 32720 34000
rect 36352 34040 36720 34049
rect 36392 34000 36434 34040
rect 36474 34000 36516 34040
rect 36556 34000 36598 34040
rect 36638 34000 36680 34040
rect 36352 33991 36720 34000
rect 40352 34040 40720 34049
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40352 33991 40720 34000
rect 44352 34040 44720 34049
rect 44392 34000 44434 34040
rect 44474 34000 44516 34040
rect 44556 34000 44598 34040
rect 44638 34000 44680 34040
rect 44352 33991 44720 34000
rect 48352 34040 48720 34049
rect 48392 34000 48434 34040
rect 48474 34000 48516 34040
rect 48556 34000 48598 34040
rect 48638 34000 48680 34040
rect 48352 33991 48720 34000
rect 52352 34040 52720 34049
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52352 33991 52720 34000
rect 56352 34040 56720 34049
rect 56392 34000 56434 34040
rect 56474 34000 56516 34040
rect 56556 34000 56598 34040
rect 56638 34000 56680 34040
rect 56352 33991 56720 34000
rect 60352 34040 60720 34049
rect 60392 34000 60434 34040
rect 60474 34000 60516 34040
rect 60556 34000 60598 34040
rect 60638 34000 60680 34040
rect 60352 33991 60720 34000
rect 64352 34040 64720 34049
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64352 33991 64720 34000
rect 68352 34040 68720 34049
rect 68392 34000 68434 34040
rect 68474 34000 68516 34040
rect 68556 34000 68598 34040
rect 68638 34000 68680 34040
rect 68352 33991 68720 34000
rect 72352 34040 72720 34049
rect 72392 34000 72434 34040
rect 72474 34000 72516 34040
rect 72556 34000 72598 34040
rect 72638 34000 72680 34040
rect 72352 33991 72720 34000
rect 76352 34040 76720 34049
rect 76392 34000 76434 34040
rect 76474 34000 76516 34040
rect 76556 34000 76598 34040
rect 76638 34000 76680 34040
rect 76352 33991 76720 34000
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 7112 33284 7480 33293
rect 7152 33244 7194 33284
rect 7234 33244 7276 33284
rect 7316 33244 7358 33284
rect 7398 33244 7440 33284
rect 7112 33235 7480 33244
rect 11112 33284 11480 33293
rect 11152 33244 11194 33284
rect 11234 33244 11276 33284
rect 11316 33244 11358 33284
rect 11398 33244 11440 33284
rect 11112 33235 11480 33244
rect 15112 33284 15480 33293
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15112 33235 15480 33244
rect 19112 33284 19480 33293
rect 19152 33244 19194 33284
rect 19234 33244 19276 33284
rect 19316 33244 19358 33284
rect 19398 33244 19440 33284
rect 19112 33235 19480 33244
rect 23112 33284 23480 33293
rect 23152 33244 23194 33284
rect 23234 33244 23276 33284
rect 23316 33244 23358 33284
rect 23398 33244 23440 33284
rect 23112 33235 23480 33244
rect 27112 33284 27480 33293
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27112 33235 27480 33244
rect 31112 33284 31480 33293
rect 31152 33244 31194 33284
rect 31234 33244 31276 33284
rect 31316 33244 31358 33284
rect 31398 33244 31440 33284
rect 31112 33235 31480 33244
rect 35112 33284 35480 33293
rect 35152 33244 35194 33284
rect 35234 33244 35276 33284
rect 35316 33244 35358 33284
rect 35398 33244 35440 33284
rect 35112 33235 35480 33244
rect 39112 33284 39480 33293
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39112 33235 39480 33244
rect 43112 33284 43480 33293
rect 43152 33244 43194 33284
rect 43234 33244 43276 33284
rect 43316 33244 43358 33284
rect 43398 33244 43440 33284
rect 43112 33235 43480 33244
rect 47112 33284 47480 33293
rect 47152 33244 47194 33284
rect 47234 33244 47276 33284
rect 47316 33244 47358 33284
rect 47398 33244 47440 33284
rect 47112 33235 47480 33244
rect 51112 33284 51480 33293
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51112 33235 51480 33244
rect 55112 33284 55480 33293
rect 55152 33244 55194 33284
rect 55234 33244 55276 33284
rect 55316 33244 55358 33284
rect 55398 33244 55440 33284
rect 55112 33235 55480 33244
rect 59112 33284 59480 33293
rect 59152 33244 59194 33284
rect 59234 33244 59276 33284
rect 59316 33244 59358 33284
rect 59398 33244 59440 33284
rect 59112 33235 59480 33244
rect 63112 33284 63480 33293
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63112 33235 63480 33244
rect 67112 33284 67480 33293
rect 67152 33244 67194 33284
rect 67234 33244 67276 33284
rect 67316 33244 67358 33284
rect 67398 33244 67440 33284
rect 67112 33235 67480 33244
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 8352 32528 8720 32537
rect 8392 32488 8434 32528
rect 8474 32488 8516 32528
rect 8556 32488 8598 32528
rect 8638 32488 8680 32528
rect 8352 32479 8720 32488
rect 12352 32528 12720 32537
rect 12392 32488 12434 32528
rect 12474 32488 12516 32528
rect 12556 32488 12598 32528
rect 12638 32488 12680 32528
rect 12352 32479 12720 32488
rect 16352 32528 16720 32537
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16352 32479 16720 32488
rect 20352 32528 20720 32537
rect 20392 32488 20434 32528
rect 20474 32488 20516 32528
rect 20556 32488 20598 32528
rect 20638 32488 20680 32528
rect 20352 32479 20720 32488
rect 24352 32528 24720 32537
rect 24392 32488 24434 32528
rect 24474 32488 24516 32528
rect 24556 32488 24598 32528
rect 24638 32488 24680 32528
rect 24352 32479 24720 32488
rect 28352 32528 28720 32537
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28352 32479 28720 32488
rect 32352 32528 32720 32537
rect 32392 32488 32434 32528
rect 32474 32488 32516 32528
rect 32556 32488 32598 32528
rect 32638 32488 32680 32528
rect 32352 32479 32720 32488
rect 36352 32528 36720 32537
rect 36392 32488 36434 32528
rect 36474 32488 36516 32528
rect 36556 32488 36598 32528
rect 36638 32488 36680 32528
rect 36352 32479 36720 32488
rect 40352 32528 40720 32537
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40352 32479 40720 32488
rect 44352 32528 44720 32537
rect 44392 32488 44434 32528
rect 44474 32488 44516 32528
rect 44556 32488 44598 32528
rect 44638 32488 44680 32528
rect 44352 32479 44720 32488
rect 48352 32528 48720 32537
rect 48392 32488 48434 32528
rect 48474 32488 48516 32528
rect 48556 32488 48598 32528
rect 48638 32488 48680 32528
rect 48352 32479 48720 32488
rect 52352 32528 52720 32537
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52352 32479 52720 32488
rect 56352 32528 56720 32537
rect 56392 32488 56434 32528
rect 56474 32488 56516 32528
rect 56556 32488 56598 32528
rect 56638 32488 56680 32528
rect 56352 32479 56720 32488
rect 60352 32528 60720 32537
rect 60392 32488 60434 32528
rect 60474 32488 60516 32528
rect 60556 32488 60598 32528
rect 60638 32488 60680 32528
rect 60352 32479 60720 32488
rect 64352 32528 64720 32537
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64352 32479 64720 32488
rect 68352 32528 68720 32537
rect 68392 32488 68434 32528
rect 68474 32488 68516 32528
rect 68556 32488 68598 32528
rect 68638 32488 68680 32528
rect 68352 32479 68720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 7112 31772 7480 31781
rect 7152 31732 7194 31772
rect 7234 31732 7276 31772
rect 7316 31732 7358 31772
rect 7398 31732 7440 31772
rect 7112 31723 7480 31732
rect 11112 31772 11480 31781
rect 11152 31732 11194 31772
rect 11234 31732 11276 31772
rect 11316 31732 11358 31772
rect 11398 31732 11440 31772
rect 11112 31723 11480 31732
rect 15112 31772 15480 31781
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15112 31723 15480 31732
rect 19112 31772 19480 31781
rect 19152 31732 19194 31772
rect 19234 31732 19276 31772
rect 19316 31732 19358 31772
rect 19398 31732 19440 31772
rect 19112 31723 19480 31732
rect 23112 31772 23480 31781
rect 23152 31732 23194 31772
rect 23234 31732 23276 31772
rect 23316 31732 23358 31772
rect 23398 31732 23440 31772
rect 23112 31723 23480 31732
rect 27112 31772 27480 31781
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27112 31723 27480 31732
rect 31112 31772 31480 31781
rect 31152 31732 31194 31772
rect 31234 31732 31276 31772
rect 31316 31732 31358 31772
rect 31398 31732 31440 31772
rect 31112 31723 31480 31732
rect 35112 31772 35480 31781
rect 35152 31732 35194 31772
rect 35234 31732 35276 31772
rect 35316 31732 35358 31772
rect 35398 31732 35440 31772
rect 35112 31723 35480 31732
rect 39112 31772 39480 31781
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39112 31723 39480 31732
rect 43112 31772 43480 31781
rect 43152 31732 43194 31772
rect 43234 31732 43276 31772
rect 43316 31732 43358 31772
rect 43398 31732 43440 31772
rect 43112 31723 43480 31732
rect 47112 31772 47480 31781
rect 47152 31732 47194 31772
rect 47234 31732 47276 31772
rect 47316 31732 47358 31772
rect 47398 31732 47440 31772
rect 47112 31723 47480 31732
rect 51112 31772 51480 31781
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51112 31723 51480 31732
rect 55112 31772 55480 31781
rect 55152 31732 55194 31772
rect 55234 31732 55276 31772
rect 55316 31732 55358 31772
rect 55398 31732 55440 31772
rect 55112 31723 55480 31732
rect 59112 31772 59480 31781
rect 59152 31732 59194 31772
rect 59234 31732 59276 31772
rect 59316 31732 59358 31772
rect 59398 31732 59440 31772
rect 59112 31723 59480 31732
rect 63112 31772 63480 31781
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63112 31723 63480 31732
rect 67112 31772 67480 31781
rect 67152 31732 67194 31772
rect 67234 31732 67276 31772
rect 67316 31732 67358 31772
rect 67398 31732 67440 31772
rect 67112 31723 67480 31732
rect 76780 31520 76820 35680
rect 85228 35720 85268 35729
rect 80352 35552 80720 35561
rect 80392 35512 80434 35552
rect 80474 35512 80516 35552
rect 80556 35512 80598 35552
rect 80638 35512 80680 35552
rect 80352 35503 80720 35512
rect 84352 35552 84720 35561
rect 84392 35512 84434 35552
rect 84474 35512 84516 35552
rect 84556 35512 84598 35552
rect 84638 35512 84680 35552
rect 84352 35503 84720 35512
rect 79112 34796 79480 34805
rect 79152 34756 79194 34796
rect 79234 34756 79276 34796
rect 79316 34756 79358 34796
rect 79398 34756 79440 34796
rect 79112 34747 79480 34756
rect 83112 34796 83480 34805
rect 83152 34756 83194 34796
rect 83234 34756 83276 34796
rect 83316 34756 83358 34796
rect 83398 34756 83440 34796
rect 83112 34747 83480 34756
rect 80236 34712 80276 34721
rect 80236 33788 80276 34672
rect 80352 34040 80720 34049
rect 80392 34000 80434 34040
rect 80474 34000 80516 34040
rect 80556 34000 80598 34040
rect 80638 34000 80680 34040
rect 80352 33991 80720 34000
rect 84352 34040 84720 34049
rect 84392 34000 84434 34040
rect 84474 34000 84516 34040
rect 84556 34000 84598 34040
rect 84638 34000 84680 34040
rect 84352 33991 84720 34000
rect 80236 33739 80276 33748
rect 76780 31471 76820 31480
rect 85228 31520 85268 35680
rect 92236 35720 92276 35729
rect 88352 35552 88720 35561
rect 88392 35512 88434 35552
rect 88474 35512 88516 35552
rect 88556 35512 88598 35552
rect 88638 35512 88680 35552
rect 88352 35503 88720 35512
rect 89932 35300 89972 35309
rect 86667 34964 86709 34973
rect 86667 34924 86668 34964
rect 86708 34924 86709 34964
rect 86667 34915 86709 34924
rect 86956 34964 86996 34973
rect 86668 34830 86708 34915
rect 85228 31471 85268 31480
rect 86860 34628 86900 34637
rect 86860 31520 86900 34588
rect 86956 31604 86996 34924
rect 87112 34796 87480 34805
rect 87152 34756 87194 34796
rect 87234 34756 87276 34796
rect 87316 34756 87358 34796
rect 87398 34756 87440 34796
rect 87112 34747 87480 34756
rect 88352 34040 88720 34049
rect 88392 34000 88434 34040
rect 88474 34000 88516 34040
rect 88556 34000 88598 34040
rect 88638 34000 88680 34040
rect 88352 33991 88720 34000
rect 86956 31555 86996 31564
rect 86860 31471 86900 31480
rect 89932 31520 89972 35260
rect 91112 34796 91480 34805
rect 91152 34756 91194 34796
rect 91234 34756 91276 34796
rect 91316 34756 91358 34796
rect 91398 34756 91440 34796
rect 91112 34747 91480 34756
rect 89932 31471 89972 31480
rect 92236 31520 92276 35680
rect 92352 35552 92720 35561
rect 92392 35512 92434 35552
rect 92474 35512 92516 35552
rect 92556 35512 92598 35552
rect 92638 35512 92680 35552
rect 92352 35503 92720 35512
rect 96352 35552 96720 35561
rect 96392 35512 96434 35552
rect 96474 35512 96516 35552
rect 96556 35512 96598 35552
rect 96638 35512 96680 35552
rect 96352 35503 96720 35512
rect 95112 34796 95480 34805
rect 95152 34756 95194 34796
rect 95234 34756 95276 34796
rect 95316 34756 95358 34796
rect 95398 34756 95440 34796
rect 95112 34747 95480 34756
rect 99112 34796 99480 34805
rect 99152 34756 99194 34796
rect 99234 34756 99276 34796
rect 99316 34756 99358 34796
rect 99398 34756 99440 34796
rect 99112 34747 99480 34756
rect 92352 34040 92720 34049
rect 92392 34000 92434 34040
rect 92474 34000 92516 34040
rect 92556 34000 92598 34040
rect 92638 34000 92680 34040
rect 92352 33991 92720 34000
rect 96352 34040 96720 34049
rect 96392 34000 96434 34040
rect 96474 34000 96516 34040
rect 96556 34000 96598 34040
rect 96638 34000 96680 34040
rect 96352 33991 96720 34000
rect 92236 31471 92276 31480
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 8352 31016 8720 31025
rect 8392 30976 8434 31016
rect 8474 30976 8516 31016
rect 8556 30976 8598 31016
rect 8638 30976 8680 31016
rect 8352 30967 8720 30976
rect 12352 31016 12720 31025
rect 12392 30976 12434 31016
rect 12474 30976 12516 31016
rect 12556 30976 12598 31016
rect 12638 30976 12680 31016
rect 12352 30967 12720 30976
rect 16352 31016 16720 31025
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16352 30967 16720 30976
rect 20352 31016 20720 31025
rect 20392 30976 20434 31016
rect 20474 30976 20516 31016
rect 20556 30976 20598 31016
rect 20638 30976 20680 31016
rect 20352 30967 20720 30976
rect 24352 31016 24720 31025
rect 24392 30976 24434 31016
rect 24474 30976 24516 31016
rect 24556 30976 24598 31016
rect 24638 30976 24680 31016
rect 24352 30967 24720 30976
rect 28352 31016 28720 31025
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28352 30967 28720 30976
rect 32352 31016 32720 31025
rect 32392 30976 32434 31016
rect 32474 30976 32516 31016
rect 32556 30976 32598 31016
rect 32638 30976 32680 31016
rect 32352 30967 32720 30976
rect 36352 31016 36720 31025
rect 36392 30976 36434 31016
rect 36474 30976 36516 31016
rect 36556 30976 36598 31016
rect 36638 30976 36680 31016
rect 36352 30967 36720 30976
rect 40352 31016 40720 31025
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40352 30967 40720 30976
rect 44352 31016 44720 31025
rect 44392 30976 44434 31016
rect 44474 30976 44516 31016
rect 44556 30976 44598 31016
rect 44638 30976 44680 31016
rect 44352 30967 44720 30976
rect 48352 31016 48720 31025
rect 48392 30976 48434 31016
rect 48474 30976 48516 31016
rect 48556 30976 48598 31016
rect 48638 30976 48680 31016
rect 48352 30967 48720 30976
rect 52352 31016 52720 31025
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52352 30967 52720 30976
rect 56352 31016 56720 31025
rect 56392 30976 56434 31016
rect 56474 30976 56516 31016
rect 56556 30976 56598 31016
rect 56638 30976 56680 31016
rect 56352 30967 56720 30976
rect 60352 31016 60720 31025
rect 60392 30976 60434 31016
rect 60474 30976 60516 31016
rect 60556 30976 60598 31016
rect 60638 30976 60680 31016
rect 60352 30967 60720 30976
rect 64352 31016 64720 31025
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64352 30967 64720 30976
rect 68352 31016 68720 31025
rect 68392 30976 68434 31016
rect 68474 30976 68516 31016
rect 68556 30976 68598 31016
rect 68638 30976 68680 31016
rect 68352 30967 68720 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 7112 30260 7480 30269
rect 7152 30220 7194 30260
rect 7234 30220 7276 30260
rect 7316 30220 7358 30260
rect 7398 30220 7440 30260
rect 7112 30211 7480 30220
rect 11112 30260 11480 30269
rect 11152 30220 11194 30260
rect 11234 30220 11276 30260
rect 11316 30220 11358 30260
rect 11398 30220 11440 30260
rect 11112 30211 11480 30220
rect 15112 30260 15480 30269
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15112 30211 15480 30220
rect 19112 30260 19480 30269
rect 19152 30220 19194 30260
rect 19234 30220 19276 30260
rect 19316 30220 19358 30260
rect 19398 30220 19440 30260
rect 19112 30211 19480 30220
rect 23112 30260 23480 30269
rect 23152 30220 23194 30260
rect 23234 30220 23276 30260
rect 23316 30220 23358 30260
rect 23398 30220 23440 30260
rect 23112 30211 23480 30220
rect 27112 30260 27480 30269
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27112 30211 27480 30220
rect 31112 30260 31480 30269
rect 31152 30220 31194 30260
rect 31234 30220 31276 30260
rect 31316 30220 31358 30260
rect 31398 30220 31440 30260
rect 31112 30211 31480 30220
rect 35112 30260 35480 30269
rect 35152 30220 35194 30260
rect 35234 30220 35276 30260
rect 35316 30220 35358 30260
rect 35398 30220 35440 30260
rect 35112 30211 35480 30220
rect 39112 30260 39480 30269
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39112 30211 39480 30220
rect 43112 30260 43480 30269
rect 43152 30220 43194 30260
rect 43234 30220 43276 30260
rect 43316 30220 43358 30260
rect 43398 30220 43440 30260
rect 43112 30211 43480 30220
rect 47112 30260 47480 30269
rect 47152 30220 47194 30260
rect 47234 30220 47276 30260
rect 47316 30220 47358 30260
rect 47398 30220 47440 30260
rect 47112 30211 47480 30220
rect 51112 30260 51480 30269
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51112 30211 51480 30220
rect 55112 30260 55480 30269
rect 55152 30220 55194 30260
rect 55234 30220 55276 30260
rect 55316 30220 55358 30260
rect 55398 30220 55440 30260
rect 55112 30211 55480 30220
rect 59112 30260 59480 30269
rect 59152 30220 59194 30260
rect 59234 30220 59276 30260
rect 59316 30220 59358 30260
rect 59398 30220 59440 30260
rect 59112 30211 59480 30220
rect 63112 30260 63480 30269
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63112 30211 63480 30220
rect 67112 30260 67480 30269
rect 67152 30220 67194 30260
rect 67234 30220 67276 30260
rect 67316 30220 67358 30260
rect 67398 30220 67440 30260
rect 67112 30211 67480 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 8352 29504 8720 29513
rect 8392 29464 8434 29504
rect 8474 29464 8516 29504
rect 8556 29464 8598 29504
rect 8638 29464 8680 29504
rect 8352 29455 8720 29464
rect 12352 29504 12720 29513
rect 12392 29464 12434 29504
rect 12474 29464 12516 29504
rect 12556 29464 12598 29504
rect 12638 29464 12680 29504
rect 12352 29455 12720 29464
rect 16352 29504 16720 29513
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16352 29455 16720 29464
rect 20352 29504 20720 29513
rect 20392 29464 20434 29504
rect 20474 29464 20516 29504
rect 20556 29464 20598 29504
rect 20638 29464 20680 29504
rect 20352 29455 20720 29464
rect 24352 29504 24720 29513
rect 24392 29464 24434 29504
rect 24474 29464 24516 29504
rect 24556 29464 24598 29504
rect 24638 29464 24680 29504
rect 24352 29455 24720 29464
rect 28352 29504 28720 29513
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28352 29455 28720 29464
rect 32352 29504 32720 29513
rect 32392 29464 32434 29504
rect 32474 29464 32516 29504
rect 32556 29464 32598 29504
rect 32638 29464 32680 29504
rect 32352 29455 32720 29464
rect 36352 29504 36720 29513
rect 36392 29464 36434 29504
rect 36474 29464 36516 29504
rect 36556 29464 36598 29504
rect 36638 29464 36680 29504
rect 36352 29455 36720 29464
rect 40352 29504 40720 29513
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40352 29455 40720 29464
rect 44352 29504 44720 29513
rect 44392 29464 44434 29504
rect 44474 29464 44516 29504
rect 44556 29464 44598 29504
rect 44638 29464 44680 29504
rect 44352 29455 44720 29464
rect 48352 29504 48720 29513
rect 48392 29464 48434 29504
rect 48474 29464 48516 29504
rect 48556 29464 48598 29504
rect 48638 29464 48680 29504
rect 48352 29455 48720 29464
rect 52352 29504 52720 29513
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52352 29455 52720 29464
rect 56352 29504 56720 29513
rect 56392 29464 56434 29504
rect 56474 29464 56516 29504
rect 56556 29464 56598 29504
rect 56638 29464 56680 29504
rect 56352 29455 56720 29464
rect 60352 29504 60720 29513
rect 60392 29464 60434 29504
rect 60474 29464 60516 29504
rect 60556 29464 60598 29504
rect 60638 29464 60680 29504
rect 60352 29455 60720 29464
rect 64352 29504 64720 29513
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64352 29455 64720 29464
rect 68352 29504 68720 29513
rect 68392 29464 68434 29504
rect 68474 29464 68516 29504
rect 68556 29464 68598 29504
rect 68638 29464 68680 29504
rect 68352 29455 68720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 7112 28748 7480 28757
rect 7152 28708 7194 28748
rect 7234 28708 7276 28748
rect 7316 28708 7358 28748
rect 7398 28708 7440 28748
rect 7112 28699 7480 28708
rect 11112 28748 11480 28757
rect 11152 28708 11194 28748
rect 11234 28708 11276 28748
rect 11316 28708 11358 28748
rect 11398 28708 11440 28748
rect 11112 28699 11480 28708
rect 15112 28748 15480 28757
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15112 28699 15480 28708
rect 19112 28748 19480 28757
rect 19152 28708 19194 28748
rect 19234 28708 19276 28748
rect 19316 28708 19358 28748
rect 19398 28708 19440 28748
rect 19112 28699 19480 28708
rect 23112 28748 23480 28757
rect 23152 28708 23194 28748
rect 23234 28708 23276 28748
rect 23316 28708 23358 28748
rect 23398 28708 23440 28748
rect 23112 28699 23480 28708
rect 27112 28748 27480 28757
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27112 28699 27480 28708
rect 31112 28748 31480 28757
rect 31152 28708 31194 28748
rect 31234 28708 31276 28748
rect 31316 28708 31358 28748
rect 31398 28708 31440 28748
rect 31112 28699 31480 28708
rect 35112 28748 35480 28757
rect 35152 28708 35194 28748
rect 35234 28708 35276 28748
rect 35316 28708 35358 28748
rect 35398 28708 35440 28748
rect 35112 28699 35480 28708
rect 39112 28748 39480 28757
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39112 28699 39480 28708
rect 43112 28748 43480 28757
rect 43152 28708 43194 28748
rect 43234 28708 43276 28748
rect 43316 28708 43358 28748
rect 43398 28708 43440 28748
rect 43112 28699 43480 28708
rect 47112 28748 47480 28757
rect 47152 28708 47194 28748
rect 47234 28708 47276 28748
rect 47316 28708 47358 28748
rect 47398 28708 47440 28748
rect 47112 28699 47480 28708
rect 51112 28748 51480 28757
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51112 28699 51480 28708
rect 55112 28748 55480 28757
rect 55152 28708 55194 28748
rect 55234 28708 55276 28748
rect 55316 28708 55358 28748
rect 55398 28708 55440 28748
rect 55112 28699 55480 28708
rect 59112 28748 59480 28757
rect 59152 28708 59194 28748
rect 59234 28708 59276 28748
rect 59316 28708 59358 28748
rect 59398 28708 59440 28748
rect 59112 28699 59480 28708
rect 63112 28748 63480 28757
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63112 28699 63480 28708
rect 67112 28748 67480 28757
rect 67152 28708 67194 28748
rect 67234 28708 67276 28748
rect 67316 28708 67358 28748
rect 67398 28708 67440 28748
rect 67112 28699 67480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 8352 27992 8720 28001
rect 8392 27952 8434 27992
rect 8474 27952 8516 27992
rect 8556 27952 8598 27992
rect 8638 27952 8680 27992
rect 8352 27943 8720 27952
rect 12352 27992 12720 28001
rect 12392 27952 12434 27992
rect 12474 27952 12516 27992
rect 12556 27952 12598 27992
rect 12638 27952 12680 27992
rect 12352 27943 12720 27952
rect 16352 27992 16720 28001
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16352 27943 16720 27952
rect 20352 27992 20720 28001
rect 20392 27952 20434 27992
rect 20474 27952 20516 27992
rect 20556 27952 20598 27992
rect 20638 27952 20680 27992
rect 20352 27943 20720 27952
rect 24352 27992 24720 28001
rect 24392 27952 24434 27992
rect 24474 27952 24516 27992
rect 24556 27952 24598 27992
rect 24638 27952 24680 27992
rect 24352 27943 24720 27952
rect 28352 27992 28720 28001
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28352 27943 28720 27952
rect 32352 27992 32720 28001
rect 32392 27952 32434 27992
rect 32474 27952 32516 27992
rect 32556 27952 32598 27992
rect 32638 27952 32680 27992
rect 32352 27943 32720 27952
rect 36352 27992 36720 28001
rect 36392 27952 36434 27992
rect 36474 27952 36516 27992
rect 36556 27952 36598 27992
rect 36638 27952 36680 27992
rect 36352 27943 36720 27952
rect 40352 27992 40720 28001
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40352 27943 40720 27952
rect 44352 27992 44720 28001
rect 44392 27952 44434 27992
rect 44474 27952 44516 27992
rect 44556 27952 44598 27992
rect 44638 27952 44680 27992
rect 44352 27943 44720 27952
rect 48352 27992 48720 28001
rect 48392 27952 48434 27992
rect 48474 27952 48516 27992
rect 48556 27952 48598 27992
rect 48638 27952 48680 27992
rect 48352 27943 48720 27952
rect 52352 27992 52720 28001
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52352 27943 52720 27952
rect 56352 27992 56720 28001
rect 56392 27952 56434 27992
rect 56474 27952 56516 27992
rect 56556 27952 56598 27992
rect 56638 27952 56680 27992
rect 56352 27943 56720 27952
rect 60352 27992 60720 28001
rect 60392 27952 60434 27992
rect 60474 27952 60516 27992
rect 60556 27952 60598 27992
rect 60638 27952 60680 27992
rect 60352 27943 60720 27952
rect 64352 27992 64720 28001
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64352 27943 64720 27952
rect 68352 27992 68720 28001
rect 68392 27952 68434 27992
rect 68474 27952 68516 27992
rect 68556 27952 68598 27992
rect 68638 27952 68680 27992
rect 68352 27943 68720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 7112 27236 7480 27245
rect 7152 27196 7194 27236
rect 7234 27196 7276 27236
rect 7316 27196 7358 27236
rect 7398 27196 7440 27236
rect 7112 27187 7480 27196
rect 11112 27236 11480 27245
rect 11152 27196 11194 27236
rect 11234 27196 11276 27236
rect 11316 27196 11358 27236
rect 11398 27196 11440 27236
rect 11112 27187 11480 27196
rect 15112 27236 15480 27245
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15112 27187 15480 27196
rect 19112 27236 19480 27245
rect 19152 27196 19194 27236
rect 19234 27196 19276 27236
rect 19316 27196 19358 27236
rect 19398 27196 19440 27236
rect 19112 27187 19480 27196
rect 23112 27236 23480 27245
rect 23152 27196 23194 27236
rect 23234 27196 23276 27236
rect 23316 27196 23358 27236
rect 23398 27196 23440 27236
rect 23112 27187 23480 27196
rect 27112 27236 27480 27245
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27112 27187 27480 27196
rect 31112 27236 31480 27245
rect 31152 27196 31194 27236
rect 31234 27196 31276 27236
rect 31316 27196 31358 27236
rect 31398 27196 31440 27236
rect 31112 27187 31480 27196
rect 35112 27236 35480 27245
rect 35152 27196 35194 27236
rect 35234 27196 35276 27236
rect 35316 27196 35358 27236
rect 35398 27196 35440 27236
rect 35112 27187 35480 27196
rect 39112 27236 39480 27245
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39112 27187 39480 27196
rect 43112 27236 43480 27245
rect 43152 27196 43194 27236
rect 43234 27196 43276 27236
rect 43316 27196 43358 27236
rect 43398 27196 43440 27236
rect 43112 27187 43480 27196
rect 47112 27236 47480 27245
rect 47152 27196 47194 27236
rect 47234 27196 47276 27236
rect 47316 27196 47358 27236
rect 47398 27196 47440 27236
rect 47112 27187 47480 27196
rect 51112 27236 51480 27245
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51112 27187 51480 27196
rect 55112 27236 55480 27245
rect 55152 27196 55194 27236
rect 55234 27196 55276 27236
rect 55316 27196 55358 27236
rect 55398 27196 55440 27236
rect 55112 27187 55480 27196
rect 59112 27236 59480 27245
rect 59152 27196 59194 27236
rect 59234 27196 59276 27236
rect 59316 27196 59358 27236
rect 59398 27196 59440 27236
rect 59112 27187 59480 27196
rect 63112 27236 63480 27245
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63112 27187 63480 27196
rect 67112 27236 67480 27245
rect 67152 27196 67194 27236
rect 67234 27196 67276 27236
rect 67316 27196 67358 27236
rect 67398 27196 67440 27236
rect 67112 27187 67480 27196
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 8352 26480 8720 26489
rect 8392 26440 8434 26480
rect 8474 26440 8516 26480
rect 8556 26440 8598 26480
rect 8638 26440 8680 26480
rect 8352 26431 8720 26440
rect 12352 26480 12720 26489
rect 12392 26440 12434 26480
rect 12474 26440 12516 26480
rect 12556 26440 12598 26480
rect 12638 26440 12680 26480
rect 12352 26431 12720 26440
rect 16352 26480 16720 26489
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16352 26431 16720 26440
rect 20352 26480 20720 26489
rect 20392 26440 20434 26480
rect 20474 26440 20516 26480
rect 20556 26440 20598 26480
rect 20638 26440 20680 26480
rect 20352 26431 20720 26440
rect 24352 26480 24720 26489
rect 24392 26440 24434 26480
rect 24474 26440 24516 26480
rect 24556 26440 24598 26480
rect 24638 26440 24680 26480
rect 24352 26431 24720 26440
rect 28352 26480 28720 26489
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28352 26431 28720 26440
rect 32352 26480 32720 26489
rect 32392 26440 32434 26480
rect 32474 26440 32516 26480
rect 32556 26440 32598 26480
rect 32638 26440 32680 26480
rect 32352 26431 32720 26440
rect 36352 26480 36720 26489
rect 36392 26440 36434 26480
rect 36474 26440 36516 26480
rect 36556 26440 36598 26480
rect 36638 26440 36680 26480
rect 36352 26431 36720 26440
rect 40352 26480 40720 26489
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40352 26431 40720 26440
rect 44352 26480 44720 26489
rect 44392 26440 44434 26480
rect 44474 26440 44516 26480
rect 44556 26440 44598 26480
rect 44638 26440 44680 26480
rect 44352 26431 44720 26440
rect 48352 26480 48720 26489
rect 48392 26440 48434 26480
rect 48474 26440 48516 26480
rect 48556 26440 48598 26480
rect 48638 26440 48680 26480
rect 48352 26431 48720 26440
rect 52352 26480 52720 26489
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52352 26431 52720 26440
rect 56352 26480 56720 26489
rect 56392 26440 56434 26480
rect 56474 26440 56516 26480
rect 56556 26440 56598 26480
rect 56638 26440 56680 26480
rect 56352 26431 56720 26440
rect 60352 26480 60720 26489
rect 60392 26440 60434 26480
rect 60474 26440 60516 26480
rect 60556 26440 60598 26480
rect 60638 26440 60680 26480
rect 60352 26431 60720 26440
rect 64352 26480 64720 26489
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64352 26431 64720 26440
rect 68352 26480 68720 26489
rect 68392 26440 68434 26480
rect 68474 26440 68516 26480
rect 68556 26440 68598 26480
rect 68638 26440 68680 26480
rect 68352 26431 68720 26440
rect 71788 26060 71828 26069
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 7112 25724 7480 25733
rect 7152 25684 7194 25724
rect 7234 25684 7276 25724
rect 7316 25684 7358 25724
rect 7398 25684 7440 25724
rect 7112 25675 7480 25684
rect 11112 25724 11480 25733
rect 11152 25684 11194 25724
rect 11234 25684 11276 25724
rect 11316 25684 11358 25724
rect 11398 25684 11440 25724
rect 11112 25675 11480 25684
rect 15112 25724 15480 25733
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15112 25675 15480 25684
rect 19112 25724 19480 25733
rect 19152 25684 19194 25724
rect 19234 25684 19276 25724
rect 19316 25684 19358 25724
rect 19398 25684 19440 25724
rect 19112 25675 19480 25684
rect 23112 25724 23480 25733
rect 23152 25684 23194 25724
rect 23234 25684 23276 25724
rect 23316 25684 23358 25724
rect 23398 25684 23440 25724
rect 23112 25675 23480 25684
rect 27112 25724 27480 25733
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27112 25675 27480 25684
rect 31112 25724 31480 25733
rect 31152 25684 31194 25724
rect 31234 25684 31276 25724
rect 31316 25684 31358 25724
rect 31398 25684 31440 25724
rect 31112 25675 31480 25684
rect 35112 25724 35480 25733
rect 35152 25684 35194 25724
rect 35234 25684 35276 25724
rect 35316 25684 35358 25724
rect 35398 25684 35440 25724
rect 35112 25675 35480 25684
rect 39112 25724 39480 25733
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39112 25675 39480 25684
rect 43112 25724 43480 25733
rect 43152 25684 43194 25724
rect 43234 25684 43276 25724
rect 43316 25684 43358 25724
rect 43398 25684 43440 25724
rect 43112 25675 43480 25684
rect 47112 25724 47480 25733
rect 47152 25684 47194 25724
rect 47234 25684 47276 25724
rect 47316 25684 47358 25724
rect 47398 25684 47440 25724
rect 47112 25675 47480 25684
rect 51112 25724 51480 25733
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51112 25675 51480 25684
rect 55112 25724 55480 25733
rect 55152 25684 55194 25724
rect 55234 25684 55276 25724
rect 55316 25684 55358 25724
rect 55398 25684 55440 25724
rect 55112 25675 55480 25684
rect 59112 25724 59480 25733
rect 59152 25684 59194 25724
rect 59234 25684 59276 25724
rect 59316 25684 59358 25724
rect 59398 25684 59440 25724
rect 59112 25675 59480 25684
rect 63112 25724 63480 25733
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63112 25675 63480 25684
rect 67112 25724 67480 25733
rect 67152 25684 67194 25724
rect 67234 25684 67276 25724
rect 67316 25684 67358 25724
rect 67398 25684 67440 25724
rect 67112 25675 67480 25684
rect 71788 25649 71828 26020
rect 71884 25976 71924 25985
rect 71884 25892 71924 25936
rect 72460 25892 72500 25901
rect 71884 25852 72460 25892
rect 72460 25843 72500 25852
rect 94924 25808 94964 25817
rect 71787 25640 71829 25649
rect 71787 25600 71788 25640
rect 71828 25600 71829 25640
rect 71787 25591 71829 25600
rect 72939 25640 72981 25649
rect 72939 25600 72940 25640
rect 72980 25600 72981 25640
rect 72939 25591 72981 25600
rect 72940 25506 72980 25591
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 8352 24968 8720 24977
rect 8392 24928 8434 24968
rect 8474 24928 8516 24968
rect 8556 24928 8598 24968
rect 8638 24928 8680 24968
rect 8352 24919 8720 24928
rect 12352 24968 12720 24977
rect 12392 24928 12434 24968
rect 12474 24928 12516 24968
rect 12556 24928 12598 24968
rect 12638 24928 12680 24968
rect 12352 24919 12720 24928
rect 16352 24968 16720 24977
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16352 24919 16720 24928
rect 20352 24968 20720 24977
rect 20392 24928 20434 24968
rect 20474 24928 20516 24968
rect 20556 24928 20598 24968
rect 20638 24928 20680 24968
rect 20352 24919 20720 24928
rect 24352 24968 24720 24977
rect 24392 24928 24434 24968
rect 24474 24928 24516 24968
rect 24556 24928 24598 24968
rect 24638 24928 24680 24968
rect 24352 24919 24720 24928
rect 28352 24968 28720 24977
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28352 24919 28720 24928
rect 32352 24968 32720 24977
rect 32392 24928 32434 24968
rect 32474 24928 32516 24968
rect 32556 24928 32598 24968
rect 32638 24928 32680 24968
rect 32352 24919 32720 24928
rect 36352 24968 36720 24977
rect 36392 24928 36434 24968
rect 36474 24928 36516 24968
rect 36556 24928 36598 24968
rect 36638 24928 36680 24968
rect 36352 24919 36720 24928
rect 40352 24968 40720 24977
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40352 24919 40720 24928
rect 44352 24968 44720 24977
rect 44392 24928 44434 24968
rect 44474 24928 44516 24968
rect 44556 24928 44598 24968
rect 44638 24928 44680 24968
rect 44352 24919 44720 24928
rect 48352 24968 48720 24977
rect 48392 24928 48434 24968
rect 48474 24928 48516 24968
rect 48556 24928 48598 24968
rect 48638 24928 48680 24968
rect 48352 24919 48720 24928
rect 52352 24968 52720 24977
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52352 24919 52720 24928
rect 56352 24968 56720 24977
rect 56392 24928 56434 24968
rect 56474 24928 56516 24968
rect 56556 24928 56598 24968
rect 56638 24928 56680 24968
rect 56352 24919 56720 24928
rect 60352 24968 60720 24977
rect 60392 24928 60434 24968
rect 60474 24928 60516 24968
rect 60556 24928 60598 24968
rect 60638 24928 60680 24968
rect 60352 24919 60720 24928
rect 64352 24968 64720 24977
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64352 24919 64720 24928
rect 68352 24968 68720 24977
rect 68392 24928 68434 24968
rect 68474 24928 68516 24968
rect 68556 24928 68598 24968
rect 68638 24928 68680 24968
rect 68352 24919 68720 24928
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 7112 24212 7480 24221
rect 7152 24172 7194 24212
rect 7234 24172 7276 24212
rect 7316 24172 7358 24212
rect 7398 24172 7440 24212
rect 7112 24163 7480 24172
rect 11112 24212 11480 24221
rect 11152 24172 11194 24212
rect 11234 24172 11276 24212
rect 11316 24172 11358 24212
rect 11398 24172 11440 24212
rect 11112 24163 11480 24172
rect 15112 24212 15480 24221
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15112 24163 15480 24172
rect 19112 24212 19480 24221
rect 19152 24172 19194 24212
rect 19234 24172 19276 24212
rect 19316 24172 19358 24212
rect 19398 24172 19440 24212
rect 19112 24163 19480 24172
rect 23112 24212 23480 24221
rect 23152 24172 23194 24212
rect 23234 24172 23276 24212
rect 23316 24172 23358 24212
rect 23398 24172 23440 24212
rect 23112 24163 23480 24172
rect 27112 24212 27480 24221
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27112 24163 27480 24172
rect 31112 24212 31480 24221
rect 31152 24172 31194 24212
rect 31234 24172 31276 24212
rect 31316 24172 31358 24212
rect 31398 24172 31440 24212
rect 31112 24163 31480 24172
rect 35112 24212 35480 24221
rect 35152 24172 35194 24212
rect 35234 24172 35276 24212
rect 35316 24172 35358 24212
rect 35398 24172 35440 24212
rect 35112 24163 35480 24172
rect 39112 24212 39480 24221
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39112 24163 39480 24172
rect 43112 24212 43480 24221
rect 43152 24172 43194 24212
rect 43234 24172 43276 24212
rect 43316 24172 43358 24212
rect 43398 24172 43440 24212
rect 43112 24163 43480 24172
rect 47112 24212 47480 24221
rect 47152 24172 47194 24212
rect 47234 24172 47276 24212
rect 47316 24172 47358 24212
rect 47398 24172 47440 24212
rect 47112 24163 47480 24172
rect 51112 24212 51480 24221
rect 51152 24172 51194 24212
rect 51234 24172 51276 24212
rect 51316 24172 51358 24212
rect 51398 24172 51440 24212
rect 51112 24163 51480 24172
rect 55112 24212 55480 24221
rect 55152 24172 55194 24212
rect 55234 24172 55276 24212
rect 55316 24172 55358 24212
rect 55398 24172 55440 24212
rect 55112 24163 55480 24172
rect 59112 24212 59480 24221
rect 59152 24172 59194 24212
rect 59234 24172 59276 24212
rect 59316 24172 59358 24212
rect 59398 24172 59440 24212
rect 59112 24163 59480 24172
rect 63112 24212 63480 24221
rect 63152 24172 63194 24212
rect 63234 24172 63276 24212
rect 63316 24172 63358 24212
rect 63398 24172 63440 24212
rect 63112 24163 63480 24172
rect 67112 24212 67480 24221
rect 67152 24172 67194 24212
rect 67234 24172 67276 24212
rect 67316 24172 67358 24212
rect 67398 24172 67440 24212
rect 67112 24163 67480 24172
rect 85420 23960 85460 23969
rect 84268 23792 84308 23801
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 8352 23456 8720 23465
rect 8392 23416 8434 23456
rect 8474 23416 8516 23456
rect 8556 23416 8598 23456
rect 8638 23416 8680 23456
rect 8352 23407 8720 23416
rect 12352 23456 12720 23465
rect 12392 23416 12434 23456
rect 12474 23416 12516 23456
rect 12556 23416 12598 23456
rect 12638 23416 12680 23456
rect 12352 23407 12720 23416
rect 16352 23456 16720 23465
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16352 23407 16720 23416
rect 20352 23456 20720 23465
rect 20392 23416 20434 23456
rect 20474 23416 20516 23456
rect 20556 23416 20598 23456
rect 20638 23416 20680 23456
rect 20352 23407 20720 23416
rect 24352 23456 24720 23465
rect 24392 23416 24434 23456
rect 24474 23416 24516 23456
rect 24556 23416 24598 23456
rect 24638 23416 24680 23456
rect 24352 23407 24720 23416
rect 28352 23456 28720 23465
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28352 23407 28720 23416
rect 32352 23456 32720 23465
rect 32392 23416 32434 23456
rect 32474 23416 32516 23456
rect 32556 23416 32598 23456
rect 32638 23416 32680 23456
rect 32352 23407 32720 23416
rect 36352 23456 36720 23465
rect 36392 23416 36434 23456
rect 36474 23416 36516 23456
rect 36556 23416 36598 23456
rect 36638 23416 36680 23456
rect 36352 23407 36720 23416
rect 40352 23456 40720 23465
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40352 23407 40720 23416
rect 44352 23456 44720 23465
rect 44392 23416 44434 23456
rect 44474 23416 44516 23456
rect 44556 23416 44598 23456
rect 44638 23416 44680 23456
rect 44352 23407 44720 23416
rect 48352 23456 48720 23465
rect 48392 23416 48434 23456
rect 48474 23416 48516 23456
rect 48556 23416 48598 23456
rect 48638 23416 48680 23456
rect 48352 23407 48720 23416
rect 52352 23456 52720 23465
rect 52392 23416 52434 23456
rect 52474 23416 52516 23456
rect 52556 23416 52598 23456
rect 52638 23416 52680 23456
rect 52352 23407 52720 23416
rect 56352 23456 56720 23465
rect 56392 23416 56434 23456
rect 56474 23416 56516 23456
rect 56556 23416 56598 23456
rect 56638 23416 56680 23456
rect 56352 23407 56720 23416
rect 60352 23456 60720 23465
rect 60392 23416 60434 23456
rect 60474 23416 60516 23456
rect 60556 23416 60598 23456
rect 60638 23416 60680 23456
rect 60352 23407 60720 23416
rect 64352 23456 64720 23465
rect 64392 23416 64434 23456
rect 64474 23416 64516 23456
rect 64556 23416 64598 23456
rect 64638 23416 64680 23456
rect 64352 23407 64720 23416
rect 68352 23456 68720 23465
rect 68392 23416 68434 23456
rect 68474 23416 68516 23456
rect 68556 23416 68598 23456
rect 68638 23416 68680 23456
rect 68352 23407 68720 23416
rect 72352 23456 72720 23465
rect 72392 23416 72434 23456
rect 72474 23416 72516 23456
rect 72556 23416 72598 23456
rect 72638 23416 72680 23456
rect 72352 23407 72720 23416
rect 76352 23456 76720 23465
rect 76392 23416 76434 23456
rect 76474 23416 76516 23456
rect 76556 23416 76598 23456
rect 76638 23416 76680 23456
rect 76352 23407 76720 23416
rect 80352 23456 80720 23465
rect 80392 23416 80434 23456
rect 80474 23416 80516 23456
rect 80556 23416 80598 23456
rect 80638 23416 80680 23456
rect 80352 23407 80720 23416
rect 83596 23288 83636 23297
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 7112 22700 7480 22709
rect 7152 22660 7194 22700
rect 7234 22660 7276 22700
rect 7316 22660 7358 22700
rect 7398 22660 7440 22700
rect 7112 22651 7480 22660
rect 11112 22700 11480 22709
rect 11152 22660 11194 22700
rect 11234 22660 11276 22700
rect 11316 22660 11358 22700
rect 11398 22660 11440 22700
rect 11112 22651 11480 22660
rect 15112 22700 15480 22709
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15112 22651 15480 22660
rect 19112 22700 19480 22709
rect 19152 22660 19194 22700
rect 19234 22660 19276 22700
rect 19316 22660 19358 22700
rect 19398 22660 19440 22700
rect 19112 22651 19480 22660
rect 23112 22700 23480 22709
rect 23152 22660 23194 22700
rect 23234 22660 23276 22700
rect 23316 22660 23358 22700
rect 23398 22660 23440 22700
rect 23112 22651 23480 22660
rect 27112 22700 27480 22709
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27112 22651 27480 22660
rect 31112 22700 31480 22709
rect 31152 22660 31194 22700
rect 31234 22660 31276 22700
rect 31316 22660 31358 22700
rect 31398 22660 31440 22700
rect 31112 22651 31480 22660
rect 35112 22700 35480 22709
rect 35152 22660 35194 22700
rect 35234 22660 35276 22700
rect 35316 22660 35358 22700
rect 35398 22660 35440 22700
rect 35112 22651 35480 22660
rect 39112 22700 39480 22709
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39112 22651 39480 22660
rect 43112 22700 43480 22709
rect 43152 22660 43194 22700
rect 43234 22660 43276 22700
rect 43316 22660 43358 22700
rect 43398 22660 43440 22700
rect 43112 22651 43480 22660
rect 47112 22700 47480 22709
rect 47152 22660 47194 22700
rect 47234 22660 47276 22700
rect 47316 22660 47358 22700
rect 47398 22660 47440 22700
rect 47112 22651 47480 22660
rect 51112 22700 51480 22709
rect 51152 22660 51194 22700
rect 51234 22660 51276 22700
rect 51316 22660 51358 22700
rect 51398 22660 51440 22700
rect 51112 22651 51480 22660
rect 55112 22700 55480 22709
rect 55152 22660 55194 22700
rect 55234 22660 55276 22700
rect 55316 22660 55358 22700
rect 55398 22660 55440 22700
rect 55112 22651 55480 22660
rect 59112 22700 59480 22709
rect 59152 22660 59194 22700
rect 59234 22660 59276 22700
rect 59316 22660 59358 22700
rect 59398 22660 59440 22700
rect 59112 22651 59480 22660
rect 63112 22700 63480 22709
rect 63152 22660 63194 22700
rect 63234 22660 63276 22700
rect 63316 22660 63358 22700
rect 63398 22660 63440 22700
rect 63112 22651 63480 22660
rect 67112 22700 67480 22709
rect 67152 22660 67194 22700
rect 67234 22660 67276 22700
rect 67316 22660 67358 22700
rect 67398 22660 67440 22700
rect 67112 22651 67480 22660
rect 71112 22700 71480 22709
rect 71152 22660 71194 22700
rect 71234 22660 71276 22700
rect 71316 22660 71358 22700
rect 71398 22660 71440 22700
rect 71112 22651 71480 22660
rect 75112 22700 75480 22709
rect 75152 22660 75194 22700
rect 75234 22660 75276 22700
rect 75316 22660 75358 22700
rect 75398 22660 75440 22700
rect 75112 22651 75480 22660
rect 79112 22700 79480 22709
rect 79152 22660 79194 22700
rect 79234 22660 79276 22700
rect 79316 22660 79358 22700
rect 79398 22660 79440 22700
rect 79112 22651 79480 22660
rect 83112 22700 83480 22709
rect 83152 22660 83194 22700
rect 83234 22660 83276 22700
rect 83316 22660 83358 22700
rect 83398 22660 83440 22700
rect 83112 22651 83480 22660
rect 83596 22364 83636 23248
rect 83596 22315 83636 22324
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 8352 21944 8720 21953
rect 8392 21904 8434 21944
rect 8474 21904 8516 21944
rect 8556 21904 8598 21944
rect 8638 21904 8680 21944
rect 8352 21895 8720 21904
rect 12352 21944 12720 21953
rect 12392 21904 12434 21944
rect 12474 21904 12516 21944
rect 12556 21904 12598 21944
rect 12638 21904 12680 21944
rect 12352 21895 12720 21904
rect 16352 21944 16720 21953
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16352 21895 16720 21904
rect 20352 21944 20720 21953
rect 20392 21904 20434 21944
rect 20474 21904 20516 21944
rect 20556 21904 20598 21944
rect 20638 21904 20680 21944
rect 20352 21895 20720 21904
rect 24352 21944 24720 21953
rect 24392 21904 24434 21944
rect 24474 21904 24516 21944
rect 24556 21904 24598 21944
rect 24638 21904 24680 21944
rect 24352 21895 24720 21904
rect 28352 21944 28720 21953
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28352 21895 28720 21904
rect 32352 21944 32720 21953
rect 32392 21904 32434 21944
rect 32474 21904 32516 21944
rect 32556 21904 32598 21944
rect 32638 21904 32680 21944
rect 32352 21895 32720 21904
rect 36352 21944 36720 21953
rect 36392 21904 36434 21944
rect 36474 21904 36516 21944
rect 36556 21904 36598 21944
rect 36638 21904 36680 21944
rect 36352 21895 36720 21904
rect 40352 21944 40720 21953
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40352 21895 40720 21904
rect 44352 21944 44720 21953
rect 44392 21904 44434 21944
rect 44474 21904 44516 21944
rect 44556 21904 44598 21944
rect 44638 21904 44680 21944
rect 44352 21895 44720 21904
rect 48352 21944 48720 21953
rect 48392 21904 48434 21944
rect 48474 21904 48516 21944
rect 48556 21904 48598 21944
rect 48638 21904 48680 21944
rect 48352 21895 48720 21904
rect 52352 21944 52720 21953
rect 52392 21904 52434 21944
rect 52474 21904 52516 21944
rect 52556 21904 52598 21944
rect 52638 21904 52680 21944
rect 52352 21895 52720 21904
rect 56352 21944 56720 21953
rect 56392 21904 56434 21944
rect 56474 21904 56516 21944
rect 56556 21904 56598 21944
rect 56638 21904 56680 21944
rect 56352 21895 56720 21904
rect 60352 21944 60720 21953
rect 60392 21904 60434 21944
rect 60474 21904 60516 21944
rect 60556 21904 60598 21944
rect 60638 21904 60680 21944
rect 60352 21895 60720 21904
rect 64352 21944 64720 21953
rect 64392 21904 64434 21944
rect 64474 21904 64516 21944
rect 64556 21904 64598 21944
rect 64638 21904 64680 21944
rect 64352 21895 64720 21904
rect 68352 21944 68720 21953
rect 68392 21904 68434 21944
rect 68474 21904 68516 21944
rect 68556 21904 68598 21944
rect 68638 21904 68680 21944
rect 68352 21895 68720 21904
rect 72352 21944 72720 21953
rect 72392 21904 72434 21944
rect 72474 21904 72516 21944
rect 72556 21904 72598 21944
rect 72638 21904 72680 21944
rect 72352 21895 72720 21904
rect 76352 21944 76720 21953
rect 76392 21904 76434 21944
rect 76474 21904 76516 21944
rect 76556 21904 76598 21944
rect 76638 21904 76680 21944
rect 76352 21895 76720 21904
rect 80352 21944 80720 21953
rect 80392 21904 80434 21944
rect 80474 21904 80516 21944
rect 80556 21904 80598 21944
rect 80638 21904 80680 21944
rect 80352 21895 80720 21904
rect 84268 21776 84308 23752
rect 84352 23456 84720 23465
rect 84392 23416 84434 23456
rect 84474 23416 84516 23456
rect 84556 23416 84598 23456
rect 84638 23416 84680 23456
rect 84352 23407 84720 23416
rect 85420 22532 85460 23920
rect 88352 23456 88720 23465
rect 88392 23416 88434 23456
rect 88474 23416 88516 23456
rect 88556 23416 88598 23456
rect 88638 23416 88680 23456
rect 88352 23407 88720 23416
rect 92352 23456 92720 23465
rect 92392 23416 92434 23456
rect 92474 23416 92516 23456
rect 92556 23416 92598 23456
rect 92638 23416 92680 23456
rect 92352 23407 92720 23416
rect 86667 23120 86709 23129
rect 86667 23080 86668 23120
rect 86708 23080 86709 23120
rect 86667 23071 86709 23080
rect 86668 22986 86708 23071
rect 87532 22868 87572 22877
rect 87112 22700 87480 22709
rect 87152 22660 87194 22700
rect 87234 22660 87276 22700
rect 87316 22660 87358 22700
rect 87398 22660 87440 22700
rect 87112 22651 87480 22660
rect 85420 22483 85460 22492
rect 87532 22196 87572 22828
rect 91112 22700 91480 22709
rect 91152 22660 91194 22700
rect 91234 22660 91276 22700
rect 91316 22660 91358 22700
rect 91398 22660 91440 22700
rect 91112 22651 91480 22660
rect 94924 22448 94964 25768
rect 94924 22399 94964 22408
rect 95020 25724 95060 25733
rect 87532 22147 87572 22156
rect 84352 21944 84720 21953
rect 84392 21904 84434 21944
rect 84474 21904 84516 21944
rect 84556 21904 84598 21944
rect 84638 21904 84680 21944
rect 84352 21895 84720 21904
rect 88352 21944 88720 21953
rect 88392 21904 88434 21944
rect 88474 21904 88516 21944
rect 88556 21904 88598 21944
rect 88638 21904 88680 21944
rect 88352 21895 88720 21904
rect 92352 21944 92720 21953
rect 92392 21904 92434 21944
rect 92474 21904 92516 21944
rect 92556 21904 92598 21944
rect 92638 21904 92680 21944
rect 92352 21895 92720 21904
rect 84268 21727 84308 21736
rect 95020 21776 95060 25684
rect 96352 23456 96720 23465
rect 96392 23416 96434 23456
rect 96474 23416 96516 23456
rect 96556 23416 96598 23456
rect 96638 23416 96680 23456
rect 96352 23407 96720 23416
rect 95112 22700 95480 22709
rect 95152 22660 95194 22700
rect 95234 22660 95276 22700
rect 95316 22660 95358 22700
rect 95398 22660 95440 22700
rect 95112 22651 95480 22660
rect 99112 22700 99480 22709
rect 99152 22660 99194 22700
rect 99234 22660 99276 22700
rect 99316 22660 99358 22700
rect 99398 22660 99440 22700
rect 99112 22651 99480 22660
rect 96352 21944 96720 21953
rect 96392 21904 96434 21944
rect 96474 21904 96516 21944
rect 96556 21904 96598 21944
rect 96638 21904 96680 21944
rect 96352 21895 96720 21904
rect 95020 21727 95060 21736
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 7112 21188 7480 21197
rect 7152 21148 7194 21188
rect 7234 21148 7276 21188
rect 7316 21148 7358 21188
rect 7398 21148 7440 21188
rect 7112 21139 7480 21148
rect 11112 21188 11480 21197
rect 11152 21148 11194 21188
rect 11234 21148 11276 21188
rect 11316 21148 11358 21188
rect 11398 21148 11440 21188
rect 11112 21139 11480 21148
rect 15112 21188 15480 21197
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15112 21139 15480 21148
rect 19112 21188 19480 21197
rect 19152 21148 19194 21188
rect 19234 21148 19276 21188
rect 19316 21148 19358 21188
rect 19398 21148 19440 21188
rect 19112 21139 19480 21148
rect 23112 21188 23480 21197
rect 23152 21148 23194 21188
rect 23234 21148 23276 21188
rect 23316 21148 23358 21188
rect 23398 21148 23440 21188
rect 23112 21139 23480 21148
rect 27112 21188 27480 21197
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27112 21139 27480 21148
rect 31112 21188 31480 21197
rect 31152 21148 31194 21188
rect 31234 21148 31276 21188
rect 31316 21148 31358 21188
rect 31398 21148 31440 21188
rect 31112 21139 31480 21148
rect 35112 21188 35480 21197
rect 35152 21148 35194 21188
rect 35234 21148 35276 21188
rect 35316 21148 35358 21188
rect 35398 21148 35440 21188
rect 35112 21139 35480 21148
rect 39112 21188 39480 21197
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39112 21139 39480 21148
rect 43112 21188 43480 21197
rect 43152 21148 43194 21188
rect 43234 21148 43276 21188
rect 43316 21148 43358 21188
rect 43398 21148 43440 21188
rect 43112 21139 43480 21148
rect 47112 21188 47480 21197
rect 47152 21148 47194 21188
rect 47234 21148 47276 21188
rect 47316 21148 47358 21188
rect 47398 21148 47440 21188
rect 47112 21139 47480 21148
rect 51112 21188 51480 21197
rect 51152 21148 51194 21188
rect 51234 21148 51276 21188
rect 51316 21148 51358 21188
rect 51398 21148 51440 21188
rect 51112 21139 51480 21148
rect 55112 21188 55480 21197
rect 55152 21148 55194 21188
rect 55234 21148 55276 21188
rect 55316 21148 55358 21188
rect 55398 21148 55440 21188
rect 55112 21139 55480 21148
rect 59112 21188 59480 21197
rect 59152 21148 59194 21188
rect 59234 21148 59276 21188
rect 59316 21148 59358 21188
rect 59398 21148 59440 21188
rect 59112 21139 59480 21148
rect 63112 21188 63480 21197
rect 63152 21148 63194 21188
rect 63234 21148 63276 21188
rect 63316 21148 63358 21188
rect 63398 21148 63440 21188
rect 63112 21139 63480 21148
rect 67112 21188 67480 21197
rect 67152 21148 67194 21188
rect 67234 21148 67276 21188
rect 67316 21148 67358 21188
rect 67398 21148 67440 21188
rect 67112 21139 67480 21148
rect 71112 21188 71480 21197
rect 71152 21148 71194 21188
rect 71234 21148 71276 21188
rect 71316 21148 71358 21188
rect 71398 21148 71440 21188
rect 71112 21139 71480 21148
rect 75112 21188 75480 21197
rect 75152 21148 75194 21188
rect 75234 21148 75276 21188
rect 75316 21148 75358 21188
rect 75398 21148 75440 21188
rect 75112 21139 75480 21148
rect 79112 21188 79480 21197
rect 79152 21148 79194 21188
rect 79234 21148 79276 21188
rect 79316 21148 79358 21188
rect 79398 21148 79440 21188
rect 79112 21139 79480 21148
rect 83112 21188 83480 21197
rect 83152 21148 83194 21188
rect 83234 21148 83276 21188
rect 83316 21148 83358 21188
rect 83398 21148 83440 21188
rect 83112 21139 83480 21148
rect 87112 21188 87480 21197
rect 87152 21148 87194 21188
rect 87234 21148 87276 21188
rect 87316 21148 87358 21188
rect 87398 21148 87440 21188
rect 87112 21139 87480 21148
rect 91112 21188 91480 21197
rect 91152 21148 91194 21188
rect 91234 21148 91276 21188
rect 91316 21148 91358 21188
rect 91398 21148 91440 21188
rect 91112 21139 91480 21148
rect 95112 21188 95480 21197
rect 95152 21148 95194 21188
rect 95234 21148 95276 21188
rect 95316 21148 95358 21188
rect 95398 21148 95440 21188
rect 95112 21139 95480 21148
rect 99112 21188 99480 21197
rect 99152 21148 99194 21188
rect 99234 21148 99276 21188
rect 99316 21148 99358 21188
rect 99398 21148 99440 21188
rect 99112 21139 99480 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 8352 20432 8720 20441
rect 8392 20392 8434 20432
rect 8474 20392 8516 20432
rect 8556 20392 8598 20432
rect 8638 20392 8680 20432
rect 8352 20383 8720 20392
rect 12352 20432 12720 20441
rect 12392 20392 12434 20432
rect 12474 20392 12516 20432
rect 12556 20392 12598 20432
rect 12638 20392 12680 20432
rect 12352 20383 12720 20392
rect 16352 20432 16720 20441
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16352 20383 16720 20392
rect 20352 20432 20720 20441
rect 20392 20392 20434 20432
rect 20474 20392 20516 20432
rect 20556 20392 20598 20432
rect 20638 20392 20680 20432
rect 20352 20383 20720 20392
rect 24352 20432 24720 20441
rect 24392 20392 24434 20432
rect 24474 20392 24516 20432
rect 24556 20392 24598 20432
rect 24638 20392 24680 20432
rect 24352 20383 24720 20392
rect 28352 20432 28720 20441
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28352 20383 28720 20392
rect 32352 20432 32720 20441
rect 32392 20392 32434 20432
rect 32474 20392 32516 20432
rect 32556 20392 32598 20432
rect 32638 20392 32680 20432
rect 32352 20383 32720 20392
rect 36352 20432 36720 20441
rect 36392 20392 36434 20432
rect 36474 20392 36516 20432
rect 36556 20392 36598 20432
rect 36638 20392 36680 20432
rect 36352 20383 36720 20392
rect 40352 20432 40720 20441
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40352 20383 40720 20392
rect 44352 20432 44720 20441
rect 44392 20392 44434 20432
rect 44474 20392 44516 20432
rect 44556 20392 44598 20432
rect 44638 20392 44680 20432
rect 44352 20383 44720 20392
rect 48352 20432 48720 20441
rect 48392 20392 48434 20432
rect 48474 20392 48516 20432
rect 48556 20392 48598 20432
rect 48638 20392 48680 20432
rect 48352 20383 48720 20392
rect 52352 20432 52720 20441
rect 52392 20392 52434 20432
rect 52474 20392 52516 20432
rect 52556 20392 52598 20432
rect 52638 20392 52680 20432
rect 52352 20383 52720 20392
rect 56352 20432 56720 20441
rect 56392 20392 56434 20432
rect 56474 20392 56516 20432
rect 56556 20392 56598 20432
rect 56638 20392 56680 20432
rect 56352 20383 56720 20392
rect 60352 20432 60720 20441
rect 60392 20392 60434 20432
rect 60474 20392 60516 20432
rect 60556 20392 60598 20432
rect 60638 20392 60680 20432
rect 60352 20383 60720 20392
rect 64352 20432 64720 20441
rect 64392 20392 64434 20432
rect 64474 20392 64516 20432
rect 64556 20392 64598 20432
rect 64638 20392 64680 20432
rect 64352 20383 64720 20392
rect 68352 20432 68720 20441
rect 68392 20392 68434 20432
rect 68474 20392 68516 20432
rect 68556 20392 68598 20432
rect 68638 20392 68680 20432
rect 68352 20383 68720 20392
rect 72352 20432 72720 20441
rect 72392 20392 72434 20432
rect 72474 20392 72516 20432
rect 72556 20392 72598 20432
rect 72638 20392 72680 20432
rect 72352 20383 72720 20392
rect 76352 20432 76720 20441
rect 76392 20392 76434 20432
rect 76474 20392 76516 20432
rect 76556 20392 76598 20432
rect 76638 20392 76680 20432
rect 76352 20383 76720 20392
rect 80352 20432 80720 20441
rect 80392 20392 80434 20432
rect 80474 20392 80516 20432
rect 80556 20392 80598 20432
rect 80638 20392 80680 20432
rect 80352 20383 80720 20392
rect 84352 20432 84720 20441
rect 84392 20392 84434 20432
rect 84474 20392 84516 20432
rect 84556 20392 84598 20432
rect 84638 20392 84680 20432
rect 84352 20383 84720 20392
rect 88352 20432 88720 20441
rect 88392 20392 88434 20432
rect 88474 20392 88516 20432
rect 88556 20392 88598 20432
rect 88638 20392 88680 20432
rect 88352 20383 88720 20392
rect 92352 20432 92720 20441
rect 92392 20392 92434 20432
rect 92474 20392 92516 20432
rect 92556 20392 92598 20432
rect 92638 20392 92680 20432
rect 92352 20383 92720 20392
rect 96352 20432 96720 20441
rect 96392 20392 96434 20432
rect 96474 20392 96516 20432
rect 96556 20392 96598 20432
rect 96638 20392 96680 20432
rect 96352 20383 96720 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 7112 19676 7480 19685
rect 7152 19636 7194 19676
rect 7234 19636 7276 19676
rect 7316 19636 7358 19676
rect 7398 19636 7440 19676
rect 7112 19627 7480 19636
rect 11112 19676 11480 19685
rect 11152 19636 11194 19676
rect 11234 19636 11276 19676
rect 11316 19636 11358 19676
rect 11398 19636 11440 19676
rect 11112 19627 11480 19636
rect 15112 19676 15480 19685
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15112 19627 15480 19636
rect 19112 19676 19480 19685
rect 19152 19636 19194 19676
rect 19234 19636 19276 19676
rect 19316 19636 19358 19676
rect 19398 19636 19440 19676
rect 19112 19627 19480 19636
rect 23112 19676 23480 19685
rect 23152 19636 23194 19676
rect 23234 19636 23276 19676
rect 23316 19636 23358 19676
rect 23398 19636 23440 19676
rect 23112 19627 23480 19636
rect 27112 19676 27480 19685
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27112 19627 27480 19636
rect 31112 19676 31480 19685
rect 31152 19636 31194 19676
rect 31234 19636 31276 19676
rect 31316 19636 31358 19676
rect 31398 19636 31440 19676
rect 31112 19627 31480 19636
rect 35112 19676 35480 19685
rect 35152 19636 35194 19676
rect 35234 19636 35276 19676
rect 35316 19636 35358 19676
rect 35398 19636 35440 19676
rect 35112 19627 35480 19636
rect 39112 19676 39480 19685
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39112 19627 39480 19636
rect 43112 19676 43480 19685
rect 43152 19636 43194 19676
rect 43234 19636 43276 19676
rect 43316 19636 43358 19676
rect 43398 19636 43440 19676
rect 43112 19627 43480 19636
rect 47112 19676 47480 19685
rect 47152 19636 47194 19676
rect 47234 19636 47276 19676
rect 47316 19636 47358 19676
rect 47398 19636 47440 19676
rect 47112 19627 47480 19636
rect 51112 19676 51480 19685
rect 51152 19636 51194 19676
rect 51234 19636 51276 19676
rect 51316 19636 51358 19676
rect 51398 19636 51440 19676
rect 51112 19627 51480 19636
rect 55112 19676 55480 19685
rect 55152 19636 55194 19676
rect 55234 19636 55276 19676
rect 55316 19636 55358 19676
rect 55398 19636 55440 19676
rect 55112 19627 55480 19636
rect 59112 19676 59480 19685
rect 59152 19636 59194 19676
rect 59234 19636 59276 19676
rect 59316 19636 59358 19676
rect 59398 19636 59440 19676
rect 59112 19627 59480 19636
rect 63112 19676 63480 19685
rect 63152 19636 63194 19676
rect 63234 19636 63276 19676
rect 63316 19636 63358 19676
rect 63398 19636 63440 19676
rect 63112 19627 63480 19636
rect 67112 19676 67480 19685
rect 67152 19636 67194 19676
rect 67234 19636 67276 19676
rect 67316 19636 67358 19676
rect 67398 19636 67440 19676
rect 67112 19627 67480 19636
rect 71112 19676 71480 19685
rect 71152 19636 71194 19676
rect 71234 19636 71276 19676
rect 71316 19636 71358 19676
rect 71398 19636 71440 19676
rect 71112 19627 71480 19636
rect 75112 19676 75480 19685
rect 75152 19636 75194 19676
rect 75234 19636 75276 19676
rect 75316 19636 75358 19676
rect 75398 19636 75440 19676
rect 75112 19627 75480 19636
rect 79112 19676 79480 19685
rect 79152 19636 79194 19676
rect 79234 19636 79276 19676
rect 79316 19636 79358 19676
rect 79398 19636 79440 19676
rect 79112 19627 79480 19636
rect 83112 19676 83480 19685
rect 83152 19636 83194 19676
rect 83234 19636 83276 19676
rect 83316 19636 83358 19676
rect 83398 19636 83440 19676
rect 83112 19627 83480 19636
rect 87112 19676 87480 19685
rect 87152 19636 87194 19676
rect 87234 19636 87276 19676
rect 87316 19636 87358 19676
rect 87398 19636 87440 19676
rect 87112 19627 87480 19636
rect 91112 19676 91480 19685
rect 91152 19636 91194 19676
rect 91234 19636 91276 19676
rect 91316 19636 91358 19676
rect 91398 19636 91440 19676
rect 91112 19627 91480 19636
rect 95112 19676 95480 19685
rect 95152 19636 95194 19676
rect 95234 19636 95276 19676
rect 95316 19636 95358 19676
rect 95398 19636 95440 19676
rect 95112 19627 95480 19636
rect 99112 19676 99480 19685
rect 99152 19636 99194 19676
rect 99234 19636 99276 19676
rect 99316 19636 99358 19676
rect 99398 19636 99440 19676
rect 99112 19627 99480 19636
rect 86763 19340 86805 19349
rect 86763 19300 86764 19340
rect 86804 19300 86805 19340
rect 86763 19291 86805 19300
rect 86764 19206 86804 19291
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 8352 18920 8720 18929
rect 8392 18880 8434 18920
rect 8474 18880 8516 18920
rect 8556 18880 8598 18920
rect 8638 18880 8680 18920
rect 8352 18871 8720 18880
rect 12352 18920 12720 18929
rect 12392 18880 12434 18920
rect 12474 18880 12516 18920
rect 12556 18880 12598 18920
rect 12638 18880 12680 18920
rect 12352 18871 12720 18880
rect 16352 18920 16720 18929
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16352 18871 16720 18880
rect 20352 18920 20720 18929
rect 20392 18880 20434 18920
rect 20474 18880 20516 18920
rect 20556 18880 20598 18920
rect 20638 18880 20680 18920
rect 20352 18871 20720 18880
rect 24352 18920 24720 18929
rect 24392 18880 24434 18920
rect 24474 18880 24516 18920
rect 24556 18880 24598 18920
rect 24638 18880 24680 18920
rect 24352 18871 24720 18880
rect 28352 18920 28720 18929
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28352 18871 28720 18880
rect 32352 18920 32720 18929
rect 32392 18880 32434 18920
rect 32474 18880 32516 18920
rect 32556 18880 32598 18920
rect 32638 18880 32680 18920
rect 32352 18871 32720 18880
rect 36352 18920 36720 18929
rect 36392 18880 36434 18920
rect 36474 18880 36516 18920
rect 36556 18880 36598 18920
rect 36638 18880 36680 18920
rect 36352 18871 36720 18880
rect 40352 18920 40720 18929
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40352 18871 40720 18880
rect 44352 18920 44720 18929
rect 44392 18880 44434 18920
rect 44474 18880 44516 18920
rect 44556 18880 44598 18920
rect 44638 18880 44680 18920
rect 44352 18871 44720 18880
rect 48352 18920 48720 18929
rect 48392 18880 48434 18920
rect 48474 18880 48516 18920
rect 48556 18880 48598 18920
rect 48638 18880 48680 18920
rect 48352 18871 48720 18880
rect 52352 18920 52720 18929
rect 52392 18880 52434 18920
rect 52474 18880 52516 18920
rect 52556 18880 52598 18920
rect 52638 18880 52680 18920
rect 52352 18871 52720 18880
rect 56352 18920 56720 18929
rect 56392 18880 56434 18920
rect 56474 18880 56516 18920
rect 56556 18880 56598 18920
rect 56638 18880 56680 18920
rect 56352 18871 56720 18880
rect 60352 18920 60720 18929
rect 60392 18880 60434 18920
rect 60474 18880 60516 18920
rect 60556 18880 60598 18920
rect 60638 18880 60680 18920
rect 60352 18871 60720 18880
rect 64352 18920 64720 18929
rect 64392 18880 64434 18920
rect 64474 18880 64516 18920
rect 64556 18880 64598 18920
rect 64638 18880 64680 18920
rect 64352 18871 64720 18880
rect 68352 18920 68720 18929
rect 68392 18880 68434 18920
rect 68474 18880 68516 18920
rect 68556 18880 68598 18920
rect 68638 18880 68680 18920
rect 68352 18871 68720 18880
rect 72352 18920 72720 18929
rect 72392 18880 72434 18920
rect 72474 18880 72516 18920
rect 72556 18880 72598 18920
rect 72638 18880 72680 18920
rect 72352 18871 72720 18880
rect 76352 18920 76720 18929
rect 76392 18880 76434 18920
rect 76474 18880 76516 18920
rect 76556 18880 76598 18920
rect 76638 18880 76680 18920
rect 76352 18871 76720 18880
rect 80352 18920 80720 18929
rect 80392 18880 80434 18920
rect 80474 18880 80516 18920
rect 80556 18880 80598 18920
rect 80638 18880 80680 18920
rect 80352 18871 80720 18880
rect 84352 18920 84720 18929
rect 84392 18880 84434 18920
rect 84474 18880 84516 18920
rect 84556 18880 84598 18920
rect 84638 18880 84680 18920
rect 84352 18871 84720 18880
rect 88352 18920 88720 18929
rect 88392 18880 88434 18920
rect 88474 18880 88516 18920
rect 88556 18880 88598 18920
rect 88638 18880 88680 18920
rect 88352 18871 88720 18880
rect 92352 18920 92720 18929
rect 92392 18880 92434 18920
rect 92474 18880 92516 18920
rect 92556 18880 92598 18920
rect 92638 18880 92680 18920
rect 92352 18871 92720 18880
rect 96352 18920 96720 18929
rect 96392 18880 96434 18920
rect 96474 18880 96516 18920
rect 96556 18880 96598 18920
rect 96638 18880 96680 18920
rect 96352 18871 96720 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 7112 18164 7480 18173
rect 7152 18124 7194 18164
rect 7234 18124 7276 18164
rect 7316 18124 7358 18164
rect 7398 18124 7440 18164
rect 7112 18115 7480 18124
rect 11112 18164 11480 18173
rect 11152 18124 11194 18164
rect 11234 18124 11276 18164
rect 11316 18124 11358 18164
rect 11398 18124 11440 18164
rect 11112 18115 11480 18124
rect 15112 18164 15480 18173
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15112 18115 15480 18124
rect 19112 18164 19480 18173
rect 19152 18124 19194 18164
rect 19234 18124 19276 18164
rect 19316 18124 19358 18164
rect 19398 18124 19440 18164
rect 19112 18115 19480 18124
rect 23112 18164 23480 18173
rect 23152 18124 23194 18164
rect 23234 18124 23276 18164
rect 23316 18124 23358 18164
rect 23398 18124 23440 18164
rect 23112 18115 23480 18124
rect 27112 18164 27480 18173
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27112 18115 27480 18124
rect 31112 18164 31480 18173
rect 31152 18124 31194 18164
rect 31234 18124 31276 18164
rect 31316 18124 31358 18164
rect 31398 18124 31440 18164
rect 31112 18115 31480 18124
rect 35112 18164 35480 18173
rect 35152 18124 35194 18164
rect 35234 18124 35276 18164
rect 35316 18124 35358 18164
rect 35398 18124 35440 18164
rect 35112 18115 35480 18124
rect 39112 18164 39480 18173
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39112 18115 39480 18124
rect 43112 18164 43480 18173
rect 43152 18124 43194 18164
rect 43234 18124 43276 18164
rect 43316 18124 43358 18164
rect 43398 18124 43440 18164
rect 43112 18115 43480 18124
rect 47112 18164 47480 18173
rect 47152 18124 47194 18164
rect 47234 18124 47276 18164
rect 47316 18124 47358 18164
rect 47398 18124 47440 18164
rect 47112 18115 47480 18124
rect 51112 18164 51480 18173
rect 51152 18124 51194 18164
rect 51234 18124 51276 18164
rect 51316 18124 51358 18164
rect 51398 18124 51440 18164
rect 51112 18115 51480 18124
rect 55112 18164 55480 18173
rect 55152 18124 55194 18164
rect 55234 18124 55276 18164
rect 55316 18124 55358 18164
rect 55398 18124 55440 18164
rect 55112 18115 55480 18124
rect 59112 18164 59480 18173
rect 59152 18124 59194 18164
rect 59234 18124 59276 18164
rect 59316 18124 59358 18164
rect 59398 18124 59440 18164
rect 59112 18115 59480 18124
rect 63112 18164 63480 18173
rect 63152 18124 63194 18164
rect 63234 18124 63276 18164
rect 63316 18124 63358 18164
rect 63398 18124 63440 18164
rect 63112 18115 63480 18124
rect 67112 18164 67480 18173
rect 67152 18124 67194 18164
rect 67234 18124 67276 18164
rect 67316 18124 67358 18164
rect 67398 18124 67440 18164
rect 67112 18115 67480 18124
rect 71112 18164 71480 18173
rect 71152 18124 71194 18164
rect 71234 18124 71276 18164
rect 71316 18124 71358 18164
rect 71398 18124 71440 18164
rect 71112 18115 71480 18124
rect 75112 18164 75480 18173
rect 75152 18124 75194 18164
rect 75234 18124 75276 18164
rect 75316 18124 75358 18164
rect 75398 18124 75440 18164
rect 75112 18115 75480 18124
rect 79112 18164 79480 18173
rect 79152 18124 79194 18164
rect 79234 18124 79276 18164
rect 79316 18124 79358 18164
rect 79398 18124 79440 18164
rect 79112 18115 79480 18124
rect 83112 18164 83480 18173
rect 83152 18124 83194 18164
rect 83234 18124 83276 18164
rect 83316 18124 83358 18164
rect 83398 18124 83440 18164
rect 83112 18115 83480 18124
rect 87112 18164 87480 18173
rect 87152 18124 87194 18164
rect 87234 18124 87276 18164
rect 87316 18124 87358 18164
rect 87398 18124 87440 18164
rect 87112 18115 87480 18124
rect 91112 18164 91480 18173
rect 91152 18124 91194 18164
rect 91234 18124 91276 18164
rect 91316 18124 91358 18164
rect 91398 18124 91440 18164
rect 91112 18115 91480 18124
rect 95112 18164 95480 18173
rect 95152 18124 95194 18164
rect 95234 18124 95276 18164
rect 95316 18124 95358 18164
rect 95398 18124 95440 18164
rect 95112 18115 95480 18124
rect 99112 18164 99480 18173
rect 99152 18124 99194 18164
rect 99234 18124 99276 18164
rect 99316 18124 99358 18164
rect 99398 18124 99440 18164
rect 99112 18115 99480 18124
rect 84268 17576 84308 17585
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 8352 17408 8720 17417
rect 8392 17368 8434 17408
rect 8474 17368 8516 17408
rect 8556 17368 8598 17408
rect 8638 17368 8680 17408
rect 8352 17359 8720 17368
rect 12352 17408 12720 17417
rect 12392 17368 12434 17408
rect 12474 17368 12516 17408
rect 12556 17368 12598 17408
rect 12638 17368 12680 17408
rect 12352 17359 12720 17368
rect 16352 17408 16720 17417
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16352 17359 16720 17368
rect 20352 17408 20720 17417
rect 20392 17368 20434 17408
rect 20474 17368 20516 17408
rect 20556 17368 20598 17408
rect 20638 17368 20680 17408
rect 20352 17359 20720 17368
rect 24352 17408 24720 17417
rect 24392 17368 24434 17408
rect 24474 17368 24516 17408
rect 24556 17368 24598 17408
rect 24638 17368 24680 17408
rect 24352 17359 24720 17368
rect 28352 17408 28720 17417
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28352 17359 28720 17368
rect 32352 17408 32720 17417
rect 32392 17368 32434 17408
rect 32474 17368 32516 17408
rect 32556 17368 32598 17408
rect 32638 17368 32680 17408
rect 32352 17359 32720 17368
rect 36352 17408 36720 17417
rect 36392 17368 36434 17408
rect 36474 17368 36516 17408
rect 36556 17368 36598 17408
rect 36638 17368 36680 17408
rect 36352 17359 36720 17368
rect 40352 17408 40720 17417
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40352 17359 40720 17368
rect 44352 17408 44720 17417
rect 44392 17368 44434 17408
rect 44474 17368 44516 17408
rect 44556 17368 44598 17408
rect 44638 17368 44680 17408
rect 44352 17359 44720 17368
rect 48352 17408 48720 17417
rect 48392 17368 48434 17408
rect 48474 17368 48516 17408
rect 48556 17368 48598 17408
rect 48638 17368 48680 17408
rect 48352 17359 48720 17368
rect 52352 17408 52720 17417
rect 52392 17368 52434 17408
rect 52474 17368 52516 17408
rect 52556 17368 52598 17408
rect 52638 17368 52680 17408
rect 52352 17359 52720 17368
rect 56352 17408 56720 17417
rect 56392 17368 56434 17408
rect 56474 17368 56516 17408
rect 56556 17368 56598 17408
rect 56638 17368 56680 17408
rect 56352 17359 56720 17368
rect 60352 17408 60720 17417
rect 60392 17368 60434 17408
rect 60474 17368 60516 17408
rect 60556 17368 60598 17408
rect 60638 17368 60680 17408
rect 60352 17359 60720 17368
rect 64352 17408 64720 17417
rect 64392 17368 64434 17408
rect 64474 17368 64516 17408
rect 64556 17368 64598 17408
rect 64638 17368 64680 17408
rect 64352 17359 64720 17368
rect 68352 17408 68720 17417
rect 68392 17368 68434 17408
rect 68474 17368 68516 17408
rect 68556 17368 68598 17408
rect 68638 17368 68680 17408
rect 68352 17359 68720 17368
rect 72352 17408 72720 17417
rect 72392 17368 72434 17408
rect 72474 17368 72516 17408
rect 72556 17368 72598 17408
rect 72638 17368 72680 17408
rect 72352 17359 72720 17368
rect 76352 17408 76720 17417
rect 76392 17368 76434 17408
rect 76474 17368 76516 17408
rect 76556 17368 76598 17408
rect 76638 17368 76680 17408
rect 76352 17359 76720 17368
rect 80352 17408 80720 17417
rect 80392 17368 80434 17408
rect 80474 17368 80516 17408
rect 80556 17368 80598 17408
rect 80638 17368 80680 17408
rect 80352 17359 80720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 7112 16652 7480 16661
rect 7152 16612 7194 16652
rect 7234 16612 7276 16652
rect 7316 16612 7358 16652
rect 7398 16612 7440 16652
rect 7112 16603 7480 16612
rect 11112 16652 11480 16661
rect 11152 16612 11194 16652
rect 11234 16612 11276 16652
rect 11316 16612 11358 16652
rect 11398 16612 11440 16652
rect 11112 16603 11480 16612
rect 15112 16652 15480 16661
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15112 16603 15480 16612
rect 19112 16652 19480 16661
rect 19152 16612 19194 16652
rect 19234 16612 19276 16652
rect 19316 16612 19358 16652
rect 19398 16612 19440 16652
rect 19112 16603 19480 16612
rect 23112 16652 23480 16661
rect 23152 16612 23194 16652
rect 23234 16612 23276 16652
rect 23316 16612 23358 16652
rect 23398 16612 23440 16652
rect 23112 16603 23480 16612
rect 27112 16652 27480 16661
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27112 16603 27480 16612
rect 31112 16652 31480 16661
rect 31152 16612 31194 16652
rect 31234 16612 31276 16652
rect 31316 16612 31358 16652
rect 31398 16612 31440 16652
rect 31112 16603 31480 16612
rect 35112 16652 35480 16661
rect 35152 16612 35194 16652
rect 35234 16612 35276 16652
rect 35316 16612 35358 16652
rect 35398 16612 35440 16652
rect 35112 16603 35480 16612
rect 39112 16652 39480 16661
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39112 16603 39480 16612
rect 43112 16652 43480 16661
rect 43152 16612 43194 16652
rect 43234 16612 43276 16652
rect 43316 16612 43358 16652
rect 43398 16612 43440 16652
rect 43112 16603 43480 16612
rect 47112 16652 47480 16661
rect 47152 16612 47194 16652
rect 47234 16612 47276 16652
rect 47316 16612 47358 16652
rect 47398 16612 47440 16652
rect 47112 16603 47480 16612
rect 51112 16652 51480 16661
rect 51152 16612 51194 16652
rect 51234 16612 51276 16652
rect 51316 16612 51358 16652
rect 51398 16612 51440 16652
rect 51112 16603 51480 16612
rect 55112 16652 55480 16661
rect 55152 16612 55194 16652
rect 55234 16612 55276 16652
rect 55316 16612 55358 16652
rect 55398 16612 55440 16652
rect 55112 16603 55480 16612
rect 59112 16652 59480 16661
rect 59152 16612 59194 16652
rect 59234 16612 59276 16652
rect 59316 16612 59358 16652
rect 59398 16612 59440 16652
rect 59112 16603 59480 16612
rect 63112 16652 63480 16661
rect 63152 16612 63194 16652
rect 63234 16612 63276 16652
rect 63316 16612 63358 16652
rect 63398 16612 63440 16652
rect 63112 16603 63480 16612
rect 67112 16652 67480 16661
rect 67152 16612 67194 16652
rect 67234 16612 67276 16652
rect 67316 16612 67358 16652
rect 67398 16612 67440 16652
rect 67112 16603 67480 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 8352 15896 8720 15905
rect 8392 15856 8434 15896
rect 8474 15856 8516 15896
rect 8556 15856 8598 15896
rect 8638 15856 8680 15896
rect 8352 15847 8720 15856
rect 12352 15896 12720 15905
rect 12392 15856 12434 15896
rect 12474 15856 12516 15896
rect 12556 15856 12598 15896
rect 12638 15856 12680 15896
rect 12352 15847 12720 15856
rect 16352 15896 16720 15905
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16352 15847 16720 15856
rect 20352 15896 20720 15905
rect 20392 15856 20434 15896
rect 20474 15856 20516 15896
rect 20556 15856 20598 15896
rect 20638 15856 20680 15896
rect 20352 15847 20720 15856
rect 24352 15896 24720 15905
rect 24392 15856 24434 15896
rect 24474 15856 24516 15896
rect 24556 15856 24598 15896
rect 24638 15856 24680 15896
rect 24352 15847 24720 15856
rect 28352 15896 28720 15905
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28352 15847 28720 15856
rect 32352 15896 32720 15905
rect 32392 15856 32434 15896
rect 32474 15856 32516 15896
rect 32556 15856 32598 15896
rect 32638 15856 32680 15896
rect 32352 15847 32720 15856
rect 36352 15896 36720 15905
rect 36392 15856 36434 15896
rect 36474 15856 36516 15896
rect 36556 15856 36598 15896
rect 36638 15856 36680 15896
rect 36352 15847 36720 15856
rect 40352 15896 40720 15905
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40352 15847 40720 15856
rect 44352 15896 44720 15905
rect 44392 15856 44434 15896
rect 44474 15856 44516 15896
rect 44556 15856 44598 15896
rect 44638 15856 44680 15896
rect 44352 15847 44720 15856
rect 48352 15896 48720 15905
rect 48392 15856 48434 15896
rect 48474 15856 48516 15896
rect 48556 15856 48598 15896
rect 48638 15856 48680 15896
rect 48352 15847 48720 15856
rect 52352 15896 52720 15905
rect 52392 15856 52434 15896
rect 52474 15856 52516 15896
rect 52556 15856 52598 15896
rect 52638 15856 52680 15896
rect 52352 15847 52720 15856
rect 56352 15896 56720 15905
rect 56392 15856 56434 15896
rect 56474 15856 56516 15896
rect 56556 15856 56598 15896
rect 56638 15856 56680 15896
rect 56352 15847 56720 15856
rect 60352 15896 60720 15905
rect 60392 15856 60434 15896
rect 60474 15856 60516 15896
rect 60556 15856 60598 15896
rect 60638 15856 60680 15896
rect 60352 15847 60720 15856
rect 64352 15896 64720 15905
rect 64392 15856 64434 15896
rect 64474 15856 64516 15896
rect 64556 15856 64598 15896
rect 64638 15856 64680 15896
rect 64352 15847 64720 15856
rect 68352 15896 68720 15905
rect 68392 15856 68434 15896
rect 68474 15856 68516 15896
rect 68556 15856 68598 15896
rect 68638 15856 68680 15896
rect 68352 15847 68720 15856
rect 71788 15560 71828 15569
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 7112 15140 7480 15149
rect 7152 15100 7194 15140
rect 7234 15100 7276 15140
rect 7316 15100 7358 15140
rect 7398 15100 7440 15140
rect 7112 15091 7480 15100
rect 11112 15140 11480 15149
rect 11152 15100 11194 15140
rect 11234 15100 11276 15140
rect 11316 15100 11358 15140
rect 11398 15100 11440 15140
rect 11112 15091 11480 15100
rect 15112 15140 15480 15149
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15112 15091 15480 15100
rect 19112 15140 19480 15149
rect 19152 15100 19194 15140
rect 19234 15100 19276 15140
rect 19316 15100 19358 15140
rect 19398 15100 19440 15140
rect 19112 15091 19480 15100
rect 23112 15140 23480 15149
rect 23152 15100 23194 15140
rect 23234 15100 23276 15140
rect 23316 15100 23358 15140
rect 23398 15100 23440 15140
rect 23112 15091 23480 15100
rect 27112 15140 27480 15149
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27112 15091 27480 15100
rect 31112 15140 31480 15149
rect 31152 15100 31194 15140
rect 31234 15100 31276 15140
rect 31316 15100 31358 15140
rect 31398 15100 31440 15140
rect 31112 15091 31480 15100
rect 35112 15140 35480 15149
rect 35152 15100 35194 15140
rect 35234 15100 35276 15140
rect 35316 15100 35358 15140
rect 35398 15100 35440 15140
rect 35112 15091 35480 15100
rect 39112 15140 39480 15149
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39112 15091 39480 15100
rect 43112 15140 43480 15149
rect 43152 15100 43194 15140
rect 43234 15100 43276 15140
rect 43316 15100 43358 15140
rect 43398 15100 43440 15140
rect 43112 15091 43480 15100
rect 47112 15140 47480 15149
rect 47152 15100 47194 15140
rect 47234 15100 47276 15140
rect 47316 15100 47358 15140
rect 47398 15100 47440 15140
rect 47112 15091 47480 15100
rect 51112 15140 51480 15149
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51112 15091 51480 15100
rect 55112 15140 55480 15149
rect 55152 15100 55194 15140
rect 55234 15100 55276 15140
rect 55316 15100 55358 15140
rect 55398 15100 55440 15140
rect 55112 15091 55480 15100
rect 59112 15140 59480 15149
rect 59152 15100 59194 15140
rect 59234 15100 59276 15140
rect 59316 15100 59358 15140
rect 59398 15100 59440 15140
rect 59112 15091 59480 15100
rect 63112 15140 63480 15149
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63112 15091 63480 15100
rect 67112 15140 67480 15149
rect 67152 15100 67194 15140
rect 67234 15100 67276 15140
rect 67316 15100 67358 15140
rect 67398 15100 67440 15140
rect 67112 15091 67480 15100
rect 71788 15056 71828 15520
rect 84268 15560 84308 17536
rect 84352 17408 84720 17417
rect 84392 17368 84434 17408
rect 84474 17368 84516 17408
rect 84556 17368 84598 17408
rect 84638 17368 84680 17408
rect 84352 17359 84720 17368
rect 88352 17408 88720 17417
rect 88392 17368 88434 17408
rect 88474 17368 88516 17408
rect 88556 17368 88598 17408
rect 88638 17368 88680 17408
rect 88352 17359 88720 17368
rect 92352 17408 92720 17417
rect 92392 17368 92434 17408
rect 92474 17368 92516 17408
rect 92556 17368 92598 17408
rect 92638 17368 92680 17408
rect 92352 17359 92720 17368
rect 96352 17408 96720 17417
rect 96392 17368 96434 17408
rect 96474 17368 96516 17408
rect 96556 17368 96598 17408
rect 96638 17368 96680 17408
rect 96352 17359 96720 17368
rect 84268 15511 84308 15520
rect 98860 15476 98900 15485
rect 71788 15007 71828 15016
rect 71884 15392 71924 15401
rect 71884 14888 71924 15352
rect 71884 14839 71924 14848
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 8352 14384 8720 14393
rect 8392 14344 8434 14384
rect 8474 14344 8516 14384
rect 8556 14344 8598 14384
rect 8638 14344 8680 14384
rect 8352 14335 8720 14344
rect 12352 14384 12720 14393
rect 12392 14344 12434 14384
rect 12474 14344 12516 14384
rect 12556 14344 12598 14384
rect 12638 14344 12680 14384
rect 12352 14335 12720 14344
rect 16352 14384 16720 14393
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16352 14335 16720 14344
rect 20352 14384 20720 14393
rect 20392 14344 20434 14384
rect 20474 14344 20516 14384
rect 20556 14344 20598 14384
rect 20638 14344 20680 14384
rect 20352 14335 20720 14344
rect 24352 14384 24720 14393
rect 24392 14344 24434 14384
rect 24474 14344 24516 14384
rect 24556 14344 24598 14384
rect 24638 14344 24680 14384
rect 24352 14335 24720 14344
rect 28352 14384 28720 14393
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28352 14335 28720 14344
rect 32352 14384 32720 14393
rect 32392 14344 32434 14384
rect 32474 14344 32516 14384
rect 32556 14344 32598 14384
rect 32638 14344 32680 14384
rect 32352 14335 32720 14344
rect 36352 14384 36720 14393
rect 36392 14344 36434 14384
rect 36474 14344 36516 14384
rect 36556 14344 36598 14384
rect 36638 14344 36680 14384
rect 36352 14335 36720 14344
rect 40352 14384 40720 14393
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40352 14335 40720 14344
rect 44352 14384 44720 14393
rect 44392 14344 44434 14384
rect 44474 14344 44516 14384
rect 44556 14344 44598 14384
rect 44638 14344 44680 14384
rect 44352 14335 44720 14344
rect 48352 14384 48720 14393
rect 48392 14344 48434 14384
rect 48474 14344 48516 14384
rect 48556 14344 48598 14384
rect 48638 14344 48680 14384
rect 48352 14335 48720 14344
rect 52352 14384 52720 14393
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52352 14335 52720 14344
rect 56352 14384 56720 14393
rect 56392 14344 56434 14384
rect 56474 14344 56516 14384
rect 56556 14344 56598 14384
rect 56638 14344 56680 14384
rect 56352 14335 56720 14344
rect 60352 14384 60720 14393
rect 60392 14344 60434 14384
rect 60474 14344 60516 14384
rect 60556 14344 60598 14384
rect 60638 14344 60680 14384
rect 60352 14335 60720 14344
rect 64352 14384 64720 14393
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64352 14335 64720 14344
rect 68352 14384 68720 14393
rect 68392 14344 68434 14384
rect 68474 14344 68516 14384
rect 68556 14344 68598 14384
rect 68638 14344 68680 14384
rect 68352 14335 68720 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 7112 13628 7480 13637
rect 7152 13588 7194 13628
rect 7234 13588 7276 13628
rect 7316 13588 7358 13628
rect 7398 13588 7440 13628
rect 7112 13579 7480 13588
rect 11112 13628 11480 13637
rect 11152 13588 11194 13628
rect 11234 13588 11276 13628
rect 11316 13588 11358 13628
rect 11398 13588 11440 13628
rect 11112 13579 11480 13588
rect 15112 13628 15480 13637
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15112 13579 15480 13588
rect 19112 13628 19480 13637
rect 19152 13588 19194 13628
rect 19234 13588 19276 13628
rect 19316 13588 19358 13628
rect 19398 13588 19440 13628
rect 19112 13579 19480 13588
rect 23112 13628 23480 13637
rect 23152 13588 23194 13628
rect 23234 13588 23276 13628
rect 23316 13588 23358 13628
rect 23398 13588 23440 13628
rect 23112 13579 23480 13588
rect 27112 13628 27480 13637
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27112 13579 27480 13588
rect 31112 13628 31480 13637
rect 31152 13588 31194 13628
rect 31234 13588 31276 13628
rect 31316 13588 31358 13628
rect 31398 13588 31440 13628
rect 31112 13579 31480 13588
rect 35112 13628 35480 13637
rect 35152 13588 35194 13628
rect 35234 13588 35276 13628
rect 35316 13588 35358 13628
rect 35398 13588 35440 13628
rect 35112 13579 35480 13588
rect 39112 13628 39480 13637
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39112 13579 39480 13588
rect 43112 13628 43480 13637
rect 43152 13588 43194 13628
rect 43234 13588 43276 13628
rect 43316 13588 43358 13628
rect 43398 13588 43440 13628
rect 43112 13579 43480 13588
rect 47112 13628 47480 13637
rect 47152 13588 47194 13628
rect 47234 13588 47276 13628
rect 47316 13588 47358 13628
rect 47398 13588 47440 13628
rect 47112 13579 47480 13588
rect 51112 13628 51480 13637
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51112 13579 51480 13588
rect 55112 13628 55480 13637
rect 55152 13588 55194 13628
rect 55234 13588 55276 13628
rect 55316 13588 55358 13628
rect 55398 13588 55440 13628
rect 55112 13579 55480 13588
rect 59112 13628 59480 13637
rect 59152 13588 59194 13628
rect 59234 13588 59276 13628
rect 59316 13588 59358 13628
rect 59398 13588 59440 13628
rect 59112 13579 59480 13588
rect 63112 13628 63480 13637
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63112 13579 63480 13588
rect 67112 13628 67480 13637
rect 67152 13588 67194 13628
rect 67234 13588 67276 13628
rect 67316 13588 67358 13628
rect 67398 13588 67440 13628
rect 67112 13579 67480 13588
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 8352 12872 8720 12881
rect 8392 12832 8434 12872
rect 8474 12832 8516 12872
rect 8556 12832 8598 12872
rect 8638 12832 8680 12872
rect 8352 12823 8720 12832
rect 12352 12872 12720 12881
rect 12392 12832 12434 12872
rect 12474 12832 12516 12872
rect 12556 12832 12598 12872
rect 12638 12832 12680 12872
rect 12352 12823 12720 12832
rect 16352 12872 16720 12881
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16352 12823 16720 12832
rect 20352 12872 20720 12881
rect 20392 12832 20434 12872
rect 20474 12832 20516 12872
rect 20556 12832 20598 12872
rect 20638 12832 20680 12872
rect 20352 12823 20720 12832
rect 24352 12872 24720 12881
rect 24392 12832 24434 12872
rect 24474 12832 24516 12872
rect 24556 12832 24598 12872
rect 24638 12832 24680 12872
rect 24352 12823 24720 12832
rect 28352 12872 28720 12881
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28352 12823 28720 12832
rect 32352 12872 32720 12881
rect 32392 12832 32434 12872
rect 32474 12832 32516 12872
rect 32556 12832 32598 12872
rect 32638 12832 32680 12872
rect 32352 12823 32720 12832
rect 36352 12872 36720 12881
rect 36392 12832 36434 12872
rect 36474 12832 36516 12872
rect 36556 12832 36598 12872
rect 36638 12832 36680 12872
rect 36352 12823 36720 12832
rect 40352 12872 40720 12881
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40352 12823 40720 12832
rect 44352 12872 44720 12881
rect 44392 12832 44434 12872
rect 44474 12832 44516 12872
rect 44556 12832 44598 12872
rect 44638 12832 44680 12872
rect 44352 12823 44720 12832
rect 48352 12872 48720 12881
rect 48392 12832 48434 12872
rect 48474 12832 48516 12872
rect 48556 12832 48598 12872
rect 48638 12832 48680 12872
rect 48352 12823 48720 12832
rect 52352 12872 52720 12881
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52352 12823 52720 12832
rect 56352 12872 56720 12881
rect 56392 12832 56434 12872
rect 56474 12832 56516 12872
rect 56556 12832 56598 12872
rect 56638 12832 56680 12872
rect 56352 12823 56720 12832
rect 60352 12872 60720 12881
rect 60392 12832 60434 12872
rect 60474 12832 60516 12872
rect 60556 12832 60598 12872
rect 60638 12832 60680 12872
rect 60352 12823 60720 12832
rect 64352 12872 64720 12881
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64352 12823 64720 12832
rect 68352 12872 68720 12881
rect 68392 12832 68434 12872
rect 68474 12832 68516 12872
rect 68556 12832 68598 12872
rect 68638 12832 68680 12872
rect 68352 12823 68720 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 7112 12116 7480 12125
rect 7152 12076 7194 12116
rect 7234 12076 7276 12116
rect 7316 12076 7358 12116
rect 7398 12076 7440 12116
rect 7112 12067 7480 12076
rect 11112 12116 11480 12125
rect 11152 12076 11194 12116
rect 11234 12076 11276 12116
rect 11316 12076 11358 12116
rect 11398 12076 11440 12116
rect 11112 12067 11480 12076
rect 15112 12116 15480 12125
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15112 12067 15480 12076
rect 19112 12116 19480 12125
rect 19152 12076 19194 12116
rect 19234 12076 19276 12116
rect 19316 12076 19358 12116
rect 19398 12076 19440 12116
rect 19112 12067 19480 12076
rect 23112 12116 23480 12125
rect 23152 12076 23194 12116
rect 23234 12076 23276 12116
rect 23316 12076 23358 12116
rect 23398 12076 23440 12116
rect 23112 12067 23480 12076
rect 27112 12116 27480 12125
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27112 12067 27480 12076
rect 31112 12116 31480 12125
rect 31152 12076 31194 12116
rect 31234 12076 31276 12116
rect 31316 12076 31358 12116
rect 31398 12076 31440 12116
rect 31112 12067 31480 12076
rect 35112 12116 35480 12125
rect 35152 12076 35194 12116
rect 35234 12076 35276 12116
rect 35316 12076 35358 12116
rect 35398 12076 35440 12116
rect 35112 12067 35480 12076
rect 39112 12116 39480 12125
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39112 12067 39480 12076
rect 43112 12116 43480 12125
rect 43152 12076 43194 12116
rect 43234 12076 43276 12116
rect 43316 12076 43358 12116
rect 43398 12076 43440 12116
rect 43112 12067 43480 12076
rect 47112 12116 47480 12125
rect 47152 12076 47194 12116
rect 47234 12076 47276 12116
rect 47316 12076 47358 12116
rect 47398 12076 47440 12116
rect 47112 12067 47480 12076
rect 51112 12116 51480 12125
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51112 12067 51480 12076
rect 55112 12116 55480 12125
rect 55152 12076 55194 12116
rect 55234 12076 55276 12116
rect 55316 12076 55358 12116
rect 55398 12076 55440 12116
rect 55112 12067 55480 12076
rect 59112 12116 59480 12125
rect 59152 12076 59194 12116
rect 59234 12076 59276 12116
rect 59316 12076 59358 12116
rect 59398 12076 59440 12116
rect 59112 12067 59480 12076
rect 63112 12116 63480 12125
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63112 12067 63480 12076
rect 67112 12116 67480 12125
rect 67152 12076 67194 12116
rect 67234 12076 67276 12116
rect 67316 12076 67358 12116
rect 67398 12076 67440 12116
rect 67112 12067 67480 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 8352 11360 8720 11369
rect 8392 11320 8434 11360
rect 8474 11320 8516 11360
rect 8556 11320 8598 11360
rect 8638 11320 8680 11360
rect 8352 11311 8720 11320
rect 12352 11360 12720 11369
rect 12392 11320 12434 11360
rect 12474 11320 12516 11360
rect 12556 11320 12598 11360
rect 12638 11320 12680 11360
rect 12352 11311 12720 11320
rect 16352 11360 16720 11369
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16352 11311 16720 11320
rect 20352 11360 20720 11369
rect 20392 11320 20434 11360
rect 20474 11320 20516 11360
rect 20556 11320 20598 11360
rect 20638 11320 20680 11360
rect 20352 11311 20720 11320
rect 24352 11360 24720 11369
rect 24392 11320 24434 11360
rect 24474 11320 24516 11360
rect 24556 11320 24598 11360
rect 24638 11320 24680 11360
rect 24352 11311 24720 11320
rect 28352 11360 28720 11369
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28352 11311 28720 11320
rect 32352 11360 32720 11369
rect 32392 11320 32434 11360
rect 32474 11320 32516 11360
rect 32556 11320 32598 11360
rect 32638 11320 32680 11360
rect 32352 11311 32720 11320
rect 36352 11360 36720 11369
rect 36392 11320 36434 11360
rect 36474 11320 36516 11360
rect 36556 11320 36598 11360
rect 36638 11320 36680 11360
rect 36352 11311 36720 11320
rect 40352 11360 40720 11369
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40352 11311 40720 11320
rect 44352 11360 44720 11369
rect 44392 11320 44434 11360
rect 44474 11320 44516 11360
rect 44556 11320 44598 11360
rect 44638 11320 44680 11360
rect 44352 11311 44720 11320
rect 48352 11360 48720 11369
rect 48392 11320 48434 11360
rect 48474 11320 48516 11360
rect 48556 11320 48598 11360
rect 48638 11320 48680 11360
rect 48352 11311 48720 11320
rect 52352 11360 52720 11369
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52352 11311 52720 11320
rect 56352 11360 56720 11369
rect 56392 11320 56434 11360
rect 56474 11320 56516 11360
rect 56556 11320 56598 11360
rect 56638 11320 56680 11360
rect 56352 11311 56720 11320
rect 60352 11360 60720 11369
rect 60392 11320 60434 11360
rect 60474 11320 60516 11360
rect 60556 11320 60598 11360
rect 60638 11320 60680 11360
rect 60352 11311 60720 11320
rect 64352 11360 64720 11369
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64352 11311 64720 11320
rect 68352 11360 68720 11369
rect 68392 11320 68434 11360
rect 68474 11320 68516 11360
rect 68556 11320 68598 11360
rect 68638 11320 68680 11360
rect 68352 11311 68720 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 7112 10604 7480 10613
rect 7152 10564 7194 10604
rect 7234 10564 7276 10604
rect 7316 10564 7358 10604
rect 7398 10564 7440 10604
rect 7112 10555 7480 10564
rect 11112 10604 11480 10613
rect 11152 10564 11194 10604
rect 11234 10564 11276 10604
rect 11316 10564 11358 10604
rect 11398 10564 11440 10604
rect 11112 10555 11480 10564
rect 15112 10604 15480 10613
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15112 10555 15480 10564
rect 19112 10604 19480 10613
rect 19152 10564 19194 10604
rect 19234 10564 19276 10604
rect 19316 10564 19358 10604
rect 19398 10564 19440 10604
rect 19112 10555 19480 10564
rect 23112 10604 23480 10613
rect 23152 10564 23194 10604
rect 23234 10564 23276 10604
rect 23316 10564 23358 10604
rect 23398 10564 23440 10604
rect 23112 10555 23480 10564
rect 27112 10604 27480 10613
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27112 10555 27480 10564
rect 31112 10604 31480 10613
rect 31152 10564 31194 10604
rect 31234 10564 31276 10604
rect 31316 10564 31358 10604
rect 31398 10564 31440 10604
rect 31112 10555 31480 10564
rect 35112 10604 35480 10613
rect 35152 10564 35194 10604
rect 35234 10564 35276 10604
rect 35316 10564 35358 10604
rect 35398 10564 35440 10604
rect 35112 10555 35480 10564
rect 39112 10604 39480 10613
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39112 10555 39480 10564
rect 43112 10604 43480 10613
rect 43152 10564 43194 10604
rect 43234 10564 43276 10604
rect 43316 10564 43358 10604
rect 43398 10564 43440 10604
rect 43112 10555 43480 10564
rect 47112 10604 47480 10613
rect 47152 10564 47194 10604
rect 47234 10564 47276 10604
rect 47316 10564 47358 10604
rect 47398 10564 47440 10604
rect 47112 10555 47480 10564
rect 51112 10604 51480 10613
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51112 10555 51480 10564
rect 55112 10604 55480 10613
rect 55152 10564 55194 10604
rect 55234 10564 55276 10604
rect 55316 10564 55358 10604
rect 55398 10564 55440 10604
rect 55112 10555 55480 10564
rect 59112 10604 59480 10613
rect 59152 10564 59194 10604
rect 59234 10564 59276 10604
rect 59316 10564 59358 10604
rect 59398 10564 59440 10604
rect 59112 10555 59480 10564
rect 63112 10604 63480 10613
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63112 10555 63480 10564
rect 67112 10604 67480 10613
rect 67152 10564 67194 10604
rect 67234 10564 67276 10604
rect 67316 10564 67358 10604
rect 67398 10564 67440 10604
rect 67112 10555 67480 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 8352 9848 8720 9857
rect 8392 9808 8434 9848
rect 8474 9808 8516 9848
rect 8556 9808 8598 9848
rect 8638 9808 8680 9848
rect 8352 9799 8720 9808
rect 12352 9848 12720 9857
rect 12392 9808 12434 9848
rect 12474 9808 12516 9848
rect 12556 9808 12598 9848
rect 12638 9808 12680 9848
rect 12352 9799 12720 9808
rect 16352 9848 16720 9857
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16352 9799 16720 9808
rect 20352 9848 20720 9857
rect 20392 9808 20434 9848
rect 20474 9808 20516 9848
rect 20556 9808 20598 9848
rect 20638 9808 20680 9848
rect 20352 9799 20720 9808
rect 24352 9848 24720 9857
rect 24392 9808 24434 9848
rect 24474 9808 24516 9848
rect 24556 9808 24598 9848
rect 24638 9808 24680 9848
rect 24352 9799 24720 9808
rect 28352 9848 28720 9857
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28352 9799 28720 9808
rect 32352 9848 32720 9857
rect 32392 9808 32434 9848
rect 32474 9808 32516 9848
rect 32556 9808 32598 9848
rect 32638 9808 32680 9848
rect 32352 9799 32720 9808
rect 36352 9848 36720 9857
rect 36392 9808 36434 9848
rect 36474 9808 36516 9848
rect 36556 9808 36598 9848
rect 36638 9808 36680 9848
rect 36352 9799 36720 9808
rect 40352 9848 40720 9857
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40352 9799 40720 9808
rect 44352 9848 44720 9857
rect 44392 9808 44434 9848
rect 44474 9808 44516 9848
rect 44556 9808 44598 9848
rect 44638 9808 44680 9848
rect 44352 9799 44720 9808
rect 48352 9848 48720 9857
rect 48392 9808 48434 9848
rect 48474 9808 48516 9848
rect 48556 9808 48598 9848
rect 48638 9808 48680 9848
rect 48352 9799 48720 9808
rect 52352 9848 52720 9857
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52352 9799 52720 9808
rect 56352 9848 56720 9857
rect 56392 9808 56434 9848
rect 56474 9808 56516 9848
rect 56556 9808 56598 9848
rect 56638 9808 56680 9848
rect 56352 9799 56720 9808
rect 60352 9848 60720 9857
rect 60392 9808 60434 9848
rect 60474 9808 60516 9848
rect 60556 9808 60598 9848
rect 60638 9808 60680 9848
rect 60352 9799 60720 9808
rect 64352 9848 64720 9857
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64352 9799 64720 9808
rect 68352 9848 68720 9857
rect 68392 9808 68434 9848
rect 68474 9808 68516 9848
rect 68556 9808 68598 9848
rect 68638 9808 68680 9848
rect 68352 9799 68720 9808
rect 80140 9764 80180 9773
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 7112 9092 7480 9101
rect 7152 9052 7194 9092
rect 7234 9052 7276 9092
rect 7316 9052 7358 9092
rect 7398 9052 7440 9092
rect 7112 9043 7480 9052
rect 11112 9092 11480 9101
rect 11152 9052 11194 9092
rect 11234 9052 11276 9092
rect 11316 9052 11358 9092
rect 11398 9052 11440 9092
rect 11112 9043 11480 9052
rect 15112 9092 15480 9101
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15112 9043 15480 9052
rect 19112 9092 19480 9101
rect 19152 9052 19194 9092
rect 19234 9052 19276 9092
rect 19316 9052 19358 9092
rect 19398 9052 19440 9092
rect 19112 9043 19480 9052
rect 23112 9092 23480 9101
rect 23152 9052 23194 9092
rect 23234 9052 23276 9092
rect 23316 9052 23358 9092
rect 23398 9052 23440 9092
rect 23112 9043 23480 9052
rect 27112 9092 27480 9101
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27112 9043 27480 9052
rect 31112 9092 31480 9101
rect 31152 9052 31194 9092
rect 31234 9052 31276 9092
rect 31316 9052 31358 9092
rect 31398 9052 31440 9092
rect 31112 9043 31480 9052
rect 35112 9092 35480 9101
rect 35152 9052 35194 9092
rect 35234 9052 35276 9092
rect 35316 9052 35358 9092
rect 35398 9052 35440 9092
rect 35112 9043 35480 9052
rect 39112 9092 39480 9101
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39112 9043 39480 9052
rect 43112 9092 43480 9101
rect 43152 9052 43194 9092
rect 43234 9052 43276 9092
rect 43316 9052 43358 9092
rect 43398 9052 43440 9092
rect 43112 9043 43480 9052
rect 47112 9092 47480 9101
rect 47152 9052 47194 9092
rect 47234 9052 47276 9092
rect 47316 9052 47358 9092
rect 47398 9052 47440 9092
rect 47112 9043 47480 9052
rect 51112 9092 51480 9101
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51112 9043 51480 9052
rect 55112 9092 55480 9101
rect 55152 9052 55194 9092
rect 55234 9052 55276 9092
rect 55316 9052 55358 9092
rect 55398 9052 55440 9092
rect 55112 9043 55480 9052
rect 59112 9092 59480 9101
rect 59152 9052 59194 9092
rect 59234 9052 59276 9092
rect 59316 9052 59358 9092
rect 59398 9052 59440 9092
rect 59112 9043 59480 9052
rect 63112 9092 63480 9101
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63112 9043 63480 9052
rect 67112 9092 67480 9101
rect 67152 9052 67194 9092
rect 67234 9052 67276 9092
rect 67316 9052 67358 9092
rect 67398 9052 67440 9092
rect 67112 9043 67480 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 8352 8336 8720 8345
rect 8392 8296 8434 8336
rect 8474 8296 8516 8336
rect 8556 8296 8598 8336
rect 8638 8296 8680 8336
rect 8352 8287 8720 8296
rect 12352 8336 12720 8345
rect 12392 8296 12434 8336
rect 12474 8296 12516 8336
rect 12556 8296 12598 8336
rect 12638 8296 12680 8336
rect 12352 8287 12720 8296
rect 16352 8336 16720 8345
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16352 8287 16720 8296
rect 20352 8336 20720 8345
rect 20392 8296 20434 8336
rect 20474 8296 20516 8336
rect 20556 8296 20598 8336
rect 20638 8296 20680 8336
rect 20352 8287 20720 8296
rect 24352 8336 24720 8345
rect 24392 8296 24434 8336
rect 24474 8296 24516 8336
rect 24556 8296 24598 8336
rect 24638 8296 24680 8336
rect 24352 8287 24720 8296
rect 28352 8336 28720 8345
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28352 8287 28720 8296
rect 32352 8336 32720 8345
rect 32392 8296 32434 8336
rect 32474 8296 32516 8336
rect 32556 8296 32598 8336
rect 32638 8296 32680 8336
rect 32352 8287 32720 8296
rect 36352 8336 36720 8345
rect 36392 8296 36434 8336
rect 36474 8296 36516 8336
rect 36556 8296 36598 8336
rect 36638 8296 36680 8336
rect 36352 8287 36720 8296
rect 40352 8336 40720 8345
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40352 8287 40720 8296
rect 44352 8336 44720 8345
rect 44392 8296 44434 8336
rect 44474 8296 44516 8336
rect 44556 8296 44598 8336
rect 44638 8296 44680 8336
rect 44352 8287 44720 8296
rect 48352 8336 48720 8345
rect 48392 8296 48434 8336
rect 48474 8296 48516 8336
rect 48556 8296 48598 8336
rect 48638 8296 48680 8336
rect 48352 8287 48720 8296
rect 52352 8336 52720 8345
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52352 8287 52720 8296
rect 56352 8336 56720 8345
rect 56392 8296 56434 8336
rect 56474 8296 56516 8336
rect 56556 8296 56598 8336
rect 56638 8296 56680 8336
rect 56352 8287 56720 8296
rect 60352 8336 60720 8345
rect 60392 8296 60434 8336
rect 60474 8296 60516 8336
rect 60556 8296 60598 8336
rect 60638 8296 60680 8336
rect 60352 8287 60720 8296
rect 64352 8336 64720 8345
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64352 8287 64720 8296
rect 68352 8336 68720 8345
rect 68392 8296 68434 8336
rect 68474 8296 68516 8336
rect 68556 8296 68598 8336
rect 68638 8296 68680 8336
rect 68352 8287 68720 8296
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 7112 7580 7480 7589
rect 7152 7540 7194 7580
rect 7234 7540 7276 7580
rect 7316 7540 7358 7580
rect 7398 7540 7440 7580
rect 7112 7531 7480 7540
rect 11112 7580 11480 7589
rect 11152 7540 11194 7580
rect 11234 7540 11276 7580
rect 11316 7540 11358 7580
rect 11398 7540 11440 7580
rect 11112 7531 11480 7540
rect 15112 7580 15480 7589
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15112 7531 15480 7540
rect 19112 7580 19480 7589
rect 19152 7540 19194 7580
rect 19234 7540 19276 7580
rect 19316 7540 19358 7580
rect 19398 7540 19440 7580
rect 19112 7531 19480 7540
rect 23112 7580 23480 7589
rect 23152 7540 23194 7580
rect 23234 7540 23276 7580
rect 23316 7540 23358 7580
rect 23398 7540 23440 7580
rect 23112 7531 23480 7540
rect 27112 7580 27480 7589
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27112 7531 27480 7540
rect 31112 7580 31480 7589
rect 31152 7540 31194 7580
rect 31234 7540 31276 7580
rect 31316 7540 31358 7580
rect 31398 7540 31440 7580
rect 31112 7531 31480 7540
rect 35112 7580 35480 7589
rect 35152 7540 35194 7580
rect 35234 7540 35276 7580
rect 35316 7540 35358 7580
rect 35398 7540 35440 7580
rect 35112 7531 35480 7540
rect 39112 7580 39480 7589
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39112 7531 39480 7540
rect 43112 7580 43480 7589
rect 43152 7540 43194 7580
rect 43234 7540 43276 7580
rect 43316 7540 43358 7580
rect 43398 7540 43440 7580
rect 43112 7531 43480 7540
rect 47112 7580 47480 7589
rect 47152 7540 47194 7580
rect 47234 7540 47276 7580
rect 47316 7540 47358 7580
rect 47398 7540 47440 7580
rect 47112 7531 47480 7540
rect 51112 7580 51480 7589
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51112 7531 51480 7540
rect 55112 7580 55480 7589
rect 55152 7540 55194 7580
rect 55234 7540 55276 7580
rect 55316 7540 55358 7580
rect 55398 7540 55440 7580
rect 55112 7531 55480 7540
rect 59112 7580 59480 7589
rect 59152 7540 59194 7580
rect 59234 7540 59276 7580
rect 59316 7540 59358 7580
rect 59398 7540 59440 7580
rect 59112 7531 59480 7540
rect 63112 7580 63480 7589
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63112 7531 63480 7540
rect 67112 7580 67480 7589
rect 67152 7540 67194 7580
rect 67234 7540 67276 7580
rect 67316 7540 67358 7580
rect 67398 7540 67440 7580
rect 67112 7531 67480 7540
rect 71112 7580 71480 7589
rect 71152 7540 71194 7580
rect 71234 7540 71276 7580
rect 71316 7540 71358 7580
rect 71398 7540 71440 7580
rect 71112 7531 71480 7540
rect 75112 7580 75480 7589
rect 75152 7540 75194 7580
rect 75234 7540 75276 7580
rect 75316 7540 75358 7580
rect 75398 7540 75440 7580
rect 75112 7531 75480 7540
rect 79112 7580 79480 7589
rect 79152 7540 79194 7580
rect 79234 7540 79276 7580
rect 79316 7540 79358 7580
rect 79398 7540 79440 7580
rect 79112 7531 79480 7540
rect 76780 7412 76820 7421
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 8352 6824 8720 6833
rect 8392 6784 8434 6824
rect 8474 6784 8516 6824
rect 8556 6784 8598 6824
rect 8638 6784 8680 6824
rect 8352 6775 8720 6784
rect 12352 6824 12720 6833
rect 12392 6784 12434 6824
rect 12474 6784 12516 6824
rect 12556 6784 12598 6824
rect 12638 6784 12680 6824
rect 12352 6775 12720 6784
rect 16352 6824 16720 6833
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16352 6775 16720 6784
rect 20352 6824 20720 6833
rect 20392 6784 20434 6824
rect 20474 6784 20516 6824
rect 20556 6784 20598 6824
rect 20638 6784 20680 6824
rect 20352 6775 20720 6784
rect 24352 6824 24720 6833
rect 24392 6784 24434 6824
rect 24474 6784 24516 6824
rect 24556 6784 24598 6824
rect 24638 6784 24680 6824
rect 24352 6775 24720 6784
rect 28352 6824 28720 6833
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28352 6775 28720 6784
rect 32352 6824 32720 6833
rect 32392 6784 32434 6824
rect 32474 6784 32516 6824
rect 32556 6784 32598 6824
rect 32638 6784 32680 6824
rect 32352 6775 32720 6784
rect 36352 6824 36720 6833
rect 36392 6784 36434 6824
rect 36474 6784 36516 6824
rect 36556 6784 36598 6824
rect 36638 6784 36680 6824
rect 36352 6775 36720 6784
rect 40352 6824 40720 6833
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40352 6775 40720 6784
rect 44352 6824 44720 6833
rect 44392 6784 44434 6824
rect 44474 6784 44516 6824
rect 44556 6784 44598 6824
rect 44638 6784 44680 6824
rect 44352 6775 44720 6784
rect 48352 6824 48720 6833
rect 48392 6784 48434 6824
rect 48474 6784 48516 6824
rect 48556 6784 48598 6824
rect 48638 6784 48680 6824
rect 48352 6775 48720 6784
rect 52352 6824 52720 6833
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52352 6775 52720 6784
rect 56352 6824 56720 6833
rect 56392 6784 56434 6824
rect 56474 6784 56516 6824
rect 56556 6784 56598 6824
rect 56638 6784 56680 6824
rect 56352 6775 56720 6784
rect 60352 6824 60720 6833
rect 60392 6784 60434 6824
rect 60474 6784 60516 6824
rect 60556 6784 60598 6824
rect 60638 6784 60680 6824
rect 60352 6775 60720 6784
rect 64352 6824 64720 6833
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64352 6775 64720 6784
rect 68352 6824 68720 6833
rect 68392 6784 68434 6824
rect 68474 6784 68516 6824
rect 68556 6784 68598 6824
rect 68638 6784 68680 6824
rect 68352 6775 68720 6784
rect 72352 6824 72720 6833
rect 72392 6784 72434 6824
rect 72474 6784 72516 6824
rect 72556 6784 72598 6824
rect 72638 6784 72680 6824
rect 72352 6775 72720 6784
rect 76352 6824 76720 6833
rect 76392 6784 76434 6824
rect 76474 6784 76516 6824
rect 76556 6784 76598 6824
rect 76638 6784 76680 6824
rect 76352 6775 76720 6784
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 7112 6068 7480 6077
rect 7152 6028 7194 6068
rect 7234 6028 7276 6068
rect 7316 6028 7358 6068
rect 7398 6028 7440 6068
rect 7112 6019 7480 6028
rect 11112 6068 11480 6077
rect 11152 6028 11194 6068
rect 11234 6028 11276 6068
rect 11316 6028 11358 6068
rect 11398 6028 11440 6068
rect 11112 6019 11480 6028
rect 15112 6068 15480 6077
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15112 6019 15480 6028
rect 19112 6068 19480 6077
rect 19152 6028 19194 6068
rect 19234 6028 19276 6068
rect 19316 6028 19358 6068
rect 19398 6028 19440 6068
rect 19112 6019 19480 6028
rect 23112 6068 23480 6077
rect 23152 6028 23194 6068
rect 23234 6028 23276 6068
rect 23316 6028 23358 6068
rect 23398 6028 23440 6068
rect 23112 6019 23480 6028
rect 27112 6068 27480 6077
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27112 6019 27480 6028
rect 31112 6068 31480 6077
rect 31152 6028 31194 6068
rect 31234 6028 31276 6068
rect 31316 6028 31358 6068
rect 31398 6028 31440 6068
rect 31112 6019 31480 6028
rect 35112 6068 35480 6077
rect 35152 6028 35194 6068
rect 35234 6028 35276 6068
rect 35316 6028 35358 6068
rect 35398 6028 35440 6068
rect 35112 6019 35480 6028
rect 39112 6068 39480 6077
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39112 6019 39480 6028
rect 43112 6068 43480 6077
rect 43152 6028 43194 6068
rect 43234 6028 43276 6068
rect 43316 6028 43358 6068
rect 43398 6028 43440 6068
rect 43112 6019 43480 6028
rect 47112 6068 47480 6077
rect 47152 6028 47194 6068
rect 47234 6028 47276 6068
rect 47316 6028 47358 6068
rect 47398 6028 47440 6068
rect 47112 6019 47480 6028
rect 51112 6068 51480 6077
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51112 6019 51480 6028
rect 55112 6068 55480 6077
rect 55152 6028 55194 6068
rect 55234 6028 55276 6068
rect 55316 6028 55358 6068
rect 55398 6028 55440 6068
rect 55112 6019 55480 6028
rect 59112 6068 59480 6077
rect 59152 6028 59194 6068
rect 59234 6028 59276 6068
rect 59316 6028 59358 6068
rect 59398 6028 59440 6068
rect 59112 6019 59480 6028
rect 63112 6068 63480 6077
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63112 6019 63480 6028
rect 67112 6068 67480 6077
rect 67152 6028 67194 6068
rect 67234 6028 67276 6068
rect 67316 6028 67358 6068
rect 67398 6028 67440 6068
rect 67112 6019 67480 6028
rect 71112 6068 71480 6077
rect 71152 6028 71194 6068
rect 71234 6028 71276 6068
rect 71316 6028 71358 6068
rect 71398 6028 71440 6068
rect 71112 6019 71480 6028
rect 75112 6068 75480 6077
rect 75152 6028 75194 6068
rect 75234 6028 75276 6068
rect 75316 6028 75358 6068
rect 75398 6028 75440 6068
rect 75112 6019 75480 6028
rect 76780 5900 76820 7372
rect 79112 6068 79480 6077
rect 79152 6028 79194 6068
rect 79234 6028 79276 6068
rect 79316 6028 79358 6068
rect 79398 6028 79440 6068
rect 79112 6019 79480 6028
rect 76780 5851 76820 5860
rect 80140 5900 80180 9724
rect 83596 9764 83636 9773
rect 82924 7916 82964 7925
rect 82924 7076 82964 7876
rect 83112 7580 83480 7589
rect 83152 7540 83194 7580
rect 83234 7540 83276 7580
rect 83316 7540 83358 7580
rect 83398 7540 83440 7580
rect 83112 7531 83480 7540
rect 82924 7027 82964 7036
rect 80352 6824 80720 6833
rect 80392 6784 80434 6824
rect 80474 6784 80516 6824
rect 80556 6784 80598 6824
rect 80638 6784 80680 6824
rect 80352 6775 80720 6784
rect 83112 6068 83480 6077
rect 83152 6028 83194 6068
rect 83234 6028 83276 6068
rect 83316 6028 83358 6068
rect 83398 6028 83440 6068
rect 83112 6019 83480 6028
rect 80140 5851 80180 5860
rect 83596 5900 83636 9724
rect 89068 9764 89108 9773
rect 85612 8840 85652 8849
rect 84352 6824 84720 6833
rect 84392 6784 84434 6824
rect 84474 6784 84516 6824
rect 84556 6784 84598 6824
rect 84638 6784 84680 6824
rect 84352 6775 84720 6784
rect 83596 5851 83636 5860
rect 85612 5900 85652 8800
rect 87112 7580 87480 7589
rect 87152 7540 87194 7580
rect 87234 7540 87276 7580
rect 87316 7540 87358 7580
rect 87398 7540 87440 7580
rect 87112 7531 87480 7540
rect 86667 7412 86709 7421
rect 86667 7372 86668 7412
rect 86708 7372 86709 7412
rect 86667 7363 86709 7372
rect 86668 7278 86708 7363
rect 88204 6992 88244 7001
rect 88204 6656 88244 6952
rect 88352 6824 88720 6833
rect 88392 6784 88434 6824
rect 88474 6784 88516 6824
rect 88556 6784 88598 6824
rect 88638 6784 88680 6824
rect 88352 6775 88720 6784
rect 88204 6607 88244 6616
rect 87112 6068 87480 6077
rect 87152 6028 87194 6068
rect 87234 6028 87276 6068
rect 87316 6028 87358 6068
rect 87398 6028 87440 6068
rect 87112 6019 87480 6028
rect 85612 5851 85652 5860
rect 89068 5900 89108 9724
rect 98860 9512 98900 15436
rect 98860 9463 98900 9472
rect 95596 7832 95636 7841
rect 91112 7580 91480 7589
rect 91152 7540 91194 7580
rect 91234 7540 91276 7580
rect 91316 7540 91358 7580
rect 91398 7540 91440 7580
rect 91112 7531 91480 7540
rect 95112 7580 95480 7589
rect 95152 7540 95194 7580
rect 95234 7540 95276 7580
rect 95316 7540 95358 7580
rect 95398 7540 95440 7580
rect 95112 7531 95480 7540
rect 92352 6824 92720 6833
rect 92392 6784 92434 6824
rect 92474 6784 92516 6824
rect 92556 6784 92598 6824
rect 92638 6784 92680 6824
rect 92352 6775 92720 6784
rect 95596 6740 95636 7792
rect 99112 7580 99480 7589
rect 99152 7540 99194 7580
rect 99234 7540 99276 7580
rect 99316 7540 99358 7580
rect 99398 7540 99440 7580
rect 99112 7531 99480 7540
rect 96352 6824 96720 6833
rect 96392 6784 96434 6824
rect 96474 6784 96516 6824
rect 96556 6784 96598 6824
rect 96638 6784 96680 6824
rect 96352 6775 96720 6784
rect 95596 6691 95636 6700
rect 91112 6068 91480 6077
rect 91152 6028 91194 6068
rect 91234 6028 91276 6068
rect 91316 6028 91358 6068
rect 91398 6028 91440 6068
rect 91112 6019 91480 6028
rect 95112 6068 95480 6077
rect 95152 6028 95194 6068
rect 95234 6028 95276 6068
rect 95316 6028 95358 6068
rect 95398 6028 95440 6068
rect 95112 6019 95480 6028
rect 99112 6068 99480 6077
rect 99152 6028 99194 6068
rect 99234 6028 99276 6068
rect 99316 6028 99358 6068
rect 99398 6028 99440 6068
rect 99112 6019 99480 6028
rect 89068 5851 89108 5860
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 8352 5312 8720 5321
rect 8392 5272 8434 5312
rect 8474 5272 8516 5312
rect 8556 5272 8598 5312
rect 8638 5272 8680 5312
rect 8352 5263 8720 5272
rect 12352 5312 12720 5321
rect 12392 5272 12434 5312
rect 12474 5272 12516 5312
rect 12556 5272 12598 5312
rect 12638 5272 12680 5312
rect 12352 5263 12720 5272
rect 16352 5312 16720 5321
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16352 5263 16720 5272
rect 20352 5312 20720 5321
rect 20392 5272 20434 5312
rect 20474 5272 20516 5312
rect 20556 5272 20598 5312
rect 20638 5272 20680 5312
rect 20352 5263 20720 5272
rect 24352 5312 24720 5321
rect 24392 5272 24434 5312
rect 24474 5272 24516 5312
rect 24556 5272 24598 5312
rect 24638 5272 24680 5312
rect 24352 5263 24720 5272
rect 28352 5312 28720 5321
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28352 5263 28720 5272
rect 32352 5312 32720 5321
rect 32392 5272 32434 5312
rect 32474 5272 32516 5312
rect 32556 5272 32598 5312
rect 32638 5272 32680 5312
rect 32352 5263 32720 5272
rect 36352 5312 36720 5321
rect 36392 5272 36434 5312
rect 36474 5272 36516 5312
rect 36556 5272 36598 5312
rect 36638 5272 36680 5312
rect 36352 5263 36720 5272
rect 40352 5312 40720 5321
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40352 5263 40720 5272
rect 44352 5312 44720 5321
rect 44392 5272 44434 5312
rect 44474 5272 44516 5312
rect 44556 5272 44598 5312
rect 44638 5272 44680 5312
rect 44352 5263 44720 5272
rect 48352 5312 48720 5321
rect 48392 5272 48434 5312
rect 48474 5272 48516 5312
rect 48556 5272 48598 5312
rect 48638 5272 48680 5312
rect 48352 5263 48720 5272
rect 52352 5312 52720 5321
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52352 5263 52720 5272
rect 56352 5312 56720 5321
rect 56392 5272 56434 5312
rect 56474 5272 56516 5312
rect 56556 5272 56598 5312
rect 56638 5272 56680 5312
rect 56352 5263 56720 5272
rect 60352 5312 60720 5321
rect 60392 5272 60434 5312
rect 60474 5272 60516 5312
rect 60556 5272 60598 5312
rect 60638 5272 60680 5312
rect 60352 5263 60720 5272
rect 64352 5312 64720 5321
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64352 5263 64720 5272
rect 68352 5312 68720 5321
rect 68392 5272 68434 5312
rect 68474 5272 68516 5312
rect 68556 5272 68598 5312
rect 68638 5272 68680 5312
rect 68352 5263 68720 5272
rect 72352 5312 72720 5321
rect 72392 5272 72434 5312
rect 72474 5272 72516 5312
rect 72556 5272 72598 5312
rect 72638 5272 72680 5312
rect 72352 5263 72720 5272
rect 76352 5312 76720 5321
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76352 5263 76720 5272
rect 80352 5312 80720 5321
rect 80392 5272 80434 5312
rect 80474 5272 80516 5312
rect 80556 5272 80598 5312
rect 80638 5272 80680 5312
rect 80352 5263 80720 5272
rect 84352 5312 84720 5321
rect 84392 5272 84434 5312
rect 84474 5272 84516 5312
rect 84556 5272 84598 5312
rect 84638 5272 84680 5312
rect 84352 5263 84720 5272
rect 88352 5312 88720 5321
rect 88392 5272 88434 5312
rect 88474 5272 88516 5312
rect 88556 5272 88598 5312
rect 88638 5272 88680 5312
rect 88352 5263 88720 5272
rect 92352 5312 92720 5321
rect 92392 5272 92434 5312
rect 92474 5272 92516 5312
rect 92556 5272 92598 5312
rect 92638 5272 92680 5312
rect 92352 5263 92720 5272
rect 96352 5312 96720 5321
rect 96392 5272 96434 5312
rect 96474 5272 96516 5312
rect 96556 5272 96598 5312
rect 96638 5272 96680 5312
rect 96352 5263 96720 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 7112 4556 7480 4565
rect 7152 4516 7194 4556
rect 7234 4516 7276 4556
rect 7316 4516 7358 4556
rect 7398 4516 7440 4556
rect 7112 4507 7480 4516
rect 11112 4556 11480 4565
rect 11152 4516 11194 4556
rect 11234 4516 11276 4556
rect 11316 4516 11358 4556
rect 11398 4516 11440 4556
rect 11112 4507 11480 4516
rect 15112 4556 15480 4565
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15112 4507 15480 4516
rect 19112 4556 19480 4565
rect 19152 4516 19194 4556
rect 19234 4516 19276 4556
rect 19316 4516 19358 4556
rect 19398 4516 19440 4556
rect 19112 4507 19480 4516
rect 23112 4556 23480 4565
rect 23152 4516 23194 4556
rect 23234 4516 23276 4556
rect 23316 4516 23358 4556
rect 23398 4516 23440 4556
rect 23112 4507 23480 4516
rect 27112 4556 27480 4565
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27112 4507 27480 4516
rect 31112 4556 31480 4565
rect 31152 4516 31194 4556
rect 31234 4516 31276 4556
rect 31316 4516 31358 4556
rect 31398 4516 31440 4556
rect 31112 4507 31480 4516
rect 35112 4556 35480 4565
rect 35152 4516 35194 4556
rect 35234 4516 35276 4556
rect 35316 4516 35358 4556
rect 35398 4516 35440 4556
rect 35112 4507 35480 4516
rect 39112 4556 39480 4565
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39112 4507 39480 4516
rect 43112 4556 43480 4565
rect 43152 4516 43194 4556
rect 43234 4516 43276 4556
rect 43316 4516 43358 4556
rect 43398 4516 43440 4556
rect 43112 4507 43480 4516
rect 47112 4556 47480 4565
rect 47152 4516 47194 4556
rect 47234 4516 47276 4556
rect 47316 4516 47358 4556
rect 47398 4516 47440 4556
rect 47112 4507 47480 4516
rect 51112 4556 51480 4565
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51112 4507 51480 4516
rect 55112 4556 55480 4565
rect 55152 4516 55194 4556
rect 55234 4516 55276 4556
rect 55316 4516 55358 4556
rect 55398 4516 55440 4556
rect 55112 4507 55480 4516
rect 59112 4556 59480 4565
rect 59152 4516 59194 4556
rect 59234 4516 59276 4556
rect 59316 4516 59358 4556
rect 59398 4516 59440 4556
rect 59112 4507 59480 4516
rect 63112 4556 63480 4565
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63112 4507 63480 4516
rect 67112 4556 67480 4565
rect 67152 4516 67194 4556
rect 67234 4516 67276 4556
rect 67316 4516 67358 4556
rect 67398 4516 67440 4556
rect 67112 4507 67480 4516
rect 71112 4556 71480 4565
rect 71152 4516 71194 4556
rect 71234 4516 71276 4556
rect 71316 4516 71358 4556
rect 71398 4516 71440 4556
rect 71112 4507 71480 4516
rect 75112 4556 75480 4565
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75112 4507 75480 4516
rect 79112 4556 79480 4565
rect 79152 4516 79194 4556
rect 79234 4516 79276 4556
rect 79316 4516 79358 4556
rect 79398 4516 79440 4556
rect 79112 4507 79480 4516
rect 83112 4556 83480 4565
rect 83152 4516 83194 4556
rect 83234 4516 83276 4556
rect 83316 4516 83358 4556
rect 83398 4516 83440 4556
rect 83112 4507 83480 4516
rect 87112 4556 87480 4565
rect 87152 4516 87194 4556
rect 87234 4516 87276 4556
rect 87316 4516 87358 4556
rect 87398 4516 87440 4556
rect 87112 4507 87480 4516
rect 91112 4556 91480 4565
rect 91152 4516 91194 4556
rect 91234 4516 91276 4556
rect 91316 4516 91358 4556
rect 91398 4516 91440 4556
rect 91112 4507 91480 4516
rect 95112 4556 95480 4565
rect 95152 4516 95194 4556
rect 95234 4516 95276 4556
rect 95316 4516 95358 4556
rect 95398 4516 95440 4556
rect 95112 4507 95480 4516
rect 99112 4556 99480 4565
rect 99152 4516 99194 4556
rect 99234 4516 99276 4556
rect 99316 4516 99358 4556
rect 99398 4516 99440 4556
rect 99112 4507 99480 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 8352 3800 8720 3809
rect 8392 3760 8434 3800
rect 8474 3760 8516 3800
rect 8556 3760 8598 3800
rect 8638 3760 8680 3800
rect 8352 3751 8720 3760
rect 12352 3800 12720 3809
rect 12392 3760 12434 3800
rect 12474 3760 12516 3800
rect 12556 3760 12598 3800
rect 12638 3760 12680 3800
rect 12352 3751 12720 3760
rect 16352 3800 16720 3809
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16352 3751 16720 3760
rect 20352 3800 20720 3809
rect 20392 3760 20434 3800
rect 20474 3760 20516 3800
rect 20556 3760 20598 3800
rect 20638 3760 20680 3800
rect 20352 3751 20720 3760
rect 24352 3800 24720 3809
rect 24392 3760 24434 3800
rect 24474 3760 24516 3800
rect 24556 3760 24598 3800
rect 24638 3760 24680 3800
rect 24352 3751 24720 3760
rect 28352 3800 28720 3809
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28352 3751 28720 3760
rect 32352 3800 32720 3809
rect 32392 3760 32434 3800
rect 32474 3760 32516 3800
rect 32556 3760 32598 3800
rect 32638 3760 32680 3800
rect 32352 3751 32720 3760
rect 36352 3800 36720 3809
rect 36392 3760 36434 3800
rect 36474 3760 36516 3800
rect 36556 3760 36598 3800
rect 36638 3760 36680 3800
rect 36352 3751 36720 3760
rect 40352 3800 40720 3809
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40352 3751 40720 3760
rect 44352 3800 44720 3809
rect 44392 3760 44434 3800
rect 44474 3760 44516 3800
rect 44556 3760 44598 3800
rect 44638 3760 44680 3800
rect 44352 3751 44720 3760
rect 48352 3800 48720 3809
rect 48392 3760 48434 3800
rect 48474 3760 48516 3800
rect 48556 3760 48598 3800
rect 48638 3760 48680 3800
rect 48352 3751 48720 3760
rect 52352 3800 52720 3809
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52352 3751 52720 3760
rect 56352 3800 56720 3809
rect 56392 3760 56434 3800
rect 56474 3760 56516 3800
rect 56556 3760 56598 3800
rect 56638 3760 56680 3800
rect 56352 3751 56720 3760
rect 60352 3800 60720 3809
rect 60392 3760 60434 3800
rect 60474 3760 60516 3800
rect 60556 3760 60598 3800
rect 60638 3760 60680 3800
rect 60352 3751 60720 3760
rect 64352 3800 64720 3809
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64352 3751 64720 3760
rect 68352 3800 68720 3809
rect 68392 3760 68434 3800
rect 68474 3760 68516 3800
rect 68556 3760 68598 3800
rect 68638 3760 68680 3800
rect 68352 3751 68720 3760
rect 72352 3800 72720 3809
rect 72392 3760 72434 3800
rect 72474 3760 72516 3800
rect 72556 3760 72598 3800
rect 72638 3760 72680 3800
rect 72352 3751 72720 3760
rect 76352 3800 76720 3809
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76352 3751 76720 3760
rect 80352 3800 80720 3809
rect 80392 3760 80434 3800
rect 80474 3760 80516 3800
rect 80556 3760 80598 3800
rect 80638 3760 80680 3800
rect 80352 3751 80720 3760
rect 84352 3800 84720 3809
rect 84392 3760 84434 3800
rect 84474 3760 84516 3800
rect 84556 3760 84598 3800
rect 84638 3760 84680 3800
rect 84352 3751 84720 3760
rect 88352 3800 88720 3809
rect 88392 3760 88434 3800
rect 88474 3760 88516 3800
rect 88556 3760 88598 3800
rect 88638 3760 88680 3800
rect 88352 3751 88720 3760
rect 92352 3800 92720 3809
rect 92392 3760 92434 3800
rect 92474 3760 92516 3800
rect 92556 3760 92598 3800
rect 92638 3760 92680 3800
rect 92352 3751 92720 3760
rect 96352 3800 96720 3809
rect 96392 3760 96434 3800
rect 96474 3760 96516 3800
rect 96556 3760 96598 3800
rect 96638 3760 96680 3800
rect 96352 3751 96720 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 7112 3044 7480 3053
rect 7152 3004 7194 3044
rect 7234 3004 7276 3044
rect 7316 3004 7358 3044
rect 7398 3004 7440 3044
rect 7112 2995 7480 3004
rect 11112 3044 11480 3053
rect 11152 3004 11194 3044
rect 11234 3004 11276 3044
rect 11316 3004 11358 3044
rect 11398 3004 11440 3044
rect 11112 2995 11480 3004
rect 15112 3044 15480 3053
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15112 2995 15480 3004
rect 19112 3044 19480 3053
rect 19152 3004 19194 3044
rect 19234 3004 19276 3044
rect 19316 3004 19358 3044
rect 19398 3004 19440 3044
rect 19112 2995 19480 3004
rect 23112 3044 23480 3053
rect 23152 3004 23194 3044
rect 23234 3004 23276 3044
rect 23316 3004 23358 3044
rect 23398 3004 23440 3044
rect 23112 2995 23480 3004
rect 27112 3044 27480 3053
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27112 2995 27480 3004
rect 31112 3044 31480 3053
rect 31152 3004 31194 3044
rect 31234 3004 31276 3044
rect 31316 3004 31358 3044
rect 31398 3004 31440 3044
rect 31112 2995 31480 3004
rect 35112 3044 35480 3053
rect 35152 3004 35194 3044
rect 35234 3004 35276 3044
rect 35316 3004 35358 3044
rect 35398 3004 35440 3044
rect 35112 2995 35480 3004
rect 39112 3044 39480 3053
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39112 2995 39480 3004
rect 43112 3044 43480 3053
rect 43152 3004 43194 3044
rect 43234 3004 43276 3044
rect 43316 3004 43358 3044
rect 43398 3004 43440 3044
rect 43112 2995 43480 3004
rect 47112 3044 47480 3053
rect 47152 3004 47194 3044
rect 47234 3004 47276 3044
rect 47316 3004 47358 3044
rect 47398 3004 47440 3044
rect 47112 2995 47480 3004
rect 51112 3044 51480 3053
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51112 2995 51480 3004
rect 55112 3044 55480 3053
rect 55152 3004 55194 3044
rect 55234 3004 55276 3044
rect 55316 3004 55358 3044
rect 55398 3004 55440 3044
rect 55112 2995 55480 3004
rect 59112 3044 59480 3053
rect 59152 3004 59194 3044
rect 59234 3004 59276 3044
rect 59316 3004 59358 3044
rect 59398 3004 59440 3044
rect 59112 2995 59480 3004
rect 63112 3044 63480 3053
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63112 2995 63480 3004
rect 67112 3044 67480 3053
rect 67152 3004 67194 3044
rect 67234 3004 67276 3044
rect 67316 3004 67358 3044
rect 67398 3004 67440 3044
rect 67112 2995 67480 3004
rect 71112 3044 71480 3053
rect 71152 3004 71194 3044
rect 71234 3004 71276 3044
rect 71316 3004 71358 3044
rect 71398 3004 71440 3044
rect 71112 2995 71480 3004
rect 75112 3044 75480 3053
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75112 2995 75480 3004
rect 79112 3044 79480 3053
rect 79152 3004 79194 3044
rect 79234 3004 79276 3044
rect 79316 3004 79358 3044
rect 79398 3004 79440 3044
rect 79112 2995 79480 3004
rect 83112 3044 83480 3053
rect 83152 3004 83194 3044
rect 83234 3004 83276 3044
rect 83316 3004 83358 3044
rect 83398 3004 83440 3044
rect 83112 2995 83480 3004
rect 87112 3044 87480 3053
rect 87152 3004 87194 3044
rect 87234 3004 87276 3044
rect 87316 3004 87358 3044
rect 87398 3004 87440 3044
rect 87112 2995 87480 3004
rect 91112 3044 91480 3053
rect 91152 3004 91194 3044
rect 91234 3004 91276 3044
rect 91316 3004 91358 3044
rect 91398 3004 91440 3044
rect 91112 2995 91480 3004
rect 95112 3044 95480 3053
rect 95152 3004 95194 3044
rect 95234 3004 95276 3044
rect 95316 3004 95358 3044
rect 95398 3004 95440 3044
rect 95112 2995 95480 3004
rect 99112 3044 99480 3053
rect 99152 3004 99194 3044
rect 99234 3004 99276 3044
rect 99316 3004 99358 3044
rect 99398 3004 99440 3044
rect 99112 2995 99480 3004
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 8352 2288 8720 2297
rect 8392 2248 8434 2288
rect 8474 2248 8516 2288
rect 8556 2248 8598 2288
rect 8638 2248 8680 2288
rect 8352 2239 8720 2248
rect 12352 2288 12720 2297
rect 12392 2248 12434 2288
rect 12474 2248 12516 2288
rect 12556 2248 12598 2288
rect 12638 2248 12680 2288
rect 12352 2239 12720 2248
rect 16352 2288 16720 2297
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16352 2239 16720 2248
rect 20352 2288 20720 2297
rect 20392 2248 20434 2288
rect 20474 2248 20516 2288
rect 20556 2248 20598 2288
rect 20638 2248 20680 2288
rect 20352 2239 20720 2248
rect 24352 2288 24720 2297
rect 24392 2248 24434 2288
rect 24474 2248 24516 2288
rect 24556 2248 24598 2288
rect 24638 2248 24680 2288
rect 24352 2239 24720 2248
rect 28352 2288 28720 2297
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28352 2239 28720 2248
rect 32352 2288 32720 2297
rect 32392 2248 32434 2288
rect 32474 2248 32516 2288
rect 32556 2248 32598 2288
rect 32638 2248 32680 2288
rect 32352 2239 32720 2248
rect 36352 2288 36720 2297
rect 36392 2248 36434 2288
rect 36474 2248 36516 2288
rect 36556 2248 36598 2288
rect 36638 2248 36680 2288
rect 36352 2239 36720 2248
rect 40352 2288 40720 2297
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40352 2239 40720 2248
rect 44352 2288 44720 2297
rect 44392 2248 44434 2288
rect 44474 2248 44516 2288
rect 44556 2248 44598 2288
rect 44638 2248 44680 2288
rect 44352 2239 44720 2248
rect 48352 2288 48720 2297
rect 48392 2248 48434 2288
rect 48474 2248 48516 2288
rect 48556 2248 48598 2288
rect 48638 2248 48680 2288
rect 48352 2239 48720 2248
rect 52352 2288 52720 2297
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52352 2239 52720 2248
rect 56352 2288 56720 2297
rect 56392 2248 56434 2288
rect 56474 2248 56516 2288
rect 56556 2248 56598 2288
rect 56638 2248 56680 2288
rect 56352 2239 56720 2248
rect 60352 2288 60720 2297
rect 60392 2248 60434 2288
rect 60474 2248 60516 2288
rect 60556 2248 60598 2288
rect 60638 2248 60680 2288
rect 60352 2239 60720 2248
rect 64352 2288 64720 2297
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64352 2239 64720 2248
rect 68352 2288 68720 2297
rect 68392 2248 68434 2288
rect 68474 2248 68516 2288
rect 68556 2248 68598 2288
rect 68638 2248 68680 2288
rect 68352 2239 68720 2248
rect 72352 2288 72720 2297
rect 72392 2248 72434 2288
rect 72474 2248 72516 2288
rect 72556 2248 72598 2288
rect 72638 2248 72680 2288
rect 72352 2239 72720 2248
rect 76352 2288 76720 2297
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76352 2239 76720 2248
rect 80352 2288 80720 2297
rect 80392 2248 80434 2288
rect 80474 2248 80516 2288
rect 80556 2248 80598 2288
rect 80638 2248 80680 2288
rect 80352 2239 80720 2248
rect 84352 2288 84720 2297
rect 84392 2248 84434 2288
rect 84474 2248 84516 2288
rect 84556 2248 84598 2288
rect 84638 2248 84680 2288
rect 84352 2239 84720 2248
rect 88352 2288 88720 2297
rect 88392 2248 88434 2288
rect 88474 2248 88516 2288
rect 88556 2248 88598 2288
rect 88638 2248 88680 2288
rect 88352 2239 88720 2248
rect 92352 2288 92720 2297
rect 92392 2248 92434 2288
rect 92474 2248 92516 2288
rect 92556 2248 92598 2288
rect 92638 2248 92680 2288
rect 92352 2239 92720 2248
rect 96352 2288 96720 2297
rect 96392 2248 96434 2288
rect 96474 2248 96516 2288
rect 96556 2248 96598 2288
rect 96638 2248 96680 2288
rect 96352 2239 96720 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 7112 1532 7480 1541
rect 7152 1492 7194 1532
rect 7234 1492 7276 1532
rect 7316 1492 7358 1532
rect 7398 1492 7440 1532
rect 7112 1483 7480 1492
rect 11112 1532 11480 1541
rect 11152 1492 11194 1532
rect 11234 1492 11276 1532
rect 11316 1492 11358 1532
rect 11398 1492 11440 1532
rect 11112 1483 11480 1492
rect 15112 1532 15480 1541
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15112 1483 15480 1492
rect 19112 1532 19480 1541
rect 19152 1492 19194 1532
rect 19234 1492 19276 1532
rect 19316 1492 19358 1532
rect 19398 1492 19440 1532
rect 19112 1483 19480 1492
rect 23112 1532 23480 1541
rect 23152 1492 23194 1532
rect 23234 1492 23276 1532
rect 23316 1492 23358 1532
rect 23398 1492 23440 1532
rect 23112 1483 23480 1492
rect 27112 1532 27480 1541
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27112 1483 27480 1492
rect 31112 1532 31480 1541
rect 31152 1492 31194 1532
rect 31234 1492 31276 1532
rect 31316 1492 31358 1532
rect 31398 1492 31440 1532
rect 31112 1483 31480 1492
rect 35112 1532 35480 1541
rect 35152 1492 35194 1532
rect 35234 1492 35276 1532
rect 35316 1492 35358 1532
rect 35398 1492 35440 1532
rect 35112 1483 35480 1492
rect 39112 1532 39480 1541
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39112 1483 39480 1492
rect 43112 1532 43480 1541
rect 43152 1492 43194 1532
rect 43234 1492 43276 1532
rect 43316 1492 43358 1532
rect 43398 1492 43440 1532
rect 43112 1483 43480 1492
rect 47112 1532 47480 1541
rect 47152 1492 47194 1532
rect 47234 1492 47276 1532
rect 47316 1492 47358 1532
rect 47398 1492 47440 1532
rect 47112 1483 47480 1492
rect 51112 1532 51480 1541
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51112 1483 51480 1492
rect 55112 1532 55480 1541
rect 55152 1492 55194 1532
rect 55234 1492 55276 1532
rect 55316 1492 55358 1532
rect 55398 1492 55440 1532
rect 55112 1483 55480 1492
rect 59112 1532 59480 1541
rect 59152 1492 59194 1532
rect 59234 1492 59276 1532
rect 59316 1492 59358 1532
rect 59398 1492 59440 1532
rect 59112 1483 59480 1492
rect 63112 1532 63480 1541
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63112 1483 63480 1492
rect 67112 1532 67480 1541
rect 67152 1492 67194 1532
rect 67234 1492 67276 1532
rect 67316 1492 67358 1532
rect 67398 1492 67440 1532
rect 67112 1483 67480 1492
rect 71112 1532 71480 1541
rect 71152 1492 71194 1532
rect 71234 1492 71276 1532
rect 71316 1492 71358 1532
rect 71398 1492 71440 1532
rect 71112 1483 71480 1492
rect 75112 1532 75480 1541
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75112 1483 75480 1492
rect 79112 1532 79480 1541
rect 79152 1492 79194 1532
rect 79234 1492 79276 1532
rect 79316 1492 79358 1532
rect 79398 1492 79440 1532
rect 79112 1483 79480 1492
rect 83112 1532 83480 1541
rect 83152 1492 83194 1532
rect 83234 1492 83276 1532
rect 83316 1492 83358 1532
rect 83398 1492 83440 1532
rect 83112 1483 83480 1492
rect 87112 1532 87480 1541
rect 87152 1492 87194 1532
rect 87234 1492 87276 1532
rect 87316 1492 87358 1532
rect 87398 1492 87440 1532
rect 87112 1483 87480 1492
rect 91112 1532 91480 1541
rect 91152 1492 91194 1532
rect 91234 1492 91276 1532
rect 91316 1492 91358 1532
rect 91398 1492 91440 1532
rect 91112 1483 91480 1492
rect 95112 1532 95480 1541
rect 95152 1492 95194 1532
rect 95234 1492 95276 1532
rect 95316 1492 95358 1532
rect 95398 1492 95440 1532
rect 95112 1483 95480 1492
rect 99112 1532 99480 1541
rect 99152 1492 99194 1532
rect 99234 1492 99276 1532
rect 99316 1492 99358 1532
rect 99398 1492 99440 1532
rect 99112 1483 99480 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 8352 776 8720 785
rect 8392 736 8434 776
rect 8474 736 8516 776
rect 8556 736 8598 776
rect 8638 736 8680 776
rect 8352 727 8720 736
rect 12352 776 12720 785
rect 12392 736 12434 776
rect 12474 736 12516 776
rect 12556 736 12598 776
rect 12638 736 12680 776
rect 12352 727 12720 736
rect 16352 776 16720 785
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16352 727 16720 736
rect 20352 776 20720 785
rect 20392 736 20434 776
rect 20474 736 20516 776
rect 20556 736 20598 776
rect 20638 736 20680 776
rect 20352 727 20720 736
rect 24352 776 24720 785
rect 24392 736 24434 776
rect 24474 736 24516 776
rect 24556 736 24598 776
rect 24638 736 24680 776
rect 24352 727 24720 736
rect 28352 776 28720 785
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28352 727 28720 736
rect 32352 776 32720 785
rect 32392 736 32434 776
rect 32474 736 32516 776
rect 32556 736 32598 776
rect 32638 736 32680 776
rect 32352 727 32720 736
rect 36352 776 36720 785
rect 36392 736 36434 776
rect 36474 736 36516 776
rect 36556 736 36598 776
rect 36638 736 36680 776
rect 36352 727 36720 736
rect 40352 776 40720 785
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40352 727 40720 736
rect 44352 776 44720 785
rect 44392 736 44434 776
rect 44474 736 44516 776
rect 44556 736 44598 776
rect 44638 736 44680 776
rect 44352 727 44720 736
rect 48352 776 48720 785
rect 48392 736 48434 776
rect 48474 736 48516 776
rect 48556 736 48598 776
rect 48638 736 48680 776
rect 48352 727 48720 736
rect 52352 776 52720 785
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52352 727 52720 736
rect 56352 776 56720 785
rect 56392 736 56434 776
rect 56474 736 56516 776
rect 56556 736 56598 776
rect 56638 736 56680 776
rect 56352 727 56720 736
rect 60352 776 60720 785
rect 60392 736 60434 776
rect 60474 736 60516 776
rect 60556 736 60598 776
rect 60638 736 60680 776
rect 60352 727 60720 736
rect 64352 776 64720 785
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64352 727 64720 736
rect 68352 776 68720 785
rect 68392 736 68434 776
rect 68474 736 68516 776
rect 68556 736 68598 776
rect 68638 736 68680 776
rect 68352 727 68720 736
rect 72352 776 72720 785
rect 72392 736 72434 776
rect 72474 736 72516 776
rect 72556 736 72598 776
rect 72638 736 72680 776
rect 72352 727 72720 736
rect 76352 776 76720 785
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76352 727 76720 736
rect 80352 776 80720 785
rect 80392 736 80434 776
rect 80474 736 80516 776
rect 80556 736 80598 776
rect 80638 736 80680 776
rect 80352 727 80720 736
rect 84352 776 84720 785
rect 84392 736 84434 776
rect 84474 736 84516 776
rect 84556 736 84598 776
rect 84638 736 84680 776
rect 84352 727 84720 736
rect 88352 776 88720 785
rect 88392 736 88434 776
rect 88474 736 88516 776
rect 88556 736 88598 776
rect 88638 736 88680 776
rect 88352 727 88720 736
rect 92352 776 92720 785
rect 92392 736 92434 776
rect 92474 736 92516 776
rect 92556 736 92598 776
rect 92638 736 92680 776
rect 92352 727 92720 736
rect 96352 776 96720 785
rect 96392 736 96434 776
rect 96474 736 96516 776
rect 96556 736 96598 776
rect 96638 736 96680 776
rect 96352 727 96720 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 8352 38536 8392 38576
rect 8434 38536 8474 38576
rect 8516 38536 8556 38576
rect 8598 38536 8638 38576
rect 8680 38536 8720 38576
rect 12352 38536 12392 38576
rect 12434 38536 12474 38576
rect 12516 38536 12556 38576
rect 12598 38536 12638 38576
rect 12680 38536 12720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 20352 38536 20392 38576
rect 20434 38536 20474 38576
rect 20516 38536 20556 38576
rect 20598 38536 20638 38576
rect 20680 38536 20720 38576
rect 24352 38536 24392 38576
rect 24434 38536 24474 38576
rect 24516 38536 24556 38576
rect 24598 38536 24638 38576
rect 24680 38536 24720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 32352 38536 32392 38576
rect 32434 38536 32474 38576
rect 32516 38536 32556 38576
rect 32598 38536 32638 38576
rect 32680 38536 32720 38576
rect 36352 38536 36392 38576
rect 36434 38536 36474 38576
rect 36516 38536 36556 38576
rect 36598 38536 36638 38576
rect 36680 38536 36720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 44352 38536 44392 38576
rect 44434 38536 44474 38576
rect 44516 38536 44556 38576
rect 44598 38536 44638 38576
rect 44680 38536 44720 38576
rect 48352 38536 48392 38576
rect 48434 38536 48474 38576
rect 48516 38536 48556 38576
rect 48598 38536 48638 38576
rect 48680 38536 48720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 56352 38536 56392 38576
rect 56434 38536 56474 38576
rect 56516 38536 56556 38576
rect 56598 38536 56638 38576
rect 56680 38536 56720 38576
rect 60352 38536 60392 38576
rect 60434 38536 60474 38576
rect 60516 38536 60556 38576
rect 60598 38536 60638 38576
rect 60680 38536 60720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 68352 38536 68392 38576
rect 68434 38536 68474 38576
rect 68516 38536 68556 38576
rect 68598 38536 68638 38576
rect 68680 38536 68720 38576
rect 72352 38536 72392 38576
rect 72434 38536 72474 38576
rect 72516 38536 72556 38576
rect 72598 38536 72638 38576
rect 72680 38536 72720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 80352 38536 80392 38576
rect 80434 38536 80474 38576
rect 80516 38536 80556 38576
rect 80598 38536 80638 38576
rect 80680 38536 80720 38576
rect 84352 38536 84392 38576
rect 84434 38536 84474 38576
rect 84516 38536 84556 38576
rect 84598 38536 84638 38576
rect 84680 38536 84720 38576
rect 88352 38536 88392 38576
rect 88434 38536 88474 38576
rect 88516 38536 88556 38576
rect 88598 38536 88638 38576
rect 88680 38536 88720 38576
rect 92352 38536 92392 38576
rect 92434 38536 92474 38576
rect 92516 38536 92556 38576
rect 92598 38536 92638 38576
rect 92680 38536 92720 38576
rect 96352 38536 96392 38576
rect 96434 38536 96474 38576
rect 96516 38536 96556 38576
rect 96598 38536 96638 38576
rect 96680 38536 96720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 7112 37780 7152 37820
rect 7194 37780 7234 37820
rect 7276 37780 7316 37820
rect 7358 37780 7398 37820
rect 7440 37780 7480 37820
rect 11112 37780 11152 37820
rect 11194 37780 11234 37820
rect 11276 37780 11316 37820
rect 11358 37780 11398 37820
rect 11440 37780 11480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 19112 37780 19152 37820
rect 19194 37780 19234 37820
rect 19276 37780 19316 37820
rect 19358 37780 19398 37820
rect 19440 37780 19480 37820
rect 23112 37780 23152 37820
rect 23194 37780 23234 37820
rect 23276 37780 23316 37820
rect 23358 37780 23398 37820
rect 23440 37780 23480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 31112 37780 31152 37820
rect 31194 37780 31234 37820
rect 31276 37780 31316 37820
rect 31358 37780 31398 37820
rect 31440 37780 31480 37820
rect 35112 37780 35152 37820
rect 35194 37780 35234 37820
rect 35276 37780 35316 37820
rect 35358 37780 35398 37820
rect 35440 37780 35480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 43112 37780 43152 37820
rect 43194 37780 43234 37820
rect 43276 37780 43316 37820
rect 43358 37780 43398 37820
rect 43440 37780 43480 37820
rect 47112 37780 47152 37820
rect 47194 37780 47234 37820
rect 47276 37780 47316 37820
rect 47358 37780 47398 37820
rect 47440 37780 47480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 55112 37780 55152 37820
rect 55194 37780 55234 37820
rect 55276 37780 55316 37820
rect 55358 37780 55398 37820
rect 55440 37780 55480 37820
rect 59112 37780 59152 37820
rect 59194 37780 59234 37820
rect 59276 37780 59316 37820
rect 59358 37780 59398 37820
rect 59440 37780 59480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 67112 37780 67152 37820
rect 67194 37780 67234 37820
rect 67276 37780 67316 37820
rect 67358 37780 67398 37820
rect 67440 37780 67480 37820
rect 71112 37780 71152 37820
rect 71194 37780 71234 37820
rect 71276 37780 71316 37820
rect 71358 37780 71398 37820
rect 71440 37780 71480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 79112 37780 79152 37820
rect 79194 37780 79234 37820
rect 79276 37780 79316 37820
rect 79358 37780 79398 37820
rect 79440 37780 79480 37820
rect 83112 37780 83152 37820
rect 83194 37780 83234 37820
rect 83276 37780 83316 37820
rect 83358 37780 83398 37820
rect 83440 37780 83480 37820
rect 87112 37780 87152 37820
rect 87194 37780 87234 37820
rect 87276 37780 87316 37820
rect 87358 37780 87398 37820
rect 87440 37780 87480 37820
rect 91112 37780 91152 37820
rect 91194 37780 91234 37820
rect 91276 37780 91316 37820
rect 91358 37780 91398 37820
rect 91440 37780 91480 37820
rect 95112 37780 95152 37820
rect 95194 37780 95234 37820
rect 95276 37780 95316 37820
rect 95358 37780 95398 37820
rect 95440 37780 95480 37820
rect 99112 37780 99152 37820
rect 99194 37780 99234 37820
rect 99276 37780 99316 37820
rect 99358 37780 99398 37820
rect 99440 37780 99480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 8352 37024 8392 37064
rect 8434 37024 8474 37064
rect 8516 37024 8556 37064
rect 8598 37024 8638 37064
rect 8680 37024 8720 37064
rect 12352 37024 12392 37064
rect 12434 37024 12474 37064
rect 12516 37024 12556 37064
rect 12598 37024 12638 37064
rect 12680 37024 12720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 20352 37024 20392 37064
rect 20434 37024 20474 37064
rect 20516 37024 20556 37064
rect 20598 37024 20638 37064
rect 20680 37024 20720 37064
rect 24352 37024 24392 37064
rect 24434 37024 24474 37064
rect 24516 37024 24556 37064
rect 24598 37024 24638 37064
rect 24680 37024 24720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 32352 37024 32392 37064
rect 32434 37024 32474 37064
rect 32516 37024 32556 37064
rect 32598 37024 32638 37064
rect 32680 37024 32720 37064
rect 36352 37024 36392 37064
rect 36434 37024 36474 37064
rect 36516 37024 36556 37064
rect 36598 37024 36638 37064
rect 36680 37024 36720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 44352 37024 44392 37064
rect 44434 37024 44474 37064
rect 44516 37024 44556 37064
rect 44598 37024 44638 37064
rect 44680 37024 44720 37064
rect 48352 37024 48392 37064
rect 48434 37024 48474 37064
rect 48516 37024 48556 37064
rect 48598 37024 48638 37064
rect 48680 37024 48720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 56352 37024 56392 37064
rect 56434 37024 56474 37064
rect 56516 37024 56556 37064
rect 56598 37024 56638 37064
rect 56680 37024 56720 37064
rect 60352 37024 60392 37064
rect 60434 37024 60474 37064
rect 60516 37024 60556 37064
rect 60598 37024 60638 37064
rect 60680 37024 60720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 68352 37024 68392 37064
rect 68434 37024 68474 37064
rect 68516 37024 68556 37064
rect 68598 37024 68638 37064
rect 68680 37024 68720 37064
rect 72352 37024 72392 37064
rect 72434 37024 72474 37064
rect 72516 37024 72556 37064
rect 72598 37024 72638 37064
rect 72680 37024 72720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 80352 37024 80392 37064
rect 80434 37024 80474 37064
rect 80516 37024 80556 37064
rect 80598 37024 80638 37064
rect 80680 37024 80720 37064
rect 84352 37024 84392 37064
rect 84434 37024 84474 37064
rect 84516 37024 84556 37064
rect 84598 37024 84638 37064
rect 84680 37024 84720 37064
rect 88352 37024 88392 37064
rect 88434 37024 88474 37064
rect 88516 37024 88556 37064
rect 88598 37024 88638 37064
rect 88680 37024 88720 37064
rect 92352 37024 92392 37064
rect 92434 37024 92474 37064
rect 92516 37024 92556 37064
rect 92598 37024 92638 37064
rect 92680 37024 92720 37064
rect 96352 37024 96392 37064
rect 96434 37024 96474 37064
rect 96516 37024 96556 37064
rect 96598 37024 96638 37064
rect 96680 37024 96720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 7112 36268 7152 36308
rect 7194 36268 7234 36308
rect 7276 36268 7316 36308
rect 7358 36268 7398 36308
rect 7440 36268 7480 36308
rect 11112 36268 11152 36308
rect 11194 36268 11234 36308
rect 11276 36268 11316 36308
rect 11358 36268 11398 36308
rect 11440 36268 11480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 19112 36268 19152 36308
rect 19194 36268 19234 36308
rect 19276 36268 19316 36308
rect 19358 36268 19398 36308
rect 19440 36268 19480 36308
rect 23112 36268 23152 36308
rect 23194 36268 23234 36308
rect 23276 36268 23316 36308
rect 23358 36268 23398 36308
rect 23440 36268 23480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 31112 36268 31152 36308
rect 31194 36268 31234 36308
rect 31276 36268 31316 36308
rect 31358 36268 31398 36308
rect 31440 36268 31480 36308
rect 35112 36268 35152 36308
rect 35194 36268 35234 36308
rect 35276 36268 35316 36308
rect 35358 36268 35398 36308
rect 35440 36268 35480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 43112 36268 43152 36308
rect 43194 36268 43234 36308
rect 43276 36268 43316 36308
rect 43358 36268 43398 36308
rect 43440 36268 43480 36308
rect 47112 36268 47152 36308
rect 47194 36268 47234 36308
rect 47276 36268 47316 36308
rect 47358 36268 47398 36308
rect 47440 36268 47480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 55112 36268 55152 36308
rect 55194 36268 55234 36308
rect 55276 36268 55316 36308
rect 55358 36268 55398 36308
rect 55440 36268 55480 36308
rect 59112 36268 59152 36308
rect 59194 36268 59234 36308
rect 59276 36268 59316 36308
rect 59358 36268 59398 36308
rect 59440 36268 59480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 67112 36268 67152 36308
rect 67194 36268 67234 36308
rect 67276 36268 67316 36308
rect 67358 36268 67398 36308
rect 67440 36268 67480 36308
rect 71112 36268 71152 36308
rect 71194 36268 71234 36308
rect 71276 36268 71316 36308
rect 71358 36268 71398 36308
rect 71440 36268 71480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 79112 36268 79152 36308
rect 79194 36268 79234 36308
rect 79276 36268 79316 36308
rect 79358 36268 79398 36308
rect 79440 36268 79480 36308
rect 83112 36268 83152 36308
rect 83194 36268 83234 36308
rect 83276 36268 83316 36308
rect 83358 36268 83398 36308
rect 83440 36268 83480 36308
rect 87112 36268 87152 36308
rect 87194 36268 87234 36308
rect 87276 36268 87316 36308
rect 87358 36268 87398 36308
rect 87440 36268 87480 36308
rect 91112 36268 91152 36308
rect 91194 36268 91234 36308
rect 91276 36268 91316 36308
rect 91358 36268 91398 36308
rect 91440 36268 91480 36308
rect 95112 36268 95152 36308
rect 95194 36268 95234 36308
rect 95276 36268 95316 36308
rect 95358 36268 95398 36308
rect 95440 36268 95480 36308
rect 99112 36268 99152 36308
rect 99194 36268 99234 36308
rect 99276 36268 99316 36308
rect 99358 36268 99398 36308
rect 99440 36268 99480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 8352 35512 8392 35552
rect 8434 35512 8474 35552
rect 8516 35512 8556 35552
rect 8598 35512 8638 35552
rect 8680 35512 8720 35552
rect 12352 35512 12392 35552
rect 12434 35512 12474 35552
rect 12516 35512 12556 35552
rect 12598 35512 12638 35552
rect 12680 35512 12720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 20352 35512 20392 35552
rect 20434 35512 20474 35552
rect 20516 35512 20556 35552
rect 20598 35512 20638 35552
rect 20680 35512 20720 35552
rect 24352 35512 24392 35552
rect 24434 35512 24474 35552
rect 24516 35512 24556 35552
rect 24598 35512 24638 35552
rect 24680 35512 24720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 32352 35512 32392 35552
rect 32434 35512 32474 35552
rect 32516 35512 32556 35552
rect 32598 35512 32638 35552
rect 32680 35512 32720 35552
rect 36352 35512 36392 35552
rect 36434 35512 36474 35552
rect 36516 35512 36556 35552
rect 36598 35512 36638 35552
rect 36680 35512 36720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 44352 35512 44392 35552
rect 44434 35512 44474 35552
rect 44516 35512 44556 35552
rect 44598 35512 44638 35552
rect 44680 35512 44720 35552
rect 48352 35512 48392 35552
rect 48434 35512 48474 35552
rect 48516 35512 48556 35552
rect 48598 35512 48638 35552
rect 48680 35512 48720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 56352 35512 56392 35552
rect 56434 35512 56474 35552
rect 56516 35512 56556 35552
rect 56598 35512 56638 35552
rect 56680 35512 56720 35552
rect 60352 35512 60392 35552
rect 60434 35512 60474 35552
rect 60516 35512 60556 35552
rect 60598 35512 60638 35552
rect 60680 35512 60720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 68352 35512 68392 35552
rect 68434 35512 68474 35552
rect 68516 35512 68556 35552
rect 68598 35512 68638 35552
rect 68680 35512 68720 35552
rect 72352 35512 72392 35552
rect 72434 35512 72474 35552
rect 72516 35512 72556 35552
rect 72598 35512 72638 35552
rect 72680 35512 72720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 7112 34756 7152 34796
rect 7194 34756 7234 34796
rect 7276 34756 7316 34796
rect 7358 34756 7398 34796
rect 7440 34756 7480 34796
rect 11112 34756 11152 34796
rect 11194 34756 11234 34796
rect 11276 34756 11316 34796
rect 11358 34756 11398 34796
rect 11440 34756 11480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 19112 34756 19152 34796
rect 19194 34756 19234 34796
rect 19276 34756 19316 34796
rect 19358 34756 19398 34796
rect 19440 34756 19480 34796
rect 23112 34756 23152 34796
rect 23194 34756 23234 34796
rect 23276 34756 23316 34796
rect 23358 34756 23398 34796
rect 23440 34756 23480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 31112 34756 31152 34796
rect 31194 34756 31234 34796
rect 31276 34756 31316 34796
rect 31358 34756 31398 34796
rect 31440 34756 31480 34796
rect 35112 34756 35152 34796
rect 35194 34756 35234 34796
rect 35276 34756 35316 34796
rect 35358 34756 35398 34796
rect 35440 34756 35480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 43112 34756 43152 34796
rect 43194 34756 43234 34796
rect 43276 34756 43316 34796
rect 43358 34756 43398 34796
rect 43440 34756 43480 34796
rect 47112 34756 47152 34796
rect 47194 34756 47234 34796
rect 47276 34756 47316 34796
rect 47358 34756 47398 34796
rect 47440 34756 47480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 55112 34756 55152 34796
rect 55194 34756 55234 34796
rect 55276 34756 55316 34796
rect 55358 34756 55398 34796
rect 55440 34756 55480 34796
rect 59112 34756 59152 34796
rect 59194 34756 59234 34796
rect 59276 34756 59316 34796
rect 59358 34756 59398 34796
rect 59440 34756 59480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 67112 34756 67152 34796
rect 67194 34756 67234 34796
rect 67276 34756 67316 34796
rect 67358 34756 67398 34796
rect 67440 34756 67480 34796
rect 71112 34756 71152 34796
rect 71194 34756 71234 34796
rect 71276 34756 71316 34796
rect 71358 34756 71398 34796
rect 71440 34756 71480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 8352 34000 8392 34040
rect 8434 34000 8474 34040
rect 8516 34000 8556 34040
rect 8598 34000 8638 34040
rect 8680 34000 8720 34040
rect 12352 34000 12392 34040
rect 12434 34000 12474 34040
rect 12516 34000 12556 34040
rect 12598 34000 12638 34040
rect 12680 34000 12720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 20352 34000 20392 34040
rect 20434 34000 20474 34040
rect 20516 34000 20556 34040
rect 20598 34000 20638 34040
rect 20680 34000 20720 34040
rect 24352 34000 24392 34040
rect 24434 34000 24474 34040
rect 24516 34000 24556 34040
rect 24598 34000 24638 34040
rect 24680 34000 24720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 32352 34000 32392 34040
rect 32434 34000 32474 34040
rect 32516 34000 32556 34040
rect 32598 34000 32638 34040
rect 32680 34000 32720 34040
rect 36352 34000 36392 34040
rect 36434 34000 36474 34040
rect 36516 34000 36556 34040
rect 36598 34000 36638 34040
rect 36680 34000 36720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 44352 34000 44392 34040
rect 44434 34000 44474 34040
rect 44516 34000 44556 34040
rect 44598 34000 44638 34040
rect 44680 34000 44720 34040
rect 48352 34000 48392 34040
rect 48434 34000 48474 34040
rect 48516 34000 48556 34040
rect 48598 34000 48638 34040
rect 48680 34000 48720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 56352 34000 56392 34040
rect 56434 34000 56474 34040
rect 56516 34000 56556 34040
rect 56598 34000 56638 34040
rect 56680 34000 56720 34040
rect 60352 34000 60392 34040
rect 60434 34000 60474 34040
rect 60516 34000 60556 34040
rect 60598 34000 60638 34040
rect 60680 34000 60720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 68352 34000 68392 34040
rect 68434 34000 68474 34040
rect 68516 34000 68556 34040
rect 68598 34000 68638 34040
rect 68680 34000 68720 34040
rect 72352 34000 72392 34040
rect 72434 34000 72474 34040
rect 72516 34000 72556 34040
rect 72598 34000 72638 34040
rect 72680 34000 72720 34040
rect 76352 34000 76392 34040
rect 76434 34000 76474 34040
rect 76516 34000 76556 34040
rect 76598 34000 76638 34040
rect 76680 34000 76720 34040
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 7112 33244 7152 33284
rect 7194 33244 7234 33284
rect 7276 33244 7316 33284
rect 7358 33244 7398 33284
rect 7440 33244 7480 33284
rect 11112 33244 11152 33284
rect 11194 33244 11234 33284
rect 11276 33244 11316 33284
rect 11358 33244 11398 33284
rect 11440 33244 11480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 19112 33244 19152 33284
rect 19194 33244 19234 33284
rect 19276 33244 19316 33284
rect 19358 33244 19398 33284
rect 19440 33244 19480 33284
rect 23112 33244 23152 33284
rect 23194 33244 23234 33284
rect 23276 33244 23316 33284
rect 23358 33244 23398 33284
rect 23440 33244 23480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 31112 33244 31152 33284
rect 31194 33244 31234 33284
rect 31276 33244 31316 33284
rect 31358 33244 31398 33284
rect 31440 33244 31480 33284
rect 35112 33244 35152 33284
rect 35194 33244 35234 33284
rect 35276 33244 35316 33284
rect 35358 33244 35398 33284
rect 35440 33244 35480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 43112 33244 43152 33284
rect 43194 33244 43234 33284
rect 43276 33244 43316 33284
rect 43358 33244 43398 33284
rect 43440 33244 43480 33284
rect 47112 33244 47152 33284
rect 47194 33244 47234 33284
rect 47276 33244 47316 33284
rect 47358 33244 47398 33284
rect 47440 33244 47480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 55112 33244 55152 33284
rect 55194 33244 55234 33284
rect 55276 33244 55316 33284
rect 55358 33244 55398 33284
rect 55440 33244 55480 33284
rect 59112 33244 59152 33284
rect 59194 33244 59234 33284
rect 59276 33244 59316 33284
rect 59358 33244 59398 33284
rect 59440 33244 59480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 67112 33244 67152 33284
rect 67194 33244 67234 33284
rect 67276 33244 67316 33284
rect 67358 33244 67398 33284
rect 67440 33244 67480 33284
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 8352 32488 8392 32528
rect 8434 32488 8474 32528
rect 8516 32488 8556 32528
rect 8598 32488 8638 32528
rect 8680 32488 8720 32528
rect 12352 32488 12392 32528
rect 12434 32488 12474 32528
rect 12516 32488 12556 32528
rect 12598 32488 12638 32528
rect 12680 32488 12720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 20352 32488 20392 32528
rect 20434 32488 20474 32528
rect 20516 32488 20556 32528
rect 20598 32488 20638 32528
rect 20680 32488 20720 32528
rect 24352 32488 24392 32528
rect 24434 32488 24474 32528
rect 24516 32488 24556 32528
rect 24598 32488 24638 32528
rect 24680 32488 24720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 32352 32488 32392 32528
rect 32434 32488 32474 32528
rect 32516 32488 32556 32528
rect 32598 32488 32638 32528
rect 32680 32488 32720 32528
rect 36352 32488 36392 32528
rect 36434 32488 36474 32528
rect 36516 32488 36556 32528
rect 36598 32488 36638 32528
rect 36680 32488 36720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 44352 32488 44392 32528
rect 44434 32488 44474 32528
rect 44516 32488 44556 32528
rect 44598 32488 44638 32528
rect 44680 32488 44720 32528
rect 48352 32488 48392 32528
rect 48434 32488 48474 32528
rect 48516 32488 48556 32528
rect 48598 32488 48638 32528
rect 48680 32488 48720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 56352 32488 56392 32528
rect 56434 32488 56474 32528
rect 56516 32488 56556 32528
rect 56598 32488 56638 32528
rect 56680 32488 56720 32528
rect 60352 32488 60392 32528
rect 60434 32488 60474 32528
rect 60516 32488 60556 32528
rect 60598 32488 60638 32528
rect 60680 32488 60720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 68352 32488 68392 32528
rect 68434 32488 68474 32528
rect 68516 32488 68556 32528
rect 68598 32488 68638 32528
rect 68680 32488 68720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 7112 31732 7152 31772
rect 7194 31732 7234 31772
rect 7276 31732 7316 31772
rect 7358 31732 7398 31772
rect 7440 31732 7480 31772
rect 11112 31732 11152 31772
rect 11194 31732 11234 31772
rect 11276 31732 11316 31772
rect 11358 31732 11398 31772
rect 11440 31732 11480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 19112 31732 19152 31772
rect 19194 31732 19234 31772
rect 19276 31732 19316 31772
rect 19358 31732 19398 31772
rect 19440 31732 19480 31772
rect 23112 31732 23152 31772
rect 23194 31732 23234 31772
rect 23276 31732 23316 31772
rect 23358 31732 23398 31772
rect 23440 31732 23480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 31112 31732 31152 31772
rect 31194 31732 31234 31772
rect 31276 31732 31316 31772
rect 31358 31732 31398 31772
rect 31440 31732 31480 31772
rect 35112 31732 35152 31772
rect 35194 31732 35234 31772
rect 35276 31732 35316 31772
rect 35358 31732 35398 31772
rect 35440 31732 35480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 43112 31732 43152 31772
rect 43194 31732 43234 31772
rect 43276 31732 43316 31772
rect 43358 31732 43398 31772
rect 43440 31732 43480 31772
rect 47112 31732 47152 31772
rect 47194 31732 47234 31772
rect 47276 31732 47316 31772
rect 47358 31732 47398 31772
rect 47440 31732 47480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 55112 31732 55152 31772
rect 55194 31732 55234 31772
rect 55276 31732 55316 31772
rect 55358 31732 55398 31772
rect 55440 31732 55480 31772
rect 59112 31732 59152 31772
rect 59194 31732 59234 31772
rect 59276 31732 59316 31772
rect 59358 31732 59398 31772
rect 59440 31732 59480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 67112 31732 67152 31772
rect 67194 31732 67234 31772
rect 67276 31732 67316 31772
rect 67358 31732 67398 31772
rect 67440 31732 67480 31772
rect 80352 35512 80392 35552
rect 80434 35512 80474 35552
rect 80516 35512 80556 35552
rect 80598 35512 80638 35552
rect 80680 35512 80720 35552
rect 84352 35512 84392 35552
rect 84434 35512 84474 35552
rect 84516 35512 84556 35552
rect 84598 35512 84638 35552
rect 84680 35512 84720 35552
rect 79112 34756 79152 34796
rect 79194 34756 79234 34796
rect 79276 34756 79316 34796
rect 79358 34756 79398 34796
rect 79440 34756 79480 34796
rect 83112 34756 83152 34796
rect 83194 34756 83234 34796
rect 83276 34756 83316 34796
rect 83358 34756 83398 34796
rect 83440 34756 83480 34796
rect 80352 34000 80392 34040
rect 80434 34000 80474 34040
rect 80516 34000 80556 34040
rect 80598 34000 80638 34040
rect 80680 34000 80720 34040
rect 84352 34000 84392 34040
rect 84434 34000 84474 34040
rect 84516 34000 84556 34040
rect 84598 34000 84638 34040
rect 84680 34000 84720 34040
rect 88352 35512 88392 35552
rect 88434 35512 88474 35552
rect 88516 35512 88556 35552
rect 88598 35512 88638 35552
rect 88680 35512 88720 35552
rect 86668 34924 86708 34964
rect 87112 34756 87152 34796
rect 87194 34756 87234 34796
rect 87276 34756 87316 34796
rect 87358 34756 87398 34796
rect 87440 34756 87480 34796
rect 88352 34000 88392 34040
rect 88434 34000 88474 34040
rect 88516 34000 88556 34040
rect 88598 34000 88638 34040
rect 88680 34000 88720 34040
rect 91112 34756 91152 34796
rect 91194 34756 91234 34796
rect 91276 34756 91316 34796
rect 91358 34756 91398 34796
rect 91440 34756 91480 34796
rect 92352 35512 92392 35552
rect 92434 35512 92474 35552
rect 92516 35512 92556 35552
rect 92598 35512 92638 35552
rect 92680 35512 92720 35552
rect 96352 35512 96392 35552
rect 96434 35512 96474 35552
rect 96516 35512 96556 35552
rect 96598 35512 96638 35552
rect 96680 35512 96720 35552
rect 95112 34756 95152 34796
rect 95194 34756 95234 34796
rect 95276 34756 95316 34796
rect 95358 34756 95398 34796
rect 95440 34756 95480 34796
rect 99112 34756 99152 34796
rect 99194 34756 99234 34796
rect 99276 34756 99316 34796
rect 99358 34756 99398 34796
rect 99440 34756 99480 34796
rect 92352 34000 92392 34040
rect 92434 34000 92474 34040
rect 92516 34000 92556 34040
rect 92598 34000 92638 34040
rect 92680 34000 92720 34040
rect 96352 34000 96392 34040
rect 96434 34000 96474 34040
rect 96516 34000 96556 34040
rect 96598 34000 96638 34040
rect 96680 34000 96720 34040
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 8352 30976 8392 31016
rect 8434 30976 8474 31016
rect 8516 30976 8556 31016
rect 8598 30976 8638 31016
rect 8680 30976 8720 31016
rect 12352 30976 12392 31016
rect 12434 30976 12474 31016
rect 12516 30976 12556 31016
rect 12598 30976 12638 31016
rect 12680 30976 12720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 20352 30976 20392 31016
rect 20434 30976 20474 31016
rect 20516 30976 20556 31016
rect 20598 30976 20638 31016
rect 20680 30976 20720 31016
rect 24352 30976 24392 31016
rect 24434 30976 24474 31016
rect 24516 30976 24556 31016
rect 24598 30976 24638 31016
rect 24680 30976 24720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 32352 30976 32392 31016
rect 32434 30976 32474 31016
rect 32516 30976 32556 31016
rect 32598 30976 32638 31016
rect 32680 30976 32720 31016
rect 36352 30976 36392 31016
rect 36434 30976 36474 31016
rect 36516 30976 36556 31016
rect 36598 30976 36638 31016
rect 36680 30976 36720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 44352 30976 44392 31016
rect 44434 30976 44474 31016
rect 44516 30976 44556 31016
rect 44598 30976 44638 31016
rect 44680 30976 44720 31016
rect 48352 30976 48392 31016
rect 48434 30976 48474 31016
rect 48516 30976 48556 31016
rect 48598 30976 48638 31016
rect 48680 30976 48720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 56352 30976 56392 31016
rect 56434 30976 56474 31016
rect 56516 30976 56556 31016
rect 56598 30976 56638 31016
rect 56680 30976 56720 31016
rect 60352 30976 60392 31016
rect 60434 30976 60474 31016
rect 60516 30976 60556 31016
rect 60598 30976 60638 31016
rect 60680 30976 60720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 68352 30976 68392 31016
rect 68434 30976 68474 31016
rect 68516 30976 68556 31016
rect 68598 30976 68638 31016
rect 68680 30976 68720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 7112 30220 7152 30260
rect 7194 30220 7234 30260
rect 7276 30220 7316 30260
rect 7358 30220 7398 30260
rect 7440 30220 7480 30260
rect 11112 30220 11152 30260
rect 11194 30220 11234 30260
rect 11276 30220 11316 30260
rect 11358 30220 11398 30260
rect 11440 30220 11480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 19112 30220 19152 30260
rect 19194 30220 19234 30260
rect 19276 30220 19316 30260
rect 19358 30220 19398 30260
rect 19440 30220 19480 30260
rect 23112 30220 23152 30260
rect 23194 30220 23234 30260
rect 23276 30220 23316 30260
rect 23358 30220 23398 30260
rect 23440 30220 23480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 31112 30220 31152 30260
rect 31194 30220 31234 30260
rect 31276 30220 31316 30260
rect 31358 30220 31398 30260
rect 31440 30220 31480 30260
rect 35112 30220 35152 30260
rect 35194 30220 35234 30260
rect 35276 30220 35316 30260
rect 35358 30220 35398 30260
rect 35440 30220 35480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 43112 30220 43152 30260
rect 43194 30220 43234 30260
rect 43276 30220 43316 30260
rect 43358 30220 43398 30260
rect 43440 30220 43480 30260
rect 47112 30220 47152 30260
rect 47194 30220 47234 30260
rect 47276 30220 47316 30260
rect 47358 30220 47398 30260
rect 47440 30220 47480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 55112 30220 55152 30260
rect 55194 30220 55234 30260
rect 55276 30220 55316 30260
rect 55358 30220 55398 30260
rect 55440 30220 55480 30260
rect 59112 30220 59152 30260
rect 59194 30220 59234 30260
rect 59276 30220 59316 30260
rect 59358 30220 59398 30260
rect 59440 30220 59480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 67112 30220 67152 30260
rect 67194 30220 67234 30260
rect 67276 30220 67316 30260
rect 67358 30220 67398 30260
rect 67440 30220 67480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 8352 29464 8392 29504
rect 8434 29464 8474 29504
rect 8516 29464 8556 29504
rect 8598 29464 8638 29504
rect 8680 29464 8720 29504
rect 12352 29464 12392 29504
rect 12434 29464 12474 29504
rect 12516 29464 12556 29504
rect 12598 29464 12638 29504
rect 12680 29464 12720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 20352 29464 20392 29504
rect 20434 29464 20474 29504
rect 20516 29464 20556 29504
rect 20598 29464 20638 29504
rect 20680 29464 20720 29504
rect 24352 29464 24392 29504
rect 24434 29464 24474 29504
rect 24516 29464 24556 29504
rect 24598 29464 24638 29504
rect 24680 29464 24720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 32352 29464 32392 29504
rect 32434 29464 32474 29504
rect 32516 29464 32556 29504
rect 32598 29464 32638 29504
rect 32680 29464 32720 29504
rect 36352 29464 36392 29504
rect 36434 29464 36474 29504
rect 36516 29464 36556 29504
rect 36598 29464 36638 29504
rect 36680 29464 36720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 44352 29464 44392 29504
rect 44434 29464 44474 29504
rect 44516 29464 44556 29504
rect 44598 29464 44638 29504
rect 44680 29464 44720 29504
rect 48352 29464 48392 29504
rect 48434 29464 48474 29504
rect 48516 29464 48556 29504
rect 48598 29464 48638 29504
rect 48680 29464 48720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 56352 29464 56392 29504
rect 56434 29464 56474 29504
rect 56516 29464 56556 29504
rect 56598 29464 56638 29504
rect 56680 29464 56720 29504
rect 60352 29464 60392 29504
rect 60434 29464 60474 29504
rect 60516 29464 60556 29504
rect 60598 29464 60638 29504
rect 60680 29464 60720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 68352 29464 68392 29504
rect 68434 29464 68474 29504
rect 68516 29464 68556 29504
rect 68598 29464 68638 29504
rect 68680 29464 68720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 7112 28708 7152 28748
rect 7194 28708 7234 28748
rect 7276 28708 7316 28748
rect 7358 28708 7398 28748
rect 7440 28708 7480 28748
rect 11112 28708 11152 28748
rect 11194 28708 11234 28748
rect 11276 28708 11316 28748
rect 11358 28708 11398 28748
rect 11440 28708 11480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 19112 28708 19152 28748
rect 19194 28708 19234 28748
rect 19276 28708 19316 28748
rect 19358 28708 19398 28748
rect 19440 28708 19480 28748
rect 23112 28708 23152 28748
rect 23194 28708 23234 28748
rect 23276 28708 23316 28748
rect 23358 28708 23398 28748
rect 23440 28708 23480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 31112 28708 31152 28748
rect 31194 28708 31234 28748
rect 31276 28708 31316 28748
rect 31358 28708 31398 28748
rect 31440 28708 31480 28748
rect 35112 28708 35152 28748
rect 35194 28708 35234 28748
rect 35276 28708 35316 28748
rect 35358 28708 35398 28748
rect 35440 28708 35480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 43112 28708 43152 28748
rect 43194 28708 43234 28748
rect 43276 28708 43316 28748
rect 43358 28708 43398 28748
rect 43440 28708 43480 28748
rect 47112 28708 47152 28748
rect 47194 28708 47234 28748
rect 47276 28708 47316 28748
rect 47358 28708 47398 28748
rect 47440 28708 47480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 55112 28708 55152 28748
rect 55194 28708 55234 28748
rect 55276 28708 55316 28748
rect 55358 28708 55398 28748
rect 55440 28708 55480 28748
rect 59112 28708 59152 28748
rect 59194 28708 59234 28748
rect 59276 28708 59316 28748
rect 59358 28708 59398 28748
rect 59440 28708 59480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 67112 28708 67152 28748
rect 67194 28708 67234 28748
rect 67276 28708 67316 28748
rect 67358 28708 67398 28748
rect 67440 28708 67480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 8352 27952 8392 27992
rect 8434 27952 8474 27992
rect 8516 27952 8556 27992
rect 8598 27952 8638 27992
rect 8680 27952 8720 27992
rect 12352 27952 12392 27992
rect 12434 27952 12474 27992
rect 12516 27952 12556 27992
rect 12598 27952 12638 27992
rect 12680 27952 12720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 20352 27952 20392 27992
rect 20434 27952 20474 27992
rect 20516 27952 20556 27992
rect 20598 27952 20638 27992
rect 20680 27952 20720 27992
rect 24352 27952 24392 27992
rect 24434 27952 24474 27992
rect 24516 27952 24556 27992
rect 24598 27952 24638 27992
rect 24680 27952 24720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 32352 27952 32392 27992
rect 32434 27952 32474 27992
rect 32516 27952 32556 27992
rect 32598 27952 32638 27992
rect 32680 27952 32720 27992
rect 36352 27952 36392 27992
rect 36434 27952 36474 27992
rect 36516 27952 36556 27992
rect 36598 27952 36638 27992
rect 36680 27952 36720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 44352 27952 44392 27992
rect 44434 27952 44474 27992
rect 44516 27952 44556 27992
rect 44598 27952 44638 27992
rect 44680 27952 44720 27992
rect 48352 27952 48392 27992
rect 48434 27952 48474 27992
rect 48516 27952 48556 27992
rect 48598 27952 48638 27992
rect 48680 27952 48720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 56352 27952 56392 27992
rect 56434 27952 56474 27992
rect 56516 27952 56556 27992
rect 56598 27952 56638 27992
rect 56680 27952 56720 27992
rect 60352 27952 60392 27992
rect 60434 27952 60474 27992
rect 60516 27952 60556 27992
rect 60598 27952 60638 27992
rect 60680 27952 60720 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 68352 27952 68392 27992
rect 68434 27952 68474 27992
rect 68516 27952 68556 27992
rect 68598 27952 68638 27992
rect 68680 27952 68720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 7112 27196 7152 27236
rect 7194 27196 7234 27236
rect 7276 27196 7316 27236
rect 7358 27196 7398 27236
rect 7440 27196 7480 27236
rect 11112 27196 11152 27236
rect 11194 27196 11234 27236
rect 11276 27196 11316 27236
rect 11358 27196 11398 27236
rect 11440 27196 11480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 19112 27196 19152 27236
rect 19194 27196 19234 27236
rect 19276 27196 19316 27236
rect 19358 27196 19398 27236
rect 19440 27196 19480 27236
rect 23112 27196 23152 27236
rect 23194 27196 23234 27236
rect 23276 27196 23316 27236
rect 23358 27196 23398 27236
rect 23440 27196 23480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 31112 27196 31152 27236
rect 31194 27196 31234 27236
rect 31276 27196 31316 27236
rect 31358 27196 31398 27236
rect 31440 27196 31480 27236
rect 35112 27196 35152 27236
rect 35194 27196 35234 27236
rect 35276 27196 35316 27236
rect 35358 27196 35398 27236
rect 35440 27196 35480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 43112 27196 43152 27236
rect 43194 27196 43234 27236
rect 43276 27196 43316 27236
rect 43358 27196 43398 27236
rect 43440 27196 43480 27236
rect 47112 27196 47152 27236
rect 47194 27196 47234 27236
rect 47276 27196 47316 27236
rect 47358 27196 47398 27236
rect 47440 27196 47480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 55112 27196 55152 27236
rect 55194 27196 55234 27236
rect 55276 27196 55316 27236
rect 55358 27196 55398 27236
rect 55440 27196 55480 27236
rect 59112 27196 59152 27236
rect 59194 27196 59234 27236
rect 59276 27196 59316 27236
rect 59358 27196 59398 27236
rect 59440 27196 59480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 67112 27196 67152 27236
rect 67194 27196 67234 27236
rect 67276 27196 67316 27236
rect 67358 27196 67398 27236
rect 67440 27196 67480 27236
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 8352 26440 8392 26480
rect 8434 26440 8474 26480
rect 8516 26440 8556 26480
rect 8598 26440 8638 26480
rect 8680 26440 8720 26480
rect 12352 26440 12392 26480
rect 12434 26440 12474 26480
rect 12516 26440 12556 26480
rect 12598 26440 12638 26480
rect 12680 26440 12720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 20352 26440 20392 26480
rect 20434 26440 20474 26480
rect 20516 26440 20556 26480
rect 20598 26440 20638 26480
rect 20680 26440 20720 26480
rect 24352 26440 24392 26480
rect 24434 26440 24474 26480
rect 24516 26440 24556 26480
rect 24598 26440 24638 26480
rect 24680 26440 24720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 32352 26440 32392 26480
rect 32434 26440 32474 26480
rect 32516 26440 32556 26480
rect 32598 26440 32638 26480
rect 32680 26440 32720 26480
rect 36352 26440 36392 26480
rect 36434 26440 36474 26480
rect 36516 26440 36556 26480
rect 36598 26440 36638 26480
rect 36680 26440 36720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 44352 26440 44392 26480
rect 44434 26440 44474 26480
rect 44516 26440 44556 26480
rect 44598 26440 44638 26480
rect 44680 26440 44720 26480
rect 48352 26440 48392 26480
rect 48434 26440 48474 26480
rect 48516 26440 48556 26480
rect 48598 26440 48638 26480
rect 48680 26440 48720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 56352 26440 56392 26480
rect 56434 26440 56474 26480
rect 56516 26440 56556 26480
rect 56598 26440 56638 26480
rect 56680 26440 56720 26480
rect 60352 26440 60392 26480
rect 60434 26440 60474 26480
rect 60516 26440 60556 26480
rect 60598 26440 60638 26480
rect 60680 26440 60720 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 68352 26440 68392 26480
rect 68434 26440 68474 26480
rect 68516 26440 68556 26480
rect 68598 26440 68638 26480
rect 68680 26440 68720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 7112 25684 7152 25724
rect 7194 25684 7234 25724
rect 7276 25684 7316 25724
rect 7358 25684 7398 25724
rect 7440 25684 7480 25724
rect 11112 25684 11152 25724
rect 11194 25684 11234 25724
rect 11276 25684 11316 25724
rect 11358 25684 11398 25724
rect 11440 25684 11480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 19112 25684 19152 25724
rect 19194 25684 19234 25724
rect 19276 25684 19316 25724
rect 19358 25684 19398 25724
rect 19440 25684 19480 25724
rect 23112 25684 23152 25724
rect 23194 25684 23234 25724
rect 23276 25684 23316 25724
rect 23358 25684 23398 25724
rect 23440 25684 23480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 31112 25684 31152 25724
rect 31194 25684 31234 25724
rect 31276 25684 31316 25724
rect 31358 25684 31398 25724
rect 31440 25684 31480 25724
rect 35112 25684 35152 25724
rect 35194 25684 35234 25724
rect 35276 25684 35316 25724
rect 35358 25684 35398 25724
rect 35440 25684 35480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 43112 25684 43152 25724
rect 43194 25684 43234 25724
rect 43276 25684 43316 25724
rect 43358 25684 43398 25724
rect 43440 25684 43480 25724
rect 47112 25684 47152 25724
rect 47194 25684 47234 25724
rect 47276 25684 47316 25724
rect 47358 25684 47398 25724
rect 47440 25684 47480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 55112 25684 55152 25724
rect 55194 25684 55234 25724
rect 55276 25684 55316 25724
rect 55358 25684 55398 25724
rect 55440 25684 55480 25724
rect 59112 25684 59152 25724
rect 59194 25684 59234 25724
rect 59276 25684 59316 25724
rect 59358 25684 59398 25724
rect 59440 25684 59480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 67112 25684 67152 25724
rect 67194 25684 67234 25724
rect 67276 25684 67316 25724
rect 67358 25684 67398 25724
rect 67440 25684 67480 25724
rect 71788 25600 71828 25640
rect 72940 25600 72980 25640
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 8352 24928 8392 24968
rect 8434 24928 8474 24968
rect 8516 24928 8556 24968
rect 8598 24928 8638 24968
rect 8680 24928 8720 24968
rect 12352 24928 12392 24968
rect 12434 24928 12474 24968
rect 12516 24928 12556 24968
rect 12598 24928 12638 24968
rect 12680 24928 12720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 20352 24928 20392 24968
rect 20434 24928 20474 24968
rect 20516 24928 20556 24968
rect 20598 24928 20638 24968
rect 20680 24928 20720 24968
rect 24352 24928 24392 24968
rect 24434 24928 24474 24968
rect 24516 24928 24556 24968
rect 24598 24928 24638 24968
rect 24680 24928 24720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 32352 24928 32392 24968
rect 32434 24928 32474 24968
rect 32516 24928 32556 24968
rect 32598 24928 32638 24968
rect 32680 24928 32720 24968
rect 36352 24928 36392 24968
rect 36434 24928 36474 24968
rect 36516 24928 36556 24968
rect 36598 24928 36638 24968
rect 36680 24928 36720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 44352 24928 44392 24968
rect 44434 24928 44474 24968
rect 44516 24928 44556 24968
rect 44598 24928 44638 24968
rect 44680 24928 44720 24968
rect 48352 24928 48392 24968
rect 48434 24928 48474 24968
rect 48516 24928 48556 24968
rect 48598 24928 48638 24968
rect 48680 24928 48720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 56352 24928 56392 24968
rect 56434 24928 56474 24968
rect 56516 24928 56556 24968
rect 56598 24928 56638 24968
rect 56680 24928 56720 24968
rect 60352 24928 60392 24968
rect 60434 24928 60474 24968
rect 60516 24928 60556 24968
rect 60598 24928 60638 24968
rect 60680 24928 60720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 68352 24928 68392 24968
rect 68434 24928 68474 24968
rect 68516 24928 68556 24968
rect 68598 24928 68638 24968
rect 68680 24928 68720 24968
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 7112 24172 7152 24212
rect 7194 24172 7234 24212
rect 7276 24172 7316 24212
rect 7358 24172 7398 24212
rect 7440 24172 7480 24212
rect 11112 24172 11152 24212
rect 11194 24172 11234 24212
rect 11276 24172 11316 24212
rect 11358 24172 11398 24212
rect 11440 24172 11480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 19112 24172 19152 24212
rect 19194 24172 19234 24212
rect 19276 24172 19316 24212
rect 19358 24172 19398 24212
rect 19440 24172 19480 24212
rect 23112 24172 23152 24212
rect 23194 24172 23234 24212
rect 23276 24172 23316 24212
rect 23358 24172 23398 24212
rect 23440 24172 23480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 31112 24172 31152 24212
rect 31194 24172 31234 24212
rect 31276 24172 31316 24212
rect 31358 24172 31398 24212
rect 31440 24172 31480 24212
rect 35112 24172 35152 24212
rect 35194 24172 35234 24212
rect 35276 24172 35316 24212
rect 35358 24172 35398 24212
rect 35440 24172 35480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 43112 24172 43152 24212
rect 43194 24172 43234 24212
rect 43276 24172 43316 24212
rect 43358 24172 43398 24212
rect 43440 24172 43480 24212
rect 47112 24172 47152 24212
rect 47194 24172 47234 24212
rect 47276 24172 47316 24212
rect 47358 24172 47398 24212
rect 47440 24172 47480 24212
rect 51112 24172 51152 24212
rect 51194 24172 51234 24212
rect 51276 24172 51316 24212
rect 51358 24172 51398 24212
rect 51440 24172 51480 24212
rect 55112 24172 55152 24212
rect 55194 24172 55234 24212
rect 55276 24172 55316 24212
rect 55358 24172 55398 24212
rect 55440 24172 55480 24212
rect 59112 24172 59152 24212
rect 59194 24172 59234 24212
rect 59276 24172 59316 24212
rect 59358 24172 59398 24212
rect 59440 24172 59480 24212
rect 63112 24172 63152 24212
rect 63194 24172 63234 24212
rect 63276 24172 63316 24212
rect 63358 24172 63398 24212
rect 63440 24172 63480 24212
rect 67112 24172 67152 24212
rect 67194 24172 67234 24212
rect 67276 24172 67316 24212
rect 67358 24172 67398 24212
rect 67440 24172 67480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 8352 23416 8392 23456
rect 8434 23416 8474 23456
rect 8516 23416 8556 23456
rect 8598 23416 8638 23456
rect 8680 23416 8720 23456
rect 12352 23416 12392 23456
rect 12434 23416 12474 23456
rect 12516 23416 12556 23456
rect 12598 23416 12638 23456
rect 12680 23416 12720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 20352 23416 20392 23456
rect 20434 23416 20474 23456
rect 20516 23416 20556 23456
rect 20598 23416 20638 23456
rect 20680 23416 20720 23456
rect 24352 23416 24392 23456
rect 24434 23416 24474 23456
rect 24516 23416 24556 23456
rect 24598 23416 24638 23456
rect 24680 23416 24720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 32352 23416 32392 23456
rect 32434 23416 32474 23456
rect 32516 23416 32556 23456
rect 32598 23416 32638 23456
rect 32680 23416 32720 23456
rect 36352 23416 36392 23456
rect 36434 23416 36474 23456
rect 36516 23416 36556 23456
rect 36598 23416 36638 23456
rect 36680 23416 36720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 44352 23416 44392 23456
rect 44434 23416 44474 23456
rect 44516 23416 44556 23456
rect 44598 23416 44638 23456
rect 44680 23416 44720 23456
rect 48352 23416 48392 23456
rect 48434 23416 48474 23456
rect 48516 23416 48556 23456
rect 48598 23416 48638 23456
rect 48680 23416 48720 23456
rect 52352 23416 52392 23456
rect 52434 23416 52474 23456
rect 52516 23416 52556 23456
rect 52598 23416 52638 23456
rect 52680 23416 52720 23456
rect 56352 23416 56392 23456
rect 56434 23416 56474 23456
rect 56516 23416 56556 23456
rect 56598 23416 56638 23456
rect 56680 23416 56720 23456
rect 60352 23416 60392 23456
rect 60434 23416 60474 23456
rect 60516 23416 60556 23456
rect 60598 23416 60638 23456
rect 60680 23416 60720 23456
rect 64352 23416 64392 23456
rect 64434 23416 64474 23456
rect 64516 23416 64556 23456
rect 64598 23416 64638 23456
rect 64680 23416 64720 23456
rect 68352 23416 68392 23456
rect 68434 23416 68474 23456
rect 68516 23416 68556 23456
rect 68598 23416 68638 23456
rect 68680 23416 68720 23456
rect 72352 23416 72392 23456
rect 72434 23416 72474 23456
rect 72516 23416 72556 23456
rect 72598 23416 72638 23456
rect 72680 23416 72720 23456
rect 76352 23416 76392 23456
rect 76434 23416 76474 23456
rect 76516 23416 76556 23456
rect 76598 23416 76638 23456
rect 76680 23416 76720 23456
rect 80352 23416 80392 23456
rect 80434 23416 80474 23456
rect 80516 23416 80556 23456
rect 80598 23416 80638 23456
rect 80680 23416 80720 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 7112 22660 7152 22700
rect 7194 22660 7234 22700
rect 7276 22660 7316 22700
rect 7358 22660 7398 22700
rect 7440 22660 7480 22700
rect 11112 22660 11152 22700
rect 11194 22660 11234 22700
rect 11276 22660 11316 22700
rect 11358 22660 11398 22700
rect 11440 22660 11480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 19112 22660 19152 22700
rect 19194 22660 19234 22700
rect 19276 22660 19316 22700
rect 19358 22660 19398 22700
rect 19440 22660 19480 22700
rect 23112 22660 23152 22700
rect 23194 22660 23234 22700
rect 23276 22660 23316 22700
rect 23358 22660 23398 22700
rect 23440 22660 23480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 31112 22660 31152 22700
rect 31194 22660 31234 22700
rect 31276 22660 31316 22700
rect 31358 22660 31398 22700
rect 31440 22660 31480 22700
rect 35112 22660 35152 22700
rect 35194 22660 35234 22700
rect 35276 22660 35316 22700
rect 35358 22660 35398 22700
rect 35440 22660 35480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 43112 22660 43152 22700
rect 43194 22660 43234 22700
rect 43276 22660 43316 22700
rect 43358 22660 43398 22700
rect 43440 22660 43480 22700
rect 47112 22660 47152 22700
rect 47194 22660 47234 22700
rect 47276 22660 47316 22700
rect 47358 22660 47398 22700
rect 47440 22660 47480 22700
rect 51112 22660 51152 22700
rect 51194 22660 51234 22700
rect 51276 22660 51316 22700
rect 51358 22660 51398 22700
rect 51440 22660 51480 22700
rect 55112 22660 55152 22700
rect 55194 22660 55234 22700
rect 55276 22660 55316 22700
rect 55358 22660 55398 22700
rect 55440 22660 55480 22700
rect 59112 22660 59152 22700
rect 59194 22660 59234 22700
rect 59276 22660 59316 22700
rect 59358 22660 59398 22700
rect 59440 22660 59480 22700
rect 63112 22660 63152 22700
rect 63194 22660 63234 22700
rect 63276 22660 63316 22700
rect 63358 22660 63398 22700
rect 63440 22660 63480 22700
rect 67112 22660 67152 22700
rect 67194 22660 67234 22700
rect 67276 22660 67316 22700
rect 67358 22660 67398 22700
rect 67440 22660 67480 22700
rect 71112 22660 71152 22700
rect 71194 22660 71234 22700
rect 71276 22660 71316 22700
rect 71358 22660 71398 22700
rect 71440 22660 71480 22700
rect 75112 22660 75152 22700
rect 75194 22660 75234 22700
rect 75276 22660 75316 22700
rect 75358 22660 75398 22700
rect 75440 22660 75480 22700
rect 79112 22660 79152 22700
rect 79194 22660 79234 22700
rect 79276 22660 79316 22700
rect 79358 22660 79398 22700
rect 79440 22660 79480 22700
rect 83112 22660 83152 22700
rect 83194 22660 83234 22700
rect 83276 22660 83316 22700
rect 83358 22660 83398 22700
rect 83440 22660 83480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 8352 21904 8392 21944
rect 8434 21904 8474 21944
rect 8516 21904 8556 21944
rect 8598 21904 8638 21944
rect 8680 21904 8720 21944
rect 12352 21904 12392 21944
rect 12434 21904 12474 21944
rect 12516 21904 12556 21944
rect 12598 21904 12638 21944
rect 12680 21904 12720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 20352 21904 20392 21944
rect 20434 21904 20474 21944
rect 20516 21904 20556 21944
rect 20598 21904 20638 21944
rect 20680 21904 20720 21944
rect 24352 21904 24392 21944
rect 24434 21904 24474 21944
rect 24516 21904 24556 21944
rect 24598 21904 24638 21944
rect 24680 21904 24720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 32352 21904 32392 21944
rect 32434 21904 32474 21944
rect 32516 21904 32556 21944
rect 32598 21904 32638 21944
rect 32680 21904 32720 21944
rect 36352 21904 36392 21944
rect 36434 21904 36474 21944
rect 36516 21904 36556 21944
rect 36598 21904 36638 21944
rect 36680 21904 36720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 44352 21904 44392 21944
rect 44434 21904 44474 21944
rect 44516 21904 44556 21944
rect 44598 21904 44638 21944
rect 44680 21904 44720 21944
rect 48352 21904 48392 21944
rect 48434 21904 48474 21944
rect 48516 21904 48556 21944
rect 48598 21904 48638 21944
rect 48680 21904 48720 21944
rect 52352 21904 52392 21944
rect 52434 21904 52474 21944
rect 52516 21904 52556 21944
rect 52598 21904 52638 21944
rect 52680 21904 52720 21944
rect 56352 21904 56392 21944
rect 56434 21904 56474 21944
rect 56516 21904 56556 21944
rect 56598 21904 56638 21944
rect 56680 21904 56720 21944
rect 60352 21904 60392 21944
rect 60434 21904 60474 21944
rect 60516 21904 60556 21944
rect 60598 21904 60638 21944
rect 60680 21904 60720 21944
rect 64352 21904 64392 21944
rect 64434 21904 64474 21944
rect 64516 21904 64556 21944
rect 64598 21904 64638 21944
rect 64680 21904 64720 21944
rect 68352 21904 68392 21944
rect 68434 21904 68474 21944
rect 68516 21904 68556 21944
rect 68598 21904 68638 21944
rect 68680 21904 68720 21944
rect 72352 21904 72392 21944
rect 72434 21904 72474 21944
rect 72516 21904 72556 21944
rect 72598 21904 72638 21944
rect 72680 21904 72720 21944
rect 76352 21904 76392 21944
rect 76434 21904 76474 21944
rect 76516 21904 76556 21944
rect 76598 21904 76638 21944
rect 76680 21904 76720 21944
rect 80352 21904 80392 21944
rect 80434 21904 80474 21944
rect 80516 21904 80556 21944
rect 80598 21904 80638 21944
rect 80680 21904 80720 21944
rect 84352 23416 84392 23456
rect 84434 23416 84474 23456
rect 84516 23416 84556 23456
rect 84598 23416 84638 23456
rect 84680 23416 84720 23456
rect 88352 23416 88392 23456
rect 88434 23416 88474 23456
rect 88516 23416 88556 23456
rect 88598 23416 88638 23456
rect 88680 23416 88720 23456
rect 92352 23416 92392 23456
rect 92434 23416 92474 23456
rect 92516 23416 92556 23456
rect 92598 23416 92638 23456
rect 92680 23416 92720 23456
rect 86668 23080 86708 23120
rect 87112 22660 87152 22700
rect 87194 22660 87234 22700
rect 87276 22660 87316 22700
rect 87358 22660 87398 22700
rect 87440 22660 87480 22700
rect 91112 22660 91152 22700
rect 91194 22660 91234 22700
rect 91276 22660 91316 22700
rect 91358 22660 91398 22700
rect 91440 22660 91480 22700
rect 84352 21904 84392 21944
rect 84434 21904 84474 21944
rect 84516 21904 84556 21944
rect 84598 21904 84638 21944
rect 84680 21904 84720 21944
rect 88352 21904 88392 21944
rect 88434 21904 88474 21944
rect 88516 21904 88556 21944
rect 88598 21904 88638 21944
rect 88680 21904 88720 21944
rect 92352 21904 92392 21944
rect 92434 21904 92474 21944
rect 92516 21904 92556 21944
rect 92598 21904 92638 21944
rect 92680 21904 92720 21944
rect 96352 23416 96392 23456
rect 96434 23416 96474 23456
rect 96516 23416 96556 23456
rect 96598 23416 96638 23456
rect 96680 23416 96720 23456
rect 95112 22660 95152 22700
rect 95194 22660 95234 22700
rect 95276 22660 95316 22700
rect 95358 22660 95398 22700
rect 95440 22660 95480 22700
rect 99112 22660 99152 22700
rect 99194 22660 99234 22700
rect 99276 22660 99316 22700
rect 99358 22660 99398 22700
rect 99440 22660 99480 22700
rect 96352 21904 96392 21944
rect 96434 21904 96474 21944
rect 96516 21904 96556 21944
rect 96598 21904 96638 21944
rect 96680 21904 96720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 7112 21148 7152 21188
rect 7194 21148 7234 21188
rect 7276 21148 7316 21188
rect 7358 21148 7398 21188
rect 7440 21148 7480 21188
rect 11112 21148 11152 21188
rect 11194 21148 11234 21188
rect 11276 21148 11316 21188
rect 11358 21148 11398 21188
rect 11440 21148 11480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 19112 21148 19152 21188
rect 19194 21148 19234 21188
rect 19276 21148 19316 21188
rect 19358 21148 19398 21188
rect 19440 21148 19480 21188
rect 23112 21148 23152 21188
rect 23194 21148 23234 21188
rect 23276 21148 23316 21188
rect 23358 21148 23398 21188
rect 23440 21148 23480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 31112 21148 31152 21188
rect 31194 21148 31234 21188
rect 31276 21148 31316 21188
rect 31358 21148 31398 21188
rect 31440 21148 31480 21188
rect 35112 21148 35152 21188
rect 35194 21148 35234 21188
rect 35276 21148 35316 21188
rect 35358 21148 35398 21188
rect 35440 21148 35480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 43112 21148 43152 21188
rect 43194 21148 43234 21188
rect 43276 21148 43316 21188
rect 43358 21148 43398 21188
rect 43440 21148 43480 21188
rect 47112 21148 47152 21188
rect 47194 21148 47234 21188
rect 47276 21148 47316 21188
rect 47358 21148 47398 21188
rect 47440 21148 47480 21188
rect 51112 21148 51152 21188
rect 51194 21148 51234 21188
rect 51276 21148 51316 21188
rect 51358 21148 51398 21188
rect 51440 21148 51480 21188
rect 55112 21148 55152 21188
rect 55194 21148 55234 21188
rect 55276 21148 55316 21188
rect 55358 21148 55398 21188
rect 55440 21148 55480 21188
rect 59112 21148 59152 21188
rect 59194 21148 59234 21188
rect 59276 21148 59316 21188
rect 59358 21148 59398 21188
rect 59440 21148 59480 21188
rect 63112 21148 63152 21188
rect 63194 21148 63234 21188
rect 63276 21148 63316 21188
rect 63358 21148 63398 21188
rect 63440 21148 63480 21188
rect 67112 21148 67152 21188
rect 67194 21148 67234 21188
rect 67276 21148 67316 21188
rect 67358 21148 67398 21188
rect 67440 21148 67480 21188
rect 71112 21148 71152 21188
rect 71194 21148 71234 21188
rect 71276 21148 71316 21188
rect 71358 21148 71398 21188
rect 71440 21148 71480 21188
rect 75112 21148 75152 21188
rect 75194 21148 75234 21188
rect 75276 21148 75316 21188
rect 75358 21148 75398 21188
rect 75440 21148 75480 21188
rect 79112 21148 79152 21188
rect 79194 21148 79234 21188
rect 79276 21148 79316 21188
rect 79358 21148 79398 21188
rect 79440 21148 79480 21188
rect 83112 21148 83152 21188
rect 83194 21148 83234 21188
rect 83276 21148 83316 21188
rect 83358 21148 83398 21188
rect 83440 21148 83480 21188
rect 87112 21148 87152 21188
rect 87194 21148 87234 21188
rect 87276 21148 87316 21188
rect 87358 21148 87398 21188
rect 87440 21148 87480 21188
rect 91112 21148 91152 21188
rect 91194 21148 91234 21188
rect 91276 21148 91316 21188
rect 91358 21148 91398 21188
rect 91440 21148 91480 21188
rect 95112 21148 95152 21188
rect 95194 21148 95234 21188
rect 95276 21148 95316 21188
rect 95358 21148 95398 21188
rect 95440 21148 95480 21188
rect 99112 21148 99152 21188
rect 99194 21148 99234 21188
rect 99276 21148 99316 21188
rect 99358 21148 99398 21188
rect 99440 21148 99480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 8352 20392 8392 20432
rect 8434 20392 8474 20432
rect 8516 20392 8556 20432
rect 8598 20392 8638 20432
rect 8680 20392 8720 20432
rect 12352 20392 12392 20432
rect 12434 20392 12474 20432
rect 12516 20392 12556 20432
rect 12598 20392 12638 20432
rect 12680 20392 12720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 20352 20392 20392 20432
rect 20434 20392 20474 20432
rect 20516 20392 20556 20432
rect 20598 20392 20638 20432
rect 20680 20392 20720 20432
rect 24352 20392 24392 20432
rect 24434 20392 24474 20432
rect 24516 20392 24556 20432
rect 24598 20392 24638 20432
rect 24680 20392 24720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 32352 20392 32392 20432
rect 32434 20392 32474 20432
rect 32516 20392 32556 20432
rect 32598 20392 32638 20432
rect 32680 20392 32720 20432
rect 36352 20392 36392 20432
rect 36434 20392 36474 20432
rect 36516 20392 36556 20432
rect 36598 20392 36638 20432
rect 36680 20392 36720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 44352 20392 44392 20432
rect 44434 20392 44474 20432
rect 44516 20392 44556 20432
rect 44598 20392 44638 20432
rect 44680 20392 44720 20432
rect 48352 20392 48392 20432
rect 48434 20392 48474 20432
rect 48516 20392 48556 20432
rect 48598 20392 48638 20432
rect 48680 20392 48720 20432
rect 52352 20392 52392 20432
rect 52434 20392 52474 20432
rect 52516 20392 52556 20432
rect 52598 20392 52638 20432
rect 52680 20392 52720 20432
rect 56352 20392 56392 20432
rect 56434 20392 56474 20432
rect 56516 20392 56556 20432
rect 56598 20392 56638 20432
rect 56680 20392 56720 20432
rect 60352 20392 60392 20432
rect 60434 20392 60474 20432
rect 60516 20392 60556 20432
rect 60598 20392 60638 20432
rect 60680 20392 60720 20432
rect 64352 20392 64392 20432
rect 64434 20392 64474 20432
rect 64516 20392 64556 20432
rect 64598 20392 64638 20432
rect 64680 20392 64720 20432
rect 68352 20392 68392 20432
rect 68434 20392 68474 20432
rect 68516 20392 68556 20432
rect 68598 20392 68638 20432
rect 68680 20392 68720 20432
rect 72352 20392 72392 20432
rect 72434 20392 72474 20432
rect 72516 20392 72556 20432
rect 72598 20392 72638 20432
rect 72680 20392 72720 20432
rect 76352 20392 76392 20432
rect 76434 20392 76474 20432
rect 76516 20392 76556 20432
rect 76598 20392 76638 20432
rect 76680 20392 76720 20432
rect 80352 20392 80392 20432
rect 80434 20392 80474 20432
rect 80516 20392 80556 20432
rect 80598 20392 80638 20432
rect 80680 20392 80720 20432
rect 84352 20392 84392 20432
rect 84434 20392 84474 20432
rect 84516 20392 84556 20432
rect 84598 20392 84638 20432
rect 84680 20392 84720 20432
rect 88352 20392 88392 20432
rect 88434 20392 88474 20432
rect 88516 20392 88556 20432
rect 88598 20392 88638 20432
rect 88680 20392 88720 20432
rect 92352 20392 92392 20432
rect 92434 20392 92474 20432
rect 92516 20392 92556 20432
rect 92598 20392 92638 20432
rect 92680 20392 92720 20432
rect 96352 20392 96392 20432
rect 96434 20392 96474 20432
rect 96516 20392 96556 20432
rect 96598 20392 96638 20432
rect 96680 20392 96720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 7112 19636 7152 19676
rect 7194 19636 7234 19676
rect 7276 19636 7316 19676
rect 7358 19636 7398 19676
rect 7440 19636 7480 19676
rect 11112 19636 11152 19676
rect 11194 19636 11234 19676
rect 11276 19636 11316 19676
rect 11358 19636 11398 19676
rect 11440 19636 11480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 19112 19636 19152 19676
rect 19194 19636 19234 19676
rect 19276 19636 19316 19676
rect 19358 19636 19398 19676
rect 19440 19636 19480 19676
rect 23112 19636 23152 19676
rect 23194 19636 23234 19676
rect 23276 19636 23316 19676
rect 23358 19636 23398 19676
rect 23440 19636 23480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 31112 19636 31152 19676
rect 31194 19636 31234 19676
rect 31276 19636 31316 19676
rect 31358 19636 31398 19676
rect 31440 19636 31480 19676
rect 35112 19636 35152 19676
rect 35194 19636 35234 19676
rect 35276 19636 35316 19676
rect 35358 19636 35398 19676
rect 35440 19636 35480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 43112 19636 43152 19676
rect 43194 19636 43234 19676
rect 43276 19636 43316 19676
rect 43358 19636 43398 19676
rect 43440 19636 43480 19676
rect 47112 19636 47152 19676
rect 47194 19636 47234 19676
rect 47276 19636 47316 19676
rect 47358 19636 47398 19676
rect 47440 19636 47480 19676
rect 51112 19636 51152 19676
rect 51194 19636 51234 19676
rect 51276 19636 51316 19676
rect 51358 19636 51398 19676
rect 51440 19636 51480 19676
rect 55112 19636 55152 19676
rect 55194 19636 55234 19676
rect 55276 19636 55316 19676
rect 55358 19636 55398 19676
rect 55440 19636 55480 19676
rect 59112 19636 59152 19676
rect 59194 19636 59234 19676
rect 59276 19636 59316 19676
rect 59358 19636 59398 19676
rect 59440 19636 59480 19676
rect 63112 19636 63152 19676
rect 63194 19636 63234 19676
rect 63276 19636 63316 19676
rect 63358 19636 63398 19676
rect 63440 19636 63480 19676
rect 67112 19636 67152 19676
rect 67194 19636 67234 19676
rect 67276 19636 67316 19676
rect 67358 19636 67398 19676
rect 67440 19636 67480 19676
rect 71112 19636 71152 19676
rect 71194 19636 71234 19676
rect 71276 19636 71316 19676
rect 71358 19636 71398 19676
rect 71440 19636 71480 19676
rect 75112 19636 75152 19676
rect 75194 19636 75234 19676
rect 75276 19636 75316 19676
rect 75358 19636 75398 19676
rect 75440 19636 75480 19676
rect 79112 19636 79152 19676
rect 79194 19636 79234 19676
rect 79276 19636 79316 19676
rect 79358 19636 79398 19676
rect 79440 19636 79480 19676
rect 83112 19636 83152 19676
rect 83194 19636 83234 19676
rect 83276 19636 83316 19676
rect 83358 19636 83398 19676
rect 83440 19636 83480 19676
rect 87112 19636 87152 19676
rect 87194 19636 87234 19676
rect 87276 19636 87316 19676
rect 87358 19636 87398 19676
rect 87440 19636 87480 19676
rect 91112 19636 91152 19676
rect 91194 19636 91234 19676
rect 91276 19636 91316 19676
rect 91358 19636 91398 19676
rect 91440 19636 91480 19676
rect 95112 19636 95152 19676
rect 95194 19636 95234 19676
rect 95276 19636 95316 19676
rect 95358 19636 95398 19676
rect 95440 19636 95480 19676
rect 99112 19636 99152 19676
rect 99194 19636 99234 19676
rect 99276 19636 99316 19676
rect 99358 19636 99398 19676
rect 99440 19636 99480 19676
rect 86764 19300 86804 19340
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 8352 18880 8392 18920
rect 8434 18880 8474 18920
rect 8516 18880 8556 18920
rect 8598 18880 8638 18920
rect 8680 18880 8720 18920
rect 12352 18880 12392 18920
rect 12434 18880 12474 18920
rect 12516 18880 12556 18920
rect 12598 18880 12638 18920
rect 12680 18880 12720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 20352 18880 20392 18920
rect 20434 18880 20474 18920
rect 20516 18880 20556 18920
rect 20598 18880 20638 18920
rect 20680 18880 20720 18920
rect 24352 18880 24392 18920
rect 24434 18880 24474 18920
rect 24516 18880 24556 18920
rect 24598 18880 24638 18920
rect 24680 18880 24720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 32352 18880 32392 18920
rect 32434 18880 32474 18920
rect 32516 18880 32556 18920
rect 32598 18880 32638 18920
rect 32680 18880 32720 18920
rect 36352 18880 36392 18920
rect 36434 18880 36474 18920
rect 36516 18880 36556 18920
rect 36598 18880 36638 18920
rect 36680 18880 36720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 44352 18880 44392 18920
rect 44434 18880 44474 18920
rect 44516 18880 44556 18920
rect 44598 18880 44638 18920
rect 44680 18880 44720 18920
rect 48352 18880 48392 18920
rect 48434 18880 48474 18920
rect 48516 18880 48556 18920
rect 48598 18880 48638 18920
rect 48680 18880 48720 18920
rect 52352 18880 52392 18920
rect 52434 18880 52474 18920
rect 52516 18880 52556 18920
rect 52598 18880 52638 18920
rect 52680 18880 52720 18920
rect 56352 18880 56392 18920
rect 56434 18880 56474 18920
rect 56516 18880 56556 18920
rect 56598 18880 56638 18920
rect 56680 18880 56720 18920
rect 60352 18880 60392 18920
rect 60434 18880 60474 18920
rect 60516 18880 60556 18920
rect 60598 18880 60638 18920
rect 60680 18880 60720 18920
rect 64352 18880 64392 18920
rect 64434 18880 64474 18920
rect 64516 18880 64556 18920
rect 64598 18880 64638 18920
rect 64680 18880 64720 18920
rect 68352 18880 68392 18920
rect 68434 18880 68474 18920
rect 68516 18880 68556 18920
rect 68598 18880 68638 18920
rect 68680 18880 68720 18920
rect 72352 18880 72392 18920
rect 72434 18880 72474 18920
rect 72516 18880 72556 18920
rect 72598 18880 72638 18920
rect 72680 18880 72720 18920
rect 76352 18880 76392 18920
rect 76434 18880 76474 18920
rect 76516 18880 76556 18920
rect 76598 18880 76638 18920
rect 76680 18880 76720 18920
rect 80352 18880 80392 18920
rect 80434 18880 80474 18920
rect 80516 18880 80556 18920
rect 80598 18880 80638 18920
rect 80680 18880 80720 18920
rect 84352 18880 84392 18920
rect 84434 18880 84474 18920
rect 84516 18880 84556 18920
rect 84598 18880 84638 18920
rect 84680 18880 84720 18920
rect 88352 18880 88392 18920
rect 88434 18880 88474 18920
rect 88516 18880 88556 18920
rect 88598 18880 88638 18920
rect 88680 18880 88720 18920
rect 92352 18880 92392 18920
rect 92434 18880 92474 18920
rect 92516 18880 92556 18920
rect 92598 18880 92638 18920
rect 92680 18880 92720 18920
rect 96352 18880 96392 18920
rect 96434 18880 96474 18920
rect 96516 18880 96556 18920
rect 96598 18880 96638 18920
rect 96680 18880 96720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 7112 18124 7152 18164
rect 7194 18124 7234 18164
rect 7276 18124 7316 18164
rect 7358 18124 7398 18164
rect 7440 18124 7480 18164
rect 11112 18124 11152 18164
rect 11194 18124 11234 18164
rect 11276 18124 11316 18164
rect 11358 18124 11398 18164
rect 11440 18124 11480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 19112 18124 19152 18164
rect 19194 18124 19234 18164
rect 19276 18124 19316 18164
rect 19358 18124 19398 18164
rect 19440 18124 19480 18164
rect 23112 18124 23152 18164
rect 23194 18124 23234 18164
rect 23276 18124 23316 18164
rect 23358 18124 23398 18164
rect 23440 18124 23480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 31112 18124 31152 18164
rect 31194 18124 31234 18164
rect 31276 18124 31316 18164
rect 31358 18124 31398 18164
rect 31440 18124 31480 18164
rect 35112 18124 35152 18164
rect 35194 18124 35234 18164
rect 35276 18124 35316 18164
rect 35358 18124 35398 18164
rect 35440 18124 35480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 43112 18124 43152 18164
rect 43194 18124 43234 18164
rect 43276 18124 43316 18164
rect 43358 18124 43398 18164
rect 43440 18124 43480 18164
rect 47112 18124 47152 18164
rect 47194 18124 47234 18164
rect 47276 18124 47316 18164
rect 47358 18124 47398 18164
rect 47440 18124 47480 18164
rect 51112 18124 51152 18164
rect 51194 18124 51234 18164
rect 51276 18124 51316 18164
rect 51358 18124 51398 18164
rect 51440 18124 51480 18164
rect 55112 18124 55152 18164
rect 55194 18124 55234 18164
rect 55276 18124 55316 18164
rect 55358 18124 55398 18164
rect 55440 18124 55480 18164
rect 59112 18124 59152 18164
rect 59194 18124 59234 18164
rect 59276 18124 59316 18164
rect 59358 18124 59398 18164
rect 59440 18124 59480 18164
rect 63112 18124 63152 18164
rect 63194 18124 63234 18164
rect 63276 18124 63316 18164
rect 63358 18124 63398 18164
rect 63440 18124 63480 18164
rect 67112 18124 67152 18164
rect 67194 18124 67234 18164
rect 67276 18124 67316 18164
rect 67358 18124 67398 18164
rect 67440 18124 67480 18164
rect 71112 18124 71152 18164
rect 71194 18124 71234 18164
rect 71276 18124 71316 18164
rect 71358 18124 71398 18164
rect 71440 18124 71480 18164
rect 75112 18124 75152 18164
rect 75194 18124 75234 18164
rect 75276 18124 75316 18164
rect 75358 18124 75398 18164
rect 75440 18124 75480 18164
rect 79112 18124 79152 18164
rect 79194 18124 79234 18164
rect 79276 18124 79316 18164
rect 79358 18124 79398 18164
rect 79440 18124 79480 18164
rect 83112 18124 83152 18164
rect 83194 18124 83234 18164
rect 83276 18124 83316 18164
rect 83358 18124 83398 18164
rect 83440 18124 83480 18164
rect 87112 18124 87152 18164
rect 87194 18124 87234 18164
rect 87276 18124 87316 18164
rect 87358 18124 87398 18164
rect 87440 18124 87480 18164
rect 91112 18124 91152 18164
rect 91194 18124 91234 18164
rect 91276 18124 91316 18164
rect 91358 18124 91398 18164
rect 91440 18124 91480 18164
rect 95112 18124 95152 18164
rect 95194 18124 95234 18164
rect 95276 18124 95316 18164
rect 95358 18124 95398 18164
rect 95440 18124 95480 18164
rect 99112 18124 99152 18164
rect 99194 18124 99234 18164
rect 99276 18124 99316 18164
rect 99358 18124 99398 18164
rect 99440 18124 99480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 8352 17368 8392 17408
rect 8434 17368 8474 17408
rect 8516 17368 8556 17408
rect 8598 17368 8638 17408
rect 8680 17368 8720 17408
rect 12352 17368 12392 17408
rect 12434 17368 12474 17408
rect 12516 17368 12556 17408
rect 12598 17368 12638 17408
rect 12680 17368 12720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 20352 17368 20392 17408
rect 20434 17368 20474 17408
rect 20516 17368 20556 17408
rect 20598 17368 20638 17408
rect 20680 17368 20720 17408
rect 24352 17368 24392 17408
rect 24434 17368 24474 17408
rect 24516 17368 24556 17408
rect 24598 17368 24638 17408
rect 24680 17368 24720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 32352 17368 32392 17408
rect 32434 17368 32474 17408
rect 32516 17368 32556 17408
rect 32598 17368 32638 17408
rect 32680 17368 32720 17408
rect 36352 17368 36392 17408
rect 36434 17368 36474 17408
rect 36516 17368 36556 17408
rect 36598 17368 36638 17408
rect 36680 17368 36720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 44352 17368 44392 17408
rect 44434 17368 44474 17408
rect 44516 17368 44556 17408
rect 44598 17368 44638 17408
rect 44680 17368 44720 17408
rect 48352 17368 48392 17408
rect 48434 17368 48474 17408
rect 48516 17368 48556 17408
rect 48598 17368 48638 17408
rect 48680 17368 48720 17408
rect 52352 17368 52392 17408
rect 52434 17368 52474 17408
rect 52516 17368 52556 17408
rect 52598 17368 52638 17408
rect 52680 17368 52720 17408
rect 56352 17368 56392 17408
rect 56434 17368 56474 17408
rect 56516 17368 56556 17408
rect 56598 17368 56638 17408
rect 56680 17368 56720 17408
rect 60352 17368 60392 17408
rect 60434 17368 60474 17408
rect 60516 17368 60556 17408
rect 60598 17368 60638 17408
rect 60680 17368 60720 17408
rect 64352 17368 64392 17408
rect 64434 17368 64474 17408
rect 64516 17368 64556 17408
rect 64598 17368 64638 17408
rect 64680 17368 64720 17408
rect 68352 17368 68392 17408
rect 68434 17368 68474 17408
rect 68516 17368 68556 17408
rect 68598 17368 68638 17408
rect 68680 17368 68720 17408
rect 72352 17368 72392 17408
rect 72434 17368 72474 17408
rect 72516 17368 72556 17408
rect 72598 17368 72638 17408
rect 72680 17368 72720 17408
rect 76352 17368 76392 17408
rect 76434 17368 76474 17408
rect 76516 17368 76556 17408
rect 76598 17368 76638 17408
rect 76680 17368 76720 17408
rect 80352 17368 80392 17408
rect 80434 17368 80474 17408
rect 80516 17368 80556 17408
rect 80598 17368 80638 17408
rect 80680 17368 80720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 7112 16612 7152 16652
rect 7194 16612 7234 16652
rect 7276 16612 7316 16652
rect 7358 16612 7398 16652
rect 7440 16612 7480 16652
rect 11112 16612 11152 16652
rect 11194 16612 11234 16652
rect 11276 16612 11316 16652
rect 11358 16612 11398 16652
rect 11440 16612 11480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 19112 16612 19152 16652
rect 19194 16612 19234 16652
rect 19276 16612 19316 16652
rect 19358 16612 19398 16652
rect 19440 16612 19480 16652
rect 23112 16612 23152 16652
rect 23194 16612 23234 16652
rect 23276 16612 23316 16652
rect 23358 16612 23398 16652
rect 23440 16612 23480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 31112 16612 31152 16652
rect 31194 16612 31234 16652
rect 31276 16612 31316 16652
rect 31358 16612 31398 16652
rect 31440 16612 31480 16652
rect 35112 16612 35152 16652
rect 35194 16612 35234 16652
rect 35276 16612 35316 16652
rect 35358 16612 35398 16652
rect 35440 16612 35480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 43112 16612 43152 16652
rect 43194 16612 43234 16652
rect 43276 16612 43316 16652
rect 43358 16612 43398 16652
rect 43440 16612 43480 16652
rect 47112 16612 47152 16652
rect 47194 16612 47234 16652
rect 47276 16612 47316 16652
rect 47358 16612 47398 16652
rect 47440 16612 47480 16652
rect 51112 16612 51152 16652
rect 51194 16612 51234 16652
rect 51276 16612 51316 16652
rect 51358 16612 51398 16652
rect 51440 16612 51480 16652
rect 55112 16612 55152 16652
rect 55194 16612 55234 16652
rect 55276 16612 55316 16652
rect 55358 16612 55398 16652
rect 55440 16612 55480 16652
rect 59112 16612 59152 16652
rect 59194 16612 59234 16652
rect 59276 16612 59316 16652
rect 59358 16612 59398 16652
rect 59440 16612 59480 16652
rect 63112 16612 63152 16652
rect 63194 16612 63234 16652
rect 63276 16612 63316 16652
rect 63358 16612 63398 16652
rect 63440 16612 63480 16652
rect 67112 16612 67152 16652
rect 67194 16612 67234 16652
rect 67276 16612 67316 16652
rect 67358 16612 67398 16652
rect 67440 16612 67480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 8352 15856 8392 15896
rect 8434 15856 8474 15896
rect 8516 15856 8556 15896
rect 8598 15856 8638 15896
rect 8680 15856 8720 15896
rect 12352 15856 12392 15896
rect 12434 15856 12474 15896
rect 12516 15856 12556 15896
rect 12598 15856 12638 15896
rect 12680 15856 12720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 20352 15856 20392 15896
rect 20434 15856 20474 15896
rect 20516 15856 20556 15896
rect 20598 15856 20638 15896
rect 20680 15856 20720 15896
rect 24352 15856 24392 15896
rect 24434 15856 24474 15896
rect 24516 15856 24556 15896
rect 24598 15856 24638 15896
rect 24680 15856 24720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 32352 15856 32392 15896
rect 32434 15856 32474 15896
rect 32516 15856 32556 15896
rect 32598 15856 32638 15896
rect 32680 15856 32720 15896
rect 36352 15856 36392 15896
rect 36434 15856 36474 15896
rect 36516 15856 36556 15896
rect 36598 15856 36638 15896
rect 36680 15856 36720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 44352 15856 44392 15896
rect 44434 15856 44474 15896
rect 44516 15856 44556 15896
rect 44598 15856 44638 15896
rect 44680 15856 44720 15896
rect 48352 15856 48392 15896
rect 48434 15856 48474 15896
rect 48516 15856 48556 15896
rect 48598 15856 48638 15896
rect 48680 15856 48720 15896
rect 52352 15856 52392 15896
rect 52434 15856 52474 15896
rect 52516 15856 52556 15896
rect 52598 15856 52638 15896
rect 52680 15856 52720 15896
rect 56352 15856 56392 15896
rect 56434 15856 56474 15896
rect 56516 15856 56556 15896
rect 56598 15856 56638 15896
rect 56680 15856 56720 15896
rect 60352 15856 60392 15896
rect 60434 15856 60474 15896
rect 60516 15856 60556 15896
rect 60598 15856 60638 15896
rect 60680 15856 60720 15896
rect 64352 15856 64392 15896
rect 64434 15856 64474 15896
rect 64516 15856 64556 15896
rect 64598 15856 64638 15896
rect 64680 15856 64720 15896
rect 68352 15856 68392 15896
rect 68434 15856 68474 15896
rect 68516 15856 68556 15896
rect 68598 15856 68638 15896
rect 68680 15856 68720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 7112 15100 7152 15140
rect 7194 15100 7234 15140
rect 7276 15100 7316 15140
rect 7358 15100 7398 15140
rect 7440 15100 7480 15140
rect 11112 15100 11152 15140
rect 11194 15100 11234 15140
rect 11276 15100 11316 15140
rect 11358 15100 11398 15140
rect 11440 15100 11480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 19112 15100 19152 15140
rect 19194 15100 19234 15140
rect 19276 15100 19316 15140
rect 19358 15100 19398 15140
rect 19440 15100 19480 15140
rect 23112 15100 23152 15140
rect 23194 15100 23234 15140
rect 23276 15100 23316 15140
rect 23358 15100 23398 15140
rect 23440 15100 23480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 31112 15100 31152 15140
rect 31194 15100 31234 15140
rect 31276 15100 31316 15140
rect 31358 15100 31398 15140
rect 31440 15100 31480 15140
rect 35112 15100 35152 15140
rect 35194 15100 35234 15140
rect 35276 15100 35316 15140
rect 35358 15100 35398 15140
rect 35440 15100 35480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 43112 15100 43152 15140
rect 43194 15100 43234 15140
rect 43276 15100 43316 15140
rect 43358 15100 43398 15140
rect 43440 15100 43480 15140
rect 47112 15100 47152 15140
rect 47194 15100 47234 15140
rect 47276 15100 47316 15140
rect 47358 15100 47398 15140
rect 47440 15100 47480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 55112 15100 55152 15140
rect 55194 15100 55234 15140
rect 55276 15100 55316 15140
rect 55358 15100 55398 15140
rect 55440 15100 55480 15140
rect 59112 15100 59152 15140
rect 59194 15100 59234 15140
rect 59276 15100 59316 15140
rect 59358 15100 59398 15140
rect 59440 15100 59480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 67112 15100 67152 15140
rect 67194 15100 67234 15140
rect 67276 15100 67316 15140
rect 67358 15100 67398 15140
rect 67440 15100 67480 15140
rect 84352 17368 84392 17408
rect 84434 17368 84474 17408
rect 84516 17368 84556 17408
rect 84598 17368 84638 17408
rect 84680 17368 84720 17408
rect 88352 17368 88392 17408
rect 88434 17368 88474 17408
rect 88516 17368 88556 17408
rect 88598 17368 88638 17408
rect 88680 17368 88720 17408
rect 92352 17368 92392 17408
rect 92434 17368 92474 17408
rect 92516 17368 92556 17408
rect 92598 17368 92638 17408
rect 92680 17368 92720 17408
rect 96352 17368 96392 17408
rect 96434 17368 96474 17408
rect 96516 17368 96556 17408
rect 96598 17368 96638 17408
rect 96680 17368 96720 17408
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 8352 14344 8392 14384
rect 8434 14344 8474 14384
rect 8516 14344 8556 14384
rect 8598 14344 8638 14384
rect 8680 14344 8720 14384
rect 12352 14344 12392 14384
rect 12434 14344 12474 14384
rect 12516 14344 12556 14384
rect 12598 14344 12638 14384
rect 12680 14344 12720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 20352 14344 20392 14384
rect 20434 14344 20474 14384
rect 20516 14344 20556 14384
rect 20598 14344 20638 14384
rect 20680 14344 20720 14384
rect 24352 14344 24392 14384
rect 24434 14344 24474 14384
rect 24516 14344 24556 14384
rect 24598 14344 24638 14384
rect 24680 14344 24720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 32352 14344 32392 14384
rect 32434 14344 32474 14384
rect 32516 14344 32556 14384
rect 32598 14344 32638 14384
rect 32680 14344 32720 14384
rect 36352 14344 36392 14384
rect 36434 14344 36474 14384
rect 36516 14344 36556 14384
rect 36598 14344 36638 14384
rect 36680 14344 36720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 44352 14344 44392 14384
rect 44434 14344 44474 14384
rect 44516 14344 44556 14384
rect 44598 14344 44638 14384
rect 44680 14344 44720 14384
rect 48352 14344 48392 14384
rect 48434 14344 48474 14384
rect 48516 14344 48556 14384
rect 48598 14344 48638 14384
rect 48680 14344 48720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 56352 14344 56392 14384
rect 56434 14344 56474 14384
rect 56516 14344 56556 14384
rect 56598 14344 56638 14384
rect 56680 14344 56720 14384
rect 60352 14344 60392 14384
rect 60434 14344 60474 14384
rect 60516 14344 60556 14384
rect 60598 14344 60638 14384
rect 60680 14344 60720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 68352 14344 68392 14384
rect 68434 14344 68474 14384
rect 68516 14344 68556 14384
rect 68598 14344 68638 14384
rect 68680 14344 68720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 7112 13588 7152 13628
rect 7194 13588 7234 13628
rect 7276 13588 7316 13628
rect 7358 13588 7398 13628
rect 7440 13588 7480 13628
rect 11112 13588 11152 13628
rect 11194 13588 11234 13628
rect 11276 13588 11316 13628
rect 11358 13588 11398 13628
rect 11440 13588 11480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 19112 13588 19152 13628
rect 19194 13588 19234 13628
rect 19276 13588 19316 13628
rect 19358 13588 19398 13628
rect 19440 13588 19480 13628
rect 23112 13588 23152 13628
rect 23194 13588 23234 13628
rect 23276 13588 23316 13628
rect 23358 13588 23398 13628
rect 23440 13588 23480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 31112 13588 31152 13628
rect 31194 13588 31234 13628
rect 31276 13588 31316 13628
rect 31358 13588 31398 13628
rect 31440 13588 31480 13628
rect 35112 13588 35152 13628
rect 35194 13588 35234 13628
rect 35276 13588 35316 13628
rect 35358 13588 35398 13628
rect 35440 13588 35480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 43112 13588 43152 13628
rect 43194 13588 43234 13628
rect 43276 13588 43316 13628
rect 43358 13588 43398 13628
rect 43440 13588 43480 13628
rect 47112 13588 47152 13628
rect 47194 13588 47234 13628
rect 47276 13588 47316 13628
rect 47358 13588 47398 13628
rect 47440 13588 47480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 55112 13588 55152 13628
rect 55194 13588 55234 13628
rect 55276 13588 55316 13628
rect 55358 13588 55398 13628
rect 55440 13588 55480 13628
rect 59112 13588 59152 13628
rect 59194 13588 59234 13628
rect 59276 13588 59316 13628
rect 59358 13588 59398 13628
rect 59440 13588 59480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 67112 13588 67152 13628
rect 67194 13588 67234 13628
rect 67276 13588 67316 13628
rect 67358 13588 67398 13628
rect 67440 13588 67480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 8352 12832 8392 12872
rect 8434 12832 8474 12872
rect 8516 12832 8556 12872
rect 8598 12832 8638 12872
rect 8680 12832 8720 12872
rect 12352 12832 12392 12872
rect 12434 12832 12474 12872
rect 12516 12832 12556 12872
rect 12598 12832 12638 12872
rect 12680 12832 12720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 20352 12832 20392 12872
rect 20434 12832 20474 12872
rect 20516 12832 20556 12872
rect 20598 12832 20638 12872
rect 20680 12832 20720 12872
rect 24352 12832 24392 12872
rect 24434 12832 24474 12872
rect 24516 12832 24556 12872
rect 24598 12832 24638 12872
rect 24680 12832 24720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 32352 12832 32392 12872
rect 32434 12832 32474 12872
rect 32516 12832 32556 12872
rect 32598 12832 32638 12872
rect 32680 12832 32720 12872
rect 36352 12832 36392 12872
rect 36434 12832 36474 12872
rect 36516 12832 36556 12872
rect 36598 12832 36638 12872
rect 36680 12832 36720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 44352 12832 44392 12872
rect 44434 12832 44474 12872
rect 44516 12832 44556 12872
rect 44598 12832 44638 12872
rect 44680 12832 44720 12872
rect 48352 12832 48392 12872
rect 48434 12832 48474 12872
rect 48516 12832 48556 12872
rect 48598 12832 48638 12872
rect 48680 12832 48720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 56352 12832 56392 12872
rect 56434 12832 56474 12872
rect 56516 12832 56556 12872
rect 56598 12832 56638 12872
rect 56680 12832 56720 12872
rect 60352 12832 60392 12872
rect 60434 12832 60474 12872
rect 60516 12832 60556 12872
rect 60598 12832 60638 12872
rect 60680 12832 60720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 68352 12832 68392 12872
rect 68434 12832 68474 12872
rect 68516 12832 68556 12872
rect 68598 12832 68638 12872
rect 68680 12832 68720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 7112 12076 7152 12116
rect 7194 12076 7234 12116
rect 7276 12076 7316 12116
rect 7358 12076 7398 12116
rect 7440 12076 7480 12116
rect 11112 12076 11152 12116
rect 11194 12076 11234 12116
rect 11276 12076 11316 12116
rect 11358 12076 11398 12116
rect 11440 12076 11480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 19112 12076 19152 12116
rect 19194 12076 19234 12116
rect 19276 12076 19316 12116
rect 19358 12076 19398 12116
rect 19440 12076 19480 12116
rect 23112 12076 23152 12116
rect 23194 12076 23234 12116
rect 23276 12076 23316 12116
rect 23358 12076 23398 12116
rect 23440 12076 23480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 31112 12076 31152 12116
rect 31194 12076 31234 12116
rect 31276 12076 31316 12116
rect 31358 12076 31398 12116
rect 31440 12076 31480 12116
rect 35112 12076 35152 12116
rect 35194 12076 35234 12116
rect 35276 12076 35316 12116
rect 35358 12076 35398 12116
rect 35440 12076 35480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 43112 12076 43152 12116
rect 43194 12076 43234 12116
rect 43276 12076 43316 12116
rect 43358 12076 43398 12116
rect 43440 12076 43480 12116
rect 47112 12076 47152 12116
rect 47194 12076 47234 12116
rect 47276 12076 47316 12116
rect 47358 12076 47398 12116
rect 47440 12076 47480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 55112 12076 55152 12116
rect 55194 12076 55234 12116
rect 55276 12076 55316 12116
rect 55358 12076 55398 12116
rect 55440 12076 55480 12116
rect 59112 12076 59152 12116
rect 59194 12076 59234 12116
rect 59276 12076 59316 12116
rect 59358 12076 59398 12116
rect 59440 12076 59480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 67112 12076 67152 12116
rect 67194 12076 67234 12116
rect 67276 12076 67316 12116
rect 67358 12076 67398 12116
rect 67440 12076 67480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 8352 11320 8392 11360
rect 8434 11320 8474 11360
rect 8516 11320 8556 11360
rect 8598 11320 8638 11360
rect 8680 11320 8720 11360
rect 12352 11320 12392 11360
rect 12434 11320 12474 11360
rect 12516 11320 12556 11360
rect 12598 11320 12638 11360
rect 12680 11320 12720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 20352 11320 20392 11360
rect 20434 11320 20474 11360
rect 20516 11320 20556 11360
rect 20598 11320 20638 11360
rect 20680 11320 20720 11360
rect 24352 11320 24392 11360
rect 24434 11320 24474 11360
rect 24516 11320 24556 11360
rect 24598 11320 24638 11360
rect 24680 11320 24720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 32352 11320 32392 11360
rect 32434 11320 32474 11360
rect 32516 11320 32556 11360
rect 32598 11320 32638 11360
rect 32680 11320 32720 11360
rect 36352 11320 36392 11360
rect 36434 11320 36474 11360
rect 36516 11320 36556 11360
rect 36598 11320 36638 11360
rect 36680 11320 36720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 44352 11320 44392 11360
rect 44434 11320 44474 11360
rect 44516 11320 44556 11360
rect 44598 11320 44638 11360
rect 44680 11320 44720 11360
rect 48352 11320 48392 11360
rect 48434 11320 48474 11360
rect 48516 11320 48556 11360
rect 48598 11320 48638 11360
rect 48680 11320 48720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 56352 11320 56392 11360
rect 56434 11320 56474 11360
rect 56516 11320 56556 11360
rect 56598 11320 56638 11360
rect 56680 11320 56720 11360
rect 60352 11320 60392 11360
rect 60434 11320 60474 11360
rect 60516 11320 60556 11360
rect 60598 11320 60638 11360
rect 60680 11320 60720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 68352 11320 68392 11360
rect 68434 11320 68474 11360
rect 68516 11320 68556 11360
rect 68598 11320 68638 11360
rect 68680 11320 68720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 7112 10564 7152 10604
rect 7194 10564 7234 10604
rect 7276 10564 7316 10604
rect 7358 10564 7398 10604
rect 7440 10564 7480 10604
rect 11112 10564 11152 10604
rect 11194 10564 11234 10604
rect 11276 10564 11316 10604
rect 11358 10564 11398 10604
rect 11440 10564 11480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 19112 10564 19152 10604
rect 19194 10564 19234 10604
rect 19276 10564 19316 10604
rect 19358 10564 19398 10604
rect 19440 10564 19480 10604
rect 23112 10564 23152 10604
rect 23194 10564 23234 10604
rect 23276 10564 23316 10604
rect 23358 10564 23398 10604
rect 23440 10564 23480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 31112 10564 31152 10604
rect 31194 10564 31234 10604
rect 31276 10564 31316 10604
rect 31358 10564 31398 10604
rect 31440 10564 31480 10604
rect 35112 10564 35152 10604
rect 35194 10564 35234 10604
rect 35276 10564 35316 10604
rect 35358 10564 35398 10604
rect 35440 10564 35480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 43112 10564 43152 10604
rect 43194 10564 43234 10604
rect 43276 10564 43316 10604
rect 43358 10564 43398 10604
rect 43440 10564 43480 10604
rect 47112 10564 47152 10604
rect 47194 10564 47234 10604
rect 47276 10564 47316 10604
rect 47358 10564 47398 10604
rect 47440 10564 47480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 55112 10564 55152 10604
rect 55194 10564 55234 10604
rect 55276 10564 55316 10604
rect 55358 10564 55398 10604
rect 55440 10564 55480 10604
rect 59112 10564 59152 10604
rect 59194 10564 59234 10604
rect 59276 10564 59316 10604
rect 59358 10564 59398 10604
rect 59440 10564 59480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 67112 10564 67152 10604
rect 67194 10564 67234 10604
rect 67276 10564 67316 10604
rect 67358 10564 67398 10604
rect 67440 10564 67480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 8352 9808 8392 9848
rect 8434 9808 8474 9848
rect 8516 9808 8556 9848
rect 8598 9808 8638 9848
rect 8680 9808 8720 9848
rect 12352 9808 12392 9848
rect 12434 9808 12474 9848
rect 12516 9808 12556 9848
rect 12598 9808 12638 9848
rect 12680 9808 12720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 20352 9808 20392 9848
rect 20434 9808 20474 9848
rect 20516 9808 20556 9848
rect 20598 9808 20638 9848
rect 20680 9808 20720 9848
rect 24352 9808 24392 9848
rect 24434 9808 24474 9848
rect 24516 9808 24556 9848
rect 24598 9808 24638 9848
rect 24680 9808 24720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 32352 9808 32392 9848
rect 32434 9808 32474 9848
rect 32516 9808 32556 9848
rect 32598 9808 32638 9848
rect 32680 9808 32720 9848
rect 36352 9808 36392 9848
rect 36434 9808 36474 9848
rect 36516 9808 36556 9848
rect 36598 9808 36638 9848
rect 36680 9808 36720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 44352 9808 44392 9848
rect 44434 9808 44474 9848
rect 44516 9808 44556 9848
rect 44598 9808 44638 9848
rect 44680 9808 44720 9848
rect 48352 9808 48392 9848
rect 48434 9808 48474 9848
rect 48516 9808 48556 9848
rect 48598 9808 48638 9848
rect 48680 9808 48720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 56352 9808 56392 9848
rect 56434 9808 56474 9848
rect 56516 9808 56556 9848
rect 56598 9808 56638 9848
rect 56680 9808 56720 9848
rect 60352 9808 60392 9848
rect 60434 9808 60474 9848
rect 60516 9808 60556 9848
rect 60598 9808 60638 9848
rect 60680 9808 60720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 68352 9808 68392 9848
rect 68434 9808 68474 9848
rect 68516 9808 68556 9848
rect 68598 9808 68638 9848
rect 68680 9808 68720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 7112 9052 7152 9092
rect 7194 9052 7234 9092
rect 7276 9052 7316 9092
rect 7358 9052 7398 9092
rect 7440 9052 7480 9092
rect 11112 9052 11152 9092
rect 11194 9052 11234 9092
rect 11276 9052 11316 9092
rect 11358 9052 11398 9092
rect 11440 9052 11480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 19112 9052 19152 9092
rect 19194 9052 19234 9092
rect 19276 9052 19316 9092
rect 19358 9052 19398 9092
rect 19440 9052 19480 9092
rect 23112 9052 23152 9092
rect 23194 9052 23234 9092
rect 23276 9052 23316 9092
rect 23358 9052 23398 9092
rect 23440 9052 23480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 31112 9052 31152 9092
rect 31194 9052 31234 9092
rect 31276 9052 31316 9092
rect 31358 9052 31398 9092
rect 31440 9052 31480 9092
rect 35112 9052 35152 9092
rect 35194 9052 35234 9092
rect 35276 9052 35316 9092
rect 35358 9052 35398 9092
rect 35440 9052 35480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 43112 9052 43152 9092
rect 43194 9052 43234 9092
rect 43276 9052 43316 9092
rect 43358 9052 43398 9092
rect 43440 9052 43480 9092
rect 47112 9052 47152 9092
rect 47194 9052 47234 9092
rect 47276 9052 47316 9092
rect 47358 9052 47398 9092
rect 47440 9052 47480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 55112 9052 55152 9092
rect 55194 9052 55234 9092
rect 55276 9052 55316 9092
rect 55358 9052 55398 9092
rect 55440 9052 55480 9092
rect 59112 9052 59152 9092
rect 59194 9052 59234 9092
rect 59276 9052 59316 9092
rect 59358 9052 59398 9092
rect 59440 9052 59480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 67112 9052 67152 9092
rect 67194 9052 67234 9092
rect 67276 9052 67316 9092
rect 67358 9052 67398 9092
rect 67440 9052 67480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 8352 8296 8392 8336
rect 8434 8296 8474 8336
rect 8516 8296 8556 8336
rect 8598 8296 8638 8336
rect 8680 8296 8720 8336
rect 12352 8296 12392 8336
rect 12434 8296 12474 8336
rect 12516 8296 12556 8336
rect 12598 8296 12638 8336
rect 12680 8296 12720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 20352 8296 20392 8336
rect 20434 8296 20474 8336
rect 20516 8296 20556 8336
rect 20598 8296 20638 8336
rect 20680 8296 20720 8336
rect 24352 8296 24392 8336
rect 24434 8296 24474 8336
rect 24516 8296 24556 8336
rect 24598 8296 24638 8336
rect 24680 8296 24720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 32352 8296 32392 8336
rect 32434 8296 32474 8336
rect 32516 8296 32556 8336
rect 32598 8296 32638 8336
rect 32680 8296 32720 8336
rect 36352 8296 36392 8336
rect 36434 8296 36474 8336
rect 36516 8296 36556 8336
rect 36598 8296 36638 8336
rect 36680 8296 36720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 44352 8296 44392 8336
rect 44434 8296 44474 8336
rect 44516 8296 44556 8336
rect 44598 8296 44638 8336
rect 44680 8296 44720 8336
rect 48352 8296 48392 8336
rect 48434 8296 48474 8336
rect 48516 8296 48556 8336
rect 48598 8296 48638 8336
rect 48680 8296 48720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 56352 8296 56392 8336
rect 56434 8296 56474 8336
rect 56516 8296 56556 8336
rect 56598 8296 56638 8336
rect 56680 8296 56720 8336
rect 60352 8296 60392 8336
rect 60434 8296 60474 8336
rect 60516 8296 60556 8336
rect 60598 8296 60638 8336
rect 60680 8296 60720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 68352 8296 68392 8336
rect 68434 8296 68474 8336
rect 68516 8296 68556 8336
rect 68598 8296 68638 8336
rect 68680 8296 68720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 7112 7540 7152 7580
rect 7194 7540 7234 7580
rect 7276 7540 7316 7580
rect 7358 7540 7398 7580
rect 7440 7540 7480 7580
rect 11112 7540 11152 7580
rect 11194 7540 11234 7580
rect 11276 7540 11316 7580
rect 11358 7540 11398 7580
rect 11440 7540 11480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 19112 7540 19152 7580
rect 19194 7540 19234 7580
rect 19276 7540 19316 7580
rect 19358 7540 19398 7580
rect 19440 7540 19480 7580
rect 23112 7540 23152 7580
rect 23194 7540 23234 7580
rect 23276 7540 23316 7580
rect 23358 7540 23398 7580
rect 23440 7540 23480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 31112 7540 31152 7580
rect 31194 7540 31234 7580
rect 31276 7540 31316 7580
rect 31358 7540 31398 7580
rect 31440 7540 31480 7580
rect 35112 7540 35152 7580
rect 35194 7540 35234 7580
rect 35276 7540 35316 7580
rect 35358 7540 35398 7580
rect 35440 7540 35480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 43112 7540 43152 7580
rect 43194 7540 43234 7580
rect 43276 7540 43316 7580
rect 43358 7540 43398 7580
rect 43440 7540 43480 7580
rect 47112 7540 47152 7580
rect 47194 7540 47234 7580
rect 47276 7540 47316 7580
rect 47358 7540 47398 7580
rect 47440 7540 47480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 55112 7540 55152 7580
rect 55194 7540 55234 7580
rect 55276 7540 55316 7580
rect 55358 7540 55398 7580
rect 55440 7540 55480 7580
rect 59112 7540 59152 7580
rect 59194 7540 59234 7580
rect 59276 7540 59316 7580
rect 59358 7540 59398 7580
rect 59440 7540 59480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 67112 7540 67152 7580
rect 67194 7540 67234 7580
rect 67276 7540 67316 7580
rect 67358 7540 67398 7580
rect 67440 7540 67480 7580
rect 71112 7540 71152 7580
rect 71194 7540 71234 7580
rect 71276 7540 71316 7580
rect 71358 7540 71398 7580
rect 71440 7540 71480 7580
rect 75112 7540 75152 7580
rect 75194 7540 75234 7580
rect 75276 7540 75316 7580
rect 75358 7540 75398 7580
rect 75440 7540 75480 7580
rect 79112 7540 79152 7580
rect 79194 7540 79234 7580
rect 79276 7540 79316 7580
rect 79358 7540 79398 7580
rect 79440 7540 79480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 8352 6784 8392 6824
rect 8434 6784 8474 6824
rect 8516 6784 8556 6824
rect 8598 6784 8638 6824
rect 8680 6784 8720 6824
rect 12352 6784 12392 6824
rect 12434 6784 12474 6824
rect 12516 6784 12556 6824
rect 12598 6784 12638 6824
rect 12680 6784 12720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 20352 6784 20392 6824
rect 20434 6784 20474 6824
rect 20516 6784 20556 6824
rect 20598 6784 20638 6824
rect 20680 6784 20720 6824
rect 24352 6784 24392 6824
rect 24434 6784 24474 6824
rect 24516 6784 24556 6824
rect 24598 6784 24638 6824
rect 24680 6784 24720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 32352 6784 32392 6824
rect 32434 6784 32474 6824
rect 32516 6784 32556 6824
rect 32598 6784 32638 6824
rect 32680 6784 32720 6824
rect 36352 6784 36392 6824
rect 36434 6784 36474 6824
rect 36516 6784 36556 6824
rect 36598 6784 36638 6824
rect 36680 6784 36720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 44352 6784 44392 6824
rect 44434 6784 44474 6824
rect 44516 6784 44556 6824
rect 44598 6784 44638 6824
rect 44680 6784 44720 6824
rect 48352 6784 48392 6824
rect 48434 6784 48474 6824
rect 48516 6784 48556 6824
rect 48598 6784 48638 6824
rect 48680 6784 48720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 56352 6784 56392 6824
rect 56434 6784 56474 6824
rect 56516 6784 56556 6824
rect 56598 6784 56638 6824
rect 56680 6784 56720 6824
rect 60352 6784 60392 6824
rect 60434 6784 60474 6824
rect 60516 6784 60556 6824
rect 60598 6784 60638 6824
rect 60680 6784 60720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 68352 6784 68392 6824
rect 68434 6784 68474 6824
rect 68516 6784 68556 6824
rect 68598 6784 68638 6824
rect 68680 6784 68720 6824
rect 72352 6784 72392 6824
rect 72434 6784 72474 6824
rect 72516 6784 72556 6824
rect 72598 6784 72638 6824
rect 72680 6784 72720 6824
rect 76352 6784 76392 6824
rect 76434 6784 76474 6824
rect 76516 6784 76556 6824
rect 76598 6784 76638 6824
rect 76680 6784 76720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 7112 6028 7152 6068
rect 7194 6028 7234 6068
rect 7276 6028 7316 6068
rect 7358 6028 7398 6068
rect 7440 6028 7480 6068
rect 11112 6028 11152 6068
rect 11194 6028 11234 6068
rect 11276 6028 11316 6068
rect 11358 6028 11398 6068
rect 11440 6028 11480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 19112 6028 19152 6068
rect 19194 6028 19234 6068
rect 19276 6028 19316 6068
rect 19358 6028 19398 6068
rect 19440 6028 19480 6068
rect 23112 6028 23152 6068
rect 23194 6028 23234 6068
rect 23276 6028 23316 6068
rect 23358 6028 23398 6068
rect 23440 6028 23480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 31112 6028 31152 6068
rect 31194 6028 31234 6068
rect 31276 6028 31316 6068
rect 31358 6028 31398 6068
rect 31440 6028 31480 6068
rect 35112 6028 35152 6068
rect 35194 6028 35234 6068
rect 35276 6028 35316 6068
rect 35358 6028 35398 6068
rect 35440 6028 35480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 43112 6028 43152 6068
rect 43194 6028 43234 6068
rect 43276 6028 43316 6068
rect 43358 6028 43398 6068
rect 43440 6028 43480 6068
rect 47112 6028 47152 6068
rect 47194 6028 47234 6068
rect 47276 6028 47316 6068
rect 47358 6028 47398 6068
rect 47440 6028 47480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 55112 6028 55152 6068
rect 55194 6028 55234 6068
rect 55276 6028 55316 6068
rect 55358 6028 55398 6068
rect 55440 6028 55480 6068
rect 59112 6028 59152 6068
rect 59194 6028 59234 6068
rect 59276 6028 59316 6068
rect 59358 6028 59398 6068
rect 59440 6028 59480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 67112 6028 67152 6068
rect 67194 6028 67234 6068
rect 67276 6028 67316 6068
rect 67358 6028 67398 6068
rect 67440 6028 67480 6068
rect 71112 6028 71152 6068
rect 71194 6028 71234 6068
rect 71276 6028 71316 6068
rect 71358 6028 71398 6068
rect 71440 6028 71480 6068
rect 75112 6028 75152 6068
rect 75194 6028 75234 6068
rect 75276 6028 75316 6068
rect 75358 6028 75398 6068
rect 75440 6028 75480 6068
rect 79112 6028 79152 6068
rect 79194 6028 79234 6068
rect 79276 6028 79316 6068
rect 79358 6028 79398 6068
rect 79440 6028 79480 6068
rect 83112 7540 83152 7580
rect 83194 7540 83234 7580
rect 83276 7540 83316 7580
rect 83358 7540 83398 7580
rect 83440 7540 83480 7580
rect 80352 6784 80392 6824
rect 80434 6784 80474 6824
rect 80516 6784 80556 6824
rect 80598 6784 80638 6824
rect 80680 6784 80720 6824
rect 83112 6028 83152 6068
rect 83194 6028 83234 6068
rect 83276 6028 83316 6068
rect 83358 6028 83398 6068
rect 83440 6028 83480 6068
rect 84352 6784 84392 6824
rect 84434 6784 84474 6824
rect 84516 6784 84556 6824
rect 84598 6784 84638 6824
rect 84680 6784 84720 6824
rect 87112 7540 87152 7580
rect 87194 7540 87234 7580
rect 87276 7540 87316 7580
rect 87358 7540 87398 7580
rect 87440 7540 87480 7580
rect 86668 7372 86708 7412
rect 88352 6784 88392 6824
rect 88434 6784 88474 6824
rect 88516 6784 88556 6824
rect 88598 6784 88638 6824
rect 88680 6784 88720 6824
rect 87112 6028 87152 6068
rect 87194 6028 87234 6068
rect 87276 6028 87316 6068
rect 87358 6028 87398 6068
rect 87440 6028 87480 6068
rect 91112 7540 91152 7580
rect 91194 7540 91234 7580
rect 91276 7540 91316 7580
rect 91358 7540 91398 7580
rect 91440 7540 91480 7580
rect 95112 7540 95152 7580
rect 95194 7540 95234 7580
rect 95276 7540 95316 7580
rect 95358 7540 95398 7580
rect 95440 7540 95480 7580
rect 92352 6784 92392 6824
rect 92434 6784 92474 6824
rect 92516 6784 92556 6824
rect 92598 6784 92638 6824
rect 92680 6784 92720 6824
rect 99112 7540 99152 7580
rect 99194 7540 99234 7580
rect 99276 7540 99316 7580
rect 99358 7540 99398 7580
rect 99440 7540 99480 7580
rect 96352 6784 96392 6824
rect 96434 6784 96474 6824
rect 96516 6784 96556 6824
rect 96598 6784 96638 6824
rect 96680 6784 96720 6824
rect 91112 6028 91152 6068
rect 91194 6028 91234 6068
rect 91276 6028 91316 6068
rect 91358 6028 91398 6068
rect 91440 6028 91480 6068
rect 95112 6028 95152 6068
rect 95194 6028 95234 6068
rect 95276 6028 95316 6068
rect 95358 6028 95398 6068
rect 95440 6028 95480 6068
rect 99112 6028 99152 6068
rect 99194 6028 99234 6068
rect 99276 6028 99316 6068
rect 99358 6028 99398 6068
rect 99440 6028 99480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 8352 5272 8392 5312
rect 8434 5272 8474 5312
rect 8516 5272 8556 5312
rect 8598 5272 8638 5312
rect 8680 5272 8720 5312
rect 12352 5272 12392 5312
rect 12434 5272 12474 5312
rect 12516 5272 12556 5312
rect 12598 5272 12638 5312
rect 12680 5272 12720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 20352 5272 20392 5312
rect 20434 5272 20474 5312
rect 20516 5272 20556 5312
rect 20598 5272 20638 5312
rect 20680 5272 20720 5312
rect 24352 5272 24392 5312
rect 24434 5272 24474 5312
rect 24516 5272 24556 5312
rect 24598 5272 24638 5312
rect 24680 5272 24720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 32352 5272 32392 5312
rect 32434 5272 32474 5312
rect 32516 5272 32556 5312
rect 32598 5272 32638 5312
rect 32680 5272 32720 5312
rect 36352 5272 36392 5312
rect 36434 5272 36474 5312
rect 36516 5272 36556 5312
rect 36598 5272 36638 5312
rect 36680 5272 36720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 44352 5272 44392 5312
rect 44434 5272 44474 5312
rect 44516 5272 44556 5312
rect 44598 5272 44638 5312
rect 44680 5272 44720 5312
rect 48352 5272 48392 5312
rect 48434 5272 48474 5312
rect 48516 5272 48556 5312
rect 48598 5272 48638 5312
rect 48680 5272 48720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 56352 5272 56392 5312
rect 56434 5272 56474 5312
rect 56516 5272 56556 5312
rect 56598 5272 56638 5312
rect 56680 5272 56720 5312
rect 60352 5272 60392 5312
rect 60434 5272 60474 5312
rect 60516 5272 60556 5312
rect 60598 5272 60638 5312
rect 60680 5272 60720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 68352 5272 68392 5312
rect 68434 5272 68474 5312
rect 68516 5272 68556 5312
rect 68598 5272 68638 5312
rect 68680 5272 68720 5312
rect 72352 5272 72392 5312
rect 72434 5272 72474 5312
rect 72516 5272 72556 5312
rect 72598 5272 72638 5312
rect 72680 5272 72720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 80352 5272 80392 5312
rect 80434 5272 80474 5312
rect 80516 5272 80556 5312
rect 80598 5272 80638 5312
rect 80680 5272 80720 5312
rect 84352 5272 84392 5312
rect 84434 5272 84474 5312
rect 84516 5272 84556 5312
rect 84598 5272 84638 5312
rect 84680 5272 84720 5312
rect 88352 5272 88392 5312
rect 88434 5272 88474 5312
rect 88516 5272 88556 5312
rect 88598 5272 88638 5312
rect 88680 5272 88720 5312
rect 92352 5272 92392 5312
rect 92434 5272 92474 5312
rect 92516 5272 92556 5312
rect 92598 5272 92638 5312
rect 92680 5272 92720 5312
rect 96352 5272 96392 5312
rect 96434 5272 96474 5312
rect 96516 5272 96556 5312
rect 96598 5272 96638 5312
rect 96680 5272 96720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 7112 4516 7152 4556
rect 7194 4516 7234 4556
rect 7276 4516 7316 4556
rect 7358 4516 7398 4556
rect 7440 4516 7480 4556
rect 11112 4516 11152 4556
rect 11194 4516 11234 4556
rect 11276 4516 11316 4556
rect 11358 4516 11398 4556
rect 11440 4516 11480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 19112 4516 19152 4556
rect 19194 4516 19234 4556
rect 19276 4516 19316 4556
rect 19358 4516 19398 4556
rect 19440 4516 19480 4556
rect 23112 4516 23152 4556
rect 23194 4516 23234 4556
rect 23276 4516 23316 4556
rect 23358 4516 23398 4556
rect 23440 4516 23480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 31112 4516 31152 4556
rect 31194 4516 31234 4556
rect 31276 4516 31316 4556
rect 31358 4516 31398 4556
rect 31440 4516 31480 4556
rect 35112 4516 35152 4556
rect 35194 4516 35234 4556
rect 35276 4516 35316 4556
rect 35358 4516 35398 4556
rect 35440 4516 35480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 43112 4516 43152 4556
rect 43194 4516 43234 4556
rect 43276 4516 43316 4556
rect 43358 4516 43398 4556
rect 43440 4516 43480 4556
rect 47112 4516 47152 4556
rect 47194 4516 47234 4556
rect 47276 4516 47316 4556
rect 47358 4516 47398 4556
rect 47440 4516 47480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 55112 4516 55152 4556
rect 55194 4516 55234 4556
rect 55276 4516 55316 4556
rect 55358 4516 55398 4556
rect 55440 4516 55480 4556
rect 59112 4516 59152 4556
rect 59194 4516 59234 4556
rect 59276 4516 59316 4556
rect 59358 4516 59398 4556
rect 59440 4516 59480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 67112 4516 67152 4556
rect 67194 4516 67234 4556
rect 67276 4516 67316 4556
rect 67358 4516 67398 4556
rect 67440 4516 67480 4556
rect 71112 4516 71152 4556
rect 71194 4516 71234 4556
rect 71276 4516 71316 4556
rect 71358 4516 71398 4556
rect 71440 4516 71480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 79112 4516 79152 4556
rect 79194 4516 79234 4556
rect 79276 4516 79316 4556
rect 79358 4516 79398 4556
rect 79440 4516 79480 4556
rect 83112 4516 83152 4556
rect 83194 4516 83234 4556
rect 83276 4516 83316 4556
rect 83358 4516 83398 4556
rect 83440 4516 83480 4556
rect 87112 4516 87152 4556
rect 87194 4516 87234 4556
rect 87276 4516 87316 4556
rect 87358 4516 87398 4556
rect 87440 4516 87480 4556
rect 91112 4516 91152 4556
rect 91194 4516 91234 4556
rect 91276 4516 91316 4556
rect 91358 4516 91398 4556
rect 91440 4516 91480 4556
rect 95112 4516 95152 4556
rect 95194 4516 95234 4556
rect 95276 4516 95316 4556
rect 95358 4516 95398 4556
rect 95440 4516 95480 4556
rect 99112 4516 99152 4556
rect 99194 4516 99234 4556
rect 99276 4516 99316 4556
rect 99358 4516 99398 4556
rect 99440 4516 99480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 8352 3760 8392 3800
rect 8434 3760 8474 3800
rect 8516 3760 8556 3800
rect 8598 3760 8638 3800
rect 8680 3760 8720 3800
rect 12352 3760 12392 3800
rect 12434 3760 12474 3800
rect 12516 3760 12556 3800
rect 12598 3760 12638 3800
rect 12680 3760 12720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 20352 3760 20392 3800
rect 20434 3760 20474 3800
rect 20516 3760 20556 3800
rect 20598 3760 20638 3800
rect 20680 3760 20720 3800
rect 24352 3760 24392 3800
rect 24434 3760 24474 3800
rect 24516 3760 24556 3800
rect 24598 3760 24638 3800
rect 24680 3760 24720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 32352 3760 32392 3800
rect 32434 3760 32474 3800
rect 32516 3760 32556 3800
rect 32598 3760 32638 3800
rect 32680 3760 32720 3800
rect 36352 3760 36392 3800
rect 36434 3760 36474 3800
rect 36516 3760 36556 3800
rect 36598 3760 36638 3800
rect 36680 3760 36720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 44352 3760 44392 3800
rect 44434 3760 44474 3800
rect 44516 3760 44556 3800
rect 44598 3760 44638 3800
rect 44680 3760 44720 3800
rect 48352 3760 48392 3800
rect 48434 3760 48474 3800
rect 48516 3760 48556 3800
rect 48598 3760 48638 3800
rect 48680 3760 48720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 56352 3760 56392 3800
rect 56434 3760 56474 3800
rect 56516 3760 56556 3800
rect 56598 3760 56638 3800
rect 56680 3760 56720 3800
rect 60352 3760 60392 3800
rect 60434 3760 60474 3800
rect 60516 3760 60556 3800
rect 60598 3760 60638 3800
rect 60680 3760 60720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 68352 3760 68392 3800
rect 68434 3760 68474 3800
rect 68516 3760 68556 3800
rect 68598 3760 68638 3800
rect 68680 3760 68720 3800
rect 72352 3760 72392 3800
rect 72434 3760 72474 3800
rect 72516 3760 72556 3800
rect 72598 3760 72638 3800
rect 72680 3760 72720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 80352 3760 80392 3800
rect 80434 3760 80474 3800
rect 80516 3760 80556 3800
rect 80598 3760 80638 3800
rect 80680 3760 80720 3800
rect 84352 3760 84392 3800
rect 84434 3760 84474 3800
rect 84516 3760 84556 3800
rect 84598 3760 84638 3800
rect 84680 3760 84720 3800
rect 88352 3760 88392 3800
rect 88434 3760 88474 3800
rect 88516 3760 88556 3800
rect 88598 3760 88638 3800
rect 88680 3760 88720 3800
rect 92352 3760 92392 3800
rect 92434 3760 92474 3800
rect 92516 3760 92556 3800
rect 92598 3760 92638 3800
rect 92680 3760 92720 3800
rect 96352 3760 96392 3800
rect 96434 3760 96474 3800
rect 96516 3760 96556 3800
rect 96598 3760 96638 3800
rect 96680 3760 96720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 7112 3004 7152 3044
rect 7194 3004 7234 3044
rect 7276 3004 7316 3044
rect 7358 3004 7398 3044
rect 7440 3004 7480 3044
rect 11112 3004 11152 3044
rect 11194 3004 11234 3044
rect 11276 3004 11316 3044
rect 11358 3004 11398 3044
rect 11440 3004 11480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 19112 3004 19152 3044
rect 19194 3004 19234 3044
rect 19276 3004 19316 3044
rect 19358 3004 19398 3044
rect 19440 3004 19480 3044
rect 23112 3004 23152 3044
rect 23194 3004 23234 3044
rect 23276 3004 23316 3044
rect 23358 3004 23398 3044
rect 23440 3004 23480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 31112 3004 31152 3044
rect 31194 3004 31234 3044
rect 31276 3004 31316 3044
rect 31358 3004 31398 3044
rect 31440 3004 31480 3044
rect 35112 3004 35152 3044
rect 35194 3004 35234 3044
rect 35276 3004 35316 3044
rect 35358 3004 35398 3044
rect 35440 3004 35480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 43112 3004 43152 3044
rect 43194 3004 43234 3044
rect 43276 3004 43316 3044
rect 43358 3004 43398 3044
rect 43440 3004 43480 3044
rect 47112 3004 47152 3044
rect 47194 3004 47234 3044
rect 47276 3004 47316 3044
rect 47358 3004 47398 3044
rect 47440 3004 47480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 55112 3004 55152 3044
rect 55194 3004 55234 3044
rect 55276 3004 55316 3044
rect 55358 3004 55398 3044
rect 55440 3004 55480 3044
rect 59112 3004 59152 3044
rect 59194 3004 59234 3044
rect 59276 3004 59316 3044
rect 59358 3004 59398 3044
rect 59440 3004 59480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 67112 3004 67152 3044
rect 67194 3004 67234 3044
rect 67276 3004 67316 3044
rect 67358 3004 67398 3044
rect 67440 3004 67480 3044
rect 71112 3004 71152 3044
rect 71194 3004 71234 3044
rect 71276 3004 71316 3044
rect 71358 3004 71398 3044
rect 71440 3004 71480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 79112 3004 79152 3044
rect 79194 3004 79234 3044
rect 79276 3004 79316 3044
rect 79358 3004 79398 3044
rect 79440 3004 79480 3044
rect 83112 3004 83152 3044
rect 83194 3004 83234 3044
rect 83276 3004 83316 3044
rect 83358 3004 83398 3044
rect 83440 3004 83480 3044
rect 87112 3004 87152 3044
rect 87194 3004 87234 3044
rect 87276 3004 87316 3044
rect 87358 3004 87398 3044
rect 87440 3004 87480 3044
rect 91112 3004 91152 3044
rect 91194 3004 91234 3044
rect 91276 3004 91316 3044
rect 91358 3004 91398 3044
rect 91440 3004 91480 3044
rect 95112 3004 95152 3044
rect 95194 3004 95234 3044
rect 95276 3004 95316 3044
rect 95358 3004 95398 3044
rect 95440 3004 95480 3044
rect 99112 3004 99152 3044
rect 99194 3004 99234 3044
rect 99276 3004 99316 3044
rect 99358 3004 99398 3044
rect 99440 3004 99480 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 8352 2248 8392 2288
rect 8434 2248 8474 2288
rect 8516 2248 8556 2288
rect 8598 2248 8638 2288
rect 8680 2248 8720 2288
rect 12352 2248 12392 2288
rect 12434 2248 12474 2288
rect 12516 2248 12556 2288
rect 12598 2248 12638 2288
rect 12680 2248 12720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 20352 2248 20392 2288
rect 20434 2248 20474 2288
rect 20516 2248 20556 2288
rect 20598 2248 20638 2288
rect 20680 2248 20720 2288
rect 24352 2248 24392 2288
rect 24434 2248 24474 2288
rect 24516 2248 24556 2288
rect 24598 2248 24638 2288
rect 24680 2248 24720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 32352 2248 32392 2288
rect 32434 2248 32474 2288
rect 32516 2248 32556 2288
rect 32598 2248 32638 2288
rect 32680 2248 32720 2288
rect 36352 2248 36392 2288
rect 36434 2248 36474 2288
rect 36516 2248 36556 2288
rect 36598 2248 36638 2288
rect 36680 2248 36720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 44352 2248 44392 2288
rect 44434 2248 44474 2288
rect 44516 2248 44556 2288
rect 44598 2248 44638 2288
rect 44680 2248 44720 2288
rect 48352 2248 48392 2288
rect 48434 2248 48474 2288
rect 48516 2248 48556 2288
rect 48598 2248 48638 2288
rect 48680 2248 48720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 56352 2248 56392 2288
rect 56434 2248 56474 2288
rect 56516 2248 56556 2288
rect 56598 2248 56638 2288
rect 56680 2248 56720 2288
rect 60352 2248 60392 2288
rect 60434 2248 60474 2288
rect 60516 2248 60556 2288
rect 60598 2248 60638 2288
rect 60680 2248 60720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 68352 2248 68392 2288
rect 68434 2248 68474 2288
rect 68516 2248 68556 2288
rect 68598 2248 68638 2288
rect 68680 2248 68720 2288
rect 72352 2248 72392 2288
rect 72434 2248 72474 2288
rect 72516 2248 72556 2288
rect 72598 2248 72638 2288
rect 72680 2248 72720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 80352 2248 80392 2288
rect 80434 2248 80474 2288
rect 80516 2248 80556 2288
rect 80598 2248 80638 2288
rect 80680 2248 80720 2288
rect 84352 2248 84392 2288
rect 84434 2248 84474 2288
rect 84516 2248 84556 2288
rect 84598 2248 84638 2288
rect 84680 2248 84720 2288
rect 88352 2248 88392 2288
rect 88434 2248 88474 2288
rect 88516 2248 88556 2288
rect 88598 2248 88638 2288
rect 88680 2248 88720 2288
rect 92352 2248 92392 2288
rect 92434 2248 92474 2288
rect 92516 2248 92556 2288
rect 92598 2248 92638 2288
rect 92680 2248 92720 2288
rect 96352 2248 96392 2288
rect 96434 2248 96474 2288
rect 96516 2248 96556 2288
rect 96598 2248 96638 2288
rect 96680 2248 96720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 7112 1492 7152 1532
rect 7194 1492 7234 1532
rect 7276 1492 7316 1532
rect 7358 1492 7398 1532
rect 7440 1492 7480 1532
rect 11112 1492 11152 1532
rect 11194 1492 11234 1532
rect 11276 1492 11316 1532
rect 11358 1492 11398 1532
rect 11440 1492 11480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 19112 1492 19152 1532
rect 19194 1492 19234 1532
rect 19276 1492 19316 1532
rect 19358 1492 19398 1532
rect 19440 1492 19480 1532
rect 23112 1492 23152 1532
rect 23194 1492 23234 1532
rect 23276 1492 23316 1532
rect 23358 1492 23398 1532
rect 23440 1492 23480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 31112 1492 31152 1532
rect 31194 1492 31234 1532
rect 31276 1492 31316 1532
rect 31358 1492 31398 1532
rect 31440 1492 31480 1532
rect 35112 1492 35152 1532
rect 35194 1492 35234 1532
rect 35276 1492 35316 1532
rect 35358 1492 35398 1532
rect 35440 1492 35480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 43112 1492 43152 1532
rect 43194 1492 43234 1532
rect 43276 1492 43316 1532
rect 43358 1492 43398 1532
rect 43440 1492 43480 1532
rect 47112 1492 47152 1532
rect 47194 1492 47234 1532
rect 47276 1492 47316 1532
rect 47358 1492 47398 1532
rect 47440 1492 47480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 55112 1492 55152 1532
rect 55194 1492 55234 1532
rect 55276 1492 55316 1532
rect 55358 1492 55398 1532
rect 55440 1492 55480 1532
rect 59112 1492 59152 1532
rect 59194 1492 59234 1532
rect 59276 1492 59316 1532
rect 59358 1492 59398 1532
rect 59440 1492 59480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 67112 1492 67152 1532
rect 67194 1492 67234 1532
rect 67276 1492 67316 1532
rect 67358 1492 67398 1532
rect 67440 1492 67480 1532
rect 71112 1492 71152 1532
rect 71194 1492 71234 1532
rect 71276 1492 71316 1532
rect 71358 1492 71398 1532
rect 71440 1492 71480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 79112 1492 79152 1532
rect 79194 1492 79234 1532
rect 79276 1492 79316 1532
rect 79358 1492 79398 1532
rect 79440 1492 79480 1532
rect 83112 1492 83152 1532
rect 83194 1492 83234 1532
rect 83276 1492 83316 1532
rect 83358 1492 83398 1532
rect 83440 1492 83480 1532
rect 87112 1492 87152 1532
rect 87194 1492 87234 1532
rect 87276 1492 87316 1532
rect 87358 1492 87398 1532
rect 87440 1492 87480 1532
rect 91112 1492 91152 1532
rect 91194 1492 91234 1532
rect 91276 1492 91316 1532
rect 91358 1492 91398 1532
rect 91440 1492 91480 1532
rect 95112 1492 95152 1532
rect 95194 1492 95234 1532
rect 95276 1492 95316 1532
rect 95358 1492 95398 1532
rect 95440 1492 95480 1532
rect 99112 1492 99152 1532
rect 99194 1492 99234 1532
rect 99276 1492 99316 1532
rect 99358 1492 99398 1532
rect 99440 1492 99480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 8352 736 8392 776
rect 8434 736 8474 776
rect 8516 736 8556 776
rect 8598 736 8638 776
rect 8680 736 8720 776
rect 12352 736 12392 776
rect 12434 736 12474 776
rect 12516 736 12556 776
rect 12598 736 12638 776
rect 12680 736 12720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 20352 736 20392 776
rect 20434 736 20474 776
rect 20516 736 20556 776
rect 20598 736 20638 776
rect 20680 736 20720 776
rect 24352 736 24392 776
rect 24434 736 24474 776
rect 24516 736 24556 776
rect 24598 736 24638 776
rect 24680 736 24720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 32352 736 32392 776
rect 32434 736 32474 776
rect 32516 736 32556 776
rect 32598 736 32638 776
rect 32680 736 32720 776
rect 36352 736 36392 776
rect 36434 736 36474 776
rect 36516 736 36556 776
rect 36598 736 36638 776
rect 36680 736 36720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 44352 736 44392 776
rect 44434 736 44474 776
rect 44516 736 44556 776
rect 44598 736 44638 776
rect 44680 736 44720 776
rect 48352 736 48392 776
rect 48434 736 48474 776
rect 48516 736 48556 776
rect 48598 736 48638 776
rect 48680 736 48720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 56352 736 56392 776
rect 56434 736 56474 776
rect 56516 736 56556 776
rect 56598 736 56638 776
rect 56680 736 56720 776
rect 60352 736 60392 776
rect 60434 736 60474 776
rect 60516 736 60556 776
rect 60598 736 60638 776
rect 60680 736 60720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 68352 736 68392 776
rect 68434 736 68474 776
rect 68516 736 68556 776
rect 68598 736 68638 776
rect 68680 736 68720 776
rect 72352 736 72392 776
rect 72434 736 72474 776
rect 72516 736 72556 776
rect 72598 736 72638 776
rect 72680 736 72720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
rect 80352 736 80392 776
rect 80434 736 80474 776
rect 80516 736 80556 776
rect 80598 736 80638 776
rect 80680 736 80720 776
rect 84352 736 84392 776
rect 84434 736 84474 776
rect 84516 736 84556 776
rect 84598 736 84638 776
rect 84680 736 84720 776
rect 88352 736 88392 776
rect 88434 736 88474 776
rect 88516 736 88556 776
rect 88598 736 88638 776
rect 88680 736 88720 776
rect 92352 736 92392 776
rect 92434 736 92474 776
rect 92516 736 92556 776
rect 92598 736 92638 776
rect 92680 736 92720 776
rect 96352 736 96392 776
rect 96434 736 96474 776
rect 96516 736 96556 776
rect 96598 736 96638 776
rect 96680 736 96720 776
<< metal5 >>
rect 4343 38599 4729 38618
rect 4343 38576 4409 38599
rect 4495 38576 4577 38599
rect 4663 38576 4729 38599
rect 4343 38536 4352 38576
rect 4392 38536 4409 38576
rect 4495 38536 4516 38576
rect 4556 38536 4577 38576
rect 4663 38536 4680 38576
rect 4720 38536 4729 38576
rect 4343 38513 4409 38536
rect 4495 38513 4577 38536
rect 4663 38513 4729 38536
rect 4343 38494 4729 38513
rect 8343 38599 8729 38618
rect 8343 38576 8409 38599
rect 8495 38576 8577 38599
rect 8663 38576 8729 38599
rect 8343 38536 8352 38576
rect 8392 38536 8409 38576
rect 8495 38536 8516 38576
rect 8556 38536 8577 38576
rect 8663 38536 8680 38576
rect 8720 38536 8729 38576
rect 8343 38513 8409 38536
rect 8495 38513 8577 38536
rect 8663 38513 8729 38536
rect 8343 38494 8729 38513
rect 12343 38599 12729 38618
rect 12343 38576 12409 38599
rect 12495 38576 12577 38599
rect 12663 38576 12729 38599
rect 12343 38536 12352 38576
rect 12392 38536 12409 38576
rect 12495 38536 12516 38576
rect 12556 38536 12577 38576
rect 12663 38536 12680 38576
rect 12720 38536 12729 38576
rect 12343 38513 12409 38536
rect 12495 38513 12577 38536
rect 12663 38513 12729 38536
rect 12343 38494 12729 38513
rect 16343 38599 16729 38618
rect 16343 38576 16409 38599
rect 16495 38576 16577 38599
rect 16663 38576 16729 38599
rect 16343 38536 16352 38576
rect 16392 38536 16409 38576
rect 16495 38536 16516 38576
rect 16556 38536 16577 38576
rect 16663 38536 16680 38576
rect 16720 38536 16729 38576
rect 16343 38513 16409 38536
rect 16495 38513 16577 38536
rect 16663 38513 16729 38536
rect 16343 38494 16729 38513
rect 20343 38599 20729 38618
rect 20343 38576 20409 38599
rect 20495 38576 20577 38599
rect 20663 38576 20729 38599
rect 20343 38536 20352 38576
rect 20392 38536 20409 38576
rect 20495 38536 20516 38576
rect 20556 38536 20577 38576
rect 20663 38536 20680 38576
rect 20720 38536 20729 38576
rect 20343 38513 20409 38536
rect 20495 38513 20577 38536
rect 20663 38513 20729 38536
rect 20343 38494 20729 38513
rect 24343 38599 24729 38618
rect 24343 38576 24409 38599
rect 24495 38576 24577 38599
rect 24663 38576 24729 38599
rect 24343 38536 24352 38576
rect 24392 38536 24409 38576
rect 24495 38536 24516 38576
rect 24556 38536 24577 38576
rect 24663 38536 24680 38576
rect 24720 38536 24729 38576
rect 24343 38513 24409 38536
rect 24495 38513 24577 38536
rect 24663 38513 24729 38536
rect 24343 38494 24729 38513
rect 28343 38599 28729 38618
rect 28343 38576 28409 38599
rect 28495 38576 28577 38599
rect 28663 38576 28729 38599
rect 28343 38536 28352 38576
rect 28392 38536 28409 38576
rect 28495 38536 28516 38576
rect 28556 38536 28577 38576
rect 28663 38536 28680 38576
rect 28720 38536 28729 38576
rect 28343 38513 28409 38536
rect 28495 38513 28577 38536
rect 28663 38513 28729 38536
rect 28343 38494 28729 38513
rect 32343 38599 32729 38618
rect 32343 38576 32409 38599
rect 32495 38576 32577 38599
rect 32663 38576 32729 38599
rect 32343 38536 32352 38576
rect 32392 38536 32409 38576
rect 32495 38536 32516 38576
rect 32556 38536 32577 38576
rect 32663 38536 32680 38576
rect 32720 38536 32729 38576
rect 32343 38513 32409 38536
rect 32495 38513 32577 38536
rect 32663 38513 32729 38536
rect 32343 38494 32729 38513
rect 36343 38599 36729 38618
rect 36343 38576 36409 38599
rect 36495 38576 36577 38599
rect 36663 38576 36729 38599
rect 36343 38536 36352 38576
rect 36392 38536 36409 38576
rect 36495 38536 36516 38576
rect 36556 38536 36577 38576
rect 36663 38536 36680 38576
rect 36720 38536 36729 38576
rect 36343 38513 36409 38536
rect 36495 38513 36577 38536
rect 36663 38513 36729 38536
rect 36343 38494 36729 38513
rect 40343 38599 40729 38618
rect 40343 38576 40409 38599
rect 40495 38576 40577 38599
rect 40663 38576 40729 38599
rect 40343 38536 40352 38576
rect 40392 38536 40409 38576
rect 40495 38536 40516 38576
rect 40556 38536 40577 38576
rect 40663 38536 40680 38576
rect 40720 38536 40729 38576
rect 40343 38513 40409 38536
rect 40495 38513 40577 38536
rect 40663 38513 40729 38536
rect 40343 38494 40729 38513
rect 44343 38599 44729 38618
rect 44343 38576 44409 38599
rect 44495 38576 44577 38599
rect 44663 38576 44729 38599
rect 44343 38536 44352 38576
rect 44392 38536 44409 38576
rect 44495 38536 44516 38576
rect 44556 38536 44577 38576
rect 44663 38536 44680 38576
rect 44720 38536 44729 38576
rect 44343 38513 44409 38536
rect 44495 38513 44577 38536
rect 44663 38513 44729 38536
rect 44343 38494 44729 38513
rect 48343 38599 48729 38618
rect 48343 38576 48409 38599
rect 48495 38576 48577 38599
rect 48663 38576 48729 38599
rect 48343 38536 48352 38576
rect 48392 38536 48409 38576
rect 48495 38536 48516 38576
rect 48556 38536 48577 38576
rect 48663 38536 48680 38576
rect 48720 38536 48729 38576
rect 48343 38513 48409 38536
rect 48495 38513 48577 38536
rect 48663 38513 48729 38536
rect 48343 38494 48729 38513
rect 52343 38599 52729 38618
rect 52343 38576 52409 38599
rect 52495 38576 52577 38599
rect 52663 38576 52729 38599
rect 52343 38536 52352 38576
rect 52392 38536 52409 38576
rect 52495 38536 52516 38576
rect 52556 38536 52577 38576
rect 52663 38536 52680 38576
rect 52720 38536 52729 38576
rect 52343 38513 52409 38536
rect 52495 38513 52577 38536
rect 52663 38513 52729 38536
rect 52343 38494 52729 38513
rect 56343 38599 56729 38618
rect 56343 38576 56409 38599
rect 56495 38576 56577 38599
rect 56663 38576 56729 38599
rect 56343 38536 56352 38576
rect 56392 38536 56409 38576
rect 56495 38536 56516 38576
rect 56556 38536 56577 38576
rect 56663 38536 56680 38576
rect 56720 38536 56729 38576
rect 56343 38513 56409 38536
rect 56495 38513 56577 38536
rect 56663 38513 56729 38536
rect 56343 38494 56729 38513
rect 60343 38599 60729 38618
rect 60343 38576 60409 38599
rect 60495 38576 60577 38599
rect 60663 38576 60729 38599
rect 60343 38536 60352 38576
rect 60392 38536 60409 38576
rect 60495 38536 60516 38576
rect 60556 38536 60577 38576
rect 60663 38536 60680 38576
rect 60720 38536 60729 38576
rect 60343 38513 60409 38536
rect 60495 38513 60577 38536
rect 60663 38513 60729 38536
rect 60343 38494 60729 38513
rect 64343 38599 64729 38618
rect 64343 38576 64409 38599
rect 64495 38576 64577 38599
rect 64663 38576 64729 38599
rect 64343 38536 64352 38576
rect 64392 38536 64409 38576
rect 64495 38536 64516 38576
rect 64556 38536 64577 38576
rect 64663 38536 64680 38576
rect 64720 38536 64729 38576
rect 64343 38513 64409 38536
rect 64495 38513 64577 38536
rect 64663 38513 64729 38536
rect 64343 38494 64729 38513
rect 68343 38599 68729 38618
rect 68343 38576 68409 38599
rect 68495 38576 68577 38599
rect 68663 38576 68729 38599
rect 68343 38536 68352 38576
rect 68392 38536 68409 38576
rect 68495 38536 68516 38576
rect 68556 38536 68577 38576
rect 68663 38536 68680 38576
rect 68720 38536 68729 38576
rect 68343 38513 68409 38536
rect 68495 38513 68577 38536
rect 68663 38513 68729 38536
rect 68343 38494 68729 38513
rect 72343 38599 72729 38618
rect 72343 38576 72409 38599
rect 72495 38576 72577 38599
rect 72663 38576 72729 38599
rect 72343 38536 72352 38576
rect 72392 38536 72409 38576
rect 72495 38536 72516 38576
rect 72556 38536 72577 38576
rect 72663 38536 72680 38576
rect 72720 38536 72729 38576
rect 72343 38513 72409 38536
rect 72495 38513 72577 38536
rect 72663 38513 72729 38536
rect 72343 38494 72729 38513
rect 76343 38599 76729 38618
rect 76343 38576 76409 38599
rect 76495 38576 76577 38599
rect 76663 38576 76729 38599
rect 76343 38536 76352 38576
rect 76392 38536 76409 38576
rect 76495 38536 76516 38576
rect 76556 38536 76577 38576
rect 76663 38536 76680 38576
rect 76720 38536 76729 38576
rect 76343 38513 76409 38536
rect 76495 38513 76577 38536
rect 76663 38513 76729 38536
rect 76343 38494 76729 38513
rect 80343 38599 80729 38618
rect 80343 38576 80409 38599
rect 80495 38576 80577 38599
rect 80663 38576 80729 38599
rect 80343 38536 80352 38576
rect 80392 38536 80409 38576
rect 80495 38536 80516 38576
rect 80556 38536 80577 38576
rect 80663 38536 80680 38576
rect 80720 38536 80729 38576
rect 80343 38513 80409 38536
rect 80495 38513 80577 38536
rect 80663 38513 80729 38536
rect 80343 38494 80729 38513
rect 84343 38599 84729 38618
rect 84343 38576 84409 38599
rect 84495 38576 84577 38599
rect 84663 38576 84729 38599
rect 84343 38536 84352 38576
rect 84392 38536 84409 38576
rect 84495 38536 84516 38576
rect 84556 38536 84577 38576
rect 84663 38536 84680 38576
rect 84720 38536 84729 38576
rect 84343 38513 84409 38536
rect 84495 38513 84577 38536
rect 84663 38513 84729 38536
rect 84343 38494 84729 38513
rect 88343 38599 88729 38618
rect 88343 38576 88409 38599
rect 88495 38576 88577 38599
rect 88663 38576 88729 38599
rect 88343 38536 88352 38576
rect 88392 38536 88409 38576
rect 88495 38536 88516 38576
rect 88556 38536 88577 38576
rect 88663 38536 88680 38576
rect 88720 38536 88729 38576
rect 88343 38513 88409 38536
rect 88495 38513 88577 38536
rect 88663 38513 88729 38536
rect 88343 38494 88729 38513
rect 92343 38599 92729 38618
rect 92343 38576 92409 38599
rect 92495 38576 92577 38599
rect 92663 38576 92729 38599
rect 92343 38536 92352 38576
rect 92392 38536 92409 38576
rect 92495 38536 92516 38576
rect 92556 38536 92577 38576
rect 92663 38536 92680 38576
rect 92720 38536 92729 38576
rect 92343 38513 92409 38536
rect 92495 38513 92577 38536
rect 92663 38513 92729 38536
rect 92343 38494 92729 38513
rect 96343 38599 96729 38618
rect 96343 38576 96409 38599
rect 96495 38576 96577 38599
rect 96663 38576 96729 38599
rect 96343 38536 96352 38576
rect 96392 38536 96409 38576
rect 96495 38536 96516 38576
rect 96556 38536 96577 38576
rect 96663 38536 96680 38576
rect 96720 38536 96729 38576
rect 96343 38513 96409 38536
rect 96495 38513 96577 38536
rect 96663 38513 96729 38536
rect 96343 38494 96729 38513
rect 3103 37843 3489 37862
rect 3103 37820 3169 37843
rect 3255 37820 3337 37843
rect 3423 37820 3489 37843
rect 3103 37780 3112 37820
rect 3152 37780 3169 37820
rect 3255 37780 3276 37820
rect 3316 37780 3337 37820
rect 3423 37780 3440 37820
rect 3480 37780 3489 37820
rect 3103 37757 3169 37780
rect 3255 37757 3337 37780
rect 3423 37757 3489 37780
rect 3103 37738 3489 37757
rect 7103 37843 7489 37862
rect 7103 37820 7169 37843
rect 7255 37820 7337 37843
rect 7423 37820 7489 37843
rect 7103 37780 7112 37820
rect 7152 37780 7169 37820
rect 7255 37780 7276 37820
rect 7316 37780 7337 37820
rect 7423 37780 7440 37820
rect 7480 37780 7489 37820
rect 7103 37757 7169 37780
rect 7255 37757 7337 37780
rect 7423 37757 7489 37780
rect 7103 37738 7489 37757
rect 11103 37843 11489 37862
rect 11103 37820 11169 37843
rect 11255 37820 11337 37843
rect 11423 37820 11489 37843
rect 11103 37780 11112 37820
rect 11152 37780 11169 37820
rect 11255 37780 11276 37820
rect 11316 37780 11337 37820
rect 11423 37780 11440 37820
rect 11480 37780 11489 37820
rect 11103 37757 11169 37780
rect 11255 37757 11337 37780
rect 11423 37757 11489 37780
rect 11103 37738 11489 37757
rect 15103 37843 15489 37862
rect 15103 37820 15169 37843
rect 15255 37820 15337 37843
rect 15423 37820 15489 37843
rect 15103 37780 15112 37820
rect 15152 37780 15169 37820
rect 15255 37780 15276 37820
rect 15316 37780 15337 37820
rect 15423 37780 15440 37820
rect 15480 37780 15489 37820
rect 15103 37757 15169 37780
rect 15255 37757 15337 37780
rect 15423 37757 15489 37780
rect 15103 37738 15489 37757
rect 19103 37843 19489 37862
rect 19103 37820 19169 37843
rect 19255 37820 19337 37843
rect 19423 37820 19489 37843
rect 19103 37780 19112 37820
rect 19152 37780 19169 37820
rect 19255 37780 19276 37820
rect 19316 37780 19337 37820
rect 19423 37780 19440 37820
rect 19480 37780 19489 37820
rect 19103 37757 19169 37780
rect 19255 37757 19337 37780
rect 19423 37757 19489 37780
rect 19103 37738 19489 37757
rect 23103 37843 23489 37862
rect 23103 37820 23169 37843
rect 23255 37820 23337 37843
rect 23423 37820 23489 37843
rect 23103 37780 23112 37820
rect 23152 37780 23169 37820
rect 23255 37780 23276 37820
rect 23316 37780 23337 37820
rect 23423 37780 23440 37820
rect 23480 37780 23489 37820
rect 23103 37757 23169 37780
rect 23255 37757 23337 37780
rect 23423 37757 23489 37780
rect 23103 37738 23489 37757
rect 27103 37843 27489 37862
rect 27103 37820 27169 37843
rect 27255 37820 27337 37843
rect 27423 37820 27489 37843
rect 27103 37780 27112 37820
rect 27152 37780 27169 37820
rect 27255 37780 27276 37820
rect 27316 37780 27337 37820
rect 27423 37780 27440 37820
rect 27480 37780 27489 37820
rect 27103 37757 27169 37780
rect 27255 37757 27337 37780
rect 27423 37757 27489 37780
rect 27103 37738 27489 37757
rect 31103 37843 31489 37862
rect 31103 37820 31169 37843
rect 31255 37820 31337 37843
rect 31423 37820 31489 37843
rect 31103 37780 31112 37820
rect 31152 37780 31169 37820
rect 31255 37780 31276 37820
rect 31316 37780 31337 37820
rect 31423 37780 31440 37820
rect 31480 37780 31489 37820
rect 31103 37757 31169 37780
rect 31255 37757 31337 37780
rect 31423 37757 31489 37780
rect 31103 37738 31489 37757
rect 35103 37843 35489 37862
rect 35103 37820 35169 37843
rect 35255 37820 35337 37843
rect 35423 37820 35489 37843
rect 35103 37780 35112 37820
rect 35152 37780 35169 37820
rect 35255 37780 35276 37820
rect 35316 37780 35337 37820
rect 35423 37780 35440 37820
rect 35480 37780 35489 37820
rect 35103 37757 35169 37780
rect 35255 37757 35337 37780
rect 35423 37757 35489 37780
rect 35103 37738 35489 37757
rect 39103 37843 39489 37862
rect 39103 37820 39169 37843
rect 39255 37820 39337 37843
rect 39423 37820 39489 37843
rect 39103 37780 39112 37820
rect 39152 37780 39169 37820
rect 39255 37780 39276 37820
rect 39316 37780 39337 37820
rect 39423 37780 39440 37820
rect 39480 37780 39489 37820
rect 39103 37757 39169 37780
rect 39255 37757 39337 37780
rect 39423 37757 39489 37780
rect 39103 37738 39489 37757
rect 43103 37843 43489 37862
rect 43103 37820 43169 37843
rect 43255 37820 43337 37843
rect 43423 37820 43489 37843
rect 43103 37780 43112 37820
rect 43152 37780 43169 37820
rect 43255 37780 43276 37820
rect 43316 37780 43337 37820
rect 43423 37780 43440 37820
rect 43480 37780 43489 37820
rect 43103 37757 43169 37780
rect 43255 37757 43337 37780
rect 43423 37757 43489 37780
rect 43103 37738 43489 37757
rect 47103 37843 47489 37862
rect 47103 37820 47169 37843
rect 47255 37820 47337 37843
rect 47423 37820 47489 37843
rect 47103 37780 47112 37820
rect 47152 37780 47169 37820
rect 47255 37780 47276 37820
rect 47316 37780 47337 37820
rect 47423 37780 47440 37820
rect 47480 37780 47489 37820
rect 47103 37757 47169 37780
rect 47255 37757 47337 37780
rect 47423 37757 47489 37780
rect 47103 37738 47489 37757
rect 51103 37843 51489 37862
rect 51103 37820 51169 37843
rect 51255 37820 51337 37843
rect 51423 37820 51489 37843
rect 51103 37780 51112 37820
rect 51152 37780 51169 37820
rect 51255 37780 51276 37820
rect 51316 37780 51337 37820
rect 51423 37780 51440 37820
rect 51480 37780 51489 37820
rect 51103 37757 51169 37780
rect 51255 37757 51337 37780
rect 51423 37757 51489 37780
rect 51103 37738 51489 37757
rect 55103 37843 55489 37862
rect 55103 37820 55169 37843
rect 55255 37820 55337 37843
rect 55423 37820 55489 37843
rect 55103 37780 55112 37820
rect 55152 37780 55169 37820
rect 55255 37780 55276 37820
rect 55316 37780 55337 37820
rect 55423 37780 55440 37820
rect 55480 37780 55489 37820
rect 55103 37757 55169 37780
rect 55255 37757 55337 37780
rect 55423 37757 55489 37780
rect 55103 37738 55489 37757
rect 59103 37843 59489 37862
rect 59103 37820 59169 37843
rect 59255 37820 59337 37843
rect 59423 37820 59489 37843
rect 59103 37780 59112 37820
rect 59152 37780 59169 37820
rect 59255 37780 59276 37820
rect 59316 37780 59337 37820
rect 59423 37780 59440 37820
rect 59480 37780 59489 37820
rect 59103 37757 59169 37780
rect 59255 37757 59337 37780
rect 59423 37757 59489 37780
rect 59103 37738 59489 37757
rect 63103 37843 63489 37862
rect 63103 37820 63169 37843
rect 63255 37820 63337 37843
rect 63423 37820 63489 37843
rect 63103 37780 63112 37820
rect 63152 37780 63169 37820
rect 63255 37780 63276 37820
rect 63316 37780 63337 37820
rect 63423 37780 63440 37820
rect 63480 37780 63489 37820
rect 63103 37757 63169 37780
rect 63255 37757 63337 37780
rect 63423 37757 63489 37780
rect 63103 37738 63489 37757
rect 67103 37843 67489 37862
rect 67103 37820 67169 37843
rect 67255 37820 67337 37843
rect 67423 37820 67489 37843
rect 67103 37780 67112 37820
rect 67152 37780 67169 37820
rect 67255 37780 67276 37820
rect 67316 37780 67337 37820
rect 67423 37780 67440 37820
rect 67480 37780 67489 37820
rect 67103 37757 67169 37780
rect 67255 37757 67337 37780
rect 67423 37757 67489 37780
rect 67103 37738 67489 37757
rect 71103 37843 71489 37862
rect 71103 37820 71169 37843
rect 71255 37820 71337 37843
rect 71423 37820 71489 37843
rect 71103 37780 71112 37820
rect 71152 37780 71169 37820
rect 71255 37780 71276 37820
rect 71316 37780 71337 37820
rect 71423 37780 71440 37820
rect 71480 37780 71489 37820
rect 71103 37757 71169 37780
rect 71255 37757 71337 37780
rect 71423 37757 71489 37780
rect 71103 37738 71489 37757
rect 75103 37843 75489 37862
rect 75103 37820 75169 37843
rect 75255 37820 75337 37843
rect 75423 37820 75489 37843
rect 75103 37780 75112 37820
rect 75152 37780 75169 37820
rect 75255 37780 75276 37820
rect 75316 37780 75337 37820
rect 75423 37780 75440 37820
rect 75480 37780 75489 37820
rect 75103 37757 75169 37780
rect 75255 37757 75337 37780
rect 75423 37757 75489 37780
rect 75103 37738 75489 37757
rect 79103 37843 79489 37862
rect 79103 37820 79169 37843
rect 79255 37820 79337 37843
rect 79423 37820 79489 37843
rect 79103 37780 79112 37820
rect 79152 37780 79169 37820
rect 79255 37780 79276 37820
rect 79316 37780 79337 37820
rect 79423 37780 79440 37820
rect 79480 37780 79489 37820
rect 79103 37757 79169 37780
rect 79255 37757 79337 37780
rect 79423 37757 79489 37780
rect 79103 37738 79489 37757
rect 83103 37843 83489 37862
rect 83103 37820 83169 37843
rect 83255 37820 83337 37843
rect 83423 37820 83489 37843
rect 83103 37780 83112 37820
rect 83152 37780 83169 37820
rect 83255 37780 83276 37820
rect 83316 37780 83337 37820
rect 83423 37780 83440 37820
rect 83480 37780 83489 37820
rect 83103 37757 83169 37780
rect 83255 37757 83337 37780
rect 83423 37757 83489 37780
rect 83103 37738 83489 37757
rect 87103 37843 87489 37862
rect 87103 37820 87169 37843
rect 87255 37820 87337 37843
rect 87423 37820 87489 37843
rect 87103 37780 87112 37820
rect 87152 37780 87169 37820
rect 87255 37780 87276 37820
rect 87316 37780 87337 37820
rect 87423 37780 87440 37820
rect 87480 37780 87489 37820
rect 87103 37757 87169 37780
rect 87255 37757 87337 37780
rect 87423 37757 87489 37780
rect 87103 37738 87489 37757
rect 91103 37843 91489 37862
rect 91103 37820 91169 37843
rect 91255 37820 91337 37843
rect 91423 37820 91489 37843
rect 91103 37780 91112 37820
rect 91152 37780 91169 37820
rect 91255 37780 91276 37820
rect 91316 37780 91337 37820
rect 91423 37780 91440 37820
rect 91480 37780 91489 37820
rect 91103 37757 91169 37780
rect 91255 37757 91337 37780
rect 91423 37757 91489 37780
rect 91103 37738 91489 37757
rect 95103 37843 95489 37862
rect 95103 37820 95169 37843
rect 95255 37820 95337 37843
rect 95423 37820 95489 37843
rect 95103 37780 95112 37820
rect 95152 37780 95169 37820
rect 95255 37780 95276 37820
rect 95316 37780 95337 37820
rect 95423 37780 95440 37820
rect 95480 37780 95489 37820
rect 95103 37757 95169 37780
rect 95255 37757 95337 37780
rect 95423 37757 95489 37780
rect 95103 37738 95489 37757
rect 99103 37843 99489 37862
rect 99103 37820 99169 37843
rect 99255 37820 99337 37843
rect 99423 37820 99489 37843
rect 99103 37780 99112 37820
rect 99152 37780 99169 37820
rect 99255 37780 99276 37820
rect 99316 37780 99337 37820
rect 99423 37780 99440 37820
rect 99480 37780 99489 37820
rect 99103 37757 99169 37780
rect 99255 37757 99337 37780
rect 99423 37757 99489 37780
rect 99103 37738 99489 37757
rect 4343 37087 4729 37106
rect 4343 37064 4409 37087
rect 4495 37064 4577 37087
rect 4663 37064 4729 37087
rect 4343 37024 4352 37064
rect 4392 37024 4409 37064
rect 4495 37024 4516 37064
rect 4556 37024 4577 37064
rect 4663 37024 4680 37064
rect 4720 37024 4729 37064
rect 4343 37001 4409 37024
rect 4495 37001 4577 37024
rect 4663 37001 4729 37024
rect 4343 36982 4729 37001
rect 8343 37087 8729 37106
rect 8343 37064 8409 37087
rect 8495 37064 8577 37087
rect 8663 37064 8729 37087
rect 8343 37024 8352 37064
rect 8392 37024 8409 37064
rect 8495 37024 8516 37064
rect 8556 37024 8577 37064
rect 8663 37024 8680 37064
rect 8720 37024 8729 37064
rect 8343 37001 8409 37024
rect 8495 37001 8577 37024
rect 8663 37001 8729 37024
rect 8343 36982 8729 37001
rect 12343 37087 12729 37106
rect 12343 37064 12409 37087
rect 12495 37064 12577 37087
rect 12663 37064 12729 37087
rect 12343 37024 12352 37064
rect 12392 37024 12409 37064
rect 12495 37024 12516 37064
rect 12556 37024 12577 37064
rect 12663 37024 12680 37064
rect 12720 37024 12729 37064
rect 12343 37001 12409 37024
rect 12495 37001 12577 37024
rect 12663 37001 12729 37024
rect 12343 36982 12729 37001
rect 16343 37087 16729 37106
rect 16343 37064 16409 37087
rect 16495 37064 16577 37087
rect 16663 37064 16729 37087
rect 16343 37024 16352 37064
rect 16392 37024 16409 37064
rect 16495 37024 16516 37064
rect 16556 37024 16577 37064
rect 16663 37024 16680 37064
rect 16720 37024 16729 37064
rect 16343 37001 16409 37024
rect 16495 37001 16577 37024
rect 16663 37001 16729 37024
rect 16343 36982 16729 37001
rect 20343 37087 20729 37106
rect 20343 37064 20409 37087
rect 20495 37064 20577 37087
rect 20663 37064 20729 37087
rect 20343 37024 20352 37064
rect 20392 37024 20409 37064
rect 20495 37024 20516 37064
rect 20556 37024 20577 37064
rect 20663 37024 20680 37064
rect 20720 37024 20729 37064
rect 20343 37001 20409 37024
rect 20495 37001 20577 37024
rect 20663 37001 20729 37024
rect 20343 36982 20729 37001
rect 24343 37087 24729 37106
rect 24343 37064 24409 37087
rect 24495 37064 24577 37087
rect 24663 37064 24729 37087
rect 24343 37024 24352 37064
rect 24392 37024 24409 37064
rect 24495 37024 24516 37064
rect 24556 37024 24577 37064
rect 24663 37024 24680 37064
rect 24720 37024 24729 37064
rect 24343 37001 24409 37024
rect 24495 37001 24577 37024
rect 24663 37001 24729 37024
rect 24343 36982 24729 37001
rect 28343 37087 28729 37106
rect 28343 37064 28409 37087
rect 28495 37064 28577 37087
rect 28663 37064 28729 37087
rect 28343 37024 28352 37064
rect 28392 37024 28409 37064
rect 28495 37024 28516 37064
rect 28556 37024 28577 37064
rect 28663 37024 28680 37064
rect 28720 37024 28729 37064
rect 28343 37001 28409 37024
rect 28495 37001 28577 37024
rect 28663 37001 28729 37024
rect 28343 36982 28729 37001
rect 32343 37087 32729 37106
rect 32343 37064 32409 37087
rect 32495 37064 32577 37087
rect 32663 37064 32729 37087
rect 32343 37024 32352 37064
rect 32392 37024 32409 37064
rect 32495 37024 32516 37064
rect 32556 37024 32577 37064
rect 32663 37024 32680 37064
rect 32720 37024 32729 37064
rect 32343 37001 32409 37024
rect 32495 37001 32577 37024
rect 32663 37001 32729 37024
rect 32343 36982 32729 37001
rect 36343 37087 36729 37106
rect 36343 37064 36409 37087
rect 36495 37064 36577 37087
rect 36663 37064 36729 37087
rect 36343 37024 36352 37064
rect 36392 37024 36409 37064
rect 36495 37024 36516 37064
rect 36556 37024 36577 37064
rect 36663 37024 36680 37064
rect 36720 37024 36729 37064
rect 36343 37001 36409 37024
rect 36495 37001 36577 37024
rect 36663 37001 36729 37024
rect 36343 36982 36729 37001
rect 40343 37087 40729 37106
rect 40343 37064 40409 37087
rect 40495 37064 40577 37087
rect 40663 37064 40729 37087
rect 40343 37024 40352 37064
rect 40392 37024 40409 37064
rect 40495 37024 40516 37064
rect 40556 37024 40577 37064
rect 40663 37024 40680 37064
rect 40720 37024 40729 37064
rect 40343 37001 40409 37024
rect 40495 37001 40577 37024
rect 40663 37001 40729 37024
rect 40343 36982 40729 37001
rect 44343 37087 44729 37106
rect 44343 37064 44409 37087
rect 44495 37064 44577 37087
rect 44663 37064 44729 37087
rect 44343 37024 44352 37064
rect 44392 37024 44409 37064
rect 44495 37024 44516 37064
rect 44556 37024 44577 37064
rect 44663 37024 44680 37064
rect 44720 37024 44729 37064
rect 44343 37001 44409 37024
rect 44495 37001 44577 37024
rect 44663 37001 44729 37024
rect 44343 36982 44729 37001
rect 48343 37087 48729 37106
rect 48343 37064 48409 37087
rect 48495 37064 48577 37087
rect 48663 37064 48729 37087
rect 48343 37024 48352 37064
rect 48392 37024 48409 37064
rect 48495 37024 48516 37064
rect 48556 37024 48577 37064
rect 48663 37024 48680 37064
rect 48720 37024 48729 37064
rect 48343 37001 48409 37024
rect 48495 37001 48577 37024
rect 48663 37001 48729 37024
rect 48343 36982 48729 37001
rect 52343 37087 52729 37106
rect 52343 37064 52409 37087
rect 52495 37064 52577 37087
rect 52663 37064 52729 37087
rect 52343 37024 52352 37064
rect 52392 37024 52409 37064
rect 52495 37024 52516 37064
rect 52556 37024 52577 37064
rect 52663 37024 52680 37064
rect 52720 37024 52729 37064
rect 52343 37001 52409 37024
rect 52495 37001 52577 37024
rect 52663 37001 52729 37024
rect 52343 36982 52729 37001
rect 56343 37087 56729 37106
rect 56343 37064 56409 37087
rect 56495 37064 56577 37087
rect 56663 37064 56729 37087
rect 56343 37024 56352 37064
rect 56392 37024 56409 37064
rect 56495 37024 56516 37064
rect 56556 37024 56577 37064
rect 56663 37024 56680 37064
rect 56720 37024 56729 37064
rect 56343 37001 56409 37024
rect 56495 37001 56577 37024
rect 56663 37001 56729 37024
rect 56343 36982 56729 37001
rect 60343 37087 60729 37106
rect 60343 37064 60409 37087
rect 60495 37064 60577 37087
rect 60663 37064 60729 37087
rect 60343 37024 60352 37064
rect 60392 37024 60409 37064
rect 60495 37024 60516 37064
rect 60556 37024 60577 37064
rect 60663 37024 60680 37064
rect 60720 37024 60729 37064
rect 60343 37001 60409 37024
rect 60495 37001 60577 37024
rect 60663 37001 60729 37024
rect 60343 36982 60729 37001
rect 64343 37087 64729 37106
rect 64343 37064 64409 37087
rect 64495 37064 64577 37087
rect 64663 37064 64729 37087
rect 64343 37024 64352 37064
rect 64392 37024 64409 37064
rect 64495 37024 64516 37064
rect 64556 37024 64577 37064
rect 64663 37024 64680 37064
rect 64720 37024 64729 37064
rect 64343 37001 64409 37024
rect 64495 37001 64577 37024
rect 64663 37001 64729 37024
rect 64343 36982 64729 37001
rect 68343 37087 68729 37106
rect 68343 37064 68409 37087
rect 68495 37064 68577 37087
rect 68663 37064 68729 37087
rect 68343 37024 68352 37064
rect 68392 37024 68409 37064
rect 68495 37024 68516 37064
rect 68556 37024 68577 37064
rect 68663 37024 68680 37064
rect 68720 37024 68729 37064
rect 68343 37001 68409 37024
rect 68495 37001 68577 37024
rect 68663 37001 68729 37024
rect 68343 36982 68729 37001
rect 72343 37087 72729 37106
rect 72343 37064 72409 37087
rect 72495 37064 72577 37087
rect 72663 37064 72729 37087
rect 72343 37024 72352 37064
rect 72392 37024 72409 37064
rect 72495 37024 72516 37064
rect 72556 37024 72577 37064
rect 72663 37024 72680 37064
rect 72720 37024 72729 37064
rect 72343 37001 72409 37024
rect 72495 37001 72577 37024
rect 72663 37001 72729 37024
rect 72343 36982 72729 37001
rect 76343 37087 76729 37106
rect 76343 37064 76409 37087
rect 76495 37064 76577 37087
rect 76663 37064 76729 37087
rect 76343 37024 76352 37064
rect 76392 37024 76409 37064
rect 76495 37024 76516 37064
rect 76556 37024 76577 37064
rect 76663 37024 76680 37064
rect 76720 37024 76729 37064
rect 76343 37001 76409 37024
rect 76495 37001 76577 37024
rect 76663 37001 76729 37024
rect 76343 36982 76729 37001
rect 80343 37087 80729 37106
rect 80343 37064 80409 37087
rect 80495 37064 80577 37087
rect 80663 37064 80729 37087
rect 80343 37024 80352 37064
rect 80392 37024 80409 37064
rect 80495 37024 80516 37064
rect 80556 37024 80577 37064
rect 80663 37024 80680 37064
rect 80720 37024 80729 37064
rect 80343 37001 80409 37024
rect 80495 37001 80577 37024
rect 80663 37001 80729 37024
rect 80343 36982 80729 37001
rect 84343 37087 84729 37106
rect 84343 37064 84409 37087
rect 84495 37064 84577 37087
rect 84663 37064 84729 37087
rect 84343 37024 84352 37064
rect 84392 37024 84409 37064
rect 84495 37024 84516 37064
rect 84556 37024 84577 37064
rect 84663 37024 84680 37064
rect 84720 37024 84729 37064
rect 84343 37001 84409 37024
rect 84495 37001 84577 37024
rect 84663 37001 84729 37024
rect 84343 36982 84729 37001
rect 88343 37087 88729 37106
rect 88343 37064 88409 37087
rect 88495 37064 88577 37087
rect 88663 37064 88729 37087
rect 88343 37024 88352 37064
rect 88392 37024 88409 37064
rect 88495 37024 88516 37064
rect 88556 37024 88577 37064
rect 88663 37024 88680 37064
rect 88720 37024 88729 37064
rect 88343 37001 88409 37024
rect 88495 37001 88577 37024
rect 88663 37001 88729 37024
rect 88343 36982 88729 37001
rect 92343 37087 92729 37106
rect 92343 37064 92409 37087
rect 92495 37064 92577 37087
rect 92663 37064 92729 37087
rect 92343 37024 92352 37064
rect 92392 37024 92409 37064
rect 92495 37024 92516 37064
rect 92556 37024 92577 37064
rect 92663 37024 92680 37064
rect 92720 37024 92729 37064
rect 92343 37001 92409 37024
rect 92495 37001 92577 37024
rect 92663 37001 92729 37024
rect 92343 36982 92729 37001
rect 96343 37087 96729 37106
rect 96343 37064 96409 37087
rect 96495 37064 96577 37087
rect 96663 37064 96729 37087
rect 96343 37024 96352 37064
rect 96392 37024 96409 37064
rect 96495 37024 96516 37064
rect 96556 37024 96577 37064
rect 96663 37024 96680 37064
rect 96720 37024 96729 37064
rect 96343 37001 96409 37024
rect 96495 37001 96577 37024
rect 96663 37001 96729 37024
rect 96343 36982 96729 37001
rect 3103 36331 3489 36350
rect 3103 36308 3169 36331
rect 3255 36308 3337 36331
rect 3423 36308 3489 36331
rect 3103 36268 3112 36308
rect 3152 36268 3169 36308
rect 3255 36268 3276 36308
rect 3316 36268 3337 36308
rect 3423 36268 3440 36308
rect 3480 36268 3489 36308
rect 3103 36245 3169 36268
rect 3255 36245 3337 36268
rect 3423 36245 3489 36268
rect 3103 36226 3489 36245
rect 7103 36331 7489 36350
rect 7103 36308 7169 36331
rect 7255 36308 7337 36331
rect 7423 36308 7489 36331
rect 7103 36268 7112 36308
rect 7152 36268 7169 36308
rect 7255 36268 7276 36308
rect 7316 36268 7337 36308
rect 7423 36268 7440 36308
rect 7480 36268 7489 36308
rect 7103 36245 7169 36268
rect 7255 36245 7337 36268
rect 7423 36245 7489 36268
rect 7103 36226 7489 36245
rect 11103 36331 11489 36350
rect 11103 36308 11169 36331
rect 11255 36308 11337 36331
rect 11423 36308 11489 36331
rect 11103 36268 11112 36308
rect 11152 36268 11169 36308
rect 11255 36268 11276 36308
rect 11316 36268 11337 36308
rect 11423 36268 11440 36308
rect 11480 36268 11489 36308
rect 11103 36245 11169 36268
rect 11255 36245 11337 36268
rect 11423 36245 11489 36268
rect 11103 36226 11489 36245
rect 15103 36331 15489 36350
rect 15103 36308 15169 36331
rect 15255 36308 15337 36331
rect 15423 36308 15489 36331
rect 15103 36268 15112 36308
rect 15152 36268 15169 36308
rect 15255 36268 15276 36308
rect 15316 36268 15337 36308
rect 15423 36268 15440 36308
rect 15480 36268 15489 36308
rect 15103 36245 15169 36268
rect 15255 36245 15337 36268
rect 15423 36245 15489 36268
rect 15103 36226 15489 36245
rect 19103 36331 19489 36350
rect 19103 36308 19169 36331
rect 19255 36308 19337 36331
rect 19423 36308 19489 36331
rect 19103 36268 19112 36308
rect 19152 36268 19169 36308
rect 19255 36268 19276 36308
rect 19316 36268 19337 36308
rect 19423 36268 19440 36308
rect 19480 36268 19489 36308
rect 19103 36245 19169 36268
rect 19255 36245 19337 36268
rect 19423 36245 19489 36268
rect 19103 36226 19489 36245
rect 23103 36331 23489 36350
rect 23103 36308 23169 36331
rect 23255 36308 23337 36331
rect 23423 36308 23489 36331
rect 23103 36268 23112 36308
rect 23152 36268 23169 36308
rect 23255 36268 23276 36308
rect 23316 36268 23337 36308
rect 23423 36268 23440 36308
rect 23480 36268 23489 36308
rect 23103 36245 23169 36268
rect 23255 36245 23337 36268
rect 23423 36245 23489 36268
rect 23103 36226 23489 36245
rect 27103 36331 27489 36350
rect 27103 36308 27169 36331
rect 27255 36308 27337 36331
rect 27423 36308 27489 36331
rect 27103 36268 27112 36308
rect 27152 36268 27169 36308
rect 27255 36268 27276 36308
rect 27316 36268 27337 36308
rect 27423 36268 27440 36308
rect 27480 36268 27489 36308
rect 27103 36245 27169 36268
rect 27255 36245 27337 36268
rect 27423 36245 27489 36268
rect 27103 36226 27489 36245
rect 31103 36331 31489 36350
rect 31103 36308 31169 36331
rect 31255 36308 31337 36331
rect 31423 36308 31489 36331
rect 31103 36268 31112 36308
rect 31152 36268 31169 36308
rect 31255 36268 31276 36308
rect 31316 36268 31337 36308
rect 31423 36268 31440 36308
rect 31480 36268 31489 36308
rect 31103 36245 31169 36268
rect 31255 36245 31337 36268
rect 31423 36245 31489 36268
rect 31103 36226 31489 36245
rect 35103 36331 35489 36350
rect 35103 36308 35169 36331
rect 35255 36308 35337 36331
rect 35423 36308 35489 36331
rect 35103 36268 35112 36308
rect 35152 36268 35169 36308
rect 35255 36268 35276 36308
rect 35316 36268 35337 36308
rect 35423 36268 35440 36308
rect 35480 36268 35489 36308
rect 35103 36245 35169 36268
rect 35255 36245 35337 36268
rect 35423 36245 35489 36268
rect 35103 36226 35489 36245
rect 39103 36331 39489 36350
rect 39103 36308 39169 36331
rect 39255 36308 39337 36331
rect 39423 36308 39489 36331
rect 39103 36268 39112 36308
rect 39152 36268 39169 36308
rect 39255 36268 39276 36308
rect 39316 36268 39337 36308
rect 39423 36268 39440 36308
rect 39480 36268 39489 36308
rect 39103 36245 39169 36268
rect 39255 36245 39337 36268
rect 39423 36245 39489 36268
rect 39103 36226 39489 36245
rect 43103 36331 43489 36350
rect 43103 36308 43169 36331
rect 43255 36308 43337 36331
rect 43423 36308 43489 36331
rect 43103 36268 43112 36308
rect 43152 36268 43169 36308
rect 43255 36268 43276 36308
rect 43316 36268 43337 36308
rect 43423 36268 43440 36308
rect 43480 36268 43489 36308
rect 43103 36245 43169 36268
rect 43255 36245 43337 36268
rect 43423 36245 43489 36268
rect 43103 36226 43489 36245
rect 47103 36331 47489 36350
rect 47103 36308 47169 36331
rect 47255 36308 47337 36331
rect 47423 36308 47489 36331
rect 47103 36268 47112 36308
rect 47152 36268 47169 36308
rect 47255 36268 47276 36308
rect 47316 36268 47337 36308
rect 47423 36268 47440 36308
rect 47480 36268 47489 36308
rect 47103 36245 47169 36268
rect 47255 36245 47337 36268
rect 47423 36245 47489 36268
rect 47103 36226 47489 36245
rect 51103 36331 51489 36350
rect 51103 36308 51169 36331
rect 51255 36308 51337 36331
rect 51423 36308 51489 36331
rect 51103 36268 51112 36308
rect 51152 36268 51169 36308
rect 51255 36268 51276 36308
rect 51316 36268 51337 36308
rect 51423 36268 51440 36308
rect 51480 36268 51489 36308
rect 51103 36245 51169 36268
rect 51255 36245 51337 36268
rect 51423 36245 51489 36268
rect 51103 36226 51489 36245
rect 55103 36331 55489 36350
rect 55103 36308 55169 36331
rect 55255 36308 55337 36331
rect 55423 36308 55489 36331
rect 55103 36268 55112 36308
rect 55152 36268 55169 36308
rect 55255 36268 55276 36308
rect 55316 36268 55337 36308
rect 55423 36268 55440 36308
rect 55480 36268 55489 36308
rect 55103 36245 55169 36268
rect 55255 36245 55337 36268
rect 55423 36245 55489 36268
rect 55103 36226 55489 36245
rect 59103 36331 59489 36350
rect 59103 36308 59169 36331
rect 59255 36308 59337 36331
rect 59423 36308 59489 36331
rect 59103 36268 59112 36308
rect 59152 36268 59169 36308
rect 59255 36268 59276 36308
rect 59316 36268 59337 36308
rect 59423 36268 59440 36308
rect 59480 36268 59489 36308
rect 59103 36245 59169 36268
rect 59255 36245 59337 36268
rect 59423 36245 59489 36268
rect 59103 36226 59489 36245
rect 63103 36331 63489 36350
rect 63103 36308 63169 36331
rect 63255 36308 63337 36331
rect 63423 36308 63489 36331
rect 63103 36268 63112 36308
rect 63152 36268 63169 36308
rect 63255 36268 63276 36308
rect 63316 36268 63337 36308
rect 63423 36268 63440 36308
rect 63480 36268 63489 36308
rect 63103 36245 63169 36268
rect 63255 36245 63337 36268
rect 63423 36245 63489 36268
rect 63103 36226 63489 36245
rect 67103 36331 67489 36350
rect 67103 36308 67169 36331
rect 67255 36308 67337 36331
rect 67423 36308 67489 36331
rect 67103 36268 67112 36308
rect 67152 36268 67169 36308
rect 67255 36268 67276 36308
rect 67316 36268 67337 36308
rect 67423 36268 67440 36308
rect 67480 36268 67489 36308
rect 67103 36245 67169 36268
rect 67255 36245 67337 36268
rect 67423 36245 67489 36268
rect 67103 36226 67489 36245
rect 71103 36331 71489 36350
rect 71103 36308 71169 36331
rect 71255 36308 71337 36331
rect 71423 36308 71489 36331
rect 71103 36268 71112 36308
rect 71152 36268 71169 36308
rect 71255 36268 71276 36308
rect 71316 36268 71337 36308
rect 71423 36268 71440 36308
rect 71480 36268 71489 36308
rect 71103 36245 71169 36268
rect 71255 36245 71337 36268
rect 71423 36245 71489 36268
rect 71103 36226 71489 36245
rect 75103 36331 75489 36350
rect 75103 36308 75169 36331
rect 75255 36308 75337 36331
rect 75423 36308 75489 36331
rect 75103 36268 75112 36308
rect 75152 36268 75169 36308
rect 75255 36268 75276 36308
rect 75316 36268 75337 36308
rect 75423 36268 75440 36308
rect 75480 36268 75489 36308
rect 75103 36245 75169 36268
rect 75255 36245 75337 36268
rect 75423 36245 75489 36268
rect 75103 36226 75489 36245
rect 79103 36331 79489 36350
rect 79103 36308 79169 36331
rect 79255 36308 79337 36331
rect 79423 36308 79489 36331
rect 79103 36268 79112 36308
rect 79152 36268 79169 36308
rect 79255 36268 79276 36308
rect 79316 36268 79337 36308
rect 79423 36268 79440 36308
rect 79480 36268 79489 36308
rect 79103 36245 79169 36268
rect 79255 36245 79337 36268
rect 79423 36245 79489 36268
rect 79103 36226 79489 36245
rect 83103 36331 83489 36350
rect 83103 36308 83169 36331
rect 83255 36308 83337 36331
rect 83423 36308 83489 36331
rect 83103 36268 83112 36308
rect 83152 36268 83169 36308
rect 83255 36268 83276 36308
rect 83316 36268 83337 36308
rect 83423 36268 83440 36308
rect 83480 36268 83489 36308
rect 83103 36245 83169 36268
rect 83255 36245 83337 36268
rect 83423 36245 83489 36268
rect 83103 36226 83489 36245
rect 87103 36331 87489 36350
rect 87103 36308 87169 36331
rect 87255 36308 87337 36331
rect 87423 36308 87489 36331
rect 87103 36268 87112 36308
rect 87152 36268 87169 36308
rect 87255 36268 87276 36308
rect 87316 36268 87337 36308
rect 87423 36268 87440 36308
rect 87480 36268 87489 36308
rect 87103 36245 87169 36268
rect 87255 36245 87337 36268
rect 87423 36245 87489 36268
rect 87103 36226 87489 36245
rect 91103 36331 91489 36350
rect 91103 36308 91169 36331
rect 91255 36308 91337 36331
rect 91423 36308 91489 36331
rect 91103 36268 91112 36308
rect 91152 36268 91169 36308
rect 91255 36268 91276 36308
rect 91316 36268 91337 36308
rect 91423 36268 91440 36308
rect 91480 36268 91489 36308
rect 91103 36245 91169 36268
rect 91255 36245 91337 36268
rect 91423 36245 91489 36268
rect 91103 36226 91489 36245
rect 95103 36331 95489 36350
rect 95103 36308 95169 36331
rect 95255 36308 95337 36331
rect 95423 36308 95489 36331
rect 95103 36268 95112 36308
rect 95152 36268 95169 36308
rect 95255 36268 95276 36308
rect 95316 36268 95337 36308
rect 95423 36268 95440 36308
rect 95480 36268 95489 36308
rect 95103 36245 95169 36268
rect 95255 36245 95337 36268
rect 95423 36245 95489 36268
rect 95103 36226 95489 36245
rect 99103 36331 99489 36350
rect 99103 36308 99169 36331
rect 99255 36308 99337 36331
rect 99423 36308 99489 36331
rect 99103 36268 99112 36308
rect 99152 36268 99169 36308
rect 99255 36268 99276 36308
rect 99316 36268 99337 36308
rect 99423 36268 99440 36308
rect 99480 36268 99489 36308
rect 99103 36245 99169 36268
rect 99255 36245 99337 36268
rect 99423 36245 99489 36268
rect 99103 36226 99489 36245
rect 4343 35575 4729 35594
rect 4343 35552 4409 35575
rect 4495 35552 4577 35575
rect 4663 35552 4729 35575
rect 4343 35512 4352 35552
rect 4392 35512 4409 35552
rect 4495 35512 4516 35552
rect 4556 35512 4577 35552
rect 4663 35512 4680 35552
rect 4720 35512 4729 35552
rect 4343 35489 4409 35512
rect 4495 35489 4577 35512
rect 4663 35489 4729 35512
rect 4343 35470 4729 35489
rect 8343 35575 8729 35594
rect 8343 35552 8409 35575
rect 8495 35552 8577 35575
rect 8663 35552 8729 35575
rect 8343 35512 8352 35552
rect 8392 35512 8409 35552
rect 8495 35512 8516 35552
rect 8556 35512 8577 35552
rect 8663 35512 8680 35552
rect 8720 35512 8729 35552
rect 8343 35489 8409 35512
rect 8495 35489 8577 35512
rect 8663 35489 8729 35512
rect 8343 35470 8729 35489
rect 12343 35575 12729 35594
rect 12343 35552 12409 35575
rect 12495 35552 12577 35575
rect 12663 35552 12729 35575
rect 12343 35512 12352 35552
rect 12392 35512 12409 35552
rect 12495 35512 12516 35552
rect 12556 35512 12577 35552
rect 12663 35512 12680 35552
rect 12720 35512 12729 35552
rect 12343 35489 12409 35512
rect 12495 35489 12577 35512
rect 12663 35489 12729 35512
rect 12343 35470 12729 35489
rect 16343 35575 16729 35594
rect 16343 35552 16409 35575
rect 16495 35552 16577 35575
rect 16663 35552 16729 35575
rect 16343 35512 16352 35552
rect 16392 35512 16409 35552
rect 16495 35512 16516 35552
rect 16556 35512 16577 35552
rect 16663 35512 16680 35552
rect 16720 35512 16729 35552
rect 16343 35489 16409 35512
rect 16495 35489 16577 35512
rect 16663 35489 16729 35512
rect 16343 35470 16729 35489
rect 20343 35575 20729 35594
rect 20343 35552 20409 35575
rect 20495 35552 20577 35575
rect 20663 35552 20729 35575
rect 20343 35512 20352 35552
rect 20392 35512 20409 35552
rect 20495 35512 20516 35552
rect 20556 35512 20577 35552
rect 20663 35512 20680 35552
rect 20720 35512 20729 35552
rect 20343 35489 20409 35512
rect 20495 35489 20577 35512
rect 20663 35489 20729 35512
rect 20343 35470 20729 35489
rect 24343 35575 24729 35594
rect 24343 35552 24409 35575
rect 24495 35552 24577 35575
rect 24663 35552 24729 35575
rect 24343 35512 24352 35552
rect 24392 35512 24409 35552
rect 24495 35512 24516 35552
rect 24556 35512 24577 35552
rect 24663 35512 24680 35552
rect 24720 35512 24729 35552
rect 24343 35489 24409 35512
rect 24495 35489 24577 35512
rect 24663 35489 24729 35512
rect 24343 35470 24729 35489
rect 28343 35575 28729 35594
rect 28343 35552 28409 35575
rect 28495 35552 28577 35575
rect 28663 35552 28729 35575
rect 28343 35512 28352 35552
rect 28392 35512 28409 35552
rect 28495 35512 28516 35552
rect 28556 35512 28577 35552
rect 28663 35512 28680 35552
rect 28720 35512 28729 35552
rect 28343 35489 28409 35512
rect 28495 35489 28577 35512
rect 28663 35489 28729 35512
rect 28343 35470 28729 35489
rect 32343 35575 32729 35594
rect 32343 35552 32409 35575
rect 32495 35552 32577 35575
rect 32663 35552 32729 35575
rect 32343 35512 32352 35552
rect 32392 35512 32409 35552
rect 32495 35512 32516 35552
rect 32556 35512 32577 35552
rect 32663 35512 32680 35552
rect 32720 35512 32729 35552
rect 32343 35489 32409 35512
rect 32495 35489 32577 35512
rect 32663 35489 32729 35512
rect 32343 35470 32729 35489
rect 36343 35575 36729 35594
rect 36343 35552 36409 35575
rect 36495 35552 36577 35575
rect 36663 35552 36729 35575
rect 36343 35512 36352 35552
rect 36392 35512 36409 35552
rect 36495 35512 36516 35552
rect 36556 35512 36577 35552
rect 36663 35512 36680 35552
rect 36720 35512 36729 35552
rect 36343 35489 36409 35512
rect 36495 35489 36577 35512
rect 36663 35489 36729 35512
rect 36343 35470 36729 35489
rect 40343 35575 40729 35594
rect 40343 35552 40409 35575
rect 40495 35552 40577 35575
rect 40663 35552 40729 35575
rect 40343 35512 40352 35552
rect 40392 35512 40409 35552
rect 40495 35512 40516 35552
rect 40556 35512 40577 35552
rect 40663 35512 40680 35552
rect 40720 35512 40729 35552
rect 40343 35489 40409 35512
rect 40495 35489 40577 35512
rect 40663 35489 40729 35512
rect 40343 35470 40729 35489
rect 44343 35575 44729 35594
rect 44343 35552 44409 35575
rect 44495 35552 44577 35575
rect 44663 35552 44729 35575
rect 44343 35512 44352 35552
rect 44392 35512 44409 35552
rect 44495 35512 44516 35552
rect 44556 35512 44577 35552
rect 44663 35512 44680 35552
rect 44720 35512 44729 35552
rect 44343 35489 44409 35512
rect 44495 35489 44577 35512
rect 44663 35489 44729 35512
rect 44343 35470 44729 35489
rect 48343 35575 48729 35594
rect 48343 35552 48409 35575
rect 48495 35552 48577 35575
rect 48663 35552 48729 35575
rect 48343 35512 48352 35552
rect 48392 35512 48409 35552
rect 48495 35512 48516 35552
rect 48556 35512 48577 35552
rect 48663 35512 48680 35552
rect 48720 35512 48729 35552
rect 48343 35489 48409 35512
rect 48495 35489 48577 35512
rect 48663 35489 48729 35512
rect 48343 35470 48729 35489
rect 52343 35575 52729 35594
rect 52343 35552 52409 35575
rect 52495 35552 52577 35575
rect 52663 35552 52729 35575
rect 52343 35512 52352 35552
rect 52392 35512 52409 35552
rect 52495 35512 52516 35552
rect 52556 35512 52577 35552
rect 52663 35512 52680 35552
rect 52720 35512 52729 35552
rect 52343 35489 52409 35512
rect 52495 35489 52577 35512
rect 52663 35489 52729 35512
rect 52343 35470 52729 35489
rect 56343 35575 56729 35594
rect 56343 35552 56409 35575
rect 56495 35552 56577 35575
rect 56663 35552 56729 35575
rect 56343 35512 56352 35552
rect 56392 35512 56409 35552
rect 56495 35512 56516 35552
rect 56556 35512 56577 35552
rect 56663 35512 56680 35552
rect 56720 35512 56729 35552
rect 56343 35489 56409 35512
rect 56495 35489 56577 35512
rect 56663 35489 56729 35512
rect 56343 35470 56729 35489
rect 60343 35575 60729 35594
rect 60343 35552 60409 35575
rect 60495 35552 60577 35575
rect 60663 35552 60729 35575
rect 60343 35512 60352 35552
rect 60392 35512 60409 35552
rect 60495 35512 60516 35552
rect 60556 35512 60577 35552
rect 60663 35512 60680 35552
rect 60720 35512 60729 35552
rect 60343 35489 60409 35512
rect 60495 35489 60577 35512
rect 60663 35489 60729 35512
rect 60343 35470 60729 35489
rect 64343 35575 64729 35594
rect 64343 35552 64409 35575
rect 64495 35552 64577 35575
rect 64663 35552 64729 35575
rect 64343 35512 64352 35552
rect 64392 35512 64409 35552
rect 64495 35512 64516 35552
rect 64556 35512 64577 35552
rect 64663 35512 64680 35552
rect 64720 35512 64729 35552
rect 64343 35489 64409 35512
rect 64495 35489 64577 35512
rect 64663 35489 64729 35512
rect 64343 35470 64729 35489
rect 68343 35575 68729 35594
rect 68343 35552 68409 35575
rect 68495 35552 68577 35575
rect 68663 35552 68729 35575
rect 68343 35512 68352 35552
rect 68392 35512 68409 35552
rect 68495 35512 68516 35552
rect 68556 35512 68577 35552
rect 68663 35512 68680 35552
rect 68720 35512 68729 35552
rect 68343 35489 68409 35512
rect 68495 35489 68577 35512
rect 68663 35489 68729 35512
rect 68343 35470 68729 35489
rect 72343 35575 72729 35594
rect 72343 35552 72409 35575
rect 72495 35552 72577 35575
rect 72663 35552 72729 35575
rect 72343 35512 72352 35552
rect 72392 35512 72409 35552
rect 72495 35512 72516 35552
rect 72556 35512 72577 35552
rect 72663 35512 72680 35552
rect 72720 35512 72729 35552
rect 72343 35489 72409 35512
rect 72495 35489 72577 35512
rect 72663 35489 72729 35512
rect 72343 35470 72729 35489
rect 76343 35575 76729 35594
rect 76343 35552 76409 35575
rect 76495 35552 76577 35575
rect 76663 35552 76729 35575
rect 76343 35512 76352 35552
rect 76392 35512 76409 35552
rect 76495 35512 76516 35552
rect 76556 35512 76577 35552
rect 76663 35512 76680 35552
rect 76720 35512 76729 35552
rect 76343 35489 76409 35512
rect 76495 35489 76577 35512
rect 76663 35489 76729 35512
rect 76343 35470 76729 35489
rect 80343 35575 80729 35594
rect 80343 35552 80409 35575
rect 80495 35552 80577 35575
rect 80663 35552 80729 35575
rect 80343 35512 80352 35552
rect 80392 35512 80409 35552
rect 80495 35512 80516 35552
rect 80556 35512 80577 35552
rect 80663 35512 80680 35552
rect 80720 35512 80729 35552
rect 80343 35489 80409 35512
rect 80495 35489 80577 35512
rect 80663 35489 80729 35512
rect 80343 35470 80729 35489
rect 84343 35575 84729 35594
rect 84343 35552 84409 35575
rect 84495 35552 84577 35575
rect 84663 35552 84729 35575
rect 84343 35512 84352 35552
rect 84392 35512 84409 35552
rect 84495 35512 84516 35552
rect 84556 35512 84577 35552
rect 84663 35512 84680 35552
rect 84720 35512 84729 35552
rect 84343 35489 84409 35512
rect 84495 35489 84577 35512
rect 84663 35489 84729 35512
rect 84343 35470 84729 35489
rect 88343 35575 88729 35594
rect 88343 35552 88409 35575
rect 88495 35552 88577 35575
rect 88663 35552 88729 35575
rect 88343 35512 88352 35552
rect 88392 35512 88409 35552
rect 88495 35512 88516 35552
rect 88556 35512 88577 35552
rect 88663 35512 88680 35552
rect 88720 35512 88729 35552
rect 88343 35489 88409 35512
rect 88495 35489 88577 35512
rect 88663 35489 88729 35512
rect 88343 35470 88729 35489
rect 92343 35575 92729 35594
rect 92343 35552 92409 35575
rect 92495 35552 92577 35575
rect 92663 35552 92729 35575
rect 92343 35512 92352 35552
rect 92392 35512 92409 35552
rect 92495 35512 92516 35552
rect 92556 35512 92577 35552
rect 92663 35512 92680 35552
rect 92720 35512 92729 35552
rect 92343 35489 92409 35512
rect 92495 35489 92577 35512
rect 92663 35489 92729 35512
rect 92343 35470 92729 35489
rect 96343 35575 96729 35594
rect 96343 35552 96409 35575
rect 96495 35552 96577 35575
rect 96663 35552 96729 35575
rect 96343 35512 96352 35552
rect 96392 35512 96409 35552
rect 96495 35512 96516 35552
rect 96556 35512 96577 35552
rect 96663 35512 96680 35552
rect 96720 35512 96729 35552
rect 96343 35489 96409 35512
rect 96495 35489 96577 35512
rect 96663 35489 96729 35512
rect 96343 35470 96729 35489
rect 86450 34987 86574 35006
rect 86450 34901 86469 34987
rect 86555 34964 86574 34987
rect 86555 34924 86668 34964
rect 86708 34924 86717 34964
rect 86555 34901 86574 34924
rect 86450 34882 86574 34901
rect 3103 34819 3489 34838
rect 3103 34796 3169 34819
rect 3255 34796 3337 34819
rect 3423 34796 3489 34819
rect 3103 34756 3112 34796
rect 3152 34756 3169 34796
rect 3255 34756 3276 34796
rect 3316 34756 3337 34796
rect 3423 34756 3440 34796
rect 3480 34756 3489 34796
rect 3103 34733 3169 34756
rect 3255 34733 3337 34756
rect 3423 34733 3489 34756
rect 3103 34714 3489 34733
rect 7103 34819 7489 34838
rect 7103 34796 7169 34819
rect 7255 34796 7337 34819
rect 7423 34796 7489 34819
rect 7103 34756 7112 34796
rect 7152 34756 7169 34796
rect 7255 34756 7276 34796
rect 7316 34756 7337 34796
rect 7423 34756 7440 34796
rect 7480 34756 7489 34796
rect 7103 34733 7169 34756
rect 7255 34733 7337 34756
rect 7423 34733 7489 34756
rect 7103 34714 7489 34733
rect 11103 34819 11489 34838
rect 11103 34796 11169 34819
rect 11255 34796 11337 34819
rect 11423 34796 11489 34819
rect 11103 34756 11112 34796
rect 11152 34756 11169 34796
rect 11255 34756 11276 34796
rect 11316 34756 11337 34796
rect 11423 34756 11440 34796
rect 11480 34756 11489 34796
rect 11103 34733 11169 34756
rect 11255 34733 11337 34756
rect 11423 34733 11489 34756
rect 11103 34714 11489 34733
rect 15103 34819 15489 34838
rect 15103 34796 15169 34819
rect 15255 34796 15337 34819
rect 15423 34796 15489 34819
rect 15103 34756 15112 34796
rect 15152 34756 15169 34796
rect 15255 34756 15276 34796
rect 15316 34756 15337 34796
rect 15423 34756 15440 34796
rect 15480 34756 15489 34796
rect 15103 34733 15169 34756
rect 15255 34733 15337 34756
rect 15423 34733 15489 34756
rect 15103 34714 15489 34733
rect 19103 34819 19489 34838
rect 19103 34796 19169 34819
rect 19255 34796 19337 34819
rect 19423 34796 19489 34819
rect 19103 34756 19112 34796
rect 19152 34756 19169 34796
rect 19255 34756 19276 34796
rect 19316 34756 19337 34796
rect 19423 34756 19440 34796
rect 19480 34756 19489 34796
rect 19103 34733 19169 34756
rect 19255 34733 19337 34756
rect 19423 34733 19489 34756
rect 19103 34714 19489 34733
rect 23103 34819 23489 34838
rect 23103 34796 23169 34819
rect 23255 34796 23337 34819
rect 23423 34796 23489 34819
rect 23103 34756 23112 34796
rect 23152 34756 23169 34796
rect 23255 34756 23276 34796
rect 23316 34756 23337 34796
rect 23423 34756 23440 34796
rect 23480 34756 23489 34796
rect 23103 34733 23169 34756
rect 23255 34733 23337 34756
rect 23423 34733 23489 34756
rect 23103 34714 23489 34733
rect 27103 34819 27489 34838
rect 27103 34796 27169 34819
rect 27255 34796 27337 34819
rect 27423 34796 27489 34819
rect 27103 34756 27112 34796
rect 27152 34756 27169 34796
rect 27255 34756 27276 34796
rect 27316 34756 27337 34796
rect 27423 34756 27440 34796
rect 27480 34756 27489 34796
rect 27103 34733 27169 34756
rect 27255 34733 27337 34756
rect 27423 34733 27489 34756
rect 27103 34714 27489 34733
rect 31103 34819 31489 34838
rect 31103 34796 31169 34819
rect 31255 34796 31337 34819
rect 31423 34796 31489 34819
rect 31103 34756 31112 34796
rect 31152 34756 31169 34796
rect 31255 34756 31276 34796
rect 31316 34756 31337 34796
rect 31423 34756 31440 34796
rect 31480 34756 31489 34796
rect 31103 34733 31169 34756
rect 31255 34733 31337 34756
rect 31423 34733 31489 34756
rect 31103 34714 31489 34733
rect 35103 34819 35489 34838
rect 35103 34796 35169 34819
rect 35255 34796 35337 34819
rect 35423 34796 35489 34819
rect 35103 34756 35112 34796
rect 35152 34756 35169 34796
rect 35255 34756 35276 34796
rect 35316 34756 35337 34796
rect 35423 34756 35440 34796
rect 35480 34756 35489 34796
rect 35103 34733 35169 34756
rect 35255 34733 35337 34756
rect 35423 34733 35489 34756
rect 35103 34714 35489 34733
rect 39103 34819 39489 34838
rect 39103 34796 39169 34819
rect 39255 34796 39337 34819
rect 39423 34796 39489 34819
rect 39103 34756 39112 34796
rect 39152 34756 39169 34796
rect 39255 34756 39276 34796
rect 39316 34756 39337 34796
rect 39423 34756 39440 34796
rect 39480 34756 39489 34796
rect 39103 34733 39169 34756
rect 39255 34733 39337 34756
rect 39423 34733 39489 34756
rect 39103 34714 39489 34733
rect 43103 34819 43489 34838
rect 43103 34796 43169 34819
rect 43255 34796 43337 34819
rect 43423 34796 43489 34819
rect 43103 34756 43112 34796
rect 43152 34756 43169 34796
rect 43255 34756 43276 34796
rect 43316 34756 43337 34796
rect 43423 34756 43440 34796
rect 43480 34756 43489 34796
rect 43103 34733 43169 34756
rect 43255 34733 43337 34756
rect 43423 34733 43489 34756
rect 43103 34714 43489 34733
rect 47103 34819 47489 34838
rect 47103 34796 47169 34819
rect 47255 34796 47337 34819
rect 47423 34796 47489 34819
rect 47103 34756 47112 34796
rect 47152 34756 47169 34796
rect 47255 34756 47276 34796
rect 47316 34756 47337 34796
rect 47423 34756 47440 34796
rect 47480 34756 47489 34796
rect 47103 34733 47169 34756
rect 47255 34733 47337 34756
rect 47423 34733 47489 34756
rect 47103 34714 47489 34733
rect 51103 34819 51489 34838
rect 51103 34796 51169 34819
rect 51255 34796 51337 34819
rect 51423 34796 51489 34819
rect 51103 34756 51112 34796
rect 51152 34756 51169 34796
rect 51255 34756 51276 34796
rect 51316 34756 51337 34796
rect 51423 34756 51440 34796
rect 51480 34756 51489 34796
rect 51103 34733 51169 34756
rect 51255 34733 51337 34756
rect 51423 34733 51489 34756
rect 51103 34714 51489 34733
rect 55103 34819 55489 34838
rect 55103 34796 55169 34819
rect 55255 34796 55337 34819
rect 55423 34796 55489 34819
rect 55103 34756 55112 34796
rect 55152 34756 55169 34796
rect 55255 34756 55276 34796
rect 55316 34756 55337 34796
rect 55423 34756 55440 34796
rect 55480 34756 55489 34796
rect 55103 34733 55169 34756
rect 55255 34733 55337 34756
rect 55423 34733 55489 34756
rect 55103 34714 55489 34733
rect 59103 34819 59489 34838
rect 59103 34796 59169 34819
rect 59255 34796 59337 34819
rect 59423 34796 59489 34819
rect 59103 34756 59112 34796
rect 59152 34756 59169 34796
rect 59255 34756 59276 34796
rect 59316 34756 59337 34796
rect 59423 34756 59440 34796
rect 59480 34756 59489 34796
rect 59103 34733 59169 34756
rect 59255 34733 59337 34756
rect 59423 34733 59489 34756
rect 59103 34714 59489 34733
rect 63103 34819 63489 34838
rect 63103 34796 63169 34819
rect 63255 34796 63337 34819
rect 63423 34796 63489 34819
rect 63103 34756 63112 34796
rect 63152 34756 63169 34796
rect 63255 34756 63276 34796
rect 63316 34756 63337 34796
rect 63423 34756 63440 34796
rect 63480 34756 63489 34796
rect 63103 34733 63169 34756
rect 63255 34733 63337 34756
rect 63423 34733 63489 34756
rect 63103 34714 63489 34733
rect 67103 34819 67489 34838
rect 67103 34796 67169 34819
rect 67255 34796 67337 34819
rect 67423 34796 67489 34819
rect 67103 34756 67112 34796
rect 67152 34756 67169 34796
rect 67255 34756 67276 34796
rect 67316 34756 67337 34796
rect 67423 34756 67440 34796
rect 67480 34756 67489 34796
rect 67103 34733 67169 34756
rect 67255 34733 67337 34756
rect 67423 34733 67489 34756
rect 67103 34714 67489 34733
rect 71103 34819 71489 34838
rect 71103 34796 71169 34819
rect 71255 34796 71337 34819
rect 71423 34796 71489 34819
rect 71103 34756 71112 34796
rect 71152 34756 71169 34796
rect 71255 34756 71276 34796
rect 71316 34756 71337 34796
rect 71423 34756 71440 34796
rect 71480 34756 71489 34796
rect 71103 34733 71169 34756
rect 71255 34733 71337 34756
rect 71423 34733 71489 34756
rect 71103 34714 71489 34733
rect 75103 34819 75489 34838
rect 75103 34796 75169 34819
rect 75255 34796 75337 34819
rect 75423 34796 75489 34819
rect 75103 34756 75112 34796
rect 75152 34756 75169 34796
rect 75255 34756 75276 34796
rect 75316 34756 75337 34796
rect 75423 34756 75440 34796
rect 75480 34756 75489 34796
rect 75103 34733 75169 34756
rect 75255 34733 75337 34756
rect 75423 34733 75489 34756
rect 75103 34714 75489 34733
rect 79103 34819 79489 34838
rect 79103 34796 79169 34819
rect 79255 34796 79337 34819
rect 79423 34796 79489 34819
rect 79103 34756 79112 34796
rect 79152 34756 79169 34796
rect 79255 34756 79276 34796
rect 79316 34756 79337 34796
rect 79423 34756 79440 34796
rect 79480 34756 79489 34796
rect 79103 34733 79169 34756
rect 79255 34733 79337 34756
rect 79423 34733 79489 34756
rect 79103 34714 79489 34733
rect 83103 34819 83489 34838
rect 83103 34796 83169 34819
rect 83255 34796 83337 34819
rect 83423 34796 83489 34819
rect 83103 34756 83112 34796
rect 83152 34756 83169 34796
rect 83255 34756 83276 34796
rect 83316 34756 83337 34796
rect 83423 34756 83440 34796
rect 83480 34756 83489 34796
rect 83103 34733 83169 34756
rect 83255 34733 83337 34756
rect 83423 34733 83489 34756
rect 83103 34714 83489 34733
rect 87103 34819 87489 34838
rect 87103 34796 87169 34819
rect 87255 34796 87337 34819
rect 87423 34796 87489 34819
rect 87103 34756 87112 34796
rect 87152 34756 87169 34796
rect 87255 34756 87276 34796
rect 87316 34756 87337 34796
rect 87423 34756 87440 34796
rect 87480 34756 87489 34796
rect 87103 34733 87169 34756
rect 87255 34733 87337 34756
rect 87423 34733 87489 34756
rect 87103 34714 87489 34733
rect 91103 34819 91489 34838
rect 91103 34796 91169 34819
rect 91255 34796 91337 34819
rect 91423 34796 91489 34819
rect 91103 34756 91112 34796
rect 91152 34756 91169 34796
rect 91255 34756 91276 34796
rect 91316 34756 91337 34796
rect 91423 34756 91440 34796
rect 91480 34756 91489 34796
rect 91103 34733 91169 34756
rect 91255 34733 91337 34756
rect 91423 34733 91489 34756
rect 91103 34714 91489 34733
rect 95103 34819 95489 34838
rect 95103 34796 95169 34819
rect 95255 34796 95337 34819
rect 95423 34796 95489 34819
rect 95103 34756 95112 34796
rect 95152 34756 95169 34796
rect 95255 34756 95276 34796
rect 95316 34756 95337 34796
rect 95423 34756 95440 34796
rect 95480 34756 95489 34796
rect 95103 34733 95169 34756
rect 95255 34733 95337 34756
rect 95423 34733 95489 34756
rect 95103 34714 95489 34733
rect 99103 34819 99489 34838
rect 99103 34796 99169 34819
rect 99255 34796 99337 34819
rect 99423 34796 99489 34819
rect 99103 34756 99112 34796
rect 99152 34756 99169 34796
rect 99255 34756 99276 34796
rect 99316 34756 99337 34796
rect 99423 34756 99440 34796
rect 99480 34756 99489 34796
rect 99103 34733 99169 34756
rect 99255 34733 99337 34756
rect 99423 34733 99489 34756
rect 99103 34714 99489 34733
rect 4343 34063 4729 34082
rect 4343 34040 4409 34063
rect 4495 34040 4577 34063
rect 4663 34040 4729 34063
rect 4343 34000 4352 34040
rect 4392 34000 4409 34040
rect 4495 34000 4516 34040
rect 4556 34000 4577 34040
rect 4663 34000 4680 34040
rect 4720 34000 4729 34040
rect 4343 33977 4409 34000
rect 4495 33977 4577 34000
rect 4663 33977 4729 34000
rect 4343 33958 4729 33977
rect 8343 34063 8729 34082
rect 8343 34040 8409 34063
rect 8495 34040 8577 34063
rect 8663 34040 8729 34063
rect 8343 34000 8352 34040
rect 8392 34000 8409 34040
rect 8495 34000 8516 34040
rect 8556 34000 8577 34040
rect 8663 34000 8680 34040
rect 8720 34000 8729 34040
rect 8343 33977 8409 34000
rect 8495 33977 8577 34000
rect 8663 33977 8729 34000
rect 8343 33958 8729 33977
rect 12343 34063 12729 34082
rect 12343 34040 12409 34063
rect 12495 34040 12577 34063
rect 12663 34040 12729 34063
rect 12343 34000 12352 34040
rect 12392 34000 12409 34040
rect 12495 34000 12516 34040
rect 12556 34000 12577 34040
rect 12663 34000 12680 34040
rect 12720 34000 12729 34040
rect 12343 33977 12409 34000
rect 12495 33977 12577 34000
rect 12663 33977 12729 34000
rect 12343 33958 12729 33977
rect 16343 34063 16729 34082
rect 16343 34040 16409 34063
rect 16495 34040 16577 34063
rect 16663 34040 16729 34063
rect 16343 34000 16352 34040
rect 16392 34000 16409 34040
rect 16495 34000 16516 34040
rect 16556 34000 16577 34040
rect 16663 34000 16680 34040
rect 16720 34000 16729 34040
rect 16343 33977 16409 34000
rect 16495 33977 16577 34000
rect 16663 33977 16729 34000
rect 16343 33958 16729 33977
rect 20343 34063 20729 34082
rect 20343 34040 20409 34063
rect 20495 34040 20577 34063
rect 20663 34040 20729 34063
rect 20343 34000 20352 34040
rect 20392 34000 20409 34040
rect 20495 34000 20516 34040
rect 20556 34000 20577 34040
rect 20663 34000 20680 34040
rect 20720 34000 20729 34040
rect 20343 33977 20409 34000
rect 20495 33977 20577 34000
rect 20663 33977 20729 34000
rect 20343 33958 20729 33977
rect 24343 34063 24729 34082
rect 24343 34040 24409 34063
rect 24495 34040 24577 34063
rect 24663 34040 24729 34063
rect 24343 34000 24352 34040
rect 24392 34000 24409 34040
rect 24495 34000 24516 34040
rect 24556 34000 24577 34040
rect 24663 34000 24680 34040
rect 24720 34000 24729 34040
rect 24343 33977 24409 34000
rect 24495 33977 24577 34000
rect 24663 33977 24729 34000
rect 24343 33958 24729 33977
rect 28343 34063 28729 34082
rect 28343 34040 28409 34063
rect 28495 34040 28577 34063
rect 28663 34040 28729 34063
rect 28343 34000 28352 34040
rect 28392 34000 28409 34040
rect 28495 34000 28516 34040
rect 28556 34000 28577 34040
rect 28663 34000 28680 34040
rect 28720 34000 28729 34040
rect 28343 33977 28409 34000
rect 28495 33977 28577 34000
rect 28663 33977 28729 34000
rect 28343 33958 28729 33977
rect 32343 34063 32729 34082
rect 32343 34040 32409 34063
rect 32495 34040 32577 34063
rect 32663 34040 32729 34063
rect 32343 34000 32352 34040
rect 32392 34000 32409 34040
rect 32495 34000 32516 34040
rect 32556 34000 32577 34040
rect 32663 34000 32680 34040
rect 32720 34000 32729 34040
rect 32343 33977 32409 34000
rect 32495 33977 32577 34000
rect 32663 33977 32729 34000
rect 32343 33958 32729 33977
rect 36343 34063 36729 34082
rect 36343 34040 36409 34063
rect 36495 34040 36577 34063
rect 36663 34040 36729 34063
rect 36343 34000 36352 34040
rect 36392 34000 36409 34040
rect 36495 34000 36516 34040
rect 36556 34000 36577 34040
rect 36663 34000 36680 34040
rect 36720 34000 36729 34040
rect 36343 33977 36409 34000
rect 36495 33977 36577 34000
rect 36663 33977 36729 34000
rect 36343 33958 36729 33977
rect 40343 34063 40729 34082
rect 40343 34040 40409 34063
rect 40495 34040 40577 34063
rect 40663 34040 40729 34063
rect 40343 34000 40352 34040
rect 40392 34000 40409 34040
rect 40495 34000 40516 34040
rect 40556 34000 40577 34040
rect 40663 34000 40680 34040
rect 40720 34000 40729 34040
rect 40343 33977 40409 34000
rect 40495 33977 40577 34000
rect 40663 33977 40729 34000
rect 40343 33958 40729 33977
rect 44343 34063 44729 34082
rect 44343 34040 44409 34063
rect 44495 34040 44577 34063
rect 44663 34040 44729 34063
rect 44343 34000 44352 34040
rect 44392 34000 44409 34040
rect 44495 34000 44516 34040
rect 44556 34000 44577 34040
rect 44663 34000 44680 34040
rect 44720 34000 44729 34040
rect 44343 33977 44409 34000
rect 44495 33977 44577 34000
rect 44663 33977 44729 34000
rect 44343 33958 44729 33977
rect 48343 34063 48729 34082
rect 48343 34040 48409 34063
rect 48495 34040 48577 34063
rect 48663 34040 48729 34063
rect 48343 34000 48352 34040
rect 48392 34000 48409 34040
rect 48495 34000 48516 34040
rect 48556 34000 48577 34040
rect 48663 34000 48680 34040
rect 48720 34000 48729 34040
rect 48343 33977 48409 34000
rect 48495 33977 48577 34000
rect 48663 33977 48729 34000
rect 48343 33958 48729 33977
rect 52343 34063 52729 34082
rect 52343 34040 52409 34063
rect 52495 34040 52577 34063
rect 52663 34040 52729 34063
rect 52343 34000 52352 34040
rect 52392 34000 52409 34040
rect 52495 34000 52516 34040
rect 52556 34000 52577 34040
rect 52663 34000 52680 34040
rect 52720 34000 52729 34040
rect 52343 33977 52409 34000
rect 52495 33977 52577 34000
rect 52663 33977 52729 34000
rect 52343 33958 52729 33977
rect 56343 34063 56729 34082
rect 56343 34040 56409 34063
rect 56495 34040 56577 34063
rect 56663 34040 56729 34063
rect 56343 34000 56352 34040
rect 56392 34000 56409 34040
rect 56495 34000 56516 34040
rect 56556 34000 56577 34040
rect 56663 34000 56680 34040
rect 56720 34000 56729 34040
rect 56343 33977 56409 34000
rect 56495 33977 56577 34000
rect 56663 33977 56729 34000
rect 56343 33958 56729 33977
rect 60343 34063 60729 34082
rect 60343 34040 60409 34063
rect 60495 34040 60577 34063
rect 60663 34040 60729 34063
rect 60343 34000 60352 34040
rect 60392 34000 60409 34040
rect 60495 34000 60516 34040
rect 60556 34000 60577 34040
rect 60663 34000 60680 34040
rect 60720 34000 60729 34040
rect 60343 33977 60409 34000
rect 60495 33977 60577 34000
rect 60663 33977 60729 34000
rect 60343 33958 60729 33977
rect 64343 34063 64729 34082
rect 64343 34040 64409 34063
rect 64495 34040 64577 34063
rect 64663 34040 64729 34063
rect 64343 34000 64352 34040
rect 64392 34000 64409 34040
rect 64495 34000 64516 34040
rect 64556 34000 64577 34040
rect 64663 34000 64680 34040
rect 64720 34000 64729 34040
rect 64343 33977 64409 34000
rect 64495 33977 64577 34000
rect 64663 33977 64729 34000
rect 64343 33958 64729 33977
rect 68343 34063 68729 34082
rect 68343 34040 68409 34063
rect 68495 34040 68577 34063
rect 68663 34040 68729 34063
rect 68343 34000 68352 34040
rect 68392 34000 68409 34040
rect 68495 34000 68516 34040
rect 68556 34000 68577 34040
rect 68663 34000 68680 34040
rect 68720 34000 68729 34040
rect 68343 33977 68409 34000
rect 68495 33977 68577 34000
rect 68663 33977 68729 34000
rect 68343 33958 68729 33977
rect 72343 34063 72729 34082
rect 72343 34040 72409 34063
rect 72495 34040 72577 34063
rect 72663 34040 72729 34063
rect 72343 34000 72352 34040
rect 72392 34000 72409 34040
rect 72495 34000 72516 34040
rect 72556 34000 72577 34040
rect 72663 34000 72680 34040
rect 72720 34000 72729 34040
rect 72343 33977 72409 34000
rect 72495 33977 72577 34000
rect 72663 33977 72729 34000
rect 72343 33958 72729 33977
rect 76343 34063 76729 34082
rect 76343 34040 76409 34063
rect 76495 34040 76577 34063
rect 76663 34040 76729 34063
rect 76343 34000 76352 34040
rect 76392 34000 76409 34040
rect 76495 34000 76516 34040
rect 76556 34000 76577 34040
rect 76663 34000 76680 34040
rect 76720 34000 76729 34040
rect 76343 33977 76409 34000
rect 76495 33977 76577 34000
rect 76663 33977 76729 34000
rect 76343 33958 76729 33977
rect 80343 34063 80729 34082
rect 80343 34040 80409 34063
rect 80495 34040 80577 34063
rect 80663 34040 80729 34063
rect 80343 34000 80352 34040
rect 80392 34000 80409 34040
rect 80495 34000 80516 34040
rect 80556 34000 80577 34040
rect 80663 34000 80680 34040
rect 80720 34000 80729 34040
rect 80343 33977 80409 34000
rect 80495 33977 80577 34000
rect 80663 33977 80729 34000
rect 80343 33958 80729 33977
rect 84343 34063 84729 34082
rect 84343 34040 84409 34063
rect 84495 34040 84577 34063
rect 84663 34040 84729 34063
rect 84343 34000 84352 34040
rect 84392 34000 84409 34040
rect 84495 34000 84516 34040
rect 84556 34000 84577 34040
rect 84663 34000 84680 34040
rect 84720 34000 84729 34040
rect 84343 33977 84409 34000
rect 84495 33977 84577 34000
rect 84663 33977 84729 34000
rect 84343 33958 84729 33977
rect 88343 34063 88729 34082
rect 88343 34040 88409 34063
rect 88495 34040 88577 34063
rect 88663 34040 88729 34063
rect 88343 34000 88352 34040
rect 88392 34000 88409 34040
rect 88495 34000 88516 34040
rect 88556 34000 88577 34040
rect 88663 34000 88680 34040
rect 88720 34000 88729 34040
rect 88343 33977 88409 34000
rect 88495 33977 88577 34000
rect 88663 33977 88729 34000
rect 88343 33958 88729 33977
rect 92343 34063 92729 34082
rect 92343 34040 92409 34063
rect 92495 34040 92577 34063
rect 92663 34040 92729 34063
rect 92343 34000 92352 34040
rect 92392 34000 92409 34040
rect 92495 34000 92516 34040
rect 92556 34000 92577 34040
rect 92663 34000 92680 34040
rect 92720 34000 92729 34040
rect 92343 33977 92409 34000
rect 92495 33977 92577 34000
rect 92663 33977 92729 34000
rect 92343 33958 92729 33977
rect 96343 34063 96729 34082
rect 96343 34040 96409 34063
rect 96495 34040 96577 34063
rect 96663 34040 96729 34063
rect 96343 34000 96352 34040
rect 96392 34000 96409 34040
rect 96495 34000 96516 34040
rect 96556 34000 96577 34040
rect 96663 34000 96680 34040
rect 96720 34000 96729 34040
rect 96343 33977 96409 34000
rect 96495 33977 96577 34000
rect 96663 33977 96729 34000
rect 96343 33958 96729 33977
rect 3103 33307 3489 33326
rect 3103 33284 3169 33307
rect 3255 33284 3337 33307
rect 3423 33284 3489 33307
rect 3103 33244 3112 33284
rect 3152 33244 3169 33284
rect 3255 33244 3276 33284
rect 3316 33244 3337 33284
rect 3423 33244 3440 33284
rect 3480 33244 3489 33284
rect 3103 33221 3169 33244
rect 3255 33221 3337 33244
rect 3423 33221 3489 33244
rect 3103 33202 3489 33221
rect 7103 33307 7489 33326
rect 7103 33284 7169 33307
rect 7255 33284 7337 33307
rect 7423 33284 7489 33307
rect 7103 33244 7112 33284
rect 7152 33244 7169 33284
rect 7255 33244 7276 33284
rect 7316 33244 7337 33284
rect 7423 33244 7440 33284
rect 7480 33244 7489 33284
rect 7103 33221 7169 33244
rect 7255 33221 7337 33244
rect 7423 33221 7489 33244
rect 7103 33202 7489 33221
rect 11103 33307 11489 33326
rect 11103 33284 11169 33307
rect 11255 33284 11337 33307
rect 11423 33284 11489 33307
rect 11103 33244 11112 33284
rect 11152 33244 11169 33284
rect 11255 33244 11276 33284
rect 11316 33244 11337 33284
rect 11423 33244 11440 33284
rect 11480 33244 11489 33284
rect 11103 33221 11169 33244
rect 11255 33221 11337 33244
rect 11423 33221 11489 33244
rect 11103 33202 11489 33221
rect 15103 33307 15489 33326
rect 15103 33284 15169 33307
rect 15255 33284 15337 33307
rect 15423 33284 15489 33307
rect 15103 33244 15112 33284
rect 15152 33244 15169 33284
rect 15255 33244 15276 33284
rect 15316 33244 15337 33284
rect 15423 33244 15440 33284
rect 15480 33244 15489 33284
rect 15103 33221 15169 33244
rect 15255 33221 15337 33244
rect 15423 33221 15489 33244
rect 15103 33202 15489 33221
rect 19103 33307 19489 33326
rect 19103 33284 19169 33307
rect 19255 33284 19337 33307
rect 19423 33284 19489 33307
rect 19103 33244 19112 33284
rect 19152 33244 19169 33284
rect 19255 33244 19276 33284
rect 19316 33244 19337 33284
rect 19423 33244 19440 33284
rect 19480 33244 19489 33284
rect 19103 33221 19169 33244
rect 19255 33221 19337 33244
rect 19423 33221 19489 33244
rect 19103 33202 19489 33221
rect 23103 33307 23489 33326
rect 23103 33284 23169 33307
rect 23255 33284 23337 33307
rect 23423 33284 23489 33307
rect 23103 33244 23112 33284
rect 23152 33244 23169 33284
rect 23255 33244 23276 33284
rect 23316 33244 23337 33284
rect 23423 33244 23440 33284
rect 23480 33244 23489 33284
rect 23103 33221 23169 33244
rect 23255 33221 23337 33244
rect 23423 33221 23489 33244
rect 23103 33202 23489 33221
rect 27103 33307 27489 33326
rect 27103 33284 27169 33307
rect 27255 33284 27337 33307
rect 27423 33284 27489 33307
rect 27103 33244 27112 33284
rect 27152 33244 27169 33284
rect 27255 33244 27276 33284
rect 27316 33244 27337 33284
rect 27423 33244 27440 33284
rect 27480 33244 27489 33284
rect 27103 33221 27169 33244
rect 27255 33221 27337 33244
rect 27423 33221 27489 33244
rect 27103 33202 27489 33221
rect 31103 33307 31489 33326
rect 31103 33284 31169 33307
rect 31255 33284 31337 33307
rect 31423 33284 31489 33307
rect 31103 33244 31112 33284
rect 31152 33244 31169 33284
rect 31255 33244 31276 33284
rect 31316 33244 31337 33284
rect 31423 33244 31440 33284
rect 31480 33244 31489 33284
rect 31103 33221 31169 33244
rect 31255 33221 31337 33244
rect 31423 33221 31489 33244
rect 31103 33202 31489 33221
rect 35103 33307 35489 33326
rect 35103 33284 35169 33307
rect 35255 33284 35337 33307
rect 35423 33284 35489 33307
rect 35103 33244 35112 33284
rect 35152 33244 35169 33284
rect 35255 33244 35276 33284
rect 35316 33244 35337 33284
rect 35423 33244 35440 33284
rect 35480 33244 35489 33284
rect 35103 33221 35169 33244
rect 35255 33221 35337 33244
rect 35423 33221 35489 33244
rect 35103 33202 35489 33221
rect 39103 33307 39489 33326
rect 39103 33284 39169 33307
rect 39255 33284 39337 33307
rect 39423 33284 39489 33307
rect 39103 33244 39112 33284
rect 39152 33244 39169 33284
rect 39255 33244 39276 33284
rect 39316 33244 39337 33284
rect 39423 33244 39440 33284
rect 39480 33244 39489 33284
rect 39103 33221 39169 33244
rect 39255 33221 39337 33244
rect 39423 33221 39489 33244
rect 39103 33202 39489 33221
rect 43103 33307 43489 33326
rect 43103 33284 43169 33307
rect 43255 33284 43337 33307
rect 43423 33284 43489 33307
rect 43103 33244 43112 33284
rect 43152 33244 43169 33284
rect 43255 33244 43276 33284
rect 43316 33244 43337 33284
rect 43423 33244 43440 33284
rect 43480 33244 43489 33284
rect 43103 33221 43169 33244
rect 43255 33221 43337 33244
rect 43423 33221 43489 33244
rect 43103 33202 43489 33221
rect 47103 33307 47489 33326
rect 47103 33284 47169 33307
rect 47255 33284 47337 33307
rect 47423 33284 47489 33307
rect 47103 33244 47112 33284
rect 47152 33244 47169 33284
rect 47255 33244 47276 33284
rect 47316 33244 47337 33284
rect 47423 33244 47440 33284
rect 47480 33244 47489 33284
rect 47103 33221 47169 33244
rect 47255 33221 47337 33244
rect 47423 33221 47489 33244
rect 47103 33202 47489 33221
rect 51103 33307 51489 33326
rect 51103 33284 51169 33307
rect 51255 33284 51337 33307
rect 51423 33284 51489 33307
rect 51103 33244 51112 33284
rect 51152 33244 51169 33284
rect 51255 33244 51276 33284
rect 51316 33244 51337 33284
rect 51423 33244 51440 33284
rect 51480 33244 51489 33284
rect 51103 33221 51169 33244
rect 51255 33221 51337 33244
rect 51423 33221 51489 33244
rect 51103 33202 51489 33221
rect 55103 33307 55489 33326
rect 55103 33284 55169 33307
rect 55255 33284 55337 33307
rect 55423 33284 55489 33307
rect 55103 33244 55112 33284
rect 55152 33244 55169 33284
rect 55255 33244 55276 33284
rect 55316 33244 55337 33284
rect 55423 33244 55440 33284
rect 55480 33244 55489 33284
rect 55103 33221 55169 33244
rect 55255 33221 55337 33244
rect 55423 33221 55489 33244
rect 55103 33202 55489 33221
rect 59103 33307 59489 33326
rect 59103 33284 59169 33307
rect 59255 33284 59337 33307
rect 59423 33284 59489 33307
rect 59103 33244 59112 33284
rect 59152 33244 59169 33284
rect 59255 33244 59276 33284
rect 59316 33244 59337 33284
rect 59423 33244 59440 33284
rect 59480 33244 59489 33284
rect 59103 33221 59169 33244
rect 59255 33221 59337 33244
rect 59423 33221 59489 33244
rect 59103 33202 59489 33221
rect 63103 33307 63489 33326
rect 63103 33284 63169 33307
rect 63255 33284 63337 33307
rect 63423 33284 63489 33307
rect 63103 33244 63112 33284
rect 63152 33244 63169 33284
rect 63255 33244 63276 33284
rect 63316 33244 63337 33284
rect 63423 33244 63440 33284
rect 63480 33244 63489 33284
rect 63103 33221 63169 33244
rect 63255 33221 63337 33244
rect 63423 33221 63489 33244
rect 63103 33202 63489 33221
rect 67103 33307 67489 33326
rect 67103 33284 67169 33307
rect 67255 33284 67337 33307
rect 67423 33284 67489 33307
rect 67103 33244 67112 33284
rect 67152 33244 67169 33284
rect 67255 33244 67276 33284
rect 67316 33244 67337 33284
rect 67423 33244 67440 33284
rect 67480 33244 67489 33284
rect 67103 33221 67169 33244
rect 67255 33221 67337 33244
rect 67423 33221 67489 33244
rect 67103 33202 67489 33221
rect 4343 32551 4729 32570
rect 4343 32528 4409 32551
rect 4495 32528 4577 32551
rect 4663 32528 4729 32551
rect 4343 32488 4352 32528
rect 4392 32488 4409 32528
rect 4495 32488 4516 32528
rect 4556 32488 4577 32528
rect 4663 32488 4680 32528
rect 4720 32488 4729 32528
rect 4343 32465 4409 32488
rect 4495 32465 4577 32488
rect 4663 32465 4729 32488
rect 4343 32446 4729 32465
rect 8343 32551 8729 32570
rect 8343 32528 8409 32551
rect 8495 32528 8577 32551
rect 8663 32528 8729 32551
rect 8343 32488 8352 32528
rect 8392 32488 8409 32528
rect 8495 32488 8516 32528
rect 8556 32488 8577 32528
rect 8663 32488 8680 32528
rect 8720 32488 8729 32528
rect 8343 32465 8409 32488
rect 8495 32465 8577 32488
rect 8663 32465 8729 32488
rect 8343 32446 8729 32465
rect 12343 32551 12729 32570
rect 12343 32528 12409 32551
rect 12495 32528 12577 32551
rect 12663 32528 12729 32551
rect 12343 32488 12352 32528
rect 12392 32488 12409 32528
rect 12495 32488 12516 32528
rect 12556 32488 12577 32528
rect 12663 32488 12680 32528
rect 12720 32488 12729 32528
rect 12343 32465 12409 32488
rect 12495 32465 12577 32488
rect 12663 32465 12729 32488
rect 12343 32446 12729 32465
rect 16343 32551 16729 32570
rect 16343 32528 16409 32551
rect 16495 32528 16577 32551
rect 16663 32528 16729 32551
rect 16343 32488 16352 32528
rect 16392 32488 16409 32528
rect 16495 32488 16516 32528
rect 16556 32488 16577 32528
rect 16663 32488 16680 32528
rect 16720 32488 16729 32528
rect 16343 32465 16409 32488
rect 16495 32465 16577 32488
rect 16663 32465 16729 32488
rect 16343 32446 16729 32465
rect 20343 32551 20729 32570
rect 20343 32528 20409 32551
rect 20495 32528 20577 32551
rect 20663 32528 20729 32551
rect 20343 32488 20352 32528
rect 20392 32488 20409 32528
rect 20495 32488 20516 32528
rect 20556 32488 20577 32528
rect 20663 32488 20680 32528
rect 20720 32488 20729 32528
rect 20343 32465 20409 32488
rect 20495 32465 20577 32488
rect 20663 32465 20729 32488
rect 20343 32446 20729 32465
rect 24343 32551 24729 32570
rect 24343 32528 24409 32551
rect 24495 32528 24577 32551
rect 24663 32528 24729 32551
rect 24343 32488 24352 32528
rect 24392 32488 24409 32528
rect 24495 32488 24516 32528
rect 24556 32488 24577 32528
rect 24663 32488 24680 32528
rect 24720 32488 24729 32528
rect 24343 32465 24409 32488
rect 24495 32465 24577 32488
rect 24663 32465 24729 32488
rect 24343 32446 24729 32465
rect 28343 32551 28729 32570
rect 28343 32528 28409 32551
rect 28495 32528 28577 32551
rect 28663 32528 28729 32551
rect 28343 32488 28352 32528
rect 28392 32488 28409 32528
rect 28495 32488 28516 32528
rect 28556 32488 28577 32528
rect 28663 32488 28680 32528
rect 28720 32488 28729 32528
rect 28343 32465 28409 32488
rect 28495 32465 28577 32488
rect 28663 32465 28729 32488
rect 28343 32446 28729 32465
rect 32343 32551 32729 32570
rect 32343 32528 32409 32551
rect 32495 32528 32577 32551
rect 32663 32528 32729 32551
rect 32343 32488 32352 32528
rect 32392 32488 32409 32528
rect 32495 32488 32516 32528
rect 32556 32488 32577 32528
rect 32663 32488 32680 32528
rect 32720 32488 32729 32528
rect 32343 32465 32409 32488
rect 32495 32465 32577 32488
rect 32663 32465 32729 32488
rect 32343 32446 32729 32465
rect 36343 32551 36729 32570
rect 36343 32528 36409 32551
rect 36495 32528 36577 32551
rect 36663 32528 36729 32551
rect 36343 32488 36352 32528
rect 36392 32488 36409 32528
rect 36495 32488 36516 32528
rect 36556 32488 36577 32528
rect 36663 32488 36680 32528
rect 36720 32488 36729 32528
rect 36343 32465 36409 32488
rect 36495 32465 36577 32488
rect 36663 32465 36729 32488
rect 36343 32446 36729 32465
rect 40343 32551 40729 32570
rect 40343 32528 40409 32551
rect 40495 32528 40577 32551
rect 40663 32528 40729 32551
rect 40343 32488 40352 32528
rect 40392 32488 40409 32528
rect 40495 32488 40516 32528
rect 40556 32488 40577 32528
rect 40663 32488 40680 32528
rect 40720 32488 40729 32528
rect 40343 32465 40409 32488
rect 40495 32465 40577 32488
rect 40663 32465 40729 32488
rect 40343 32446 40729 32465
rect 44343 32551 44729 32570
rect 44343 32528 44409 32551
rect 44495 32528 44577 32551
rect 44663 32528 44729 32551
rect 44343 32488 44352 32528
rect 44392 32488 44409 32528
rect 44495 32488 44516 32528
rect 44556 32488 44577 32528
rect 44663 32488 44680 32528
rect 44720 32488 44729 32528
rect 44343 32465 44409 32488
rect 44495 32465 44577 32488
rect 44663 32465 44729 32488
rect 44343 32446 44729 32465
rect 48343 32551 48729 32570
rect 48343 32528 48409 32551
rect 48495 32528 48577 32551
rect 48663 32528 48729 32551
rect 48343 32488 48352 32528
rect 48392 32488 48409 32528
rect 48495 32488 48516 32528
rect 48556 32488 48577 32528
rect 48663 32488 48680 32528
rect 48720 32488 48729 32528
rect 48343 32465 48409 32488
rect 48495 32465 48577 32488
rect 48663 32465 48729 32488
rect 48343 32446 48729 32465
rect 52343 32551 52729 32570
rect 52343 32528 52409 32551
rect 52495 32528 52577 32551
rect 52663 32528 52729 32551
rect 52343 32488 52352 32528
rect 52392 32488 52409 32528
rect 52495 32488 52516 32528
rect 52556 32488 52577 32528
rect 52663 32488 52680 32528
rect 52720 32488 52729 32528
rect 52343 32465 52409 32488
rect 52495 32465 52577 32488
rect 52663 32465 52729 32488
rect 52343 32446 52729 32465
rect 56343 32551 56729 32570
rect 56343 32528 56409 32551
rect 56495 32528 56577 32551
rect 56663 32528 56729 32551
rect 56343 32488 56352 32528
rect 56392 32488 56409 32528
rect 56495 32488 56516 32528
rect 56556 32488 56577 32528
rect 56663 32488 56680 32528
rect 56720 32488 56729 32528
rect 56343 32465 56409 32488
rect 56495 32465 56577 32488
rect 56663 32465 56729 32488
rect 56343 32446 56729 32465
rect 60343 32551 60729 32570
rect 60343 32528 60409 32551
rect 60495 32528 60577 32551
rect 60663 32528 60729 32551
rect 60343 32488 60352 32528
rect 60392 32488 60409 32528
rect 60495 32488 60516 32528
rect 60556 32488 60577 32528
rect 60663 32488 60680 32528
rect 60720 32488 60729 32528
rect 60343 32465 60409 32488
rect 60495 32465 60577 32488
rect 60663 32465 60729 32488
rect 60343 32446 60729 32465
rect 64343 32551 64729 32570
rect 64343 32528 64409 32551
rect 64495 32528 64577 32551
rect 64663 32528 64729 32551
rect 64343 32488 64352 32528
rect 64392 32488 64409 32528
rect 64495 32488 64516 32528
rect 64556 32488 64577 32528
rect 64663 32488 64680 32528
rect 64720 32488 64729 32528
rect 64343 32465 64409 32488
rect 64495 32465 64577 32488
rect 64663 32465 64729 32488
rect 64343 32446 64729 32465
rect 68343 32551 68729 32570
rect 68343 32528 68409 32551
rect 68495 32528 68577 32551
rect 68663 32528 68729 32551
rect 68343 32488 68352 32528
rect 68392 32488 68409 32528
rect 68495 32488 68516 32528
rect 68556 32488 68577 32528
rect 68663 32488 68680 32528
rect 68720 32488 68729 32528
rect 68343 32465 68409 32488
rect 68495 32465 68577 32488
rect 68663 32465 68729 32488
rect 68343 32446 68729 32465
rect 3103 31795 3489 31814
rect 3103 31772 3169 31795
rect 3255 31772 3337 31795
rect 3423 31772 3489 31795
rect 3103 31732 3112 31772
rect 3152 31732 3169 31772
rect 3255 31732 3276 31772
rect 3316 31732 3337 31772
rect 3423 31732 3440 31772
rect 3480 31732 3489 31772
rect 3103 31709 3169 31732
rect 3255 31709 3337 31732
rect 3423 31709 3489 31732
rect 3103 31690 3489 31709
rect 7103 31795 7489 31814
rect 7103 31772 7169 31795
rect 7255 31772 7337 31795
rect 7423 31772 7489 31795
rect 7103 31732 7112 31772
rect 7152 31732 7169 31772
rect 7255 31732 7276 31772
rect 7316 31732 7337 31772
rect 7423 31732 7440 31772
rect 7480 31732 7489 31772
rect 7103 31709 7169 31732
rect 7255 31709 7337 31732
rect 7423 31709 7489 31732
rect 7103 31690 7489 31709
rect 11103 31795 11489 31814
rect 11103 31772 11169 31795
rect 11255 31772 11337 31795
rect 11423 31772 11489 31795
rect 11103 31732 11112 31772
rect 11152 31732 11169 31772
rect 11255 31732 11276 31772
rect 11316 31732 11337 31772
rect 11423 31732 11440 31772
rect 11480 31732 11489 31772
rect 11103 31709 11169 31732
rect 11255 31709 11337 31732
rect 11423 31709 11489 31732
rect 11103 31690 11489 31709
rect 15103 31795 15489 31814
rect 15103 31772 15169 31795
rect 15255 31772 15337 31795
rect 15423 31772 15489 31795
rect 15103 31732 15112 31772
rect 15152 31732 15169 31772
rect 15255 31732 15276 31772
rect 15316 31732 15337 31772
rect 15423 31732 15440 31772
rect 15480 31732 15489 31772
rect 15103 31709 15169 31732
rect 15255 31709 15337 31732
rect 15423 31709 15489 31732
rect 15103 31690 15489 31709
rect 19103 31795 19489 31814
rect 19103 31772 19169 31795
rect 19255 31772 19337 31795
rect 19423 31772 19489 31795
rect 19103 31732 19112 31772
rect 19152 31732 19169 31772
rect 19255 31732 19276 31772
rect 19316 31732 19337 31772
rect 19423 31732 19440 31772
rect 19480 31732 19489 31772
rect 19103 31709 19169 31732
rect 19255 31709 19337 31732
rect 19423 31709 19489 31732
rect 19103 31690 19489 31709
rect 23103 31795 23489 31814
rect 23103 31772 23169 31795
rect 23255 31772 23337 31795
rect 23423 31772 23489 31795
rect 23103 31732 23112 31772
rect 23152 31732 23169 31772
rect 23255 31732 23276 31772
rect 23316 31732 23337 31772
rect 23423 31732 23440 31772
rect 23480 31732 23489 31772
rect 23103 31709 23169 31732
rect 23255 31709 23337 31732
rect 23423 31709 23489 31732
rect 23103 31690 23489 31709
rect 27103 31795 27489 31814
rect 27103 31772 27169 31795
rect 27255 31772 27337 31795
rect 27423 31772 27489 31795
rect 27103 31732 27112 31772
rect 27152 31732 27169 31772
rect 27255 31732 27276 31772
rect 27316 31732 27337 31772
rect 27423 31732 27440 31772
rect 27480 31732 27489 31772
rect 27103 31709 27169 31732
rect 27255 31709 27337 31732
rect 27423 31709 27489 31732
rect 27103 31690 27489 31709
rect 31103 31795 31489 31814
rect 31103 31772 31169 31795
rect 31255 31772 31337 31795
rect 31423 31772 31489 31795
rect 31103 31732 31112 31772
rect 31152 31732 31169 31772
rect 31255 31732 31276 31772
rect 31316 31732 31337 31772
rect 31423 31732 31440 31772
rect 31480 31732 31489 31772
rect 31103 31709 31169 31732
rect 31255 31709 31337 31732
rect 31423 31709 31489 31732
rect 31103 31690 31489 31709
rect 35103 31795 35489 31814
rect 35103 31772 35169 31795
rect 35255 31772 35337 31795
rect 35423 31772 35489 31795
rect 35103 31732 35112 31772
rect 35152 31732 35169 31772
rect 35255 31732 35276 31772
rect 35316 31732 35337 31772
rect 35423 31732 35440 31772
rect 35480 31732 35489 31772
rect 35103 31709 35169 31732
rect 35255 31709 35337 31732
rect 35423 31709 35489 31732
rect 35103 31690 35489 31709
rect 39103 31795 39489 31814
rect 39103 31772 39169 31795
rect 39255 31772 39337 31795
rect 39423 31772 39489 31795
rect 39103 31732 39112 31772
rect 39152 31732 39169 31772
rect 39255 31732 39276 31772
rect 39316 31732 39337 31772
rect 39423 31732 39440 31772
rect 39480 31732 39489 31772
rect 39103 31709 39169 31732
rect 39255 31709 39337 31732
rect 39423 31709 39489 31732
rect 39103 31690 39489 31709
rect 43103 31795 43489 31814
rect 43103 31772 43169 31795
rect 43255 31772 43337 31795
rect 43423 31772 43489 31795
rect 43103 31732 43112 31772
rect 43152 31732 43169 31772
rect 43255 31732 43276 31772
rect 43316 31732 43337 31772
rect 43423 31732 43440 31772
rect 43480 31732 43489 31772
rect 43103 31709 43169 31732
rect 43255 31709 43337 31732
rect 43423 31709 43489 31732
rect 43103 31690 43489 31709
rect 47103 31795 47489 31814
rect 47103 31772 47169 31795
rect 47255 31772 47337 31795
rect 47423 31772 47489 31795
rect 47103 31732 47112 31772
rect 47152 31732 47169 31772
rect 47255 31732 47276 31772
rect 47316 31732 47337 31772
rect 47423 31732 47440 31772
rect 47480 31732 47489 31772
rect 47103 31709 47169 31732
rect 47255 31709 47337 31732
rect 47423 31709 47489 31732
rect 47103 31690 47489 31709
rect 51103 31795 51489 31814
rect 51103 31772 51169 31795
rect 51255 31772 51337 31795
rect 51423 31772 51489 31795
rect 51103 31732 51112 31772
rect 51152 31732 51169 31772
rect 51255 31732 51276 31772
rect 51316 31732 51337 31772
rect 51423 31732 51440 31772
rect 51480 31732 51489 31772
rect 51103 31709 51169 31732
rect 51255 31709 51337 31732
rect 51423 31709 51489 31732
rect 51103 31690 51489 31709
rect 55103 31795 55489 31814
rect 55103 31772 55169 31795
rect 55255 31772 55337 31795
rect 55423 31772 55489 31795
rect 55103 31732 55112 31772
rect 55152 31732 55169 31772
rect 55255 31732 55276 31772
rect 55316 31732 55337 31772
rect 55423 31732 55440 31772
rect 55480 31732 55489 31772
rect 55103 31709 55169 31732
rect 55255 31709 55337 31732
rect 55423 31709 55489 31732
rect 55103 31690 55489 31709
rect 59103 31795 59489 31814
rect 59103 31772 59169 31795
rect 59255 31772 59337 31795
rect 59423 31772 59489 31795
rect 59103 31732 59112 31772
rect 59152 31732 59169 31772
rect 59255 31732 59276 31772
rect 59316 31732 59337 31772
rect 59423 31732 59440 31772
rect 59480 31732 59489 31772
rect 59103 31709 59169 31732
rect 59255 31709 59337 31732
rect 59423 31709 59489 31732
rect 59103 31690 59489 31709
rect 63103 31795 63489 31814
rect 63103 31772 63169 31795
rect 63255 31772 63337 31795
rect 63423 31772 63489 31795
rect 63103 31732 63112 31772
rect 63152 31732 63169 31772
rect 63255 31732 63276 31772
rect 63316 31732 63337 31772
rect 63423 31732 63440 31772
rect 63480 31732 63489 31772
rect 63103 31709 63169 31732
rect 63255 31709 63337 31732
rect 63423 31709 63489 31732
rect 63103 31690 63489 31709
rect 67103 31795 67489 31814
rect 67103 31772 67169 31795
rect 67255 31772 67337 31795
rect 67423 31772 67489 31795
rect 67103 31732 67112 31772
rect 67152 31732 67169 31772
rect 67255 31732 67276 31772
rect 67316 31732 67337 31772
rect 67423 31732 67440 31772
rect 67480 31732 67489 31772
rect 67103 31709 67169 31732
rect 67255 31709 67337 31732
rect 67423 31709 67489 31732
rect 67103 31690 67489 31709
rect 72316 31122 72756 31252
rect 4343 31039 4729 31058
rect 4343 31016 4409 31039
rect 4495 31016 4577 31039
rect 4663 31016 4729 31039
rect 4343 30976 4352 31016
rect 4392 30976 4409 31016
rect 4495 30976 4516 31016
rect 4556 30976 4577 31016
rect 4663 30976 4680 31016
rect 4720 30976 4729 31016
rect 4343 30953 4409 30976
rect 4495 30953 4577 30976
rect 4663 30953 4729 30976
rect 4343 30934 4729 30953
rect 8343 31039 8729 31058
rect 8343 31016 8409 31039
rect 8495 31016 8577 31039
rect 8663 31016 8729 31039
rect 8343 30976 8352 31016
rect 8392 30976 8409 31016
rect 8495 30976 8516 31016
rect 8556 30976 8577 31016
rect 8663 30976 8680 31016
rect 8720 30976 8729 31016
rect 8343 30953 8409 30976
rect 8495 30953 8577 30976
rect 8663 30953 8729 30976
rect 8343 30934 8729 30953
rect 12343 31039 12729 31058
rect 12343 31016 12409 31039
rect 12495 31016 12577 31039
rect 12663 31016 12729 31039
rect 12343 30976 12352 31016
rect 12392 30976 12409 31016
rect 12495 30976 12516 31016
rect 12556 30976 12577 31016
rect 12663 30976 12680 31016
rect 12720 30976 12729 31016
rect 12343 30953 12409 30976
rect 12495 30953 12577 30976
rect 12663 30953 12729 30976
rect 12343 30934 12729 30953
rect 16343 31039 16729 31058
rect 16343 31016 16409 31039
rect 16495 31016 16577 31039
rect 16663 31016 16729 31039
rect 16343 30976 16352 31016
rect 16392 30976 16409 31016
rect 16495 30976 16516 31016
rect 16556 30976 16577 31016
rect 16663 30976 16680 31016
rect 16720 30976 16729 31016
rect 16343 30953 16409 30976
rect 16495 30953 16577 30976
rect 16663 30953 16729 30976
rect 16343 30934 16729 30953
rect 20343 31039 20729 31058
rect 20343 31016 20409 31039
rect 20495 31016 20577 31039
rect 20663 31016 20729 31039
rect 20343 30976 20352 31016
rect 20392 30976 20409 31016
rect 20495 30976 20516 31016
rect 20556 30976 20577 31016
rect 20663 30976 20680 31016
rect 20720 30976 20729 31016
rect 20343 30953 20409 30976
rect 20495 30953 20577 30976
rect 20663 30953 20729 30976
rect 20343 30934 20729 30953
rect 24343 31039 24729 31058
rect 24343 31016 24409 31039
rect 24495 31016 24577 31039
rect 24663 31016 24729 31039
rect 24343 30976 24352 31016
rect 24392 30976 24409 31016
rect 24495 30976 24516 31016
rect 24556 30976 24577 31016
rect 24663 30976 24680 31016
rect 24720 30976 24729 31016
rect 24343 30953 24409 30976
rect 24495 30953 24577 30976
rect 24663 30953 24729 30976
rect 24343 30934 24729 30953
rect 28343 31039 28729 31058
rect 28343 31016 28409 31039
rect 28495 31016 28577 31039
rect 28663 31016 28729 31039
rect 28343 30976 28352 31016
rect 28392 30976 28409 31016
rect 28495 30976 28516 31016
rect 28556 30976 28577 31016
rect 28663 30976 28680 31016
rect 28720 30976 28729 31016
rect 28343 30953 28409 30976
rect 28495 30953 28577 30976
rect 28663 30953 28729 30976
rect 28343 30934 28729 30953
rect 32343 31039 32729 31058
rect 32343 31016 32409 31039
rect 32495 31016 32577 31039
rect 32663 31016 32729 31039
rect 32343 30976 32352 31016
rect 32392 30976 32409 31016
rect 32495 30976 32516 31016
rect 32556 30976 32577 31016
rect 32663 30976 32680 31016
rect 32720 30976 32729 31016
rect 32343 30953 32409 30976
rect 32495 30953 32577 30976
rect 32663 30953 32729 30976
rect 32343 30934 32729 30953
rect 36343 31039 36729 31058
rect 36343 31016 36409 31039
rect 36495 31016 36577 31039
rect 36663 31016 36729 31039
rect 36343 30976 36352 31016
rect 36392 30976 36409 31016
rect 36495 30976 36516 31016
rect 36556 30976 36577 31016
rect 36663 30976 36680 31016
rect 36720 30976 36729 31016
rect 36343 30953 36409 30976
rect 36495 30953 36577 30976
rect 36663 30953 36729 30976
rect 36343 30934 36729 30953
rect 40343 31039 40729 31058
rect 40343 31016 40409 31039
rect 40495 31016 40577 31039
rect 40663 31016 40729 31039
rect 40343 30976 40352 31016
rect 40392 30976 40409 31016
rect 40495 30976 40516 31016
rect 40556 30976 40577 31016
rect 40663 30976 40680 31016
rect 40720 30976 40729 31016
rect 40343 30953 40409 30976
rect 40495 30953 40577 30976
rect 40663 30953 40729 30976
rect 40343 30934 40729 30953
rect 44343 31039 44729 31058
rect 44343 31016 44409 31039
rect 44495 31016 44577 31039
rect 44663 31016 44729 31039
rect 44343 30976 44352 31016
rect 44392 30976 44409 31016
rect 44495 30976 44516 31016
rect 44556 30976 44577 31016
rect 44663 30976 44680 31016
rect 44720 30976 44729 31016
rect 44343 30953 44409 30976
rect 44495 30953 44577 30976
rect 44663 30953 44729 30976
rect 44343 30934 44729 30953
rect 48343 31039 48729 31058
rect 48343 31016 48409 31039
rect 48495 31016 48577 31039
rect 48663 31016 48729 31039
rect 48343 30976 48352 31016
rect 48392 30976 48409 31016
rect 48495 30976 48516 31016
rect 48556 30976 48577 31016
rect 48663 30976 48680 31016
rect 48720 30976 48729 31016
rect 48343 30953 48409 30976
rect 48495 30953 48577 30976
rect 48663 30953 48729 30976
rect 48343 30934 48729 30953
rect 52343 31039 52729 31058
rect 52343 31016 52409 31039
rect 52495 31016 52577 31039
rect 52663 31016 52729 31039
rect 52343 30976 52352 31016
rect 52392 30976 52409 31016
rect 52495 30976 52516 31016
rect 52556 30976 52577 31016
rect 52663 30976 52680 31016
rect 52720 30976 52729 31016
rect 52343 30953 52409 30976
rect 52495 30953 52577 30976
rect 52663 30953 52729 30976
rect 52343 30934 52729 30953
rect 56343 31039 56729 31058
rect 56343 31016 56409 31039
rect 56495 31016 56577 31039
rect 56663 31016 56729 31039
rect 56343 30976 56352 31016
rect 56392 30976 56409 31016
rect 56495 30976 56516 31016
rect 56556 30976 56577 31016
rect 56663 30976 56680 31016
rect 56720 30976 56729 31016
rect 56343 30953 56409 30976
rect 56495 30953 56577 30976
rect 56663 30953 56729 30976
rect 56343 30934 56729 30953
rect 60343 31039 60729 31058
rect 60343 31016 60409 31039
rect 60495 31016 60577 31039
rect 60663 31016 60729 31039
rect 60343 30976 60352 31016
rect 60392 30976 60409 31016
rect 60495 30976 60516 31016
rect 60556 30976 60577 31016
rect 60663 30976 60680 31016
rect 60720 30976 60729 31016
rect 60343 30953 60409 30976
rect 60495 30953 60577 30976
rect 60663 30953 60729 30976
rect 60343 30934 60729 30953
rect 64343 31039 64729 31058
rect 64343 31016 64409 31039
rect 64495 31016 64577 31039
rect 64663 31016 64729 31039
rect 64343 30976 64352 31016
rect 64392 30976 64409 31016
rect 64495 30976 64516 31016
rect 64556 30976 64577 31016
rect 64663 30976 64680 31016
rect 64720 30976 64729 31016
rect 64343 30953 64409 30976
rect 64495 30953 64577 30976
rect 64663 30953 64729 30976
rect 64343 30934 64729 30953
rect 68343 31039 68729 31058
rect 68343 31016 68409 31039
rect 68495 31016 68577 31039
rect 68663 31016 68729 31039
rect 68343 30976 68352 31016
rect 68392 30976 68409 31016
rect 68495 30976 68516 31016
rect 68556 30976 68577 31016
rect 68663 30976 68680 31016
rect 68720 30976 68729 31016
rect 68343 30953 68409 30976
rect 68495 30953 68577 30976
rect 68663 30953 68729 30976
rect 68343 30934 68729 30953
rect 72316 31036 72409 31122
rect 72495 31036 72577 31122
rect 72663 31036 72756 31122
rect 72316 30954 72756 31036
rect 72316 30868 72409 30954
rect 72495 30868 72577 30954
rect 72663 30868 72756 30954
rect 72316 30786 72756 30868
rect 72316 30700 72409 30786
rect 72495 30700 72577 30786
rect 72663 30700 72756 30786
rect 72316 30618 72756 30700
rect 72316 30532 72409 30618
rect 72495 30532 72577 30618
rect 72663 30532 72756 30618
rect 72316 30450 72756 30532
rect 72316 30364 72409 30450
rect 72495 30364 72577 30450
rect 72663 30364 72756 30450
rect 3103 30283 3489 30302
rect 3103 30260 3169 30283
rect 3255 30260 3337 30283
rect 3423 30260 3489 30283
rect 3103 30220 3112 30260
rect 3152 30220 3169 30260
rect 3255 30220 3276 30260
rect 3316 30220 3337 30260
rect 3423 30220 3440 30260
rect 3480 30220 3489 30260
rect 3103 30197 3169 30220
rect 3255 30197 3337 30220
rect 3423 30197 3489 30220
rect 3103 30178 3489 30197
rect 7103 30283 7489 30302
rect 7103 30260 7169 30283
rect 7255 30260 7337 30283
rect 7423 30260 7489 30283
rect 7103 30220 7112 30260
rect 7152 30220 7169 30260
rect 7255 30220 7276 30260
rect 7316 30220 7337 30260
rect 7423 30220 7440 30260
rect 7480 30220 7489 30260
rect 7103 30197 7169 30220
rect 7255 30197 7337 30220
rect 7423 30197 7489 30220
rect 7103 30178 7489 30197
rect 11103 30283 11489 30302
rect 11103 30260 11169 30283
rect 11255 30260 11337 30283
rect 11423 30260 11489 30283
rect 11103 30220 11112 30260
rect 11152 30220 11169 30260
rect 11255 30220 11276 30260
rect 11316 30220 11337 30260
rect 11423 30220 11440 30260
rect 11480 30220 11489 30260
rect 11103 30197 11169 30220
rect 11255 30197 11337 30220
rect 11423 30197 11489 30220
rect 11103 30178 11489 30197
rect 15103 30283 15489 30302
rect 15103 30260 15169 30283
rect 15255 30260 15337 30283
rect 15423 30260 15489 30283
rect 15103 30220 15112 30260
rect 15152 30220 15169 30260
rect 15255 30220 15276 30260
rect 15316 30220 15337 30260
rect 15423 30220 15440 30260
rect 15480 30220 15489 30260
rect 15103 30197 15169 30220
rect 15255 30197 15337 30220
rect 15423 30197 15489 30220
rect 15103 30178 15489 30197
rect 19103 30283 19489 30302
rect 19103 30260 19169 30283
rect 19255 30260 19337 30283
rect 19423 30260 19489 30283
rect 19103 30220 19112 30260
rect 19152 30220 19169 30260
rect 19255 30220 19276 30260
rect 19316 30220 19337 30260
rect 19423 30220 19440 30260
rect 19480 30220 19489 30260
rect 19103 30197 19169 30220
rect 19255 30197 19337 30220
rect 19423 30197 19489 30220
rect 19103 30178 19489 30197
rect 23103 30283 23489 30302
rect 23103 30260 23169 30283
rect 23255 30260 23337 30283
rect 23423 30260 23489 30283
rect 23103 30220 23112 30260
rect 23152 30220 23169 30260
rect 23255 30220 23276 30260
rect 23316 30220 23337 30260
rect 23423 30220 23440 30260
rect 23480 30220 23489 30260
rect 23103 30197 23169 30220
rect 23255 30197 23337 30220
rect 23423 30197 23489 30220
rect 23103 30178 23489 30197
rect 27103 30283 27489 30302
rect 27103 30260 27169 30283
rect 27255 30260 27337 30283
rect 27423 30260 27489 30283
rect 27103 30220 27112 30260
rect 27152 30220 27169 30260
rect 27255 30220 27276 30260
rect 27316 30220 27337 30260
rect 27423 30220 27440 30260
rect 27480 30220 27489 30260
rect 27103 30197 27169 30220
rect 27255 30197 27337 30220
rect 27423 30197 27489 30220
rect 27103 30178 27489 30197
rect 31103 30283 31489 30302
rect 31103 30260 31169 30283
rect 31255 30260 31337 30283
rect 31423 30260 31489 30283
rect 31103 30220 31112 30260
rect 31152 30220 31169 30260
rect 31255 30220 31276 30260
rect 31316 30220 31337 30260
rect 31423 30220 31440 30260
rect 31480 30220 31489 30260
rect 31103 30197 31169 30220
rect 31255 30197 31337 30220
rect 31423 30197 31489 30220
rect 31103 30178 31489 30197
rect 35103 30283 35489 30302
rect 35103 30260 35169 30283
rect 35255 30260 35337 30283
rect 35423 30260 35489 30283
rect 35103 30220 35112 30260
rect 35152 30220 35169 30260
rect 35255 30220 35276 30260
rect 35316 30220 35337 30260
rect 35423 30220 35440 30260
rect 35480 30220 35489 30260
rect 35103 30197 35169 30220
rect 35255 30197 35337 30220
rect 35423 30197 35489 30220
rect 35103 30178 35489 30197
rect 39103 30283 39489 30302
rect 39103 30260 39169 30283
rect 39255 30260 39337 30283
rect 39423 30260 39489 30283
rect 39103 30220 39112 30260
rect 39152 30220 39169 30260
rect 39255 30220 39276 30260
rect 39316 30220 39337 30260
rect 39423 30220 39440 30260
rect 39480 30220 39489 30260
rect 39103 30197 39169 30220
rect 39255 30197 39337 30220
rect 39423 30197 39489 30220
rect 39103 30178 39489 30197
rect 43103 30283 43489 30302
rect 43103 30260 43169 30283
rect 43255 30260 43337 30283
rect 43423 30260 43489 30283
rect 43103 30220 43112 30260
rect 43152 30220 43169 30260
rect 43255 30220 43276 30260
rect 43316 30220 43337 30260
rect 43423 30220 43440 30260
rect 43480 30220 43489 30260
rect 43103 30197 43169 30220
rect 43255 30197 43337 30220
rect 43423 30197 43489 30220
rect 43103 30178 43489 30197
rect 47103 30283 47489 30302
rect 47103 30260 47169 30283
rect 47255 30260 47337 30283
rect 47423 30260 47489 30283
rect 47103 30220 47112 30260
rect 47152 30220 47169 30260
rect 47255 30220 47276 30260
rect 47316 30220 47337 30260
rect 47423 30220 47440 30260
rect 47480 30220 47489 30260
rect 47103 30197 47169 30220
rect 47255 30197 47337 30220
rect 47423 30197 47489 30220
rect 47103 30178 47489 30197
rect 51103 30283 51489 30302
rect 51103 30260 51169 30283
rect 51255 30260 51337 30283
rect 51423 30260 51489 30283
rect 51103 30220 51112 30260
rect 51152 30220 51169 30260
rect 51255 30220 51276 30260
rect 51316 30220 51337 30260
rect 51423 30220 51440 30260
rect 51480 30220 51489 30260
rect 51103 30197 51169 30220
rect 51255 30197 51337 30220
rect 51423 30197 51489 30220
rect 51103 30178 51489 30197
rect 55103 30283 55489 30302
rect 55103 30260 55169 30283
rect 55255 30260 55337 30283
rect 55423 30260 55489 30283
rect 55103 30220 55112 30260
rect 55152 30220 55169 30260
rect 55255 30220 55276 30260
rect 55316 30220 55337 30260
rect 55423 30220 55440 30260
rect 55480 30220 55489 30260
rect 55103 30197 55169 30220
rect 55255 30197 55337 30220
rect 55423 30197 55489 30220
rect 55103 30178 55489 30197
rect 59103 30283 59489 30302
rect 59103 30260 59169 30283
rect 59255 30260 59337 30283
rect 59423 30260 59489 30283
rect 59103 30220 59112 30260
rect 59152 30220 59169 30260
rect 59255 30220 59276 30260
rect 59316 30220 59337 30260
rect 59423 30220 59440 30260
rect 59480 30220 59489 30260
rect 59103 30197 59169 30220
rect 59255 30197 59337 30220
rect 59423 30197 59489 30220
rect 59103 30178 59489 30197
rect 63103 30283 63489 30302
rect 63103 30260 63169 30283
rect 63255 30260 63337 30283
rect 63423 30260 63489 30283
rect 63103 30220 63112 30260
rect 63152 30220 63169 30260
rect 63255 30220 63276 30260
rect 63316 30220 63337 30260
rect 63423 30220 63440 30260
rect 63480 30220 63489 30260
rect 63103 30197 63169 30220
rect 63255 30197 63337 30220
rect 63423 30197 63489 30220
rect 63103 30178 63489 30197
rect 67103 30283 67489 30302
rect 67103 30260 67169 30283
rect 67255 30260 67337 30283
rect 67423 30260 67489 30283
rect 67103 30220 67112 30260
rect 67152 30220 67169 30260
rect 67255 30220 67276 30260
rect 67316 30220 67337 30260
rect 67423 30220 67440 30260
rect 67480 30220 67489 30260
rect 67103 30197 67169 30220
rect 67255 30197 67337 30220
rect 67423 30197 67489 30220
rect 67103 30178 67489 30197
rect 72316 30282 72756 30364
rect 72316 30196 72409 30282
rect 72495 30196 72577 30282
rect 72663 30196 72756 30282
rect 72316 30114 72756 30196
rect 72316 30028 72409 30114
rect 72495 30028 72577 30114
rect 72663 30028 72756 30114
rect 72316 29946 72756 30028
rect 72316 29860 72409 29946
rect 72495 29860 72577 29946
rect 72663 29860 72756 29946
rect 72316 29778 72756 29860
rect 72316 29692 72409 29778
rect 72495 29692 72577 29778
rect 72663 29692 72756 29778
rect 72316 29610 72756 29692
rect 4343 29527 4729 29546
rect 4343 29504 4409 29527
rect 4495 29504 4577 29527
rect 4663 29504 4729 29527
rect 4343 29464 4352 29504
rect 4392 29464 4409 29504
rect 4495 29464 4516 29504
rect 4556 29464 4577 29504
rect 4663 29464 4680 29504
rect 4720 29464 4729 29504
rect 4343 29441 4409 29464
rect 4495 29441 4577 29464
rect 4663 29441 4729 29464
rect 4343 29422 4729 29441
rect 8343 29527 8729 29546
rect 8343 29504 8409 29527
rect 8495 29504 8577 29527
rect 8663 29504 8729 29527
rect 8343 29464 8352 29504
rect 8392 29464 8409 29504
rect 8495 29464 8516 29504
rect 8556 29464 8577 29504
rect 8663 29464 8680 29504
rect 8720 29464 8729 29504
rect 8343 29441 8409 29464
rect 8495 29441 8577 29464
rect 8663 29441 8729 29464
rect 8343 29422 8729 29441
rect 12343 29527 12729 29546
rect 12343 29504 12409 29527
rect 12495 29504 12577 29527
rect 12663 29504 12729 29527
rect 12343 29464 12352 29504
rect 12392 29464 12409 29504
rect 12495 29464 12516 29504
rect 12556 29464 12577 29504
rect 12663 29464 12680 29504
rect 12720 29464 12729 29504
rect 12343 29441 12409 29464
rect 12495 29441 12577 29464
rect 12663 29441 12729 29464
rect 12343 29422 12729 29441
rect 16343 29527 16729 29546
rect 16343 29504 16409 29527
rect 16495 29504 16577 29527
rect 16663 29504 16729 29527
rect 16343 29464 16352 29504
rect 16392 29464 16409 29504
rect 16495 29464 16516 29504
rect 16556 29464 16577 29504
rect 16663 29464 16680 29504
rect 16720 29464 16729 29504
rect 16343 29441 16409 29464
rect 16495 29441 16577 29464
rect 16663 29441 16729 29464
rect 16343 29422 16729 29441
rect 20343 29527 20729 29546
rect 20343 29504 20409 29527
rect 20495 29504 20577 29527
rect 20663 29504 20729 29527
rect 20343 29464 20352 29504
rect 20392 29464 20409 29504
rect 20495 29464 20516 29504
rect 20556 29464 20577 29504
rect 20663 29464 20680 29504
rect 20720 29464 20729 29504
rect 20343 29441 20409 29464
rect 20495 29441 20577 29464
rect 20663 29441 20729 29464
rect 20343 29422 20729 29441
rect 24343 29527 24729 29546
rect 24343 29504 24409 29527
rect 24495 29504 24577 29527
rect 24663 29504 24729 29527
rect 24343 29464 24352 29504
rect 24392 29464 24409 29504
rect 24495 29464 24516 29504
rect 24556 29464 24577 29504
rect 24663 29464 24680 29504
rect 24720 29464 24729 29504
rect 24343 29441 24409 29464
rect 24495 29441 24577 29464
rect 24663 29441 24729 29464
rect 24343 29422 24729 29441
rect 28343 29527 28729 29546
rect 28343 29504 28409 29527
rect 28495 29504 28577 29527
rect 28663 29504 28729 29527
rect 28343 29464 28352 29504
rect 28392 29464 28409 29504
rect 28495 29464 28516 29504
rect 28556 29464 28577 29504
rect 28663 29464 28680 29504
rect 28720 29464 28729 29504
rect 28343 29441 28409 29464
rect 28495 29441 28577 29464
rect 28663 29441 28729 29464
rect 28343 29422 28729 29441
rect 32343 29527 32729 29546
rect 32343 29504 32409 29527
rect 32495 29504 32577 29527
rect 32663 29504 32729 29527
rect 32343 29464 32352 29504
rect 32392 29464 32409 29504
rect 32495 29464 32516 29504
rect 32556 29464 32577 29504
rect 32663 29464 32680 29504
rect 32720 29464 32729 29504
rect 32343 29441 32409 29464
rect 32495 29441 32577 29464
rect 32663 29441 32729 29464
rect 32343 29422 32729 29441
rect 36343 29527 36729 29546
rect 36343 29504 36409 29527
rect 36495 29504 36577 29527
rect 36663 29504 36729 29527
rect 36343 29464 36352 29504
rect 36392 29464 36409 29504
rect 36495 29464 36516 29504
rect 36556 29464 36577 29504
rect 36663 29464 36680 29504
rect 36720 29464 36729 29504
rect 36343 29441 36409 29464
rect 36495 29441 36577 29464
rect 36663 29441 36729 29464
rect 36343 29422 36729 29441
rect 40343 29527 40729 29546
rect 40343 29504 40409 29527
rect 40495 29504 40577 29527
rect 40663 29504 40729 29527
rect 40343 29464 40352 29504
rect 40392 29464 40409 29504
rect 40495 29464 40516 29504
rect 40556 29464 40577 29504
rect 40663 29464 40680 29504
rect 40720 29464 40729 29504
rect 40343 29441 40409 29464
rect 40495 29441 40577 29464
rect 40663 29441 40729 29464
rect 40343 29422 40729 29441
rect 44343 29527 44729 29546
rect 44343 29504 44409 29527
rect 44495 29504 44577 29527
rect 44663 29504 44729 29527
rect 44343 29464 44352 29504
rect 44392 29464 44409 29504
rect 44495 29464 44516 29504
rect 44556 29464 44577 29504
rect 44663 29464 44680 29504
rect 44720 29464 44729 29504
rect 44343 29441 44409 29464
rect 44495 29441 44577 29464
rect 44663 29441 44729 29464
rect 44343 29422 44729 29441
rect 48343 29527 48729 29546
rect 48343 29504 48409 29527
rect 48495 29504 48577 29527
rect 48663 29504 48729 29527
rect 48343 29464 48352 29504
rect 48392 29464 48409 29504
rect 48495 29464 48516 29504
rect 48556 29464 48577 29504
rect 48663 29464 48680 29504
rect 48720 29464 48729 29504
rect 48343 29441 48409 29464
rect 48495 29441 48577 29464
rect 48663 29441 48729 29464
rect 48343 29422 48729 29441
rect 52343 29527 52729 29546
rect 52343 29504 52409 29527
rect 52495 29504 52577 29527
rect 52663 29504 52729 29527
rect 52343 29464 52352 29504
rect 52392 29464 52409 29504
rect 52495 29464 52516 29504
rect 52556 29464 52577 29504
rect 52663 29464 52680 29504
rect 52720 29464 52729 29504
rect 52343 29441 52409 29464
rect 52495 29441 52577 29464
rect 52663 29441 52729 29464
rect 52343 29422 52729 29441
rect 56343 29527 56729 29546
rect 56343 29504 56409 29527
rect 56495 29504 56577 29527
rect 56663 29504 56729 29527
rect 56343 29464 56352 29504
rect 56392 29464 56409 29504
rect 56495 29464 56516 29504
rect 56556 29464 56577 29504
rect 56663 29464 56680 29504
rect 56720 29464 56729 29504
rect 56343 29441 56409 29464
rect 56495 29441 56577 29464
rect 56663 29441 56729 29464
rect 56343 29422 56729 29441
rect 60343 29527 60729 29546
rect 60343 29504 60409 29527
rect 60495 29504 60577 29527
rect 60663 29504 60729 29527
rect 60343 29464 60352 29504
rect 60392 29464 60409 29504
rect 60495 29464 60516 29504
rect 60556 29464 60577 29504
rect 60663 29464 60680 29504
rect 60720 29464 60729 29504
rect 60343 29441 60409 29464
rect 60495 29441 60577 29464
rect 60663 29441 60729 29464
rect 60343 29422 60729 29441
rect 64343 29527 64729 29546
rect 64343 29504 64409 29527
rect 64495 29504 64577 29527
rect 64663 29504 64729 29527
rect 64343 29464 64352 29504
rect 64392 29464 64409 29504
rect 64495 29464 64516 29504
rect 64556 29464 64577 29504
rect 64663 29464 64680 29504
rect 64720 29464 64729 29504
rect 64343 29441 64409 29464
rect 64495 29441 64577 29464
rect 64663 29441 64729 29464
rect 64343 29422 64729 29441
rect 68343 29527 68729 29546
rect 68343 29504 68409 29527
rect 68495 29504 68577 29527
rect 68663 29504 68729 29527
rect 68343 29464 68352 29504
rect 68392 29464 68409 29504
rect 68495 29464 68516 29504
rect 68556 29464 68577 29504
rect 68663 29464 68680 29504
rect 68720 29464 68729 29504
rect 68343 29441 68409 29464
rect 68495 29441 68577 29464
rect 68663 29441 68729 29464
rect 68343 29422 68729 29441
rect 72316 29524 72409 29610
rect 72495 29524 72577 29610
rect 72663 29524 72756 29610
rect 72316 29442 72756 29524
rect 72316 29356 72409 29442
rect 72495 29356 72577 29442
rect 72663 29356 72756 29442
rect 72316 29274 72756 29356
rect 72316 29188 72409 29274
rect 72495 29188 72577 29274
rect 72663 29188 72756 29274
rect 72316 29106 72756 29188
rect 72316 29020 72409 29106
rect 72495 29020 72577 29106
rect 72663 29020 72756 29106
rect 72316 28890 72756 29020
rect 76316 31122 76756 31252
rect 76316 31036 76409 31122
rect 76495 31036 76577 31122
rect 76663 31036 76756 31122
rect 76316 30954 76756 31036
rect 76316 30868 76409 30954
rect 76495 30868 76577 30954
rect 76663 30868 76756 30954
rect 76316 30786 76756 30868
rect 76316 30700 76409 30786
rect 76495 30700 76577 30786
rect 76663 30700 76756 30786
rect 76316 30618 76756 30700
rect 76316 30532 76409 30618
rect 76495 30532 76577 30618
rect 76663 30532 76756 30618
rect 76316 30450 76756 30532
rect 76316 30364 76409 30450
rect 76495 30364 76577 30450
rect 76663 30364 76756 30450
rect 76316 30282 76756 30364
rect 76316 30196 76409 30282
rect 76495 30196 76577 30282
rect 76663 30196 76756 30282
rect 76316 30114 76756 30196
rect 76316 30028 76409 30114
rect 76495 30028 76577 30114
rect 76663 30028 76756 30114
rect 76316 29946 76756 30028
rect 76316 29860 76409 29946
rect 76495 29860 76577 29946
rect 76663 29860 76756 29946
rect 76316 29778 76756 29860
rect 76316 29692 76409 29778
rect 76495 29692 76577 29778
rect 76663 29692 76756 29778
rect 76316 29610 76756 29692
rect 76316 29524 76409 29610
rect 76495 29524 76577 29610
rect 76663 29524 76756 29610
rect 76316 29442 76756 29524
rect 76316 29356 76409 29442
rect 76495 29356 76577 29442
rect 76663 29356 76756 29442
rect 76316 29274 76756 29356
rect 76316 29188 76409 29274
rect 76495 29188 76577 29274
rect 76663 29188 76756 29274
rect 76316 29106 76756 29188
rect 76316 29020 76409 29106
rect 76495 29020 76577 29106
rect 76663 29020 76756 29106
rect 76316 28890 76756 29020
rect 80316 31122 80756 31252
rect 80316 31036 80409 31122
rect 80495 31036 80577 31122
rect 80663 31036 80756 31122
rect 80316 30954 80756 31036
rect 80316 30868 80409 30954
rect 80495 30868 80577 30954
rect 80663 30868 80756 30954
rect 80316 30786 80756 30868
rect 80316 30700 80409 30786
rect 80495 30700 80577 30786
rect 80663 30700 80756 30786
rect 80316 30618 80756 30700
rect 80316 30532 80409 30618
rect 80495 30532 80577 30618
rect 80663 30532 80756 30618
rect 80316 30450 80756 30532
rect 80316 30364 80409 30450
rect 80495 30364 80577 30450
rect 80663 30364 80756 30450
rect 80316 30282 80756 30364
rect 80316 30196 80409 30282
rect 80495 30196 80577 30282
rect 80663 30196 80756 30282
rect 80316 30114 80756 30196
rect 80316 30028 80409 30114
rect 80495 30028 80577 30114
rect 80663 30028 80756 30114
rect 80316 29946 80756 30028
rect 80316 29860 80409 29946
rect 80495 29860 80577 29946
rect 80663 29860 80756 29946
rect 80316 29778 80756 29860
rect 80316 29692 80409 29778
rect 80495 29692 80577 29778
rect 80663 29692 80756 29778
rect 80316 29610 80756 29692
rect 80316 29524 80409 29610
rect 80495 29524 80577 29610
rect 80663 29524 80756 29610
rect 80316 29442 80756 29524
rect 80316 29356 80409 29442
rect 80495 29356 80577 29442
rect 80663 29356 80756 29442
rect 80316 29274 80756 29356
rect 80316 29188 80409 29274
rect 80495 29188 80577 29274
rect 80663 29188 80756 29274
rect 80316 29106 80756 29188
rect 80316 29020 80409 29106
rect 80495 29020 80577 29106
rect 80663 29020 80756 29106
rect 80316 28890 80756 29020
rect 84316 31122 84756 31252
rect 84316 31036 84409 31122
rect 84495 31036 84577 31122
rect 84663 31036 84756 31122
rect 84316 30954 84756 31036
rect 84316 30868 84409 30954
rect 84495 30868 84577 30954
rect 84663 30868 84756 30954
rect 84316 30786 84756 30868
rect 84316 30700 84409 30786
rect 84495 30700 84577 30786
rect 84663 30700 84756 30786
rect 84316 30618 84756 30700
rect 84316 30532 84409 30618
rect 84495 30532 84577 30618
rect 84663 30532 84756 30618
rect 84316 30450 84756 30532
rect 84316 30364 84409 30450
rect 84495 30364 84577 30450
rect 84663 30364 84756 30450
rect 84316 30282 84756 30364
rect 84316 30196 84409 30282
rect 84495 30196 84577 30282
rect 84663 30196 84756 30282
rect 84316 30114 84756 30196
rect 84316 30028 84409 30114
rect 84495 30028 84577 30114
rect 84663 30028 84756 30114
rect 84316 29946 84756 30028
rect 84316 29860 84409 29946
rect 84495 29860 84577 29946
rect 84663 29860 84756 29946
rect 84316 29778 84756 29860
rect 84316 29692 84409 29778
rect 84495 29692 84577 29778
rect 84663 29692 84756 29778
rect 84316 29610 84756 29692
rect 84316 29524 84409 29610
rect 84495 29524 84577 29610
rect 84663 29524 84756 29610
rect 84316 29442 84756 29524
rect 84316 29356 84409 29442
rect 84495 29356 84577 29442
rect 84663 29356 84756 29442
rect 84316 29274 84756 29356
rect 84316 29188 84409 29274
rect 84495 29188 84577 29274
rect 84663 29188 84756 29274
rect 84316 29106 84756 29188
rect 84316 29020 84409 29106
rect 84495 29020 84577 29106
rect 84663 29020 84756 29106
rect 84316 28890 84756 29020
rect 88316 31122 88756 31252
rect 88316 31036 88409 31122
rect 88495 31036 88577 31122
rect 88663 31036 88756 31122
rect 88316 30954 88756 31036
rect 88316 30868 88409 30954
rect 88495 30868 88577 30954
rect 88663 30868 88756 30954
rect 88316 30786 88756 30868
rect 88316 30700 88409 30786
rect 88495 30700 88577 30786
rect 88663 30700 88756 30786
rect 88316 30618 88756 30700
rect 88316 30532 88409 30618
rect 88495 30532 88577 30618
rect 88663 30532 88756 30618
rect 88316 30450 88756 30532
rect 88316 30364 88409 30450
rect 88495 30364 88577 30450
rect 88663 30364 88756 30450
rect 88316 30282 88756 30364
rect 88316 30196 88409 30282
rect 88495 30196 88577 30282
rect 88663 30196 88756 30282
rect 88316 30114 88756 30196
rect 88316 30028 88409 30114
rect 88495 30028 88577 30114
rect 88663 30028 88756 30114
rect 88316 29946 88756 30028
rect 88316 29860 88409 29946
rect 88495 29860 88577 29946
rect 88663 29860 88756 29946
rect 88316 29778 88756 29860
rect 88316 29692 88409 29778
rect 88495 29692 88577 29778
rect 88663 29692 88756 29778
rect 88316 29610 88756 29692
rect 88316 29524 88409 29610
rect 88495 29524 88577 29610
rect 88663 29524 88756 29610
rect 88316 29442 88756 29524
rect 88316 29356 88409 29442
rect 88495 29356 88577 29442
rect 88663 29356 88756 29442
rect 88316 29274 88756 29356
rect 88316 29188 88409 29274
rect 88495 29188 88577 29274
rect 88663 29188 88756 29274
rect 88316 29106 88756 29188
rect 88316 29020 88409 29106
rect 88495 29020 88577 29106
rect 88663 29020 88756 29106
rect 88316 28890 88756 29020
rect 92316 31122 92756 31252
rect 92316 31036 92409 31122
rect 92495 31036 92577 31122
rect 92663 31036 92756 31122
rect 92316 30954 92756 31036
rect 92316 30868 92409 30954
rect 92495 30868 92577 30954
rect 92663 30868 92756 30954
rect 92316 30786 92756 30868
rect 92316 30700 92409 30786
rect 92495 30700 92577 30786
rect 92663 30700 92756 30786
rect 92316 30618 92756 30700
rect 92316 30532 92409 30618
rect 92495 30532 92577 30618
rect 92663 30532 92756 30618
rect 92316 30450 92756 30532
rect 92316 30364 92409 30450
rect 92495 30364 92577 30450
rect 92663 30364 92756 30450
rect 92316 30282 92756 30364
rect 92316 30196 92409 30282
rect 92495 30196 92577 30282
rect 92663 30196 92756 30282
rect 92316 30114 92756 30196
rect 92316 30028 92409 30114
rect 92495 30028 92577 30114
rect 92663 30028 92756 30114
rect 92316 29946 92756 30028
rect 92316 29860 92409 29946
rect 92495 29860 92577 29946
rect 92663 29860 92756 29946
rect 92316 29778 92756 29860
rect 92316 29692 92409 29778
rect 92495 29692 92577 29778
rect 92663 29692 92756 29778
rect 92316 29610 92756 29692
rect 92316 29524 92409 29610
rect 92495 29524 92577 29610
rect 92663 29524 92756 29610
rect 92316 29442 92756 29524
rect 92316 29356 92409 29442
rect 92495 29356 92577 29442
rect 92663 29356 92756 29442
rect 92316 29274 92756 29356
rect 92316 29188 92409 29274
rect 92495 29188 92577 29274
rect 92663 29188 92756 29274
rect 92316 29106 92756 29188
rect 92316 29020 92409 29106
rect 92495 29020 92577 29106
rect 92663 29020 92756 29106
rect 92316 28890 92756 29020
rect 96316 31122 96756 31252
rect 96316 31036 96409 31122
rect 96495 31036 96577 31122
rect 96663 31036 96756 31122
rect 96316 30954 96756 31036
rect 96316 30868 96409 30954
rect 96495 30868 96577 30954
rect 96663 30868 96756 30954
rect 96316 30786 96756 30868
rect 96316 30700 96409 30786
rect 96495 30700 96577 30786
rect 96663 30700 96756 30786
rect 96316 30618 96756 30700
rect 96316 30532 96409 30618
rect 96495 30532 96577 30618
rect 96663 30532 96756 30618
rect 96316 30450 96756 30532
rect 96316 30364 96409 30450
rect 96495 30364 96577 30450
rect 96663 30364 96756 30450
rect 96316 30282 96756 30364
rect 96316 30196 96409 30282
rect 96495 30196 96577 30282
rect 96663 30196 96756 30282
rect 96316 30114 96756 30196
rect 96316 30028 96409 30114
rect 96495 30028 96577 30114
rect 96663 30028 96756 30114
rect 96316 29946 96756 30028
rect 96316 29860 96409 29946
rect 96495 29860 96577 29946
rect 96663 29860 96756 29946
rect 96316 29778 96756 29860
rect 96316 29692 96409 29778
rect 96495 29692 96577 29778
rect 96663 29692 96756 29778
rect 96316 29610 96756 29692
rect 96316 29524 96409 29610
rect 96495 29524 96577 29610
rect 96663 29524 96756 29610
rect 96316 29442 96756 29524
rect 96316 29356 96409 29442
rect 96495 29356 96577 29442
rect 96663 29356 96756 29442
rect 96316 29274 96756 29356
rect 96316 29188 96409 29274
rect 96495 29188 96577 29274
rect 96663 29188 96756 29274
rect 96316 29106 96756 29188
rect 96316 29020 96409 29106
rect 96495 29020 96577 29106
rect 96663 29020 96756 29106
rect 96316 28890 96756 29020
rect 3103 28771 3489 28790
rect 3103 28748 3169 28771
rect 3255 28748 3337 28771
rect 3423 28748 3489 28771
rect 3103 28708 3112 28748
rect 3152 28708 3169 28748
rect 3255 28708 3276 28748
rect 3316 28708 3337 28748
rect 3423 28708 3440 28748
rect 3480 28708 3489 28748
rect 3103 28685 3169 28708
rect 3255 28685 3337 28708
rect 3423 28685 3489 28708
rect 3103 28666 3489 28685
rect 7103 28771 7489 28790
rect 7103 28748 7169 28771
rect 7255 28748 7337 28771
rect 7423 28748 7489 28771
rect 7103 28708 7112 28748
rect 7152 28708 7169 28748
rect 7255 28708 7276 28748
rect 7316 28708 7337 28748
rect 7423 28708 7440 28748
rect 7480 28708 7489 28748
rect 7103 28685 7169 28708
rect 7255 28685 7337 28708
rect 7423 28685 7489 28708
rect 7103 28666 7489 28685
rect 11103 28771 11489 28790
rect 11103 28748 11169 28771
rect 11255 28748 11337 28771
rect 11423 28748 11489 28771
rect 11103 28708 11112 28748
rect 11152 28708 11169 28748
rect 11255 28708 11276 28748
rect 11316 28708 11337 28748
rect 11423 28708 11440 28748
rect 11480 28708 11489 28748
rect 11103 28685 11169 28708
rect 11255 28685 11337 28708
rect 11423 28685 11489 28708
rect 11103 28666 11489 28685
rect 15103 28771 15489 28790
rect 15103 28748 15169 28771
rect 15255 28748 15337 28771
rect 15423 28748 15489 28771
rect 15103 28708 15112 28748
rect 15152 28708 15169 28748
rect 15255 28708 15276 28748
rect 15316 28708 15337 28748
rect 15423 28708 15440 28748
rect 15480 28708 15489 28748
rect 15103 28685 15169 28708
rect 15255 28685 15337 28708
rect 15423 28685 15489 28708
rect 15103 28666 15489 28685
rect 19103 28771 19489 28790
rect 19103 28748 19169 28771
rect 19255 28748 19337 28771
rect 19423 28748 19489 28771
rect 19103 28708 19112 28748
rect 19152 28708 19169 28748
rect 19255 28708 19276 28748
rect 19316 28708 19337 28748
rect 19423 28708 19440 28748
rect 19480 28708 19489 28748
rect 19103 28685 19169 28708
rect 19255 28685 19337 28708
rect 19423 28685 19489 28708
rect 19103 28666 19489 28685
rect 23103 28771 23489 28790
rect 23103 28748 23169 28771
rect 23255 28748 23337 28771
rect 23423 28748 23489 28771
rect 23103 28708 23112 28748
rect 23152 28708 23169 28748
rect 23255 28708 23276 28748
rect 23316 28708 23337 28748
rect 23423 28708 23440 28748
rect 23480 28708 23489 28748
rect 23103 28685 23169 28708
rect 23255 28685 23337 28708
rect 23423 28685 23489 28708
rect 23103 28666 23489 28685
rect 27103 28771 27489 28790
rect 27103 28748 27169 28771
rect 27255 28748 27337 28771
rect 27423 28748 27489 28771
rect 27103 28708 27112 28748
rect 27152 28708 27169 28748
rect 27255 28708 27276 28748
rect 27316 28708 27337 28748
rect 27423 28708 27440 28748
rect 27480 28708 27489 28748
rect 27103 28685 27169 28708
rect 27255 28685 27337 28708
rect 27423 28685 27489 28708
rect 27103 28666 27489 28685
rect 31103 28771 31489 28790
rect 31103 28748 31169 28771
rect 31255 28748 31337 28771
rect 31423 28748 31489 28771
rect 31103 28708 31112 28748
rect 31152 28708 31169 28748
rect 31255 28708 31276 28748
rect 31316 28708 31337 28748
rect 31423 28708 31440 28748
rect 31480 28708 31489 28748
rect 31103 28685 31169 28708
rect 31255 28685 31337 28708
rect 31423 28685 31489 28708
rect 31103 28666 31489 28685
rect 35103 28771 35489 28790
rect 35103 28748 35169 28771
rect 35255 28748 35337 28771
rect 35423 28748 35489 28771
rect 35103 28708 35112 28748
rect 35152 28708 35169 28748
rect 35255 28708 35276 28748
rect 35316 28708 35337 28748
rect 35423 28708 35440 28748
rect 35480 28708 35489 28748
rect 35103 28685 35169 28708
rect 35255 28685 35337 28708
rect 35423 28685 35489 28708
rect 35103 28666 35489 28685
rect 39103 28771 39489 28790
rect 39103 28748 39169 28771
rect 39255 28748 39337 28771
rect 39423 28748 39489 28771
rect 39103 28708 39112 28748
rect 39152 28708 39169 28748
rect 39255 28708 39276 28748
rect 39316 28708 39337 28748
rect 39423 28708 39440 28748
rect 39480 28708 39489 28748
rect 39103 28685 39169 28708
rect 39255 28685 39337 28708
rect 39423 28685 39489 28708
rect 39103 28666 39489 28685
rect 43103 28771 43489 28790
rect 43103 28748 43169 28771
rect 43255 28748 43337 28771
rect 43423 28748 43489 28771
rect 43103 28708 43112 28748
rect 43152 28708 43169 28748
rect 43255 28708 43276 28748
rect 43316 28708 43337 28748
rect 43423 28708 43440 28748
rect 43480 28708 43489 28748
rect 43103 28685 43169 28708
rect 43255 28685 43337 28708
rect 43423 28685 43489 28708
rect 43103 28666 43489 28685
rect 47103 28771 47489 28790
rect 47103 28748 47169 28771
rect 47255 28748 47337 28771
rect 47423 28748 47489 28771
rect 47103 28708 47112 28748
rect 47152 28708 47169 28748
rect 47255 28708 47276 28748
rect 47316 28708 47337 28748
rect 47423 28708 47440 28748
rect 47480 28708 47489 28748
rect 47103 28685 47169 28708
rect 47255 28685 47337 28708
rect 47423 28685 47489 28708
rect 47103 28666 47489 28685
rect 51103 28771 51489 28790
rect 51103 28748 51169 28771
rect 51255 28748 51337 28771
rect 51423 28748 51489 28771
rect 51103 28708 51112 28748
rect 51152 28708 51169 28748
rect 51255 28708 51276 28748
rect 51316 28708 51337 28748
rect 51423 28708 51440 28748
rect 51480 28708 51489 28748
rect 51103 28685 51169 28708
rect 51255 28685 51337 28708
rect 51423 28685 51489 28708
rect 51103 28666 51489 28685
rect 55103 28771 55489 28790
rect 55103 28748 55169 28771
rect 55255 28748 55337 28771
rect 55423 28748 55489 28771
rect 55103 28708 55112 28748
rect 55152 28708 55169 28748
rect 55255 28708 55276 28748
rect 55316 28708 55337 28748
rect 55423 28708 55440 28748
rect 55480 28708 55489 28748
rect 55103 28685 55169 28708
rect 55255 28685 55337 28708
rect 55423 28685 55489 28708
rect 55103 28666 55489 28685
rect 59103 28771 59489 28790
rect 59103 28748 59169 28771
rect 59255 28748 59337 28771
rect 59423 28748 59489 28771
rect 59103 28708 59112 28748
rect 59152 28708 59169 28748
rect 59255 28708 59276 28748
rect 59316 28708 59337 28748
rect 59423 28708 59440 28748
rect 59480 28708 59489 28748
rect 59103 28685 59169 28708
rect 59255 28685 59337 28708
rect 59423 28685 59489 28708
rect 59103 28666 59489 28685
rect 63103 28771 63489 28790
rect 63103 28748 63169 28771
rect 63255 28748 63337 28771
rect 63423 28748 63489 28771
rect 63103 28708 63112 28748
rect 63152 28708 63169 28748
rect 63255 28708 63276 28748
rect 63316 28708 63337 28748
rect 63423 28708 63440 28748
rect 63480 28708 63489 28748
rect 63103 28685 63169 28708
rect 63255 28685 63337 28708
rect 63423 28685 63489 28708
rect 63103 28666 63489 28685
rect 67103 28771 67489 28790
rect 67103 28748 67169 28771
rect 67255 28748 67337 28771
rect 67423 28748 67489 28771
rect 67103 28708 67112 28748
rect 67152 28708 67169 28748
rect 67255 28708 67276 28748
rect 67316 28708 67337 28748
rect 67423 28708 67440 28748
rect 67480 28708 67489 28748
rect 67103 28685 67169 28708
rect 67255 28685 67337 28708
rect 67423 28685 67489 28708
rect 67103 28666 67489 28685
rect 75076 28246 75516 28376
rect 75076 28160 75169 28246
rect 75255 28160 75337 28246
rect 75423 28160 75516 28246
rect 75076 28078 75516 28160
rect 4343 28015 4729 28034
rect 4343 27992 4409 28015
rect 4495 27992 4577 28015
rect 4663 27992 4729 28015
rect 4343 27952 4352 27992
rect 4392 27952 4409 27992
rect 4495 27952 4516 27992
rect 4556 27952 4577 27992
rect 4663 27952 4680 27992
rect 4720 27952 4729 27992
rect 4343 27929 4409 27952
rect 4495 27929 4577 27952
rect 4663 27929 4729 27952
rect 4343 27910 4729 27929
rect 8343 28015 8729 28034
rect 8343 27992 8409 28015
rect 8495 27992 8577 28015
rect 8663 27992 8729 28015
rect 8343 27952 8352 27992
rect 8392 27952 8409 27992
rect 8495 27952 8516 27992
rect 8556 27952 8577 27992
rect 8663 27952 8680 27992
rect 8720 27952 8729 27992
rect 8343 27929 8409 27952
rect 8495 27929 8577 27952
rect 8663 27929 8729 27952
rect 8343 27910 8729 27929
rect 12343 28015 12729 28034
rect 12343 27992 12409 28015
rect 12495 27992 12577 28015
rect 12663 27992 12729 28015
rect 12343 27952 12352 27992
rect 12392 27952 12409 27992
rect 12495 27952 12516 27992
rect 12556 27952 12577 27992
rect 12663 27952 12680 27992
rect 12720 27952 12729 27992
rect 12343 27929 12409 27952
rect 12495 27929 12577 27952
rect 12663 27929 12729 27952
rect 12343 27910 12729 27929
rect 16343 28015 16729 28034
rect 16343 27992 16409 28015
rect 16495 27992 16577 28015
rect 16663 27992 16729 28015
rect 16343 27952 16352 27992
rect 16392 27952 16409 27992
rect 16495 27952 16516 27992
rect 16556 27952 16577 27992
rect 16663 27952 16680 27992
rect 16720 27952 16729 27992
rect 16343 27929 16409 27952
rect 16495 27929 16577 27952
rect 16663 27929 16729 27952
rect 16343 27910 16729 27929
rect 20343 28015 20729 28034
rect 20343 27992 20409 28015
rect 20495 27992 20577 28015
rect 20663 27992 20729 28015
rect 20343 27952 20352 27992
rect 20392 27952 20409 27992
rect 20495 27952 20516 27992
rect 20556 27952 20577 27992
rect 20663 27952 20680 27992
rect 20720 27952 20729 27992
rect 20343 27929 20409 27952
rect 20495 27929 20577 27952
rect 20663 27929 20729 27952
rect 20343 27910 20729 27929
rect 24343 28015 24729 28034
rect 24343 27992 24409 28015
rect 24495 27992 24577 28015
rect 24663 27992 24729 28015
rect 24343 27952 24352 27992
rect 24392 27952 24409 27992
rect 24495 27952 24516 27992
rect 24556 27952 24577 27992
rect 24663 27952 24680 27992
rect 24720 27952 24729 27992
rect 24343 27929 24409 27952
rect 24495 27929 24577 27952
rect 24663 27929 24729 27952
rect 24343 27910 24729 27929
rect 28343 28015 28729 28034
rect 28343 27992 28409 28015
rect 28495 27992 28577 28015
rect 28663 27992 28729 28015
rect 28343 27952 28352 27992
rect 28392 27952 28409 27992
rect 28495 27952 28516 27992
rect 28556 27952 28577 27992
rect 28663 27952 28680 27992
rect 28720 27952 28729 27992
rect 28343 27929 28409 27952
rect 28495 27929 28577 27952
rect 28663 27929 28729 27952
rect 28343 27910 28729 27929
rect 32343 28015 32729 28034
rect 32343 27992 32409 28015
rect 32495 27992 32577 28015
rect 32663 27992 32729 28015
rect 32343 27952 32352 27992
rect 32392 27952 32409 27992
rect 32495 27952 32516 27992
rect 32556 27952 32577 27992
rect 32663 27952 32680 27992
rect 32720 27952 32729 27992
rect 32343 27929 32409 27952
rect 32495 27929 32577 27952
rect 32663 27929 32729 27952
rect 32343 27910 32729 27929
rect 36343 28015 36729 28034
rect 36343 27992 36409 28015
rect 36495 27992 36577 28015
rect 36663 27992 36729 28015
rect 36343 27952 36352 27992
rect 36392 27952 36409 27992
rect 36495 27952 36516 27992
rect 36556 27952 36577 27992
rect 36663 27952 36680 27992
rect 36720 27952 36729 27992
rect 36343 27929 36409 27952
rect 36495 27929 36577 27952
rect 36663 27929 36729 27952
rect 36343 27910 36729 27929
rect 40343 28015 40729 28034
rect 40343 27992 40409 28015
rect 40495 27992 40577 28015
rect 40663 27992 40729 28015
rect 40343 27952 40352 27992
rect 40392 27952 40409 27992
rect 40495 27952 40516 27992
rect 40556 27952 40577 27992
rect 40663 27952 40680 27992
rect 40720 27952 40729 27992
rect 40343 27929 40409 27952
rect 40495 27929 40577 27952
rect 40663 27929 40729 27952
rect 40343 27910 40729 27929
rect 44343 28015 44729 28034
rect 44343 27992 44409 28015
rect 44495 27992 44577 28015
rect 44663 27992 44729 28015
rect 44343 27952 44352 27992
rect 44392 27952 44409 27992
rect 44495 27952 44516 27992
rect 44556 27952 44577 27992
rect 44663 27952 44680 27992
rect 44720 27952 44729 27992
rect 44343 27929 44409 27952
rect 44495 27929 44577 27952
rect 44663 27929 44729 27952
rect 44343 27910 44729 27929
rect 48343 28015 48729 28034
rect 48343 27992 48409 28015
rect 48495 27992 48577 28015
rect 48663 27992 48729 28015
rect 48343 27952 48352 27992
rect 48392 27952 48409 27992
rect 48495 27952 48516 27992
rect 48556 27952 48577 27992
rect 48663 27952 48680 27992
rect 48720 27952 48729 27992
rect 48343 27929 48409 27952
rect 48495 27929 48577 27952
rect 48663 27929 48729 27952
rect 48343 27910 48729 27929
rect 52343 28015 52729 28034
rect 52343 27992 52409 28015
rect 52495 27992 52577 28015
rect 52663 27992 52729 28015
rect 52343 27952 52352 27992
rect 52392 27952 52409 27992
rect 52495 27952 52516 27992
rect 52556 27952 52577 27992
rect 52663 27952 52680 27992
rect 52720 27952 52729 27992
rect 52343 27929 52409 27952
rect 52495 27929 52577 27952
rect 52663 27929 52729 27952
rect 52343 27910 52729 27929
rect 56343 28015 56729 28034
rect 56343 27992 56409 28015
rect 56495 27992 56577 28015
rect 56663 27992 56729 28015
rect 56343 27952 56352 27992
rect 56392 27952 56409 27992
rect 56495 27952 56516 27992
rect 56556 27952 56577 27992
rect 56663 27952 56680 27992
rect 56720 27952 56729 27992
rect 56343 27929 56409 27952
rect 56495 27929 56577 27952
rect 56663 27929 56729 27952
rect 56343 27910 56729 27929
rect 60343 28015 60729 28034
rect 60343 27992 60409 28015
rect 60495 27992 60577 28015
rect 60663 27992 60729 28015
rect 60343 27952 60352 27992
rect 60392 27952 60409 27992
rect 60495 27952 60516 27992
rect 60556 27952 60577 27992
rect 60663 27952 60680 27992
rect 60720 27952 60729 27992
rect 60343 27929 60409 27952
rect 60495 27929 60577 27952
rect 60663 27929 60729 27952
rect 60343 27910 60729 27929
rect 64343 28015 64729 28034
rect 64343 27992 64409 28015
rect 64495 27992 64577 28015
rect 64663 27992 64729 28015
rect 64343 27952 64352 27992
rect 64392 27952 64409 27992
rect 64495 27952 64516 27992
rect 64556 27952 64577 27992
rect 64663 27952 64680 27992
rect 64720 27952 64729 27992
rect 64343 27929 64409 27952
rect 64495 27929 64577 27952
rect 64663 27929 64729 27952
rect 64343 27910 64729 27929
rect 68343 28015 68729 28034
rect 68343 27992 68409 28015
rect 68495 27992 68577 28015
rect 68663 27992 68729 28015
rect 68343 27952 68352 27992
rect 68392 27952 68409 27992
rect 68495 27952 68516 27992
rect 68556 27952 68577 27992
rect 68663 27952 68680 27992
rect 68720 27952 68729 27992
rect 68343 27929 68409 27952
rect 68495 27929 68577 27952
rect 68663 27929 68729 27952
rect 68343 27910 68729 27929
rect 75076 27992 75169 28078
rect 75255 27992 75337 28078
rect 75423 27992 75516 28078
rect 75076 27910 75516 27992
rect 75076 27824 75169 27910
rect 75255 27824 75337 27910
rect 75423 27824 75516 27910
rect 75076 27742 75516 27824
rect 75076 27656 75169 27742
rect 75255 27656 75337 27742
rect 75423 27656 75516 27742
rect 75076 27574 75516 27656
rect 75076 27488 75169 27574
rect 75255 27488 75337 27574
rect 75423 27488 75516 27574
rect 75076 27406 75516 27488
rect 75076 27320 75169 27406
rect 75255 27320 75337 27406
rect 75423 27320 75516 27406
rect 3103 27259 3489 27278
rect 3103 27236 3169 27259
rect 3255 27236 3337 27259
rect 3423 27236 3489 27259
rect 3103 27196 3112 27236
rect 3152 27196 3169 27236
rect 3255 27196 3276 27236
rect 3316 27196 3337 27236
rect 3423 27196 3440 27236
rect 3480 27196 3489 27236
rect 3103 27173 3169 27196
rect 3255 27173 3337 27196
rect 3423 27173 3489 27196
rect 3103 27154 3489 27173
rect 7103 27259 7489 27278
rect 7103 27236 7169 27259
rect 7255 27236 7337 27259
rect 7423 27236 7489 27259
rect 7103 27196 7112 27236
rect 7152 27196 7169 27236
rect 7255 27196 7276 27236
rect 7316 27196 7337 27236
rect 7423 27196 7440 27236
rect 7480 27196 7489 27236
rect 7103 27173 7169 27196
rect 7255 27173 7337 27196
rect 7423 27173 7489 27196
rect 7103 27154 7489 27173
rect 11103 27259 11489 27278
rect 11103 27236 11169 27259
rect 11255 27236 11337 27259
rect 11423 27236 11489 27259
rect 11103 27196 11112 27236
rect 11152 27196 11169 27236
rect 11255 27196 11276 27236
rect 11316 27196 11337 27236
rect 11423 27196 11440 27236
rect 11480 27196 11489 27236
rect 11103 27173 11169 27196
rect 11255 27173 11337 27196
rect 11423 27173 11489 27196
rect 11103 27154 11489 27173
rect 15103 27259 15489 27278
rect 15103 27236 15169 27259
rect 15255 27236 15337 27259
rect 15423 27236 15489 27259
rect 15103 27196 15112 27236
rect 15152 27196 15169 27236
rect 15255 27196 15276 27236
rect 15316 27196 15337 27236
rect 15423 27196 15440 27236
rect 15480 27196 15489 27236
rect 15103 27173 15169 27196
rect 15255 27173 15337 27196
rect 15423 27173 15489 27196
rect 15103 27154 15489 27173
rect 19103 27259 19489 27278
rect 19103 27236 19169 27259
rect 19255 27236 19337 27259
rect 19423 27236 19489 27259
rect 19103 27196 19112 27236
rect 19152 27196 19169 27236
rect 19255 27196 19276 27236
rect 19316 27196 19337 27236
rect 19423 27196 19440 27236
rect 19480 27196 19489 27236
rect 19103 27173 19169 27196
rect 19255 27173 19337 27196
rect 19423 27173 19489 27196
rect 19103 27154 19489 27173
rect 23103 27259 23489 27278
rect 23103 27236 23169 27259
rect 23255 27236 23337 27259
rect 23423 27236 23489 27259
rect 23103 27196 23112 27236
rect 23152 27196 23169 27236
rect 23255 27196 23276 27236
rect 23316 27196 23337 27236
rect 23423 27196 23440 27236
rect 23480 27196 23489 27236
rect 23103 27173 23169 27196
rect 23255 27173 23337 27196
rect 23423 27173 23489 27196
rect 23103 27154 23489 27173
rect 27103 27259 27489 27278
rect 27103 27236 27169 27259
rect 27255 27236 27337 27259
rect 27423 27236 27489 27259
rect 27103 27196 27112 27236
rect 27152 27196 27169 27236
rect 27255 27196 27276 27236
rect 27316 27196 27337 27236
rect 27423 27196 27440 27236
rect 27480 27196 27489 27236
rect 27103 27173 27169 27196
rect 27255 27173 27337 27196
rect 27423 27173 27489 27196
rect 27103 27154 27489 27173
rect 31103 27259 31489 27278
rect 31103 27236 31169 27259
rect 31255 27236 31337 27259
rect 31423 27236 31489 27259
rect 31103 27196 31112 27236
rect 31152 27196 31169 27236
rect 31255 27196 31276 27236
rect 31316 27196 31337 27236
rect 31423 27196 31440 27236
rect 31480 27196 31489 27236
rect 31103 27173 31169 27196
rect 31255 27173 31337 27196
rect 31423 27173 31489 27196
rect 31103 27154 31489 27173
rect 35103 27259 35489 27278
rect 35103 27236 35169 27259
rect 35255 27236 35337 27259
rect 35423 27236 35489 27259
rect 35103 27196 35112 27236
rect 35152 27196 35169 27236
rect 35255 27196 35276 27236
rect 35316 27196 35337 27236
rect 35423 27196 35440 27236
rect 35480 27196 35489 27236
rect 35103 27173 35169 27196
rect 35255 27173 35337 27196
rect 35423 27173 35489 27196
rect 35103 27154 35489 27173
rect 39103 27259 39489 27278
rect 39103 27236 39169 27259
rect 39255 27236 39337 27259
rect 39423 27236 39489 27259
rect 39103 27196 39112 27236
rect 39152 27196 39169 27236
rect 39255 27196 39276 27236
rect 39316 27196 39337 27236
rect 39423 27196 39440 27236
rect 39480 27196 39489 27236
rect 39103 27173 39169 27196
rect 39255 27173 39337 27196
rect 39423 27173 39489 27196
rect 39103 27154 39489 27173
rect 43103 27259 43489 27278
rect 43103 27236 43169 27259
rect 43255 27236 43337 27259
rect 43423 27236 43489 27259
rect 43103 27196 43112 27236
rect 43152 27196 43169 27236
rect 43255 27196 43276 27236
rect 43316 27196 43337 27236
rect 43423 27196 43440 27236
rect 43480 27196 43489 27236
rect 43103 27173 43169 27196
rect 43255 27173 43337 27196
rect 43423 27173 43489 27196
rect 43103 27154 43489 27173
rect 47103 27259 47489 27278
rect 47103 27236 47169 27259
rect 47255 27236 47337 27259
rect 47423 27236 47489 27259
rect 47103 27196 47112 27236
rect 47152 27196 47169 27236
rect 47255 27196 47276 27236
rect 47316 27196 47337 27236
rect 47423 27196 47440 27236
rect 47480 27196 47489 27236
rect 47103 27173 47169 27196
rect 47255 27173 47337 27196
rect 47423 27173 47489 27196
rect 47103 27154 47489 27173
rect 51103 27259 51489 27278
rect 51103 27236 51169 27259
rect 51255 27236 51337 27259
rect 51423 27236 51489 27259
rect 51103 27196 51112 27236
rect 51152 27196 51169 27236
rect 51255 27196 51276 27236
rect 51316 27196 51337 27236
rect 51423 27196 51440 27236
rect 51480 27196 51489 27236
rect 51103 27173 51169 27196
rect 51255 27173 51337 27196
rect 51423 27173 51489 27196
rect 51103 27154 51489 27173
rect 55103 27259 55489 27278
rect 55103 27236 55169 27259
rect 55255 27236 55337 27259
rect 55423 27236 55489 27259
rect 55103 27196 55112 27236
rect 55152 27196 55169 27236
rect 55255 27196 55276 27236
rect 55316 27196 55337 27236
rect 55423 27196 55440 27236
rect 55480 27196 55489 27236
rect 55103 27173 55169 27196
rect 55255 27173 55337 27196
rect 55423 27173 55489 27196
rect 55103 27154 55489 27173
rect 59103 27259 59489 27278
rect 59103 27236 59169 27259
rect 59255 27236 59337 27259
rect 59423 27236 59489 27259
rect 59103 27196 59112 27236
rect 59152 27196 59169 27236
rect 59255 27196 59276 27236
rect 59316 27196 59337 27236
rect 59423 27196 59440 27236
rect 59480 27196 59489 27236
rect 59103 27173 59169 27196
rect 59255 27173 59337 27196
rect 59423 27173 59489 27196
rect 59103 27154 59489 27173
rect 63103 27259 63489 27278
rect 63103 27236 63169 27259
rect 63255 27236 63337 27259
rect 63423 27236 63489 27259
rect 63103 27196 63112 27236
rect 63152 27196 63169 27236
rect 63255 27196 63276 27236
rect 63316 27196 63337 27236
rect 63423 27196 63440 27236
rect 63480 27196 63489 27236
rect 63103 27173 63169 27196
rect 63255 27173 63337 27196
rect 63423 27173 63489 27196
rect 63103 27154 63489 27173
rect 67103 27259 67489 27278
rect 67103 27236 67169 27259
rect 67255 27236 67337 27259
rect 67423 27236 67489 27259
rect 67103 27196 67112 27236
rect 67152 27196 67169 27236
rect 67255 27196 67276 27236
rect 67316 27196 67337 27236
rect 67423 27196 67440 27236
rect 67480 27196 67489 27236
rect 67103 27173 67169 27196
rect 67255 27173 67337 27196
rect 67423 27173 67489 27196
rect 67103 27154 67489 27173
rect 75076 27238 75516 27320
rect 75076 27152 75169 27238
rect 75255 27152 75337 27238
rect 75423 27152 75516 27238
rect 75076 27070 75516 27152
rect 75076 26984 75169 27070
rect 75255 26984 75337 27070
rect 75423 26984 75516 27070
rect 75076 26902 75516 26984
rect 75076 26816 75169 26902
rect 75255 26816 75337 26902
rect 75423 26816 75516 26902
rect 75076 26734 75516 26816
rect 75076 26648 75169 26734
rect 75255 26648 75337 26734
rect 75423 26648 75516 26734
rect 75076 26566 75516 26648
rect 4343 26503 4729 26522
rect 4343 26480 4409 26503
rect 4495 26480 4577 26503
rect 4663 26480 4729 26503
rect 4343 26440 4352 26480
rect 4392 26440 4409 26480
rect 4495 26440 4516 26480
rect 4556 26440 4577 26480
rect 4663 26440 4680 26480
rect 4720 26440 4729 26480
rect 4343 26417 4409 26440
rect 4495 26417 4577 26440
rect 4663 26417 4729 26440
rect 4343 26398 4729 26417
rect 8343 26503 8729 26522
rect 8343 26480 8409 26503
rect 8495 26480 8577 26503
rect 8663 26480 8729 26503
rect 8343 26440 8352 26480
rect 8392 26440 8409 26480
rect 8495 26440 8516 26480
rect 8556 26440 8577 26480
rect 8663 26440 8680 26480
rect 8720 26440 8729 26480
rect 8343 26417 8409 26440
rect 8495 26417 8577 26440
rect 8663 26417 8729 26440
rect 8343 26398 8729 26417
rect 12343 26503 12729 26522
rect 12343 26480 12409 26503
rect 12495 26480 12577 26503
rect 12663 26480 12729 26503
rect 12343 26440 12352 26480
rect 12392 26440 12409 26480
rect 12495 26440 12516 26480
rect 12556 26440 12577 26480
rect 12663 26440 12680 26480
rect 12720 26440 12729 26480
rect 12343 26417 12409 26440
rect 12495 26417 12577 26440
rect 12663 26417 12729 26440
rect 12343 26398 12729 26417
rect 16343 26503 16729 26522
rect 16343 26480 16409 26503
rect 16495 26480 16577 26503
rect 16663 26480 16729 26503
rect 16343 26440 16352 26480
rect 16392 26440 16409 26480
rect 16495 26440 16516 26480
rect 16556 26440 16577 26480
rect 16663 26440 16680 26480
rect 16720 26440 16729 26480
rect 16343 26417 16409 26440
rect 16495 26417 16577 26440
rect 16663 26417 16729 26440
rect 16343 26398 16729 26417
rect 20343 26503 20729 26522
rect 20343 26480 20409 26503
rect 20495 26480 20577 26503
rect 20663 26480 20729 26503
rect 20343 26440 20352 26480
rect 20392 26440 20409 26480
rect 20495 26440 20516 26480
rect 20556 26440 20577 26480
rect 20663 26440 20680 26480
rect 20720 26440 20729 26480
rect 20343 26417 20409 26440
rect 20495 26417 20577 26440
rect 20663 26417 20729 26440
rect 20343 26398 20729 26417
rect 24343 26503 24729 26522
rect 24343 26480 24409 26503
rect 24495 26480 24577 26503
rect 24663 26480 24729 26503
rect 24343 26440 24352 26480
rect 24392 26440 24409 26480
rect 24495 26440 24516 26480
rect 24556 26440 24577 26480
rect 24663 26440 24680 26480
rect 24720 26440 24729 26480
rect 24343 26417 24409 26440
rect 24495 26417 24577 26440
rect 24663 26417 24729 26440
rect 24343 26398 24729 26417
rect 28343 26503 28729 26522
rect 28343 26480 28409 26503
rect 28495 26480 28577 26503
rect 28663 26480 28729 26503
rect 28343 26440 28352 26480
rect 28392 26440 28409 26480
rect 28495 26440 28516 26480
rect 28556 26440 28577 26480
rect 28663 26440 28680 26480
rect 28720 26440 28729 26480
rect 28343 26417 28409 26440
rect 28495 26417 28577 26440
rect 28663 26417 28729 26440
rect 28343 26398 28729 26417
rect 32343 26503 32729 26522
rect 32343 26480 32409 26503
rect 32495 26480 32577 26503
rect 32663 26480 32729 26503
rect 32343 26440 32352 26480
rect 32392 26440 32409 26480
rect 32495 26440 32516 26480
rect 32556 26440 32577 26480
rect 32663 26440 32680 26480
rect 32720 26440 32729 26480
rect 32343 26417 32409 26440
rect 32495 26417 32577 26440
rect 32663 26417 32729 26440
rect 32343 26398 32729 26417
rect 36343 26503 36729 26522
rect 36343 26480 36409 26503
rect 36495 26480 36577 26503
rect 36663 26480 36729 26503
rect 36343 26440 36352 26480
rect 36392 26440 36409 26480
rect 36495 26440 36516 26480
rect 36556 26440 36577 26480
rect 36663 26440 36680 26480
rect 36720 26440 36729 26480
rect 36343 26417 36409 26440
rect 36495 26417 36577 26440
rect 36663 26417 36729 26440
rect 36343 26398 36729 26417
rect 40343 26503 40729 26522
rect 40343 26480 40409 26503
rect 40495 26480 40577 26503
rect 40663 26480 40729 26503
rect 40343 26440 40352 26480
rect 40392 26440 40409 26480
rect 40495 26440 40516 26480
rect 40556 26440 40577 26480
rect 40663 26440 40680 26480
rect 40720 26440 40729 26480
rect 40343 26417 40409 26440
rect 40495 26417 40577 26440
rect 40663 26417 40729 26440
rect 40343 26398 40729 26417
rect 44343 26503 44729 26522
rect 44343 26480 44409 26503
rect 44495 26480 44577 26503
rect 44663 26480 44729 26503
rect 44343 26440 44352 26480
rect 44392 26440 44409 26480
rect 44495 26440 44516 26480
rect 44556 26440 44577 26480
rect 44663 26440 44680 26480
rect 44720 26440 44729 26480
rect 44343 26417 44409 26440
rect 44495 26417 44577 26440
rect 44663 26417 44729 26440
rect 44343 26398 44729 26417
rect 48343 26503 48729 26522
rect 48343 26480 48409 26503
rect 48495 26480 48577 26503
rect 48663 26480 48729 26503
rect 48343 26440 48352 26480
rect 48392 26440 48409 26480
rect 48495 26440 48516 26480
rect 48556 26440 48577 26480
rect 48663 26440 48680 26480
rect 48720 26440 48729 26480
rect 48343 26417 48409 26440
rect 48495 26417 48577 26440
rect 48663 26417 48729 26440
rect 48343 26398 48729 26417
rect 52343 26503 52729 26522
rect 52343 26480 52409 26503
rect 52495 26480 52577 26503
rect 52663 26480 52729 26503
rect 52343 26440 52352 26480
rect 52392 26440 52409 26480
rect 52495 26440 52516 26480
rect 52556 26440 52577 26480
rect 52663 26440 52680 26480
rect 52720 26440 52729 26480
rect 52343 26417 52409 26440
rect 52495 26417 52577 26440
rect 52663 26417 52729 26440
rect 52343 26398 52729 26417
rect 56343 26503 56729 26522
rect 56343 26480 56409 26503
rect 56495 26480 56577 26503
rect 56663 26480 56729 26503
rect 56343 26440 56352 26480
rect 56392 26440 56409 26480
rect 56495 26440 56516 26480
rect 56556 26440 56577 26480
rect 56663 26440 56680 26480
rect 56720 26440 56729 26480
rect 56343 26417 56409 26440
rect 56495 26417 56577 26440
rect 56663 26417 56729 26440
rect 56343 26398 56729 26417
rect 60343 26503 60729 26522
rect 60343 26480 60409 26503
rect 60495 26480 60577 26503
rect 60663 26480 60729 26503
rect 60343 26440 60352 26480
rect 60392 26440 60409 26480
rect 60495 26440 60516 26480
rect 60556 26440 60577 26480
rect 60663 26440 60680 26480
rect 60720 26440 60729 26480
rect 60343 26417 60409 26440
rect 60495 26417 60577 26440
rect 60663 26417 60729 26440
rect 60343 26398 60729 26417
rect 64343 26503 64729 26522
rect 64343 26480 64409 26503
rect 64495 26480 64577 26503
rect 64663 26480 64729 26503
rect 64343 26440 64352 26480
rect 64392 26440 64409 26480
rect 64495 26440 64516 26480
rect 64556 26440 64577 26480
rect 64663 26440 64680 26480
rect 64720 26440 64729 26480
rect 64343 26417 64409 26440
rect 64495 26417 64577 26440
rect 64663 26417 64729 26440
rect 64343 26398 64729 26417
rect 68343 26503 68729 26522
rect 68343 26480 68409 26503
rect 68495 26480 68577 26503
rect 68663 26480 68729 26503
rect 68343 26440 68352 26480
rect 68392 26440 68409 26480
rect 68495 26440 68516 26480
rect 68556 26440 68577 26480
rect 68663 26440 68680 26480
rect 68720 26440 68729 26480
rect 68343 26417 68409 26440
rect 68495 26417 68577 26440
rect 68663 26417 68729 26440
rect 68343 26398 68729 26417
rect 75076 26480 75169 26566
rect 75255 26480 75337 26566
rect 75423 26480 75516 26566
rect 75076 26398 75516 26480
rect 75076 26312 75169 26398
rect 75255 26312 75337 26398
rect 75423 26312 75516 26398
rect 75076 26230 75516 26312
rect 75076 26144 75169 26230
rect 75255 26144 75337 26230
rect 75423 26144 75516 26230
rect 75076 26014 75516 26144
rect 79076 28246 79516 28376
rect 79076 28160 79169 28246
rect 79255 28160 79337 28246
rect 79423 28160 79516 28246
rect 79076 28078 79516 28160
rect 79076 27992 79169 28078
rect 79255 27992 79337 28078
rect 79423 27992 79516 28078
rect 79076 27910 79516 27992
rect 79076 27824 79169 27910
rect 79255 27824 79337 27910
rect 79423 27824 79516 27910
rect 79076 27742 79516 27824
rect 79076 27656 79169 27742
rect 79255 27656 79337 27742
rect 79423 27656 79516 27742
rect 79076 27574 79516 27656
rect 79076 27488 79169 27574
rect 79255 27488 79337 27574
rect 79423 27488 79516 27574
rect 79076 27406 79516 27488
rect 79076 27320 79169 27406
rect 79255 27320 79337 27406
rect 79423 27320 79516 27406
rect 79076 27238 79516 27320
rect 79076 27152 79169 27238
rect 79255 27152 79337 27238
rect 79423 27152 79516 27238
rect 79076 27070 79516 27152
rect 79076 26984 79169 27070
rect 79255 26984 79337 27070
rect 79423 26984 79516 27070
rect 79076 26902 79516 26984
rect 79076 26816 79169 26902
rect 79255 26816 79337 26902
rect 79423 26816 79516 26902
rect 79076 26734 79516 26816
rect 79076 26648 79169 26734
rect 79255 26648 79337 26734
rect 79423 26648 79516 26734
rect 79076 26566 79516 26648
rect 79076 26480 79169 26566
rect 79255 26480 79337 26566
rect 79423 26480 79516 26566
rect 79076 26398 79516 26480
rect 79076 26312 79169 26398
rect 79255 26312 79337 26398
rect 79423 26312 79516 26398
rect 79076 26230 79516 26312
rect 79076 26144 79169 26230
rect 79255 26144 79337 26230
rect 79423 26144 79516 26230
rect 79076 26014 79516 26144
rect 83076 28246 83516 28376
rect 83076 28160 83169 28246
rect 83255 28160 83337 28246
rect 83423 28160 83516 28246
rect 83076 28078 83516 28160
rect 83076 27992 83169 28078
rect 83255 27992 83337 28078
rect 83423 27992 83516 28078
rect 83076 27910 83516 27992
rect 83076 27824 83169 27910
rect 83255 27824 83337 27910
rect 83423 27824 83516 27910
rect 83076 27742 83516 27824
rect 83076 27656 83169 27742
rect 83255 27656 83337 27742
rect 83423 27656 83516 27742
rect 83076 27574 83516 27656
rect 83076 27488 83169 27574
rect 83255 27488 83337 27574
rect 83423 27488 83516 27574
rect 83076 27406 83516 27488
rect 83076 27320 83169 27406
rect 83255 27320 83337 27406
rect 83423 27320 83516 27406
rect 83076 27238 83516 27320
rect 83076 27152 83169 27238
rect 83255 27152 83337 27238
rect 83423 27152 83516 27238
rect 83076 27070 83516 27152
rect 83076 26984 83169 27070
rect 83255 26984 83337 27070
rect 83423 26984 83516 27070
rect 83076 26902 83516 26984
rect 83076 26816 83169 26902
rect 83255 26816 83337 26902
rect 83423 26816 83516 26902
rect 83076 26734 83516 26816
rect 83076 26648 83169 26734
rect 83255 26648 83337 26734
rect 83423 26648 83516 26734
rect 83076 26566 83516 26648
rect 83076 26480 83169 26566
rect 83255 26480 83337 26566
rect 83423 26480 83516 26566
rect 83076 26398 83516 26480
rect 83076 26312 83169 26398
rect 83255 26312 83337 26398
rect 83423 26312 83516 26398
rect 83076 26230 83516 26312
rect 83076 26144 83169 26230
rect 83255 26144 83337 26230
rect 83423 26144 83516 26230
rect 83076 26014 83516 26144
rect 87076 28246 87516 28376
rect 87076 28160 87169 28246
rect 87255 28160 87337 28246
rect 87423 28160 87516 28246
rect 87076 28078 87516 28160
rect 87076 27992 87169 28078
rect 87255 27992 87337 28078
rect 87423 27992 87516 28078
rect 87076 27910 87516 27992
rect 87076 27824 87169 27910
rect 87255 27824 87337 27910
rect 87423 27824 87516 27910
rect 87076 27742 87516 27824
rect 87076 27656 87169 27742
rect 87255 27656 87337 27742
rect 87423 27656 87516 27742
rect 87076 27574 87516 27656
rect 87076 27488 87169 27574
rect 87255 27488 87337 27574
rect 87423 27488 87516 27574
rect 87076 27406 87516 27488
rect 87076 27320 87169 27406
rect 87255 27320 87337 27406
rect 87423 27320 87516 27406
rect 87076 27238 87516 27320
rect 87076 27152 87169 27238
rect 87255 27152 87337 27238
rect 87423 27152 87516 27238
rect 87076 27070 87516 27152
rect 87076 26984 87169 27070
rect 87255 26984 87337 27070
rect 87423 26984 87516 27070
rect 87076 26902 87516 26984
rect 87076 26816 87169 26902
rect 87255 26816 87337 26902
rect 87423 26816 87516 26902
rect 87076 26734 87516 26816
rect 87076 26648 87169 26734
rect 87255 26648 87337 26734
rect 87423 26648 87516 26734
rect 87076 26566 87516 26648
rect 87076 26480 87169 26566
rect 87255 26480 87337 26566
rect 87423 26480 87516 26566
rect 87076 26398 87516 26480
rect 87076 26312 87169 26398
rect 87255 26312 87337 26398
rect 87423 26312 87516 26398
rect 87076 26230 87516 26312
rect 87076 26144 87169 26230
rect 87255 26144 87337 26230
rect 87423 26144 87516 26230
rect 87076 26014 87516 26144
rect 91076 28246 91516 28376
rect 91076 28160 91169 28246
rect 91255 28160 91337 28246
rect 91423 28160 91516 28246
rect 91076 28078 91516 28160
rect 91076 27992 91169 28078
rect 91255 27992 91337 28078
rect 91423 27992 91516 28078
rect 91076 27910 91516 27992
rect 91076 27824 91169 27910
rect 91255 27824 91337 27910
rect 91423 27824 91516 27910
rect 91076 27742 91516 27824
rect 91076 27656 91169 27742
rect 91255 27656 91337 27742
rect 91423 27656 91516 27742
rect 91076 27574 91516 27656
rect 91076 27488 91169 27574
rect 91255 27488 91337 27574
rect 91423 27488 91516 27574
rect 91076 27406 91516 27488
rect 91076 27320 91169 27406
rect 91255 27320 91337 27406
rect 91423 27320 91516 27406
rect 91076 27238 91516 27320
rect 91076 27152 91169 27238
rect 91255 27152 91337 27238
rect 91423 27152 91516 27238
rect 91076 27070 91516 27152
rect 91076 26984 91169 27070
rect 91255 26984 91337 27070
rect 91423 26984 91516 27070
rect 91076 26902 91516 26984
rect 91076 26816 91169 26902
rect 91255 26816 91337 26902
rect 91423 26816 91516 26902
rect 91076 26734 91516 26816
rect 91076 26648 91169 26734
rect 91255 26648 91337 26734
rect 91423 26648 91516 26734
rect 91076 26566 91516 26648
rect 91076 26480 91169 26566
rect 91255 26480 91337 26566
rect 91423 26480 91516 26566
rect 91076 26398 91516 26480
rect 91076 26312 91169 26398
rect 91255 26312 91337 26398
rect 91423 26312 91516 26398
rect 91076 26230 91516 26312
rect 91076 26144 91169 26230
rect 91255 26144 91337 26230
rect 91423 26144 91516 26230
rect 91076 26014 91516 26144
rect 95076 28246 95516 28376
rect 95076 28160 95169 28246
rect 95255 28160 95337 28246
rect 95423 28160 95516 28246
rect 95076 28078 95516 28160
rect 95076 27992 95169 28078
rect 95255 27992 95337 28078
rect 95423 27992 95516 28078
rect 95076 27910 95516 27992
rect 95076 27824 95169 27910
rect 95255 27824 95337 27910
rect 95423 27824 95516 27910
rect 95076 27742 95516 27824
rect 95076 27656 95169 27742
rect 95255 27656 95337 27742
rect 95423 27656 95516 27742
rect 95076 27574 95516 27656
rect 95076 27488 95169 27574
rect 95255 27488 95337 27574
rect 95423 27488 95516 27574
rect 95076 27406 95516 27488
rect 95076 27320 95169 27406
rect 95255 27320 95337 27406
rect 95423 27320 95516 27406
rect 95076 27238 95516 27320
rect 95076 27152 95169 27238
rect 95255 27152 95337 27238
rect 95423 27152 95516 27238
rect 95076 27070 95516 27152
rect 95076 26984 95169 27070
rect 95255 26984 95337 27070
rect 95423 26984 95516 27070
rect 95076 26902 95516 26984
rect 95076 26816 95169 26902
rect 95255 26816 95337 26902
rect 95423 26816 95516 26902
rect 95076 26734 95516 26816
rect 95076 26648 95169 26734
rect 95255 26648 95337 26734
rect 95423 26648 95516 26734
rect 95076 26566 95516 26648
rect 95076 26480 95169 26566
rect 95255 26480 95337 26566
rect 95423 26480 95516 26566
rect 95076 26398 95516 26480
rect 95076 26312 95169 26398
rect 95255 26312 95337 26398
rect 95423 26312 95516 26398
rect 95076 26230 95516 26312
rect 95076 26144 95169 26230
rect 95255 26144 95337 26230
rect 95423 26144 95516 26230
rect 95076 26014 95516 26144
rect 3103 25747 3489 25766
rect 3103 25724 3169 25747
rect 3255 25724 3337 25747
rect 3423 25724 3489 25747
rect 3103 25684 3112 25724
rect 3152 25684 3169 25724
rect 3255 25684 3276 25724
rect 3316 25684 3337 25724
rect 3423 25684 3440 25724
rect 3480 25684 3489 25724
rect 3103 25661 3169 25684
rect 3255 25661 3337 25684
rect 3423 25661 3489 25684
rect 3103 25642 3489 25661
rect 7103 25747 7489 25766
rect 7103 25724 7169 25747
rect 7255 25724 7337 25747
rect 7423 25724 7489 25747
rect 7103 25684 7112 25724
rect 7152 25684 7169 25724
rect 7255 25684 7276 25724
rect 7316 25684 7337 25724
rect 7423 25684 7440 25724
rect 7480 25684 7489 25724
rect 7103 25661 7169 25684
rect 7255 25661 7337 25684
rect 7423 25661 7489 25684
rect 7103 25642 7489 25661
rect 11103 25747 11489 25766
rect 11103 25724 11169 25747
rect 11255 25724 11337 25747
rect 11423 25724 11489 25747
rect 11103 25684 11112 25724
rect 11152 25684 11169 25724
rect 11255 25684 11276 25724
rect 11316 25684 11337 25724
rect 11423 25684 11440 25724
rect 11480 25684 11489 25724
rect 11103 25661 11169 25684
rect 11255 25661 11337 25684
rect 11423 25661 11489 25684
rect 11103 25642 11489 25661
rect 15103 25747 15489 25766
rect 15103 25724 15169 25747
rect 15255 25724 15337 25747
rect 15423 25724 15489 25747
rect 15103 25684 15112 25724
rect 15152 25684 15169 25724
rect 15255 25684 15276 25724
rect 15316 25684 15337 25724
rect 15423 25684 15440 25724
rect 15480 25684 15489 25724
rect 15103 25661 15169 25684
rect 15255 25661 15337 25684
rect 15423 25661 15489 25684
rect 15103 25642 15489 25661
rect 19103 25747 19489 25766
rect 19103 25724 19169 25747
rect 19255 25724 19337 25747
rect 19423 25724 19489 25747
rect 19103 25684 19112 25724
rect 19152 25684 19169 25724
rect 19255 25684 19276 25724
rect 19316 25684 19337 25724
rect 19423 25684 19440 25724
rect 19480 25684 19489 25724
rect 19103 25661 19169 25684
rect 19255 25661 19337 25684
rect 19423 25661 19489 25684
rect 19103 25642 19489 25661
rect 23103 25747 23489 25766
rect 23103 25724 23169 25747
rect 23255 25724 23337 25747
rect 23423 25724 23489 25747
rect 23103 25684 23112 25724
rect 23152 25684 23169 25724
rect 23255 25684 23276 25724
rect 23316 25684 23337 25724
rect 23423 25684 23440 25724
rect 23480 25684 23489 25724
rect 23103 25661 23169 25684
rect 23255 25661 23337 25684
rect 23423 25661 23489 25684
rect 23103 25642 23489 25661
rect 27103 25747 27489 25766
rect 27103 25724 27169 25747
rect 27255 25724 27337 25747
rect 27423 25724 27489 25747
rect 27103 25684 27112 25724
rect 27152 25684 27169 25724
rect 27255 25684 27276 25724
rect 27316 25684 27337 25724
rect 27423 25684 27440 25724
rect 27480 25684 27489 25724
rect 27103 25661 27169 25684
rect 27255 25661 27337 25684
rect 27423 25661 27489 25684
rect 27103 25642 27489 25661
rect 31103 25747 31489 25766
rect 31103 25724 31169 25747
rect 31255 25724 31337 25747
rect 31423 25724 31489 25747
rect 31103 25684 31112 25724
rect 31152 25684 31169 25724
rect 31255 25684 31276 25724
rect 31316 25684 31337 25724
rect 31423 25684 31440 25724
rect 31480 25684 31489 25724
rect 31103 25661 31169 25684
rect 31255 25661 31337 25684
rect 31423 25661 31489 25684
rect 31103 25642 31489 25661
rect 35103 25747 35489 25766
rect 35103 25724 35169 25747
rect 35255 25724 35337 25747
rect 35423 25724 35489 25747
rect 35103 25684 35112 25724
rect 35152 25684 35169 25724
rect 35255 25684 35276 25724
rect 35316 25684 35337 25724
rect 35423 25684 35440 25724
rect 35480 25684 35489 25724
rect 35103 25661 35169 25684
rect 35255 25661 35337 25684
rect 35423 25661 35489 25684
rect 35103 25642 35489 25661
rect 39103 25747 39489 25766
rect 39103 25724 39169 25747
rect 39255 25724 39337 25747
rect 39423 25724 39489 25747
rect 39103 25684 39112 25724
rect 39152 25684 39169 25724
rect 39255 25684 39276 25724
rect 39316 25684 39337 25724
rect 39423 25684 39440 25724
rect 39480 25684 39489 25724
rect 39103 25661 39169 25684
rect 39255 25661 39337 25684
rect 39423 25661 39489 25684
rect 39103 25642 39489 25661
rect 43103 25747 43489 25766
rect 43103 25724 43169 25747
rect 43255 25724 43337 25747
rect 43423 25724 43489 25747
rect 43103 25684 43112 25724
rect 43152 25684 43169 25724
rect 43255 25684 43276 25724
rect 43316 25684 43337 25724
rect 43423 25684 43440 25724
rect 43480 25684 43489 25724
rect 43103 25661 43169 25684
rect 43255 25661 43337 25684
rect 43423 25661 43489 25684
rect 43103 25642 43489 25661
rect 47103 25747 47489 25766
rect 47103 25724 47169 25747
rect 47255 25724 47337 25747
rect 47423 25724 47489 25747
rect 47103 25684 47112 25724
rect 47152 25684 47169 25724
rect 47255 25684 47276 25724
rect 47316 25684 47337 25724
rect 47423 25684 47440 25724
rect 47480 25684 47489 25724
rect 47103 25661 47169 25684
rect 47255 25661 47337 25684
rect 47423 25661 47489 25684
rect 47103 25642 47489 25661
rect 51103 25747 51489 25766
rect 51103 25724 51169 25747
rect 51255 25724 51337 25747
rect 51423 25724 51489 25747
rect 51103 25684 51112 25724
rect 51152 25684 51169 25724
rect 51255 25684 51276 25724
rect 51316 25684 51337 25724
rect 51423 25684 51440 25724
rect 51480 25684 51489 25724
rect 51103 25661 51169 25684
rect 51255 25661 51337 25684
rect 51423 25661 51489 25684
rect 51103 25642 51489 25661
rect 55103 25747 55489 25766
rect 55103 25724 55169 25747
rect 55255 25724 55337 25747
rect 55423 25724 55489 25747
rect 55103 25684 55112 25724
rect 55152 25684 55169 25724
rect 55255 25684 55276 25724
rect 55316 25684 55337 25724
rect 55423 25684 55440 25724
rect 55480 25684 55489 25724
rect 55103 25661 55169 25684
rect 55255 25661 55337 25684
rect 55423 25661 55489 25684
rect 55103 25642 55489 25661
rect 59103 25747 59489 25766
rect 59103 25724 59169 25747
rect 59255 25724 59337 25747
rect 59423 25724 59489 25747
rect 59103 25684 59112 25724
rect 59152 25684 59169 25724
rect 59255 25684 59276 25724
rect 59316 25684 59337 25724
rect 59423 25684 59440 25724
rect 59480 25684 59489 25724
rect 59103 25661 59169 25684
rect 59255 25661 59337 25684
rect 59423 25661 59489 25684
rect 59103 25642 59489 25661
rect 63103 25747 63489 25766
rect 63103 25724 63169 25747
rect 63255 25724 63337 25747
rect 63423 25724 63489 25747
rect 63103 25684 63112 25724
rect 63152 25684 63169 25724
rect 63255 25684 63276 25724
rect 63316 25684 63337 25724
rect 63423 25684 63440 25724
rect 63480 25684 63489 25724
rect 63103 25661 63169 25684
rect 63255 25661 63337 25684
rect 63423 25661 63489 25684
rect 63103 25642 63489 25661
rect 67103 25747 67489 25766
rect 67103 25724 67169 25747
rect 67255 25724 67337 25747
rect 67423 25724 67489 25747
rect 67103 25684 67112 25724
rect 67152 25684 67169 25724
rect 67255 25684 67276 25724
rect 67316 25684 67337 25724
rect 67423 25684 67440 25724
rect 67480 25684 67489 25724
rect 67103 25661 67169 25684
rect 67255 25661 67337 25684
rect 67423 25661 67489 25684
rect 67103 25642 67489 25661
rect 71779 25600 71788 25640
rect 71828 25600 72940 25640
rect 72980 25600 72989 25640
rect 4343 24991 4729 25010
rect 4343 24968 4409 24991
rect 4495 24968 4577 24991
rect 4663 24968 4729 24991
rect 4343 24928 4352 24968
rect 4392 24928 4409 24968
rect 4495 24928 4516 24968
rect 4556 24928 4577 24968
rect 4663 24928 4680 24968
rect 4720 24928 4729 24968
rect 4343 24905 4409 24928
rect 4495 24905 4577 24928
rect 4663 24905 4729 24928
rect 4343 24886 4729 24905
rect 8343 24991 8729 25010
rect 8343 24968 8409 24991
rect 8495 24968 8577 24991
rect 8663 24968 8729 24991
rect 8343 24928 8352 24968
rect 8392 24928 8409 24968
rect 8495 24928 8516 24968
rect 8556 24928 8577 24968
rect 8663 24928 8680 24968
rect 8720 24928 8729 24968
rect 8343 24905 8409 24928
rect 8495 24905 8577 24928
rect 8663 24905 8729 24928
rect 8343 24886 8729 24905
rect 12343 24991 12729 25010
rect 12343 24968 12409 24991
rect 12495 24968 12577 24991
rect 12663 24968 12729 24991
rect 12343 24928 12352 24968
rect 12392 24928 12409 24968
rect 12495 24928 12516 24968
rect 12556 24928 12577 24968
rect 12663 24928 12680 24968
rect 12720 24928 12729 24968
rect 12343 24905 12409 24928
rect 12495 24905 12577 24928
rect 12663 24905 12729 24928
rect 12343 24886 12729 24905
rect 16343 24991 16729 25010
rect 16343 24968 16409 24991
rect 16495 24968 16577 24991
rect 16663 24968 16729 24991
rect 16343 24928 16352 24968
rect 16392 24928 16409 24968
rect 16495 24928 16516 24968
rect 16556 24928 16577 24968
rect 16663 24928 16680 24968
rect 16720 24928 16729 24968
rect 16343 24905 16409 24928
rect 16495 24905 16577 24928
rect 16663 24905 16729 24928
rect 16343 24886 16729 24905
rect 20343 24991 20729 25010
rect 20343 24968 20409 24991
rect 20495 24968 20577 24991
rect 20663 24968 20729 24991
rect 20343 24928 20352 24968
rect 20392 24928 20409 24968
rect 20495 24928 20516 24968
rect 20556 24928 20577 24968
rect 20663 24928 20680 24968
rect 20720 24928 20729 24968
rect 20343 24905 20409 24928
rect 20495 24905 20577 24928
rect 20663 24905 20729 24928
rect 20343 24886 20729 24905
rect 24343 24991 24729 25010
rect 24343 24968 24409 24991
rect 24495 24968 24577 24991
rect 24663 24968 24729 24991
rect 24343 24928 24352 24968
rect 24392 24928 24409 24968
rect 24495 24928 24516 24968
rect 24556 24928 24577 24968
rect 24663 24928 24680 24968
rect 24720 24928 24729 24968
rect 24343 24905 24409 24928
rect 24495 24905 24577 24928
rect 24663 24905 24729 24928
rect 24343 24886 24729 24905
rect 28343 24991 28729 25010
rect 28343 24968 28409 24991
rect 28495 24968 28577 24991
rect 28663 24968 28729 24991
rect 28343 24928 28352 24968
rect 28392 24928 28409 24968
rect 28495 24928 28516 24968
rect 28556 24928 28577 24968
rect 28663 24928 28680 24968
rect 28720 24928 28729 24968
rect 28343 24905 28409 24928
rect 28495 24905 28577 24928
rect 28663 24905 28729 24928
rect 28343 24886 28729 24905
rect 32343 24991 32729 25010
rect 32343 24968 32409 24991
rect 32495 24968 32577 24991
rect 32663 24968 32729 24991
rect 32343 24928 32352 24968
rect 32392 24928 32409 24968
rect 32495 24928 32516 24968
rect 32556 24928 32577 24968
rect 32663 24928 32680 24968
rect 32720 24928 32729 24968
rect 32343 24905 32409 24928
rect 32495 24905 32577 24928
rect 32663 24905 32729 24928
rect 32343 24886 32729 24905
rect 36343 24991 36729 25010
rect 36343 24968 36409 24991
rect 36495 24968 36577 24991
rect 36663 24968 36729 24991
rect 36343 24928 36352 24968
rect 36392 24928 36409 24968
rect 36495 24928 36516 24968
rect 36556 24928 36577 24968
rect 36663 24928 36680 24968
rect 36720 24928 36729 24968
rect 36343 24905 36409 24928
rect 36495 24905 36577 24928
rect 36663 24905 36729 24928
rect 36343 24886 36729 24905
rect 40343 24991 40729 25010
rect 40343 24968 40409 24991
rect 40495 24968 40577 24991
rect 40663 24968 40729 24991
rect 40343 24928 40352 24968
rect 40392 24928 40409 24968
rect 40495 24928 40516 24968
rect 40556 24928 40577 24968
rect 40663 24928 40680 24968
rect 40720 24928 40729 24968
rect 40343 24905 40409 24928
rect 40495 24905 40577 24928
rect 40663 24905 40729 24928
rect 40343 24886 40729 24905
rect 44343 24991 44729 25010
rect 44343 24968 44409 24991
rect 44495 24968 44577 24991
rect 44663 24968 44729 24991
rect 44343 24928 44352 24968
rect 44392 24928 44409 24968
rect 44495 24928 44516 24968
rect 44556 24928 44577 24968
rect 44663 24928 44680 24968
rect 44720 24928 44729 24968
rect 44343 24905 44409 24928
rect 44495 24905 44577 24928
rect 44663 24905 44729 24928
rect 44343 24886 44729 24905
rect 48343 24991 48729 25010
rect 48343 24968 48409 24991
rect 48495 24968 48577 24991
rect 48663 24968 48729 24991
rect 48343 24928 48352 24968
rect 48392 24928 48409 24968
rect 48495 24928 48516 24968
rect 48556 24928 48577 24968
rect 48663 24928 48680 24968
rect 48720 24928 48729 24968
rect 48343 24905 48409 24928
rect 48495 24905 48577 24928
rect 48663 24905 48729 24928
rect 48343 24886 48729 24905
rect 52343 24991 52729 25010
rect 52343 24968 52409 24991
rect 52495 24968 52577 24991
rect 52663 24968 52729 24991
rect 52343 24928 52352 24968
rect 52392 24928 52409 24968
rect 52495 24928 52516 24968
rect 52556 24928 52577 24968
rect 52663 24928 52680 24968
rect 52720 24928 52729 24968
rect 52343 24905 52409 24928
rect 52495 24905 52577 24928
rect 52663 24905 52729 24928
rect 52343 24886 52729 24905
rect 56343 24991 56729 25010
rect 56343 24968 56409 24991
rect 56495 24968 56577 24991
rect 56663 24968 56729 24991
rect 56343 24928 56352 24968
rect 56392 24928 56409 24968
rect 56495 24928 56516 24968
rect 56556 24928 56577 24968
rect 56663 24928 56680 24968
rect 56720 24928 56729 24968
rect 56343 24905 56409 24928
rect 56495 24905 56577 24928
rect 56663 24905 56729 24928
rect 56343 24886 56729 24905
rect 60343 24991 60729 25010
rect 60343 24968 60409 24991
rect 60495 24968 60577 24991
rect 60663 24968 60729 24991
rect 60343 24928 60352 24968
rect 60392 24928 60409 24968
rect 60495 24928 60516 24968
rect 60556 24928 60577 24968
rect 60663 24928 60680 24968
rect 60720 24928 60729 24968
rect 60343 24905 60409 24928
rect 60495 24905 60577 24928
rect 60663 24905 60729 24928
rect 60343 24886 60729 24905
rect 64343 24991 64729 25010
rect 64343 24968 64409 24991
rect 64495 24968 64577 24991
rect 64663 24968 64729 24991
rect 64343 24928 64352 24968
rect 64392 24928 64409 24968
rect 64495 24928 64516 24968
rect 64556 24928 64577 24968
rect 64663 24928 64680 24968
rect 64720 24928 64729 24968
rect 64343 24905 64409 24928
rect 64495 24905 64577 24928
rect 64663 24905 64729 24928
rect 64343 24886 64729 24905
rect 68343 24991 68729 25010
rect 68343 24968 68409 24991
rect 68495 24968 68577 24991
rect 68663 24968 68729 24991
rect 68343 24928 68352 24968
rect 68392 24928 68409 24968
rect 68495 24928 68516 24968
rect 68556 24928 68577 24968
rect 68663 24928 68680 24968
rect 68720 24928 68729 24968
rect 68343 24905 68409 24928
rect 68495 24905 68577 24928
rect 68663 24905 68729 24928
rect 68343 24886 68729 24905
rect 3103 24235 3489 24254
rect 3103 24212 3169 24235
rect 3255 24212 3337 24235
rect 3423 24212 3489 24235
rect 3103 24172 3112 24212
rect 3152 24172 3169 24212
rect 3255 24172 3276 24212
rect 3316 24172 3337 24212
rect 3423 24172 3440 24212
rect 3480 24172 3489 24212
rect 3103 24149 3169 24172
rect 3255 24149 3337 24172
rect 3423 24149 3489 24172
rect 3103 24130 3489 24149
rect 7103 24235 7489 24254
rect 7103 24212 7169 24235
rect 7255 24212 7337 24235
rect 7423 24212 7489 24235
rect 7103 24172 7112 24212
rect 7152 24172 7169 24212
rect 7255 24172 7276 24212
rect 7316 24172 7337 24212
rect 7423 24172 7440 24212
rect 7480 24172 7489 24212
rect 7103 24149 7169 24172
rect 7255 24149 7337 24172
rect 7423 24149 7489 24172
rect 7103 24130 7489 24149
rect 11103 24235 11489 24254
rect 11103 24212 11169 24235
rect 11255 24212 11337 24235
rect 11423 24212 11489 24235
rect 11103 24172 11112 24212
rect 11152 24172 11169 24212
rect 11255 24172 11276 24212
rect 11316 24172 11337 24212
rect 11423 24172 11440 24212
rect 11480 24172 11489 24212
rect 11103 24149 11169 24172
rect 11255 24149 11337 24172
rect 11423 24149 11489 24172
rect 11103 24130 11489 24149
rect 15103 24235 15489 24254
rect 15103 24212 15169 24235
rect 15255 24212 15337 24235
rect 15423 24212 15489 24235
rect 15103 24172 15112 24212
rect 15152 24172 15169 24212
rect 15255 24172 15276 24212
rect 15316 24172 15337 24212
rect 15423 24172 15440 24212
rect 15480 24172 15489 24212
rect 15103 24149 15169 24172
rect 15255 24149 15337 24172
rect 15423 24149 15489 24172
rect 15103 24130 15489 24149
rect 19103 24235 19489 24254
rect 19103 24212 19169 24235
rect 19255 24212 19337 24235
rect 19423 24212 19489 24235
rect 19103 24172 19112 24212
rect 19152 24172 19169 24212
rect 19255 24172 19276 24212
rect 19316 24172 19337 24212
rect 19423 24172 19440 24212
rect 19480 24172 19489 24212
rect 19103 24149 19169 24172
rect 19255 24149 19337 24172
rect 19423 24149 19489 24172
rect 19103 24130 19489 24149
rect 23103 24235 23489 24254
rect 23103 24212 23169 24235
rect 23255 24212 23337 24235
rect 23423 24212 23489 24235
rect 23103 24172 23112 24212
rect 23152 24172 23169 24212
rect 23255 24172 23276 24212
rect 23316 24172 23337 24212
rect 23423 24172 23440 24212
rect 23480 24172 23489 24212
rect 23103 24149 23169 24172
rect 23255 24149 23337 24172
rect 23423 24149 23489 24172
rect 23103 24130 23489 24149
rect 27103 24235 27489 24254
rect 27103 24212 27169 24235
rect 27255 24212 27337 24235
rect 27423 24212 27489 24235
rect 27103 24172 27112 24212
rect 27152 24172 27169 24212
rect 27255 24172 27276 24212
rect 27316 24172 27337 24212
rect 27423 24172 27440 24212
rect 27480 24172 27489 24212
rect 27103 24149 27169 24172
rect 27255 24149 27337 24172
rect 27423 24149 27489 24172
rect 27103 24130 27489 24149
rect 31103 24235 31489 24254
rect 31103 24212 31169 24235
rect 31255 24212 31337 24235
rect 31423 24212 31489 24235
rect 31103 24172 31112 24212
rect 31152 24172 31169 24212
rect 31255 24172 31276 24212
rect 31316 24172 31337 24212
rect 31423 24172 31440 24212
rect 31480 24172 31489 24212
rect 31103 24149 31169 24172
rect 31255 24149 31337 24172
rect 31423 24149 31489 24172
rect 31103 24130 31489 24149
rect 35103 24235 35489 24254
rect 35103 24212 35169 24235
rect 35255 24212 35337 24235
rect 35423 24212 35489 24235
rect 35103 24172 35112 24212
rect 35152 24172 35169 24212
rect 35255 24172 35276 24212
rect 35316 24172 35337 24212
rect 35423 24172 35440 24212
rect 35480 24172 35489 24212
rect 35103 24149 35169 24172
rect 35255 24149 35337 24172
rect 35423 24149 35489 24172
rect 35103 24130 35489 24149
rect 39103 24235 39489 24254
rect 39103 24212 39169 24235
rect 39255 24212 39337 24235
rect 39423 24212 39489 24235
rect 39103 24172 39112 24212
rect 39152 24172 39169 24212
rect 39255 24172 39276 24212
rect 39316 24172 39337 24212
rect 39423 24172 39440 24212
rect 39480 24172 39489 24212
rect 39103 24149 39169 24172
rect 39255 24149 39337 24172
rect 39423 24149 39489 24172
rect 39103 24130 39489 24149
rect 43103 24235 43489 24254
rect 43103 24212 43169 24235
rect 43255 24212 43337 24235
rect 43423 24212 43489 24235
rect 43103 24172 43112 24212
rect 43152 24172 43169 24212
rect 43255 24172 43276 24212
rect 43316 24172 43337 24212
rect 43423 24172 43440 24212
rect 43480 24172 43489 24212
rect 43103 24149 43169 24172
rect 43255 24149 43337 24172
rect 43423 24149 43489 24172
rect 43103 24130 43489 24149
rect 47103 24235 47489 24254
rect 47103 24212 47169 24235
rect 47255 24212 47337 24235
rect 47423 24212 47489 24235
rect 47103 24172 47112 24212
rect 47152 24172 47169 24212
rect 47255 24172 47276 24212
rect 47316 24172 47337 24212
rect 47423 24172 47440 24212
rect 47480 24172 47489 24212
rect 47103 24149 47169 24172
rect 47255 24149 47337 24172
rect 47423 24149 47489 24172
rect 47103 24130 47489 24149
rect 51103 24235 51489 24254
rect 51103 24212 51169 24235
rect 51255 24212 51337 24235
rect 51423 24212 51489 24235
rect 51103 24172 51112 24212
rect 51152 24172 51169 24212
rect 51255 24172 51276 24212
rect 51316 24172 51337 24212
rect 51423 24172 51440 24212
rect 51480 24172 51489 24212
rect 51103 24149 51169 24172
rect 51255 24149 51337 24172
rect 51423 24149 51489 24172
rect 51103 24130 51489 24149
rect 55103 24235 55489 24254
rect 55103 24212 55169 24235
rect 55255 24212 55337 24235
rect 55423 24212 55489 24235
rect 55103 24172 55112 24212
rect 55152 24172 55169 24212
rect 55255 24172 55276 24212
rect 55316 24172 55337 24212
rect 55423 24172 55440 24212
rect 55480 24172 55489 24212
rect 55103 24149 55169 24172
rect 55255 24149 55337 24172
rect 55423 24149 55489 24172
rect 55103 24130 55489 24149
rect 59103 24235 59489 24254
rect 59103 24212 59169 24235
rect 59255 24212 59337 24235
rect 59423 24212 59489 24235
rect 59103 24172 59112 24212
rect 59152 24172 59169 24212
rect 59255 24172 59276 24212
rect 59316 24172 59337 24212
rect 59423 24172 59440 24212
rect 59480 24172 59489 24212
rect 59103 24149 59169 24172
rect 59255 24149 59337 24172
rect 59423 24149 59489 24172
rect 59103 24130 59489 24149
rect 63103 24235 63489 24254
rect 63103 24212 63169 24235
rect 63255 24212 63337 24235
rect 63423 24212 63489 24235
rect 63103 24172 63112 24212
rect 63152 24172 63169 24212
rect 63255 24172 63276 24212
rect 63316 24172 63337 24212
rect 63423 24172 63440 24212
rect 63480 24172 63489 24212
rect 63103 24149 63169 24172
rect 63255 24149 63337 24172
rect 63423 24149 63489 24172
rect 63103 24130 63489 24149
rect 67103 24235 67489 24254
rect 67103 24212 67169 24235
rect 67255 24212 67337 24235
rect 67423 24212 67489 24235
rect 67103 24172 67112 24212
rect 67152 24172 67169 24212
rect 67255 24172 67276 24212
rect 67316 24172 67337 24212
rect 67423 24172 67440 24212
rect 67480 24172 67489 24212
rect 67103 24149 67169 24172
rect 67255 24149 67337 24172
rect 67423 24149 67489 24172
rect 67103 24130 67489 24149
rect 4343 23479 4729 23498
rect 4343 23456 4409 23479
rect 4495 23456 4577 23479
rect 4663 23456 4729 23479
rect 4343 23416 4352 23456
rect 4392 23416 4409 23456
rect 4495 23416 4516 23456
rect 4556 23416 4577 23456
rect 4663 23416 4680 23456
rect 4720 23416 4729 23456
rect 4343 23393 4409 23416
rect 4495 23393 4577 23416
rect 4663 23393 4729 23416
rect 4343 23374 4729 23393
rect 8343 23479 8729 23498
rect 8343 23456 8409 23479
rect 8495 23456 8577 23479
rect 8663 23456 8729 23479
rect 8343 23416 8352 23456
rect 8392 23416 8409 23456
rect 8495 23416 8516 23456
rect 8556 23416 8577 23456
rect 8663 23416 8680 23456
rect 8720 23416 8729 23456
rect 8343 23393 8409 23416
rect 8495 23393 8577 23416
rect 8663 23393 8729 23416
rect 8343 23374 8729 23393
rect 12343 23479 12729 23498
rect 12343 23456 12409 23479
rect 12495 23456 12577 23479
rect 12663 23456 12729 23479
rect 12343 23416 12352 23456
rect 12392 23416 12409 23456
rect 12495 23416 12516 23456
rect 12556 23416 12577 23456
rect 12663 23416 12680 23456
rect 12720 23416 12729 23456
rect 12343 23393 12409 23416
rect 12495 23393 12577 23416
rect 12663 23393 12729 23416
rect 12343 23374 12729 23393
rect 16343 23479 16729 23498
rect 16343 23456 16409 23479
rect 16495 23456 16577 23479
rect 16663 23456 16729 23479
rect 16343 23416 16352 23456
rect 16392 23416 16409 23456
rect 16495 23416 16516 23456
rect 16556 23416 16577 23456
rect 16663 23416 16680 23456
rect 16720 23416 16729 23456
rect 16343 23393 16409 23416
rect 16495 23393 16577 23416
rect 16663 23393 16729 23416
rect 16343 23374 16729 23393
rect 20343 23479 20729 23498
rect 20343 23456 20409 23479
rect 20495 23456 20577 23479
rect 20663 23456 20729 23479
rect 20343 23416 20352 23456
rect 20392 23416 20409 23456
rect 20495 23416 20516 23456
rect 20556 23416 20577 23456
rect 20663 23416 20680 23456
rect 20720 23416 20729 23456
rect 20343 23393 20409 23416
rect 20495 23393 20577 23416
rect 20663 23393 20729 23416
rect 20343 23374 20729 23393
rect 24343 23479 24729 23498
rect 24343 23456 24409 23479
rect 24495 23456 24577 23479
rect 24663 23456 24729 23479
rect 24343 23416 24352 23456
rect 24392 23416 24409 23456
rect 24495 23416 24516 23456
rect 24556 23416 24577 23456
rect 24663 23416 24680 23456
rect 24720 23416 24729 23456
rect 24343 23393 24409 23416
rect 24495 23393 24577 23416
rect 24663 23393 24729 23416
rect 24343 23374 24729 23393
rect 28343 23479 28729 23498
rect 28343 23456 28409 23479
rect 28495 23456 28577 23479
rect 28663 23456 28729 23479
rect 28343 23416 28352 23456
rect 28392 23416 28409 23456
rect 28495 23416 28516 23456
rect 28556 23416 28577 23456
rect 28663 23416 28680 23456
rect 28720 23416 28729 23456
rect 28343 23393 28409 23416
rect 28495 23393 28577 23416
rect 28663 23393 28729 23416
rect 28343 23374 28729 23393
rect 32343 23479 32729 23498
rect 32343 23456 32409 23479
rect 32495 23456 32577 23479
rect 32663 23456 32729 23479
rect 32343 23416 32352 23456
rect 32392 23416 32409 23456
rect 32495 23416 32516 23456
rect 32556 23416 32577 23456
rect 32663 23416 32680 23456
rect 32720 23416 32729 23456
rect 32343 23393 32409 23416
rect 32495 23393 32577 23416
rect 32663 23393 32729 23416
rect 32343 23374 32729 23393
rect 36343 23479 36729 23498
rect 36343 23456 36409 23479
rect 36495 23456 36577 23479
rect 36663 23456 36729 23479
rect 36343 23416 36352 23456
rect 36392 23416 36409 23456
rect 36495 23416 36516 23456
rect 36556 23416 36577 23456
rect 36663 23416 36680 23456
rect 36720 23416 36729 23456
rect 36343 23393 36409 23416
rect 36495 23393 36577 23416
rect 36663 23393 36729 23416
rect 36343 23374 36729 23393
rect 40343 23479 40729 23498
rect 40343 23456 40409 23479
rect 40495 23456 40577 23479
rect 40663 23456 40729 23479
rect 40343 23416 40352 23456
rect 40392 23416 40409 23456
rect 40495 23416 40516 23456
rect 40556 23416 40577 23456
rect 40663 23416 40680 23456
rect 40720 23416 40729 23456
rect 40343 23393 40409 23416
rect 40495 23393 40577 23416
rect 40663 23393 40729 23416
rect 40343 23374 40729 23393
rect 44343 23479 44729 23498
rect 44343 23456 44409 23479
rect 44495 23456 44577 23479
rect 44663 23456 44729 23479
rect 44343 23416 44352 23456
rect 44392 23416 44409 23456
rect 44495 23416 44516 23456
rect 44556 23416 44577 23456
rect 44663 23416 44680 23456
rect 44720 23416 44729 23456
rect 44343 23393 44409 23416
rect 44495 23393 44577 23416
rect 44663 23393 44729 23416
rect 44343 23374 44729 23393
rect 48343 23479 48729 23498
rect 48343 23456 48409 23479
rect 48495 23456 48577 23479
rect 48663 23456 48729 23479
rect 48343 23416 48352 23456
rect 48392 23416 48409 23456
rect 48495 23416 48516 23456
rect 48556 23416 48577 23456
rect 48663 23416 48680 23456
rect 48720 23416 48729 23456
rect 48343 23393 48409 23416
rect 48495 23393 48577 23416
rect 48663 23393 48729 23416
rect 48343 23374 48729 23393
rect 52343 23479 52729 23498
rect 52343 23456 52409 23479
rect 52495 23456 52577 23479
rect 52663 23456 52729 23479
rect 52343 23416 52352 23456
rect 52392 23416 52409 23456
rect 52495 23416 52516 23456
rect 52556 23416 52577 23456
rect 52663 23416 52680 23456
rect 52720 23416 52729 23456
rect 52343 23393 52409 23416
rect 52495 23393 52577 23416
rect 52663 23393 52729 23416
rect 52343 23374 52729 23393
rect 56343 23479 56729 23498
rect 56343 23456 56409 23479
rect 56495 23456 56577 23479
rect 56663 23456 56729 23479
rect 56343 23416 56352 23456
rect 56392 23416 56409 23456
rect 56495 23416 56516 23456
rect 56556 23416 56577 23456
rect 56663 23416 56680 23456
rect 56720 23416 56729 23456
rect 56343 23393 56409 23416
rect 56495 23393 56577 23416
rect 56663 23393 56729 23416
rect 56343 23374 56729 23393
rect 60343 23479 60729 23498
rect 60343 23456 60409 23479
rect 60495 23456 60577 23479
rect 60663 23456 60729 23479
rect 60343 23416 60352 23456
rect 60392 23416 60409 23456
rect 60495 23416 60516 23456
rect 60556 23416 60577 23456
rect 60663 23416 60680 23456
rect 60720 23416 60729 23456
rect 60343 23393 60409 23416
rect 60495 23393 60577 23416
rect 60663 23393 60729 23416
rect 60343 23374 60729 23393
rect 64343 23479 64729 23498
rect 64343 23456 64409 23479
rect 64495 23456 64577 23479
rect 64663 23456 64729 23479
rect 64343 23416 64352 23456
rect 64392 23416 64409 23456
rect 64495 23416 64516 23456
rect 64556 23416 64577 23456
rect 64663 23416 64680 23456
rect 64720 23416 64729 23456
rect 64343 23393 64409 23416
rect 64495 23393 64577 23416
rect 64663 23393 64729 23416
rect 64343 23374 64729 23393
rect 68343 23479 68729 23498
rect 68343 23456 68409 23479
rect 68495 23456 68577 23479
rect 68663 23456 68729 23479
rect 68343 23416 68352 23456
rect 68392 23416 68409 23456
rect 68495 23416 68516 23456
rect 68556 23416 68577 23456
rect 68663 23416 68680 23456
rect 68720 23416 68729 23456
rect 68343 23393 68409 23416
rect 68495 23393 68577 23416
rect 68663 23393 68729 23416
rect 68343 23374 68729 23393
rect 72343 23479 72729 23498
rect 72343 23456 72409 23479
rect 72495 23456 72577 23479
rect 72663 23456 72729 23479
rect 72343 23416 72352 23456
rect 72392 23416 72409 23456
rect 72495 23416 72516 23456
rect 72556 23416 72577 23456
rect 72663 23416 72680 23456
rect 72720 23416 72729 23456
rect 72343 23393 72409 23416
rect 72495 23393 72577 23416
rect 72663 23393 72729 23416
rect 72343 23374 72729 23393
rect 76343 23479 76729 23498
rect 76343 23456 76409 23479
rect 76495 23456 76577 23479
rect 76663 23456 76729 23479
rect 76343 23416 76352 23456
rect 76392 23416 76409 23456
rect 76495 23416 76516 23456
rect 76556 23416 76577 23456
rect 76663 23416 76680 23456
rect 76720 23416 76729 23456
rect 76343 23393 76409 23416
rect 76495 23393 76577 23416
rect 76663 23393 76729 23416
rect 76343 23374 76729 23393
rect 80343 23479 80729 23498
rect 80343 23456 80409 23479
rect 80495 23456 80577 23479
rect 80663 23456 80729 23479
rect 80343 23416 80352 23456
rect 80392 23416 80409 23456
rect 80495 23416 80516 23456
rect 80556 23416 80577 23456
rect 80663 23416 80680 23456
rect 80720 23416 80729 23456
rect 80343 23393 80409 23416
rect 80495 23393 80577 23416
rect 80663 23393 80729 23416
rect 80343 23374 80729 23393
rect 84343 23479 84729 23498
rect 84343 23456 84409 23479
rect 84495 23456 84577 23479
rect 84663 23456 84729 23479
rect 84343 23416 84352 23456
rect 84392 23416 84409 23456
rect 84495 23416 84516 23456
rect 84556 23416 84577 23456
rect 84663 23416 84680 23456
rect 84720 23416 84729 23456
rect 84343 23393 84409 23416
rect 84495 23393 84577 23416
rect 84663 23393 84729 23416
rect 84343 23374 84729 23393
rect 88343 23479 88729 23498
rect 88343 23456 88409 23479
rect 88495 23456 88577 23479
rect 88663 23456 88729 23479
rect 88343 23416 88352 23456
rect 88392 23416 88409 23456
rect 88495 23416 88516 23456
rect 88556 23416 88577 23456
rect 88663 23416 88680 23456
rect 88720 23416 88729 23456
rect 88343 23393 88409 23416
rect 88495 23393 88577 23416
rect 88663 23393 88729 23416
rect 88343 23374 88729 23393
rect 92343 23479 92729 23498
rect 92343 23456 92409 23479
rect 92495 23456 92577 23479
rect 92663 23456 92729 23479
rect 92343 23416 92352 23456
rect 92392 23416 92409 23456
rect 92495 23416 92516 23456
rect 92556 23416 92577 23456
rect 92663 23416 92680 23456
rect 92720 23416 92729 23456
rect 92343 23393 92409 23416
rect 92495 23393 92577 23416
rect 92663 23393 92729 23416
rect 92343 23374 92729 23393
rect 96343 23479 96729 23498
rect 96343 23456 96409 23479
rect 96495 23456 96577 23479
rect 96663 23456 96729 23479
rect 96343 23416 96352 23456
rect 96392 23416 96409 23456
rect 96495 23416 96516 23456
rect 96556 23416 96577 23456
rect 96663 23416 96680 23456
rect 96720 23416 96729 23456
rect 96343 23393 96409 23416
rect 96495 23393 96577 23416
rect 96663 23393 96729 23416
rect 96343 23374 96729 23393
rect 86450 23143 86574 23162
rect 86450 23057 86469 23143
rect 86555 23120 86574 23143
rect 86555 23080 86668 23120
rect 86708 23080 86717 23120
rect 86555 23057 86574 23080
rect 86450 23038 86574 23057
rect 3103 22723 3489 22742
rect 3103 22700 3169 22723
rect 3255 22700 3337 22723
rect 3423 22700 3489 22723
rect 3103 22660 3112 22700
rect 3152 22660 3169 22700
rect 3255 22660 3276 22700
rect 3316 22660 3337 22700
rect 3423 22660 3440 22700
rect 3480 22660 3489 22700
rect 3103 22637 3169 22660
rect 3255 22637 3337 22660
rect 3423 22637 3489 22660
rect 3103 22618 3489 22637
rect 7103 22723 7489 22742
rect 7103 22700 7169 22723
rect 7255 22700 7337 22723
rect 7423 22700 7489 22723
rect 7103 22660 7112 22700
rect 7152 22660 7169 22700
rect 7255 22660 7276 22700
rect 7316 22660 7337 22700
rect 7423 22660 7440 22700
rect 7480 22660 7489 22700
rect 7103 22637 7169 22660
rect 7255 22637 7337 22660
rect 7423 22637 7489 22660
rect 7103 22618 7489 22637
rect 11103 22723 11489 22742
rect 11103 22700 11169 22723
rect 11255 22700 11337 22723
rect 11423 22700 11489 22723
rect 11103 22660 11112 22700
rect 11152 22660 11169 22700
rect 11255 22660 11276 22700
rect 11316 22660 11337 22700
rect 11423 22660 11440 22700
rect 11480 22660 11489 22700
rect 11103 22637 11169 22660
rect 11255 22637 11337 22660
rect 11423 22637 11489 22660
rect 11103 22618 11489 22637
rect 15103 22723 15489 22742
rect 15103 22700 15169 22723
rect 15255 22700 15337 22723
rect 15423 22700 15489 22723
rect 15103 22660 15112 22700
rect 15152 22660 15169 22700
rect 15255 22660 15276 22700
rect 15316 22660 15337 22700
rect 15423 22660 15440 22700
rect 15480 22660 15489 22700
rect 15103 22637 15169 22660
rect 15255 22637 15337 22660
rect 15423 22637 15489 22660
rect 15103 22618 15489 22637
rect 19103 22723 19489 22742
rect 19103 22700 19169 22723
rect 19255 22700 19337 22723
rect 19423 22700 19489 22723
rect 19103 22660 19112 22700
rect 19152 22660 19169 22700
rect 19255 22660 19276 22700
rect 19316 22660 19337 22700
rect 19423 22660 19440 22700
rect 19480 22660 19489 22700
rect 19103 22637 19169 22660
rect 19255 22637 19337 22660
rect 19423 22637 19489 22660
rect 19103 22618 19489 22637
rect 23103 22723 23489 22742
rect 23103 22700 23169 22723
rect 23255 22700 23337 22723
rect 23423 22700 23489 22723
rect 23103 22660 23112 22700
rect 23152 22660 23169 22700
rect 23255 22660 23276 22700
rect 23316 22660 23337 22700
rect 23423 22660 23440 22700
rect 23480 22660 23489 22700
rect 23103 22637 23169 22660
rect 23255 22637 23337 22660
rect 23423 22637 23489 22660
rect 23103 22618 23489 22637
rect 27103 22723 27489 22742
rect 27103 22700 27169 22723
rect 27255 22700 27337 22723
rect 27423 22700 27489 22723
rect 27103 22660 27112 22700
rect 27152 22660 27169 22700
rect 27255 22660 27276 22700
rect 27316 22660 27337 22700
rect 27423 22660 27440 22700
rect 27480 22660 27489 22700
rect 27103 22637 27169 22660
rect 27255 22637 27337 22660
rect 27423 22637 27489 22660
rect 27103 22618 27489 22637
rect 31103 22723 31489 22742
rect 31103 22700 31169 22723
rect 31255 22700 31337 22723
rect 31423 22700 31489 22723
rect 31103 22660 31112 22700
rect 31152 22660 31169 22700
rect 31255 22660 31276 22700
rect 31316 22660 31337 22700
rect 31423 22660 31440 22700
rect 31480 22660 31489 22700
rect 31103 22637 31169 22660
rect 31255 22637 31337 22660
rect 31423 22637 31489 22660
rect 31103 22618 31489 22637
rect 35103 22723 35489 22742
rect 35103 22700 35169 22723
rect 35255 22700 35337 22723
rect 35423 22700 35489 22723
rect 35103 22660 35112 22700
rect 35152 22660 35169 22700
rect 35255 22660 35276 22700
rect 35316 22660 35337 22700
rect 35423 22660 35440 22700
rect 35480 22660 35489 22700
rect 35103 22637 35169 22660
rect 35255 22637 35337 22660
rect 35423 22637 35489 22660
rect 35103 22618 35489 22637
rect 39103 22723 39489 22742
rect 39103 22700 39169 22723
rect 39255 22700 39337 22723
rect 39423 22700 39489 22723
rect 39103 22660 39112 22700
rect 39152 22660 39169 22700
rect 39255 22660 39276 22700
rect 39316 22660 39337 22700
rect 39423 22660 39440 22700
rect 39480 22660 39489 22700
rect 39103 22637 39169 22660
rect 39255 22637 39337 22660
rect 39423 22637 39489 22660
rect 39103 22618 39489 22637
rect 43103 22723 43489 22742
rect 43103 22700 43169 22723
rect 43255 22700 43337 22723
rect 43423 22700 43489 22723
rect 43103 22660 43112 22700
rect 43152 22660 43169 22700
rect 43255 22660 43276 22700
rect 43316 22660 43337 22700
rect 43423 22660 43440 22700
rect 43480 22660 43489 22700
rect 43103 22637 43169 22660
rect 43255 22637 43337 22660
rect 43423 22637 43489 22660
rect 43103 22618 43489 22637
rect 47103 22723 47489 22742
rect 47103 22700 47169 22723
rect 47255 22700 47337 22723
rect 47423 22700 47489 22723
rect 47103 22660 47112 22700
rect 47152 22660 47169 22700
rect 47255 22660 47276 22700
rect 47316 22660 47337 22700
rect 47423 22660 47440 22700
rect 47480 22660 47489 22700
rect 47103 22637 47169 22660
rect 47255 22637 47337 22660
rect 47423 22637 47489 22660
rect 47103 22618 47489 22637
rect 51103 22723 51489 22742
rect 51103 22700 51169 22723
rect 51255 22700 51337 22723
rect 51423 22700 51489 22723
rect 51103 22660 51112 22700
rect 51152 22660 51169 22700
rect 51255 22660 51276 22700
rect 51316 22660 51337 22700
rect 51423 22660 51440 22700
rect 51480 22660 51489 22700
rect 51103 22637 51169 22660
rect 51255 22637 51337 22660
rect 51423 22637 51489 22660
rect 51103 22618 51489 22637
rect 55103 22723 55489 22742
rect 55103 22700 55169 22723
rect 55255 22700 55337 22723
rect 55423 22700 55489 22723
rect 55103 22660 55112 22700
rect 55152 22660 55169 22700
rect 55255 22660 55276 22700
rect 55316 22660 55337 22700
rect 55423 22660 55440 22700
rect 55480 22660 55489 22700
rect 55103 22637 55169 22660
rect 55255 22637 55337 22660
rect 55423 22637 55489 22660
rect 55103 22618 55489 22637
rect 59103 22723 59489 22742
rect 59103 22700 59169 22723
rect 59255 22700 59337 22723
rect 59423 22700 59489 22723
rect 59103 22660 59112 22700
rect 59152 22660 59169 22700
rect 59255 22660 59276 22700
rect 59316 22660 59337 22700
rect 59423 22660 59440 22700
rect 59480 22660 59489 22700
rect 59103 22637 59169 22660
rect 59255 22637 59337 22660
rect 59423 22637 59489 22660
rect 59103 22618 59489 22637
rect 63103 22723 63489 22742
rect 63103 22700 63169 22723
rect 63255 22700 63337 22723
rect 63423 22700 63489 22723
rect 63103 22660 63112 22700
rect 63152 22660 63169 22700
rect 63255 22660 63276 22700
rect 63316 22660 63337 22700
rect 63423 22660 63440 22700
rect 63480 22660 63489 22700
rect 63103 22637 63169 22660
rect 63255 22637 63337 22660
rect 63423 22637 63489 22660
rect 63103 22618 63489 22637
rect 67103 22723 67489 22742
rect 67103 22700 67169 22723
rect 67255 22700 67337 22723
rect 67423 22700 67489 22723
rect 67103 22660 67112 22700
rect 67152 22660 67169 22700
rect 67255 22660 67276 22700
rect 67316 22660 67337 22700
rect 67423 22660 67440 22700
rect 67480 22660 67489 22700
rect 67103 22637 67169 22660
rect 67255 22637 67337 22660
rect 67423 22637 67489 22660
rect 67103 22618 67489 22637
rect 71103 22723 71489 22742
rect 71103 22700 71169 22723
rect 71255 22700 71337 22723
rect 71423 22700 71489 22723
rect 71103 22660 71112 22700
rect 71152 22660 71169 22700
rect 71255 22660 71276 22700
rect 71316 22660 71337 22700
rect 71423 22660 71440 22700
rect 71480 22660 71489 22700
rect 71103 22637 71169 22660
rect 71255 22637 71337 22660
rect 71423 22637 71489 22660
rect 71103 22618 71489 22637
rect 75103 22723 75489 22742
rect 75103 22700 75169 22723
rect 75255 22700 75337 22723
rect 75423 22700 75489 22723
rect 75103 22660 75112 22700
rect 75152 22660 75169 22700
rect 75255 22660 75276 22700
rect 75316 22660 75337 22700
rect 75423 22660 75440 22700
rect 75480 22660 75489 22700
rect 75103 22637 75169 22660
rect 75255 22637 75337 22660
rect 75423 22637 75489 22660
rect 75103 22618 75489 22637
rect 79103 22723 79489 22742
rect 79103 22700 79169 22723
rect 79255 22700 79337 22723
rect 79423 22700 79489 22723
rect 79103 22660 79112 22700
rect 79152 22660 79169 22700
rect 79255 22660 79276 22700
rect 79316 22660 79337 22700
rect 79423 22660 79440 22700
rect 79480 22660 79489 22700
rect 79103 22637 79169 22660
rect 79255 22637 79337 22660
rect 79423 22637 79489 22660
rect 79103 22618 79489 22637
rect 83103 22723 83489 22742
rect 83103 22700 83169 22723
rect 83255 22700 83337 22723
rect 83423 22700 83489 22723
rect 83103 22660 83112 22700
rect 83152 22660 83169 22700
rect 83255 22660 83276 22700
rect 83316 22660 83337 22700
rect 83423 22660 83440 22700
rect 83480 22660 83489 22700
rect 83103 22637 83169 22660
rect 83255 22637 83337 22660
rect 83423 22637 83489 22660
rect 83103 22618 83489 22637
rect 87103 22723 87489 22742
rect 87103 22700 87169 22723
rect 87255 22700 87337 22723
rect 87423 22700 87489 22723
rect 87103 22660 87112 22700
rect 87152 22660 87169 22700
rect 87255 22660 87276 22700
rect 87316 22660 87337 22700
rect 87423 22660 87440 22700
rect 87480 22660 87489 22700
rect 87103 22637 87169 22660
rect 87255 22637 87337 22660
rect 87423 22637 87489 22660
rect 87103 22618 87489 22637
rect 91103 22723 91489 22742
rect 91103 22700 91169 22723
rect 91255 22700 91337 22723
rect 91423 22700 91489 22723
rect 91103 22660 91112 22700
rect 91152 22660 91169 22700
rect 91255 22660 91276 22700
rect 91316 22660 91337 22700
rect 91423 22660 91440 22700
rect 91480 22660 91489 22700
rect 91103 22637 91169 22660
rect 91255 22637 91337 22660
rect 91423 22637 91489 22660
rect 91103 22618 91489 22637
rect 95103 22723 95489 22742
rect 95103 22700 95169 22723
rect 95255 22700 95337 22723
rect 95423 22700 95489 22723
rect 95103 22660 95112 22700
rect 95152 22660 95169 22700
rect 95255 22660 95276 22700
rect 95316 22660 95337 22700
rect 95423 22660 95440 22700
rect 95480 22660 95489 22700
rect 95103 22637 95169 22660
rect 95255 22637 95337 22660
rect 95423 22637 95489 22660
rect 95103 22618 95489 22637
rect 99103 22723 99489 22742
rect 99103 22700 99169 22723
rect 99255 22700 99337 22723
rect 99423 22700 99489 22723
rect 99103 22660 99112 22700
rect 99152 22660 99169 22700
rect 99255 22660 99276 22700
rect 99316 22660 99337 22700
rect 99423 22660 99440 22700
rect 99480 22660 99489 22700
rect 99103 22637 99169 22660
rect 99255 22637 99337 22660
rect 99423 22637 99489 22660
rect 99103 22618 99489 22637
rect 4343 21967 4729 21986
rect 4343 21944 4409 21967
rect 4495 21944 4577 21967
rect 4663 21944 4729 21967
rect 4343 21904 4352 21944
rect 4392 21904 4409 21944
rect 4495 21904 4516 21944
rect 4556 21904 4577 21944
rect 4663 21904 4680 21944
rect 4720 21904 4729 21944
rect 4343 21881 4409 21904
rect 4495 21881 4577 21904
rect 4663 21881 4729 21904
rect 4343 21862 4729 21881
rect 8343 21967 8729 21986
rect 8343 21944 8409 21967
rect 8495 21944 8577 21967
rect 8663 21944 8729 21967
rect 8343 21904 8352 21944
rect 8392 21904 8409 21944
rect 8495 21904 8516 21944
rect 8556 21904 8577 21944
rect 8663 21904 8680 21944
rect 8720 21904 8729 21944
rect 8343 21881 8409 21904
rect 8495 21881 8577 21904
rect 8663 21881 8729 21904
rect 8343 21862 8729 21881
rect 12343 21967 12729 21986
rect 12343 21944 12409 21967
rect 12495 21944 12577 21967
rect 12663 21944 12729 21967
rect 12343 21904 12352 21944
rect 12392 21904 12409 21944
rect 12495 21904 12516 21944
rect 12556 21904 12577 21944
rect 12663 21904 12680 21944
rect 12720 21904 12729 21944
rect 12343 21881 12409 21904
rect 12495 21881 12577 21904
rect 12663 21881 12729 21904
rect 12343 21862 12729 21881
rect 16343 21967 16729 21986
rect 16343 21944 16409 21967
rect 16495 21944 16577 21967
rect 16663 21944 16729 21967
rect 16343 21904 16352 21944
rect 16392 21904 16409 21944
rect 16495 21904 16516 21944
rect 16556 21904 16577 21944
rect 16663 21904 16680 21944
rect 16720 21904 16729 21944
rect 16343 21881 16409 21904
rect 16495 21881 16577 21904
rect 16663 21881 16729 21904
rect 16343 21862 16729 21881
rect 20343 21967 20729 21986
rect 20343 21944 20409 21967
rect 20495 21944 20577 21967
rect 20663 21944 20729 21967
rect 20343 21904 20352 21944
rect 20392 21904 20409 21944
rect 20495 21904 20516 21944
rect 20556 21904 20577 21944
rect 20663 21904 20680 21944
rect 20720 21904 20729 21944
rect 20343 21881 20409 21904
rect 20495 21881 20577 21904
rect 20663 21881 20729 21904
rect 20343 21862 20729 21881
rect 24343 21967 24729 21986
rect 24343 21944 24409 21967
rect 24495 21944 24577 21967
rect 24663 21944 24729 21967
rect 24343 21904 24352 21944
rect 24392 21904 24409 21944
rect 24495 21904 24516 21944
rect 24556 21904 24577 21944
rect 24663 21904 24680 21944
rect 24720 21904 24729 21944
rect 24343 21881 24409 21904
rect 24495 21881 24577 21904
rect 24663 21881 24729 21904
rect 24343 21862 24729 21881
rect 28343 21967 28729 21986
rect 28343 21944 28409 21967
rect 28495 21944 28577 21967
rect 28663 21944 28729 21967
rect 28343 21904 28352 21944
rect 28392 21904 28409 21944
rect 28495 21904 28516 21944
rect 28556 21904 28577 21944
rect 28663 21904 28680 21944
rect 28720 21904 28729 21944
rect 28343 21881 28409 21904
rect 28495 21881 28577 21904
rect 28663 21881 28729 21904
rect 28343 21862 28729 21881
rect 32343 21967 32729 21986
rect 32343 21944 32409 21967
rect 32495 21944 32577 21967
rect 32663 21944 32729 21967
rect 32343 21904 32352 21944
rect 32392 21904 32409 21944
rect 32495 21904 32516 21944
rect 32556 21904 32577 21944
rect 32663 21904 32680 21944
rect 32720 21904 32729 21944
rect 32343 21881 32409 21904
rect 32495 21881 32577 21904
rect 32663 21881 32729 21904
rect 32343 21862 32729 21881
rect 36343 21967 36729 21986
rect 36343 21944 36409 21967
rect 36495 21944 36577 21967
rect 36663 21944 36729 21967
rect 36343 21904 36352 21944
rect 36392 21904 36409 21944
rect 36495 21904 36516 21944
rect 36556 21904 36577 21944
rect 36663 21904 36680 21944
rect 36720 21904 36729 21944
rect 36343 21881 36409 21904
rect 36495 21881 36577 21904
rect 36663 21881 36729 21904
rect 36343 21862 36729 21881
rect 40343 21967 40729 21986
rect 40343 21944 40409 21967
rect 40495 21944 40577 21967
rect 40663 21944 40729 21967
rect 40343 21904 40352 21944
rect 40392 21904 40409 21944
rect 40495 21904 40516 21944
rect 40556 21904 40577 21944
rect 40663 21904 40680 21944
rect 40720 21904 40729 21944
rect 40343 21881 40409 21904
rect 40495 21881 40577 21904
rect 40663 21881 40729 21904
rect 40343 21862 40729 21881
rect 44343 21967 44729 21986
rect 44343 21944 44409 21967
rect 44495 21944 44577 21967
rect 44663 21944 44729 21967
rect 44343 21904 44352 21944
rect 44392 21904 44409 21944
rect 44495 21904 44516 21944
rect 44556 21904 44577 21944
rect 44663 21904 44680 21944
rect 44720 21904 44729 21944
rect 44343 21881 44409 21904
rect 44495 21881 44577 21904
rect 44663 21881 44729 21904
rect 44343 21862 44729 21881
rect 48343 21967 48729 21986
rect 48343 21944 48409 21967
rect 48495 21944 48577 21967
rect 48663 21944 48729 21967
rect 48343 21904 48352 21944
rect 48392 21904 48409 21944
rect 48495 21904 48516 21944
rect 48556 21904 48577 21944
rect 48663 21904 48680 21944
rect 48720 21904 48729 21944
rect 48343 21881 48409 21904
rect 48495 21881 48577 21904
rect 48663 21881 48729 21904
rect 48343 21862 48729 21881
rect 52343 21967 52729 21986
rect 52343 21944 52409 21967
rect 52495 21944 52577 21967
rect 52663 21944 52729 21967
rect 52343 21904 52352 21944
rect 52392 21904 52409 21944
rect 52495 21904 52516 21944
rect 52556 21904 52577 21944
rect 52663 21904 52680 21944
rect 52720 21904 52729 21944
rect 52343 21881 52409 21904
rect 52495 21881 52577 21904
rect 52663 21881 52729 21904
rect 52343 21862 52729 21881
rect 56343 21967 56729 21986
rect 56343 21944 56409 21967
rect 56495 21944 56577 21967
rect 56663 21944 56729 21967
rect 56343 21904 56352 21944
rect 56392 21904 56409 21944
rect 56495 21904 56516 21944
rect 56556 21904 56577 21944
rect 56663 21904 56680 21944
rect 56720 21904 56729 21944
rect 56343 21881 56409 21904
rect 56495 21881 56577 21904
rect 56663 21881 56729 21904
rect 56343 21862 56729 21881
rect 60343 21967 60729 21986
rect 60343 21944 60409 21967
rect 60495 21944 60577 21967
rect 60663 21944 60729 21967
rect 60343 21904 60352 21944
rect 60392 21904 60409 21944
rect 60495 21904 60516 21944
rect 60556 21904 60577 21944
rect 60663 21904 60680 21944
rect 60720 21904 60729 21944
rect 60343 21881 60409 21904
rect 60495 21881 60577 21904
rect 60663 21881 60729 21904
rect 60343 21862 60729 21881
rect 64343 21967 64729 21986
rect 64343 21944 64409 21967
rect 64495 21944 64577 21967
rect 64663 21944 64729 21967
rect 64343 21904 64352 21944
rect 64392 21904 64409 21944
rect 64495 21904 64516 21944
rect 64556 21904 64577 21944
rect 64663 21904 64680 21944
rect 64720 21904 64729 21944
rect 64343 21881 64409 21904
rect 64495 21881 64577 21904
rect 64663 21881 64729 21904
rect 64343 21862 64729 21881
rect 68343 21967 68729 21986
rect 68343 21944 68409 21967
rect 68495 21944 68577 21967
rect 68663 21944 68729 21967
rect 68343 21904 68352 21944
rect 68392 21904 68409 21944
rect 68495 21904 68516 21944
rect 68556 21904 68577 21944
rect 68663 21904 68680 21944
rect 68720 21904 68729 21944
rect 68343 21881 68409 21904
rect 68495 21881 68577 21904
rect 68663 21881 68729 21904
rect 68343 21862 68729 21881
rect 72343 21967 72729 21986
rect 72343 21944 72409 21967
rect 72495 21944 72577 21967
rect 72663 21944 72729 21967
rect 72343 21904 72352 21944
rect 72392 21904 72409 21944
rect 72495 21904 72516 21944
rect 72556 21904 72577 21944
rect 72663 21904 72680 21944
rect 72720 21904 72729 21944
rect 72343 21881 72409 21904
rect 72495 21881 72577 21904
rect 72663 21881 72729 21904
rect 72343 21862 72729 21881
rect 76343 21967 76729 21986
rect 76343 21944 76409 21967
rect 76495 21944 76577 21967
rect 76663 21944 76729 21967
rect 76343 21904 76352 21944
rect 76392 21904 76409 21944
rect 76495 21904 76516 21944
rect 76556 21904 76577 21944
rect 76663 21904 76680 21944
rect 76720 21904 76729 21944
rect 76343 21881 76409 21904
rect 76495 21881 76577 21904
rect 76663 21881 76729 21904
rect 76343 21862 76729 21881
rect 80343 21967 80729 21986
rect 80343 21944 80409 21967
rect 80495 21944 80577 21967
rect 80663 21944 80729 21967
rect 80343 21904 80352 21944
rect 80392 21904 80409 21944
rect 80495 21904 80516 21944
rect 80556 21904 80577 21944
rect 80663 21904 80680 21944
rect 80720 21904 80729 21944
rect 80343 21881 80409 21904
rect 80495 21881 80577 21904
rect 80663 21881 80729 21904
rect 80343 21862 80729 21881
rect 84343 21967 84729 21986
rect 84343 21944 84409 21967
rect 84495 21944 84577 21967
rect 84663 21944 84729 21967
rect 84343 21904 84352 21944
rect 84392 21904 84409 21944
rect 84495 21904 84516 21944
rect 84556 21904 84577 21944
rect 84663 21904 84680 21944
rect 84720 21904 84729 21944
rect 84343 21881 84409 21904
rect 84495 21881 84577 21904
rect 84663 21881 84729 21904
rect 84343 21862 84729 21881
rect 88343 21967 88729 21986
rect 88343 21944 88409 21967
rect 88495 21944 88577 21967
rect 88663 21944 88729 21967
rect 88343 21904 88352 21944
rect 88392 21904 88409 21944
rect 88495 21904 88516 21944
rect 88556 21904 88577 21944
rect 88663 21904 88680 21944
rect 88720 21904 88729 21944
rect 88343 21881 88409 21904
rect 88495 21881 88577 21904
rect 88663 21881 88729 21904
rect 88343 21862 88729 21881
rect 92343 21967 92729 21986
rect 92343 21944 92409 21967
rect 92495 21944 92577 21967
rect 92663 21944 92729 21967
rect 92343 21904 92352 21944
rect 92392 21904 92409 21944
rect 92495 21904 92516 21944
rect 92556 21904 92577 21944
rect 92663 21904 92680 21944
rect 92720 21904 92729 21944
rect 92343 21881 92409 21904
rect 92495 21881 92577 21904
rect 92663 21881 92729 21904
rect 92343 21862 92729 21881
rect 96343 21967 96729 21986
rect 96343 21944 96409 21967
rect 96495 21944 96577 21967
rect 96663 21944 96729 21967
rect 96343 21904 96352 21944
rect 96392 21904 96409 21944
rect 96495 21904 96516 21944
rect 96556 21904 96577 21944
rect 96663 21904 96680 21944
rect 96720 21904 96729 21944
rect 96343 21881 96409 21904
rect 96495 21881 96577 21904
rect 96663 21881 96729 21904
rect 96343 21862 96729 21881
rect 3103 21211 3489 21230
rect 3103 21188 3169 21211
rect 3255 21188 3337 21211
rect 3423 21188 3489 21211
rect 3103 21148 3112 21188
rect 3152 21148 3169 21188
rect 3255 21148 3276 21188
rect 3316 21148 3337 21188
rect 3423 21148 3440 21188
rect 3480 21148 3489 21188
rect 3103 21125 3169 21148
rect 3255 21125 3337 21148
rect 3423 21125 3489 21148
rect 3103 21106 3489 21125
rect 7103 21211 7489 21230
rect 7103 21188 7169 21211
rect 7255 21188 7337 21211
rect 7423 21188 7489 21211
rect 7103 21148 7112 21188
rect 7152 21148 7169 21188
rect 7255 21148 7276 21188
rect 7316 21148 7337 21188
rect 7423 21148 7440 21188
rect 7480 21148 7489 21188
rect 7103 21125 7169 21148
rect 7255 21125 7337 21148
rect 7423 21125 7489 21148
rect 7103 21106 7489 21125
rect 11103 21211 11489 21230
rect 11103 21188 11169 21211
rect 11255 21188 11337 21211
rect 11423 21188 11489 21211
rect 11103 21148 11112 21188
rect 11152 21148 11169 21188
rect 11255 21148 11276 21188
rect 11316 21148 11337 21188
rect 11423 21148 11440 21188
rect 11480 21148 11489 21188
rect 11103 21125 11169 21148
rect 11255 21125 11337 21148
rect 11423 21125 11489 21148
rect 11103 21106 11489 21125
rect 15103 21211 15489 21230
rect 15103 21188 15169 21211
rect 15255 21188 15337 21211
rect 15423 21188 15489 21211
rect 15103 21148 15112 21188
rect 15152 21148 15169 21188
rect 15255 21148 15276 21188
rect 15316 21148 15337 21188
rect 15423 21148 15440 21188
rect 15480 21148 15489 21188
rect 15103 21125 15169 21148
rect 15255 21125 15337 21148
rect 15423 21125 15489 21148
rect 15103 21106 15489 21125
rect 19103 21211 19489 21230
rect 19103 21188 19169 21211
rect 19255 21188 19337 21211
rect 19423 21188 19489 21211
rect 19103 21148 19112 21188
rect 19152 21148 19169 21188
rect 19255 21148 19276 21188
rect 19316 21148 19337 21188
rect 19423 21148 19440 21188
rect 19480 21148 19489 21188
rect 19103 21125 19169 21148
rect 19255 21125 19337 21148
rect 19423 21125 19489 21148
rect 19103 21106 19489 21125
rect 23103 21211 23489 21230
rect 23103 21188 23169 21211
rect 23255 21188 23337 21211
rect 23423 21188 23489 21211
rect 23103 21148 23112 21188
rect 23152 21148 23169 21188
rect 23255 21148 23276 21188
rect 23316 21148 23337 21188
rect 23423 21148 23440 21188
rect 23480 21148 23489 21188
rect 23103 21125 23169 21148
rect 23255 21125 23337 21148
rect 23423 21125 23489 21148
rect 23103 21106 23489 21125
rect 27103 21211 27489 21230
rect 27103 21188 27169 21211
rect 27255 21188 27337 21211
rect 27423 21188 27489 21211
rect 27103 21148 27112 21188
rect 27152 21148 27169 21188
rect 27255 21148 27276 21188
rect 27316 21148 27337 21188
rect 27423 21148 27440 21188
rect 27480 21148 27489 21188
rect 27103 21125 27169 21148
rect 27255 21125 27337 21148
rect 27423 21125 27489 21148
rect 27103 21106 27489 21125
rect 31103 21211 31489 21230
rect 31103 21188 31169 21211
rect 31255 21188 31337 21211
rect 31423 21188 31489 21211
rect 31103 21148 31112 21188
rect 31152 21148 31169 21188
rect 31255 21148 31276 21188
rect 31316 21148 31337 21188
rect 31423 21148 31440 21188
rect 31480 21148 31489 21188
rect 31103 21125 31169 21148
rect 31255 21125 31337 21148
rect 31423 21125 31489 21148
rect 31103 21106 31489 21125
rect 35103 21211 35489 21230
rect 35103 21188 35169 21211
rect 35255 21188 35337 21211
rect 35423 21188 35489 21211
rect 35103 21148 35112 21188
rect 35152 21148 35169 21188
rect 35255 21148 35276 21188
rect 35316 21148 35337 21188
rect 35423 21148 35440 21188
rect 35480 21148 35489 21188
rect 35103 21125 35169 21148
rect 35255 21125 35337 21148
rect 35423 21125 35489 21148
rect 35103 21106 35489 21125
rect 39103 21211 39489 21230
rect 39103 21188 39169 21211
rect 39255 21188 39337 21211
rect 39423 21188 39489 21211
rect 39103 21148 39112 21188
rect 39152 21148 39169 21188
rect 39255 21148 39276 21188
rect 39316 21148 39337 21188
rect 39423 21148 39440 21188
rect 39480 21148 39489 21188
rect 39103 21125 39169 21148
rect 39255 21125 39337 21148
rect 39423 21125 39489 21148
rect 39103 21106 39489 21125
rect 43103 21211 43489 21230
rect 43103 21188 43169 21211
rect 43255 21188 43337 21211
rect 43423 21188 43489 21211
rect 43103 21148 43112 21188
rect 43152 21148 43169 21188
rect 43255 21148 43276 21188
rect 43316 21148 43337 21188
rect 43423 21148 43440 21188
rect 43480 21148 43489 21188
rect 43103 21125 43169 21148
rect 43255 21125 43337 21148
rect 43423 21125 43489 21148
rect 43103 21106 43489 21125
rect 47103 21211 47489 21230
rect 47103 21188 47169 21211
rect 47255 21188 47337 21211
rect 47423 21188 47489 21211
rect 47103 21148 47112 21188
rect 47152 21148 47169 21188
rect 47255 21148 47276 21188
rect 47316 21148 47337 21188
rect 47423 21148 47440 21188
rect 47480 21148 47489 21188
rect 47103 21125 47169 21148
rect 47255 21125 47337 21148
rect 47423 21125 47489 21148
rect 47103 21106 47489 21125
rect 51103 21211 51489 21230
rect 51103 21188 51169 21211
rect 51255 21188 51337 21211
rect 51423 21188 51489 21211
rect 51103 21148 51112 21188
rect 51152 21148 51169 21188
rect 51255 21148 51276 21188
rect 51316 21148 51337 21188
rect 51423 21148 51440 21188
rect 51480 21148 51489 21188
rect 51103 21125 51169 21148
rect 51255 21125 51337 21148
rect 51423 21125 51489 21148
rect 51103 21106 51489 21125
rect 55103 21211 55489 21230
rect 55103 21188 55169 21211
rect 55255 21188 55337 21211
rect 55423 21188 55489 21211
rect 55103 21148 55112 21188
rect 55152 21148 55169 21188
rect 55255 21148 55276 21188
rect 55316 21148 55337 21188
rect 55423 21148 55440 21188
rect 55480 21148 55489 21188
rect 55103 21125 55169 21148
rect 55255 21125 55337 21148
rect 55423 21125 55489 21148
rect 55103 21106 55489 21125
rect 59103 21211 59489 21230
rect 59103 21188 59169 21211
rect 59255 21188 59337 21211
rect 59423 21188 59489 21211
rect 59103 21148 59112 21188
rect 59152 21148 59169 21188
rect 59255 21148 59276 21188
rect 59316 21148 59337 21188
rect 59423 21148 59440 21188
rect 59480 21148 59489 21188
rect 59103 21125 59169 21148
rect 59255 21125 59337 21148
rect 59423 21125 59489 21148
rect 59103 21106 59489 21125
rect 63103 21211 63489 21230
rect 63103 21188 63169 21211
rect 63255 21188 63337 21211
rect 63423 21188 63489 21211
rect 63103 21148 63112 21188
rect 63152 21148 63169 21188
rect 63255 21148 63276 21188
rect 63316 21148 63337 21188
rect 63423 21148 63440 21188
rect 63480 21148 63489 21188
rect 63103 21125 63169 21148
rect 63255 21125 63337 21148
rect 63423 21125 63489 21148
rect 63103 21106 63489 21125
rect 67103 21211 67489 21230
rect 67103 21188 67169 21211
rect 67255 21188 67337 21211
rect 67423 21188 67489 21211
rect 67103 21148 67112 21188
rect 67152 21148 67169 21188
rect 67255 21148 67276 21188
rect 67316 21148 67337 21188
rect 67423 21148 67440 21188
rect 67480 21148 67489 21188
rect 67103 21125 67169 21148
rect 67255 21125 67337 21148
rect 67423 21125 67489 21148
rect 67103 21106 67489 21125
rect 71103 21211 71489 21230
rect 71103 21188 71169 21211
rect 71255 21188 71337 21211
rect 71423 21188 71489 21211
rect 71103 21148 71112 21188
rect 71152 21148 71169 21188
rect 71255 21148 71276 21188
rect 71316 21148 71337 21188
rect 71423 21148 71440 21188
rect 71480 21148 71489 21188
rect 71103 21125 71169 21148
rect 71255 21125 71337 21148
rect 71423 21125 71489 21148
rect 71103 21106 71489 21125
rect 75103 21211 75489 21230
rect 75103 21188 75169 21211
rect 75255 21188 75337 21211
rect 75423 21188 75489 21211
rect 75103 21148 75112 21188
rect 75152 21148 75169 21188
rect 75255 21148 75276 21188
rect 75316 21148 75337 21188
rect 75423 21148 75440 21188
rect 75480 21148 75489 21188
rect 75103 21125 75169 21148
rect 75255 21125 75337 21148
rect 75423 21125 75489 21148
rect 75103 21106 75489 21125
rect 79103 21211 79489 21230
rect 79103 21188 79169 21211
rect 79255 21188 79337 21211
rect 79423 21188 79489 21211
rect 79103 21148 79112 21188
rect 79152 21148 79169 21188
rect 79255 21148 79276 21188
rect 79316 21148 79337 21188
rect 79423 21148 79440 21188
rect 79480 21148 79489 21188
rect 79103 21125 79169 21148
rect 79255 21125 79337 21148
rect 79423 21125 79489 21148
rect 79103 21106 79489 21125
rect 83103 21211 83489 21230
rect 83103 21188 83169 21211
rect 83255 21188 83337 21211
rect 83423 21188 83489 21211
rect 83103 21148 83112 21188
rect 83152 21148 83169 21188
rect 83255 21148 83276 21188
rect 83316 21148 83337 21188
rect 83423 21148 83440 21188
rect 83480 21148 83489 21188
rect 83103 21125 83169 21148
rect 83255 21125 83337 21148
rect 83423 21125 83489 21148
rect 83103 21106 83489 21125
rect 87103 21211 87489 21230
rect 87103 21188 87169 21211
rect 87255 21188 87337 21211
rect 87423 21188 87489 21211
rect 87103 21148 87112 21188
rect 87152 21148 87169 21188
rect 87255 21148 87276 21188
rect 87316 21148 87337 21188
rect 87423 21148 87440 21188
rect 87480 21148 87489 21188
rect 87103 21125 87169 21148
rect 87255 21125 87337 21148
rect 87423 21125 87489 21148
rect 87103 21106 87489 21125
rect 91103 21211 91489 21230
rect 91103 21188 91169 21211
rect 91255 21188 91337 21211
rect 91423 21188 91489 21211
rect 91103 21148 91112 21188
rect 91152 21148 91169 21188
rect 91255 21148 91276 21188
rect 91316 21148 91337 21188
rect 91423 21148 91440 21188
rect 91480 21148 91489 21188
rect 91103 21125 91169 21148
rect 91255 21125 91337 21148
rect 91423 21125 91489 21148
rect 91103 21106 91489 21125
rect 95103 21211 95489 21230
rect 95103 21188 95169 21211
rect 95255 21188 95337 21211
rect 95423 21188 95489 21211
rect 95103 21148 95112 21188
rect 95152 21148 95169 21188
rect 95255 21148 95276 21188
rect 95316 21148 95337 21188
rect 95423 21148 95440 21188
rect 95480 21148 95489 21188
rect 95103 21125 95169 21148
rect 95255 21125 95337 21148
rect 95423 21125 95489 21148
rect 95103 21106 95489 21125
rect 99103 21211 99489 21230
rect 99103 21188 99169 21211
rect 99255 21188 99337 21211
rect 99423 21188 99489 21211
rect 99103 21148 99112 21188
rect 99152 21148 99169 21188
rect 99255 21148 99276 21188
rect 99316 21148 99337 21188
rect 99423 21148 99440 21188
rect 99480 21148 99489 21188
rect 99103 21125 99169 21148
rect 99255 21125 99337 21148
rect 99423 21125 99489 21148
rect 99103 21106 99489 21125
rect 4343 20455 4729 20474
rect 4343 20432 4409 20455
rect 4495 20432 4577 20455
rect 4663 20432 4729 20455
rect 4343 20392 4352 20432
rect 4392 20392 4409 20432
rect 4495 20392 4516 20432
rect 4556 20392 4577 20432
rect 4663 20392 4680 20432
rect 4720 20392 4729 20432
rect 4343 20369 4409 20392
rect 4495 20369 4577 20392
rect 4663 20369 4729 20392
rect 4343 20350 4729 20369
rect 8343 20455 8729 20474
rect 8343 20432 8409 20455
rect 8495 20432 8577 20455
rect 8663 20432 8729 20455
rect 8343 20392 8352 20432
rect 8392 20392 8409 20432
rect 8495 20392 8516 20432
rect 8556 20392 8577 20432
rect 8663 20392 8680 20432
rect 8720 20392 8729 20432
rect 8343 20369 8409 20392
rect 8495 20369 8577 20392
rect 8663 20369 8729 20392
rect 8343 20350 8729 20369
rect 12343 20455 12729 20474
rect 12343 20432 12409 20455
rect 12495 20432 12577 20455
rect 12663 20432 12729 20455
rect 12343 20392 12352 20432
rect 12392 20392 12409 20432
rect 12495 20392 12516 20432
rect 12556 20392 12577 20432
rect 12663 20392 12680 20432
rect 12720 20392 12729 20432
rect 12343 20369 12409 20392
rect 12495 20369 12577 20392
rect 12663 20369 12729 20392
rect 12343 20350 12729 20369
rect 16343 20455 16729 20474
rect 16343 20432 16409 20455
rect 16495 20432 16577 20455
rect 16663 20432 16729 20455
rect 16343 20392 16352 20432
rect 16392 20392 16409 20432
rect 16495 20392 16516 20432
rect 16556 20392 16577 20432
rect 16663 20392 16680 20432
rect 16720 20392 16729 20432
rect 16343 20369 16409 20392
rect 16495 20369 16577 20392
rect 16663 20369 16729 20392
rect 16343 20350 16729 20369
rect 20343 20455 20729 20474
rect 20343 20432 20409 20455
rect 20495 20432 20577 20455
rect 20663 20432 20729 20455
rect 20343 20392 20352 20432
rect 20392 20392 20409 20432
rect 20495 20392 20516 20432
rect 20556 20392 20577 20432
rect 20663 20392 20680 20432
rect 20720 20392 20729 20432
rect 20343 20369 20409 20392
rect 20495 20369 20577 20392
rect 20663 20369 20729 20392
rect 20343 20350 20729 20369
rect 24343 20455 24729 20474
rect 24343 20432 24409 20455
rect 24495 20432 24577 20455
rect 24663 20432 24729 20455
rect 24343 20392 24352 20432
rect 24392 20392 24409 20432
rect 24495 20392 24516 20432
rect 24556 20392 24577 20432
rect 24663 20392 24680 20432
rect 24720 20392 24729 20432
rect 24343 20369 24409 20392
rect 24495 20369 24577 20392
rect 24663 20369 24729 20392
rect 24343 20350 24729 20369
rect 28343 20455 28729 20474
rect 28343 20432 28409 20455
rect 28495 20432 28577 20455
rect 28663 20432 28729 20455
rect 28343 20392 28352 20432
rect 28392 20392 28409 20432
rect 28495 20392 28516 20432
rect 28556 20392 28577 20432
rect 28663 20392 28680 20432
rect 28720 20392 28729 20432
rect 28343 20369 28409 20392
rect 28495 20369 28577 20392
rect 28663 20369 28729 20392
rect 28343 20350 28729 20369
rect 32343 20455 32729 20474
rect 32343 20432 32409 20455
rect 32495 20432 32577 20455
rect 32663 20432 32729 20455
rect 32343 20392 32352 20432
rect 32392 20392 32409 20432
rect 32495 20392 32516 20432
rect 32556 20392 32577 20432
rect 32663 20392 32680 20432
rect 32720 20392 32729 20432
rect 32343 20369 32409 20392
rect 32495 20369 32577 20392
rect 32663 20369 32729 20392
rect 32343 20350 32729 20369
rect 36343 20455 36729 20474
rect 36343 20432 36409 20455
rect 36495 20432 36577 20455
rect 36663 20432 36729 20455
rect 36343 20392 36352 20432
rect 36392 20392 36409 20432
rect 36495 20392 36516 20432
rect 36556 20392 36577 20432
rect 36663 20392 36680 20432
rect 36720 20392 36729 20432
rect 36343 20369 36409 20392
rect 36495 20369 36577 20392
rect 36663 20369 36729 20392
rect 36343 20350 36729 20369
rect 40343 20455 40729 20474
rect 40343 20432 40409 20455
rect 40495 20432 40577 20455
rect 40663 20432 40729 20455
rect 40343 20392 40352 20432
rect 40392 20392 40409 20432
rect 40495 20392 40516 20432
rect 40556 20392 40577 20432
rect 40663 20392 40680 20432
rect 40720 20392 40729 20432
rect 40343 20369 40409 20392
rect 40495 20369 40577 20392
rect 40663 20369 40729 20392
rect 40343 20350 40729 20369
rect 44343 20455 44729 20474
rect 44343 20432 44409 20455
rect 44495 20432 44577 20455
rect 44663 20432 44729 20455
rect 44343 20392 44352 20432
rect 44392 20392 44409 20432
rect 44495 20392 44516 20432
rect 44556 20392 44577 20432
rect 44663 20392 44680 20432
rect 44720 20392 44729 20432
rect 44343 20369 44409 20392
rect 44495 20369 44577 20392
rect 44663 20369 44729 20392
rect 44343 20350 44729 20369
rect 48343 20455 48729 20474
rect 48343 20432 48409 20455
rect 48495 20432 48577 20455
rect 48663 20432 48729 20455
rect 48343 20392 48352 20432
rect 48392 20392 48409 20432
rect 48495 20392 48516 20432
rect 48556 20392 48577 20432
rect 48663 20392 48680 20432
rect 48720 20392 48729 20432
rect 48343 20369 48409 20392
rect 48495 20369 48577 20392
rect 48663 20369 48729 20392
rect 48343 20350 48729 20369
rect 52343 20455 52729 20474
rect 52343 20432 52409 20455
rect 52495 20432 52577 20455
rect 52663 20432 52729 20455
rect 52343 20392 52352 20432
rect 52392 20392 52409 20432
rect 52495 20392 52516 20432
rect 52556 20392 52577 20432
rect 52663 20392 52680 20432
rect 52720 20392 52729 20432
rect 52343 20369 52409 20392
rect 52495 20369 52577 20392
rect 52663 20369 52729 20392
rect 52343 20350 52729 20369
rect 56343 20455 56729 20474
rect 56343 20432 56409 20455
rect 56495 20432 56577 20455
rect 56663 20432 56729 20455
rect 56343 20392 56352 20432
rect 56392 20392 56409 20432
rect 56495 20392 56516 20432
rect 56556 20392 56577 20432
rect 56663 20392 56680 20432
rect 56720 20392 56729 20432
rect 56343 20369 56409 20392
rect 56495 20369 56577 20392
rect 56663 20369 56729 20392
rect 56343 20350 56729 20369
rect 60343 20455 60729 20474
rect 60343 20432 60409 20455
rect 60495 20432 60577 20455
rect 60663 20432 60729 20455
rect 60343 20392 60352 20432
rect 60392 20392 60409 20432
rect 60495 20392 60516 20432
rect 60556 20392 60577 20432
rect 60663 20392 60680 20432
rect 60720 20392 60729 20432
rect 60343 20369 60409 20392
rect 60495 20369 60577 20392
rect 60663 20369 60729 20392
rect 60343 20350 60729 20369
rect 64343 20455 64729 20474
rect 64343 20432 64409 20455
rect 64495 20432 64577 20455
rect 64663 20432 64729 20455
rect 64343 20392 64352 20432
rect 64392 20392 64409 20432
rect 64495 20392 64516 20432
rect 64556 20392 64577 20432
rect 64663 20392 64680 20432
rect 64720 20392 64729 20432
rect 64343 20369 64409 20392
rect 64495 20369 64577 20392
rect 64663 20369 64729 20392
rect 64343 20350 64729 20369
rect 68343 20455 68729 20474
rect 68343 20432 68409 20455
rect 68495 20432 68577 20455
rect 68663 20432 68729 20455
rect 68343 20392 68352 20432
rect 68392 20392 68409 20432
rect 68495 20392 68516 20432
rect 68556 20392 68577 20432
rect 68663 20392 68680 20432
rect 68720 20392 68729 20432
rect 68343 20369 68409 20392
rect 68495 20369 68577 20392
rect 68663 20369 68729 20392
rect 68343 20350 68729 20369
rect 72343 20455 72729 20474
rect 72343 20432 72409 20455
rect 72495 20432 72577 20455
rect 72663 20432 72729 20455
rect 72343 20392 72352 20432
rect 72392 20392 72409 20432
rect 72495 20392 72516 20432
rect 72556 20392 72577 20432
rect 72663 20392 72680 20432
rect 72720 20392 72729 20432
rect 72343 20369 72409 20392
rect 72495 20369 72577 20392
rect 72663 20369 72729 20392
rect 72343 20350 72729 20369
rect 76343 20455 76729 20474
rect 76343 20432 76409 20455
rect 76495 20432 76577 20455
rect 76663 20432 76729 20455
rect 76343 20392 76352 20432
rect 76392 20392 76409 20432
rect 76495 20392 76516 20432
rect 76556 20392 76577 20432
rect 76663 20392 76680 20432
rect 76720 20392 76729 20432
rect 76343 20369 76409 20392
rect 76495 20369 76577 20392
rect 76663 20369 76729 20392
rect 76343 20350 76729 20369
rect 80343 20455 80729 20474
rect 80343 20432 80409 20455
rect 80495 20432 80577 20455
rect 80663 20432 80729 20455
rect 80343 20392 80352 20432
rect 80392 20392 80409 20432
rect 80495 20392 80516 20432
rect 80556 20392 80577 20432
rect 80663 20392 80680 20432
rect 80720 20392 80729 20432
rect 80343 20369 80409 20392
rect 80495 20369 80577 20392
rect 80663 20369 80729 20392
rect 80343 20350 80729 20369
rect 84343 20455 84729 20474
rect 84343 20432 84409 20455
rect 84495 20432 84577 20455
rect 84663 20432 84729 20455
rect 84343 20392 84352 20432
rect 84392 20392 84409 20432
rect 84495 20392 84516 20432
rect 84556 20392 84577 20432
rect 84663 20392 84680 20432
rect 84720 20392 84729 20432
rect 84343 20369 84409 20392
rect 84495 20369 84577 20392
rect 84663 20369 84729 20392
rect 84343 20350 84729 20369
rect 88343 20455 88729 20474
rect 88343 20432 88409 20455
rect 88495 20432 88577 20455
rect 88663 20432 88729 20455
rect 88343 20392 88352 20432
rect 88392 20392 88409 20432
rect 88495 20392 88516 20432
rect 88556 20392 88577 20432
rect 88663 20392 88680 20432
rect 88720 20392 88729 20432
rect 88343 20369 88409 20392
rect 88495 20369 88577 20392
rect 88663 20369 88729 20392
rect 88343 20350 88729 20369
rect 92343 20455 92729 20474
rect 92343 20432 92409 20455
rect 92495 20432 92577 20455
rect 92663 20432 92729 20455
rect 92343 20392 92352 20432
rect 92392 20392 92409 20432
rect 92495 20392 92516 20432
rect 92556 20392 92577 20432
rect 92663 20392 92680 20432
rect 92720 20392 92729 20432
rect 92343 20369 92409 20392
rect 92495 20369 92577 20392
rect 92663 20369 92729 20392
rect 92343 20350 92729 20369
rect 96343 20455 96729 20474
rect 96343 20432 96409 20455
rect 96495 20432 96577 20455
rect 96663 20432 96729 20455
rect 96343 20392 96352 20432
rect 96392 20392 96409 20432
rect 96495 20392 96516 20432
rect 96556 20392 96577 20432
rect 96663 20392 96680 20432
rect 96720 20392 96729 20432
rect 96343 20369 96409 20392
rect 96495 20369 96577 20392
rect 96663 20369 96729 20392
rect 96343 20350 96729 20369
rect 3103 19699 3489 19718
rect 3103 19676 3169 19699
rect 3255 19676 3337 19699
rect 3423 19676 3489 19699
rect 3103 19636 3112 19676
rect 3152 19636 3169 19676
rect 3255 19636 3276 19676
rect 3316 19636 3337 19676
rect 3423 19636 3440 19676
rect 3480 19636 3489 19676
rect 3103 19613 3169 19636
rect 3255 19613 3337 19636
rect 3423 19613 3489 19636
rect 3103 19594 3489 19613
rect 7103 19699 7489 19718
rect 7103 19676 7169 19699
rect 7255 19676 7337 19699
rect 7423 19676 7489 19699
rect 7103 19636 7112 19676
rect 7152 19636 7169 19676
rect 7255 19636 7276 19676
rect 7316 19636 7337 19676
rect 7423 19636 7440 19676
rect 7480 19636 7489 19676
rect 7103 19613 7169 19636
rect 7255 19613 7337 19636
rect 7423 19613 7489 19636
rect 7103 19594 7489 19613
rect 11103 19699 11489 19718
rect 11103 19676 11169 19699
rect 11255 19676 11337 19699
rect 11423 19676 11489 19699
rect 11103 19636 11112 19676
rect 11152 19636 11169 19676
rect 11255 19636 11276 19676
rect 11316 19636 11337 19676
rect 11423 19636 11440 19676
rect 11480 19636 11489 19676
rect 11103 19613 11169 19636
rect 11255 19613 11337 19636
rect 11423 19613 11489 19636
rect 11103 19594 11489 19613
rect 15103 19699 15489 19718
rect 15103 19676 15169 19699
rect 15255 19676 15337 19699
rect 15423 19676 15489 19699
rect 15103 19636 15112 19676
rect 15152 19636 15169 19676
rect 15255 19636 15276 19676
rect 15316 19636 15337 19676
rect 15423 19636 15440 19676
rect 15480 19636 15489 19676
rect 15103 19613 15169 19636
rect 15255 19613 15337 19636
rect 15423 19613 15489 19636
rect 15103 19594 15489 19613
rect 19103 19699 19489 19718
rect 19103 19676 19169 19699
rect 19255 19676 19337 19699
rect 19423 19676 19489 19699
rect 19103 19636 19112 19676
rect 19152 19636 19169 19676
rect 19255 19636 19276 19676
rect 19316 19636 19337 19676
rect 19423 19636 19440 19676
rect 19480 19636 19489 19676
rect 19103 19613 19169 19636
rect 19255 19613 19337 19636
rect 19423 19613 19489 19636
rect 19103 19594 19489 19613
rect 23103 19699 23489 19718
rect 23103 19676 23169 19699
rect 23255 19676 23337 19699
rect 23423 19676 23489 19699
rect 23103 19636 23112 19676
rect 23152 19636 23169 19676
rect 23255 19636 23276 19676
rect 23316 19636 23337 19676
rect 23423 19636 23440 19676
rect 23480 19636 23489 19676
rect 23103 19613 23169 19636
rect 23255 19613 23337 19636
rect 23423 19613 23489 19636
rect 23103 19594 23489 19613
rect 27103 19699 27489 19718
rect 27103 19676 27169 19699
rect 27255 19676 27337 19699
rect 27423 19676 27489 19699
rect 27103 19636 27112 19676
rect 27152 19636 27169 19676
rect 27255 19636 27276 19676
rect 27316 19636 27337 19676
rect 27423 19636 27440 19676
rect 27480 19636 27489 19676
rect 27103 19613 27169 19636
rect 27255 19613 27337 19636
rect 27423 19613 27489 19636
rect 27103 19594 27489 19613
rect 31103 19699 31489 19718
rect 31103 19676 31169 19699
rect 31255 19676 31337 19699
rect 31423 19676 31489 19699
rect 31103 19636 31112 19676
rect 31152 19636 31169 19676
rect 31255 19636 31276 19676
rect 31316 19636 31337 19676
rect 31423 19636 31440 19676
rect 31480 19636 31489 19676
rect 31103 19613 31169 19636
rect 31255 19613 31337 19636
rect 31423 19613 31489 19636
rect 31103 19594 31489 19613
rect 35103 19699 35489 19718
rect 35103 19676 35169 19699
rect 35255 19676 35337 19699
rect 35423 19676 35489 19699
rect 35103 19636 35112 19676
rect 35152 19636 35169 19676
rect 35255 19636 35276 19676
rect 35316 19636 35337 19676
rect 35423 19636 35440 19676
rect 35480 19636 35489 19676
rect 35103 19613 35169 19636
rect 35255 19613 35337 19636
rect 35423 19613 35489 19636
rect 35103 19594 35489 19613
rect 39103 19699 39489 19718
rect 39103 19676 39169 19699
rect 39255 19676 39337 19699
rect 39423 19676 39489 19699
rect 39103 19636 39112 19676
rect 39152 19636 39169 19676
rect 39255 19636 39276 19676
rect 39316 19636 39337 19676
rect 39423 19636 39440 19676
rect 39480 19636 39489 19676
rect 39103 19613 39169 19636
rect 39255 19613 39337 19636
rect 39423 19613 39489 19636
rect 39103 19594 39489 19613
rect 43103 19699 43489 19718
rect 43103 19676 43169 19699
rect 43255 19676 43337 19699
rect 43423 19676 43489 19699
rect 43103 19636 43112 19676
rect 43152 19636 43169 19676
rect 43255 19636 43276 19676
rect 43316 19636 43337 19676
rect 43423 19636 43440 19676
rect 43480 19636 43489 19676
rect 43103 19613 43169 19636
rect 43255 19613 43337 19636
rect 43423 19613 43489 19636
rect 43103 19594 43489 19613
rect 47103 19699 47489 19718
rect 47103 19676 47169 19699
rect 47255 19676 47337 19699
rect 47423 19676 47489 19699
rect 47103 19636 47112 19676
rect 47152 19636 47169 19676
rect 47255 19636 47276 19676
rect 47316 19636 47337 19676
rect 47423 19636 47440 19676
rect 47480 19636 47489 19676
rect 47103 19613 47169 19636
rect 47255 19613 47337 19636
rect 47423 19613 47489 19636
rect 47103 19594 47489 19613
rect 51103 19699 51489 19718
rect 51103 19676 51169 19699
rect 51255 19676 51337 19699
rect 51423 19676 51489 19699
rect 51103 19636 51112 19676
rect 51152 19636 51169 19676
rect 51255 19636 51276 19676
rect 51316 19636 51337 19676
rect 51423 19636 51440 19676
rect 51480 19636 51489 19676
rect 51103 19613 51169 19636
rect 51255 19613 51337 19636
rect 51423 19613 51489 19636
rect 51103 19594 51489 19613
rect 55103 19699 55489 19718
rect 55103 19676 55169 19699
rect 55255 19676 55337 19699
rect 55423 19676 55489 19699
rect 55103 19636 55112 19676
rect 55152 19636 55169 19676
rect 55255 19636 55276 19676
rect 55316 19636 55337 19676
rect 55423 19636 55440 19676
rect 55480 19636 55489 19676
rect 55103 19613 55169 19636
rect 55255 19613 55337 19636
rect 55423 19613 55489 19636
rect 55103 19594 55489 19613
rect 59103 19699 59489 19718
rect 59103 19676 59169 19699
rect 59255 19676 59337 19699
rect 59423 19676 59489 19699
rect 59103 19636 59112 19676
rect 59152 19636 59169 19676
rect 59255 19636 59276 19676
rect 59316 19636 59337 19676
rect 59423 19636 59440 19676
rect 59480 19636 59489 19676
rect 59103 19613 59169 19636
rect 59255 19613 59337 19636
rect 59423 19613 59489 19636
rect 59103 19594 59489 19613
rect 63103 19699 63489 19718
rect 63103 19676 63169 19699
rect 63255 19676 63337 19699
rect 63423 19676 63489 19699
rect 63103 19636 63112 19676
rect 63152 19636 63169 19676
rect 63255 19636 63276 19676
rect 63316 19636 63337 19676
rect 63423 19636 63440 19676
rect 63480 19636 63489 19676
rect 63103 19613 63169 19636
rect 63255 19613 63337 19636
rect 63423 19613 63489 19636
rect 63103 19594 63489 19613
rect 67103 19699 67489 19718
rect 67103 19676 67169 19699
rect 67255 19676 67337 19699
rect 67423 19676 67489 19699
rect 67103 19636 67112 19676
rect 67152 19636 67169 19676
rect 67255 19636 67276 19676
rect 67316 19636 67337 19676
rect 67423 19636 67440 19676
rect 67480 19636 67489 19676
rect 67103 19613 67169 19636
rect 67255 19613 67337 19636
rect 67423 19613 67489 19636
rect 67103 19594 67489 19613
rect 71103 19699 71489 19718
rect 71103 19676 71169 19699
rect 71255 19676 71337 19699
rect 71423 19676 71489 19699
rect 71103 19636 71112 19676
rect 71152 19636 71169 19676
rect 71255 19636 71276 19676
rect 71316 19636 71337 19676
rect 71423 19636 71440 19676
rect 71480 19636 71489 19676
rect 71103 19613 71169 19636
rect 71255 19613 71337 19636
rect 71423 19613 71489 19636
rect 71103 19594 71489 19613
rect 75103 19699 75489 19718
rect 75103 19676 75169 19699
rect 75255 19676 75337 19699
rect 75423 19676 75489 19699
rect 75103 19636 75112 19676
rect 75152 19636 75169 19676
rect 75255 19636 75276 19676
rect 75316 19636 75337 19676
rect 75423 19636 75440 19676
rect 75480 19636 75489 19676
rect 75103 19613 75169 19636
rect 75255 19613 75337 19636
rect 75423 19613 75489 19636
rect 75103 19594 75489 19613
rect 79103 19699 79489 19718
rect 79103 19676 79169 19699
rect 79255 19676 79337 19699
rect 79423 19676 79489 19699
rect 79103 19636 79112 19676
rect 79152 19636 79169 19676
rect 79255 19636 79276 19676
rect 79316 19636 79337 19676
rect 79423 19636 79440 19676
rect 79480 19636 79489 19676
rect 79103 19613 79169 19636
rect 79255 19613 79337 19636
rect 79423 19613 79489 19636
rect 79103 19594 79489 19613
rect 83103 19699 83489 19718
rect 83103 19676 83169 19699
rect 83255 19676 83337 19699
rect 83423 19676 83489 19699
rect 83103 19636 83112 19676
rect 83152 19636 83169 19676
rect 83255 19636 83276 19676
rect 83316 19636 83337 19676
rect 83423 19636 83440 19676
rect 83480 19636 83489 19676
rect 83103 19613 83169 19636
rect 83255 19613 83337 19636
rect 83423 19613 83489 19636
rect 83103 19594 83489 19613
rect 87103 19699 87489 19718
rect 87103 19676 87169 19699
rect 87255 19676 87337 19699
rect 87423 19676 87489 19699
rect 87103 19636 87112 19676
rect 87152 19636 87169 19676
rect 87255 19636 87276 19676
rect 87316 19636 87337 19676
rect 87423 19636 87440 19676
rect 87480 19636 87489 19676
rect 87103 19613 87169 19636
rect 87255 19613 87337 19636
rect 87423 19613 87489 19636
rect 87103 19594 87489 19613
rect 91103 19699 91489 19718
rect 91103 19676 91169 19699
rect 91255 19676 91337 19699
rect 91423 19676 91489 19699
rect 91103 19636 91112 19676
rect 91152 19636 91169 19676
rect 91255 19636 91276 19676
rect 91316 19636 91337 19676
rect 91423 19636 91440 19676
rect 91480 19636 91489 19676
rect 91103 19613 91169 19636
rect 91255 19613 91337 19636
rect 91423 19613 91489 19636
rect 91103 19594 91489 19613
rect 95103 19699 95489 19718
rect 95103 19676 95169 19699
rect 95255 19676 95337 19699
rect 95423 19676 95489 19699
rect 95103 19636 95112 19676
rect 95152 19636 95169 19676
rect 95255 19636 95276 19676
rect 95316 19636 95337 19676
rect 95423 19636 95440 19676
rect 95480 19636 95489 19676
rect 95103 19613 95169 19636
rect 95255 19613 95337 19636
rect 95423 19613 95489 19636
rect 95103 19594 95489 19613
rect 99103 19699 99489 19718
rect 99103 19676 99169 19699
rect 99255 19676 99337 19699
rect 99423 19676 99489 19699
rect 99103 19636 99112 19676
rect 99152 19636 99169 19676
rect 99255 19636 99276 19676
rect 99316 19636 99337 19676
rect 99423 19636 99440 19676
rect 99480 19636 99489 19676
rect 99103 19613 99169 19636
rect 99255 19613 99337 19636
rect 99423 19613 99489 19636
rect 99103 19594 99489 19613
rect 86450 19363 86574 19382
rect 86450 19277 86469 19363
rect 86555 19340 86574 19363
rect 86555 19300 86764 19340
rect 86804 19300 86813 19340
rect 86555 19277 86574 19300
rect 86450 19258 86574 19277
rect 4343 18943 4729 18962
rect 4343 18920 4409 18943
rect 4495 18920 4577 18943
rect 4663 18920 4729 18943
rect 4343 18880 4352 18920
rect 4392 18880 4409 18920
rect 4495 18880 4516 18920
rect 4556 18880 4577 18920
rect 4663 18880 4680 18920
rect 4720 18880 4729 18920
rect 4343 18857 4409 18880
rect 4495 18857 4577 18880
rect 4663 18857 4729 18880
rect 4343 18838 4729 18857
rect 8343 18943 8729 18962
rect 8343 18920 8409 18943
rect 8495 18920 8577 18943
rect 8663 18920 8729 18943
rect 8343 18880 8352 18920
rect 8392 18880 8409 18920
rect 8495 18880 8516 18920
rect 8556 18880 8577 18920
rect 8663 18880 8680 18920
rect 8720 18880 8729 18920
rect 8343 18857 8409 18880
rect 8495 18857 8577 18880
rect 8663 18857 8729 18880
rect 8343 18838 8729 18857
rect 12343 18943 12729 18962
rect 12343 18920 12409 18943
rect 12495 18920 12577 18943
rect 12663 18920 12729 18943
rect 12343 18880 12352 18920
rect 12392 18880 12409 18920
rect 12495 18880 12516 18920
rect 12556 18880 12577 18920
rect 12663 18880 12680 18920
rect 12720 18880 12729 18920
rect 12343 18857 12409 18880
rect 12495 18857 12577 18880
rect 12663 18857 12729 18880
rect 12343 18838 12729 18857
rect 16343 18943 16729 18962
rect 16343 18920 16409 18943
rect 16495 18920 16577 18943
rect 16663 18920 16729 18943
rect 16343 18880 16352 18920
rect 16392 18880 16409 18920
rect 16495 18880 16516 18920
rect 16556 18880 16577 18920
rect 16663 18880 16680 18920
rect 16720 18880 16729 18920
rect 16343 18857 16409 18880
rect 16495 18857 16577 18880
rect 16663 18857 16729 18880
rect 16343 18838 16729 18857
rect 20343 18943 20729 18962
rect 20343 18920 20409 18943
rect 20495 18920 20577 18943
rect 20663 18920 20729 18943
rect 20343 18880 20352 18920
rect 20392 18880 20409 18920
rect 20495 18880 20516 18920
rect 20556 18880 20577 18920
rect 20663 18880 20680 18920
rect 20720 18880 20729 18920
rect 20343 18857 20409 18880
rect 20495 18857 20577 18880
rect 20663 18857 20729 18880
rect 20343 18838 20729 18857
rect 24343 18943 24729 18962
rect 24343 18920 24409 18943
rect 24495 18920 24577 18943
rect 24663 18920 24729 18943
rect 24343 18880 24352 18920
rect 24392 18880 24409 18920
rect 24495 18880 24516 18920
rect 24556 18880 24577 18920
rect 24663 18880 24680 18920
rect 24720 18880 24729 18920
rect 24343 18857 24409 18880
rect 24495 18857 24577 18880
rect 24663 18857 24729 18880
rect 24343 18838 24729 18857
rect 28343 18943 28729 18962
rect 28343 18920 28409 18943
rect 28495 18920 28577 18943
rect 28663 18920 28729 18943
rect 28343 18880 28352 18920
rect 28392 18880 28409 18920
rect 28495 18880 28516 18920
rect 28556 18880 28577 18920
rect 28663 18880 28680 18920
rect 28720 18880 28729 18920
rect 28343 18857 28409 18880
rect 28495 18857 28577 18880
rect 28663 18857 28729 18880
rect 28343 18838 28729 18857
rect 32343 18943 32729 18962
rect 32343 18920 32409 18943
rect 32495 18920 32577 18943
rect 32663 18920 32729 18943
rect 32343 18880 32352 18920
rect 32392 18880 32409 18920
rect 32495 18880 32516 18920
rect 32556 18880 32577 18920
rect 32663 18880 32680 18920
rect 32720 18880 32729 18920
rect 32343 18857 32409 18880
rect 32495 18857 32577 18880
rect 32663 18857 32729 18880
rect 32343 18838 32729 18857
rect 36343 18943 36729 18962
rect 36343 18920 36409 18943
rect 36495 18920 36577 18943
rect 36663 18920 36729 18943
rect 36343 18880 36352 18920
rect 36392 18880 36409 18920
rect 36495 18880 36516 18920
rect 36556 18880 36577 18920
rect 36663 18880 36680 18920
rect 36720 18880 36729 18920
rect 36343 18857 36409 18880
rect 36495 18857 36577 18880
rect 36663 18857 36729 18880
rect 36343 18838 36729 18857
rect 40343 18943 40729 18962
rect 40343 18920 40409 18943
rect 40495 18920 40577 18943
rect 40663 18920 40729 18943
rect 40343 18880 40352 18920
rect 40392 18880 40409 18920
rect 40495 18880 40516 18920
rect 40556 18880 40577 18920
rect 40663 18880 40680 18920
rect 40720 18880 40729 18920
rect 40343 18857 40409 18880
rect 40495 18857 40577 18880
rect 40663 18857 40729 18880
rect 40343 18838 40729 18857
rect 44343 18943 44729 18962
rect 44343 18920 44409 18943
rect 44495 18920 44577 18943
rect 44663 18920 44729 18943
rect 44343 18880 44352 18920
rect 44392 18880 44409 18920
rect 44495 18880 44516 18920
rect 44556 18880 44577 18920
rect 44663 18880 44680 18920
rect 44720 18880 44729 18920
rect 44343 18857 44409 18880
rect 44495 18857 44577 18880
rect 44663 18857 44729 18880
rect 44343 18838 44729 18857
rect 48343 18943 48729 18962
rect 48343 18920 48409 18943
rect 48495 18920 48577 18943
rect 48663 18920 48729 18943
rect 48343 18880 48352 18920
rect 48392 18880 48409 18920
rect 48495 18880 48516 18920
rect 48556 18880 48577 18920
rect 48663 18880 48680 18920
rect 48720 18880 48729 18920
rect 48343 18857 48409 18880
rect 48495 18857 48577 18880
rect 48663 18857 48729 18880
rect 48343 18838 48729 18857
rect 52343 18943 52729 18962
rect 52343 18920 52409 18943
rect 52495 18920 52577 18943
rect 52663 18920 52729 18943
rect 52343 18880 52352 18920
rect 52392 18880 52409 18920
rect 52495 18880 52516 18920
rect 52556 18880 52577 18920
rect 52663 18880 52680 18920
rect 52720 18880 52729 18920
rect 52343 18857 52409 18880
rect 52495 18857 52577 18880
rect 52663 18857 52729 18880
rect 52343 18838 52729 18857
rect 56343 18943 56729 18962
rect 56343 18920 56409 18943
rect 56495 18920 56577 18943
rect 56663 18920 56729 18943
rect 56343 18880 56352 18920
rect 56392 18880 56409 18920
rect 56495 18880 56516 18920
rect 56556 18880 56577 18920
rect 56663 18880 56680 18920
rect 56720 18880 56729 18920
rect 56343 18857 56409 18880
rect 56495 18857 56577 18880
rect 56663 18857 56729 18880
rect 56343 18838 56729 18857
rect 60343 18943 60729 18962
rect 60343 18920 60409 18943
rect 60495 18920 60577 18943
rect 60663 18920 60729 18943
rect 60343 18880 60352 18920
rect 60392 18880 60409 18920
rect 60495 18880 60516 18920
rect 60556 18880 60577 18920
rect 60663 18880 60680 18920
rect 60720 18880 60729 18920
rect 60343 18857 60409 18880
rect 60495 18857 60577 18880
rect 60663 18857 60729 18880
rect 60343 18838 60729 18857
rect 64343 18943 64729 18962
rect 64343 18920 64409 18943
rect 64495 18920 64577 18943
rect 64663 18920 64729 18943
rect 64343 18880 64352 18920
rect 64392 18880 64409 18920
rect 64495 18880 64516 18920
rect 64556 18880 64577 18920
rect 64663 18880 64680 18920
rect 64720 18880 64729 18920
rect 64343 18857 64409 18880
rect 64495 18857 64577 18880
rect 64663 18857 64729 18880
rect 64343 18838 64729 18857
rect 68343 18943 68729 18962
rect 68343 18920 68409 18943
rect 68495 18920 68577 18943
rect 68663 18920 68729 18943
rect 68343 18880 68352 18920
rect 68392 18880 68409 18920
rect 68495 18880 68516 18920
rect 68556 18880 68577 18920
rect 68663 18880 68680 18920
rect 68720 18880 68729 18920
rect 68343 18857 68409 18880
rect 68495 18857 68577 18880
rect 68663 18857 68729 18880
rect 68343 18838 68729 18857
rect 72343 18943 72729 18962
rect 72343 18920 72409 18943
rect 72495 18920 72577 18943
rect 72663 18920 72729 18943
rect 72343 18880 72352 18920
rect 72392 18880 72409 18920
rect 72495 18880 72516 18920
rect 72556 18880 72577 18920
rect 72663 18880 72680 18920
rect 72720 18880 72729 18920
rect 72343 18857 72409 18880
rect 72495 18857 72577 18880
rect 72663 18857 72729 18880
rect 72343 18838 72729 18857
rect 76343 18943 76729 18962
rect 76343 18920 76409 18943
rect 76495 18920 76577 18943
rect 76663 18920 76729 18943
rect 76343 18880 76352 18920
rect 76392 18880 76409 18920
rect 76495 18880 76516 18920
rect 76556 18880 76577 18920
rect 76663 18880 76680 18920
rect 76720 18880 76729 18920
rect 76343 18857 76409 18880
rect 76495 18857 76577 18880
rect 76663 18857 76729 18880
rect 76343 18838 76729 18857
rect 80343 18943 80729 18962
rect 80343 18920 80409 18943
rect 80495 18920 80577 18943
rect 80663 18920 80729 18943
rect 80343 18880 80352 18920
rect 80392 18880 80409 18920
rect 80495 18880 80516 18920
rect 80556 18880 80577 18920
rect 80663 18880 80680 18920
rect 80720 18880 80729 18920
rect 80343 18857 80409 18880
rect 80495 18857 80577 18880
rect 80663 18857 80729 18880
rect 80343 18838 80729 18857
rect 84343 18943 84729 18962
rect 84343 18920 84409 18943
rect 84495 18920 84577 18943
rect 84663 18920 84729 18943
rect 84343 18880 84352 18920
rect 84392 18880 84409 18920
rect 84495 18880 84516 18920
rect 84556 18880 84577 18920
rect 84663 18880 84680 18920
rect 84720 18880 84729 18920
rect 84343 18857 84409 18880
rect 84495 18857 84577 18880
rect 84663 18857 84729 18880
rect 84343 18838 84729 18857
rect 88343 18943 88729 18962
rect 88343 18920 88409 18943
rect 88495 18920 88577 18943
rect 88663 18920 88729 18943
rect 88343 18880 88352 18920
rect 88392 18880 88409 18920
rect 88495 18880 88516 18920
rect 88556 18880 88577 18920
rect 88663 18880 88680 18920
rect 88720 18880 88729 18920
rect 88343 18857 88409 18880
rect 88495 18857 88577 18880
rect 88663 18857 88729 18880
rect 88343 18838 88729 18857
rect 92343 18943 92729 18962
rect 92343 18920 92409 18943
rect 92495 18920 92577 18943
rect 92663 18920 92729 18943
rect 92343 18880 92352 18920
rect 92392 18880 92409 18920
rect 92495 18880 92516 18920
rect 92556 18880 92577 18920
rect 92663 18880 92680 18920
rect 92720 18880 92729 18920
rect 92343 18857 92409 18880
rect 92495 18857 92577 18880
rect 92663 18857 92729 18880
rect 92343 18838 92729 18857
rect 96343 18943 96729 18962
rect 96343 18920 96409 18943
rect 96495 18920 96577 18943
rect 96663 18920 96729 18943
rect 96343 18880 96352 18920
rect 96392 18880 96409 18920
rect 96495 18880 96516 18920
rect 96556 18880 96577 18920
rect 96663 18880 96680 18920
rect 96720 18880 96729 18920
rect 96343 18857 96409 18880
rect 96495 18857 96577 18880
rect 96663 18857 96729 18880
rect 96343 18838 96729 18857
rect 3103 18187 3489 18206
rect 3103 18164 3169 18187
rect 3255 18164 3337 18187
rect 3423 18164 3489 18187
rect 3103 18124 3112 18164
rect 3152 18124 3169 18164
rect 3255 18124 3276 18164
rect 3316 18124 3337 18164
rect 3423 18124 3440 18164
rect 3480 18124 3489 18164
rect 3103 18101 3169 18124
rect 3255 18101 3337 18124
rect 3423 18101 3489 18124
rect 3103 18082 3489 18101
rect 7103 18187 7489 18206
rect 7103 18164 7169 18187
rect 7255 18164 7337 18187
rect 7423 18164 7489 18187
rect 7103 18124 7112 18164
rect 7152 18124 7169 18164
rect 7255 18124 7276 18164
rect 7316 18124 7337 18164
rect 7423 18124 7440 18164
rect 7480 18124 7489 18164
rect 7103 18101 7169 18124
rect 7255 18101 7337 18124
rect 7423 18101 7489 18124
rect 7103 18082 7489 18101
rect 11103 18187 11489 18206
rect 11103 18164 11169 18187
rect 11255 18164 11337 18187
rect 11423 18164 11489 18187
rect 11103 18124 11112 18164
rect 11152 18124 11169 18164
rect 11255 18124 11276 18164
rect 11316 18124 11337 18164
rect 11423 18124 11440 18164
rect 11480 18124 11489 18164
rect 11103 18101 11169 18124
rect 11255 18101 11337 18124
rect 11423 18101 11489 18124
rect 11103 18082 11489 18101
rect 15103 18187 15489 18206
rect 15103 18164 15169 18187
rect 15255 18164 15337 18187
rect 15423 18164 15489 18187
rect 15103 18124 15112 18164
rect 15152 18124 15169 18164
rect 15255 18124 15276 18164
rect 15316 18124 15337 18164
rect 15423 18124 15440 18164
rect 15480 18124 15489 18164
rect 15103 18101 15169 18124
rect 15255 18101 15337 18124
rect 15423 18101 15489 18124
rect 15103 18082 15489 18101
rect 19103 18187 19489 18206
rect 19103 18164 19169 18187
rect 19255 18164 19337 18187
rect 19423 18164 19489 18187
rect 19103 18124 19112 18164
rect 19152 18124 19169 18164
rect 19255 18124 19276 18164
rect 19316 18124 19337 18164
rect 19423 18124 19440 18164
rect 19480 18124 19489 18164
rect 19103 18101 19169 18124
rect 19255 18101 19337 18124
rect 19423 18101 19489 18124
rect 19103 18082 19489 18101
rect 23103 18187 23489 18206
rect 23103 18164 23169 18187
rect 23255 18164 23337 18187
rect 23423 18164 23489 18187
rect 23103 18124 23112 18164
rect 23152 18124 23169 18164
rect 23255 18124 23276 18164
rect 23316 18124 23337 18164
rect 23423 18124 23440 18164
rect 23480 18124 23489 18164
rect 23103 18101 23169 18124
rect 23255 18101 23337 18124
rect 23423 18101 23489 18124
rect 23103 18082 23489 18101
rect 27103 18187 27489 18206
rect 27103 18164 27169 18187
rect 27255 18164 27337 18187
rect 27423 18164 27489 18187
rect 27103 18124 27112 18164
rect 27152 18124 27169 18164
rect 27255 18124 27276 18164
rect 27316 18124 27337 18164
rect 27423 18124 27440 18164
rect 27480 18124 27489 18164
rect 27103 18101 27169 18124
rect 27255 18101 27337 18124
rect 27423 18101 27489 18124
rect 27103 18082 27489 18101
rect 31103 18187 31489 18206
rect 31103 18164 31169 18187
rect 31255 18164 31337 18187
rect 31423 18164 31489 18187
rect 31103 18124 31112 18164
rect 31152 18124 31169 18164
rect 31255 18124 31276 18164
rect 31316 18124 31337 18164
rect 31423 18124 31440 18164
rect 31480 18124 31489 18164
rect 31103 18101 31169 18124
rect 31255 18101 31337 18124
rect 31423 18101 31489 18124
rect 31103 18082 31489 18101
rect 35103 18187 35489 18206
rect 35103 18164 35169 18187
rect 35255 18164 35337 18187
rect 35423 18164 35489 18187
rect 35103 18124 35112 18164
rect 35152 18124 35169 18164
rect 35255 18124 35276 18164
rect 35316 18124 35337 18164
rect 35423 18124 35440 18164
rect 35480 18124 35489 18164
rect 35103 18101 35169 18124
rect 35255 18101 35337 18124
rect 35423 18101 35489 18124
rect 35103 18082 35489 18101
rect 39103 18187 39489 18206
rect 39103 18164 39169 18187
rect 39255 18164 39337 18187
rect 39423 18164 39489 18187
rect 39103 18124 39112 18164
rect 39152 18124 39169 18164
rect 39255 18124 39276 18164
rect 39316 18124 39337 18164
rect 39423 18124 39440 18164
rect 39480 18124 39489 18164
rect 39103 18101 39169 18124
rect 39255 18101 39337 18124
rect 39423 18101 39489 18124
rect 39103 18082 39489 18101
rect 43103 18187 43489 18206
rect 43103 18164 43169 18187
rect 43255 18164 43337 18187
rect 43423 18164 43489 18187
rect 43103 18124 43112 18164
rect 43152 18124 43169 18164
rect 43255 18124 43276 18164
rect 43316 18124 43337 18164
rect 43423 18124 43440 18164
rect 43480 18124 43489 18164
rect 43103 18101 43169 18124
rect 43255 18101 43337 18124
rect 43423 18101 43489 18124
rect 43103 18082 43489 18101
rect 47103 18187 47489 18206
rect 47103 18164 47169 18187
rect 47255 18164 47337 18187
rect 47423 18164 47489 18187
rect 47103 18124 47112 18164
rect 47152 18124 47169 18164
rect 47255 18124 47276 18164
rect 47316 18124 47337 18164
rect 47423 18124 47440 18164
rect 47480 18124 47489 18164
rect 47103 18101 47169 18124
rect 47255 18101 47337 18124
rect 47423 18101 47489 18124
rect 47103 18082 47489 18101
rect 51103 18187 51489 18206
rect 51103 18164 51169 18187
rect 51255 18164 51337 18187
rect 51423 18164 51489 18187
rect 51103 18124 51112 18164
rect 51152 18124 51169 18164
rect 51255 18124 51276 18164
rect 51316 18124 51337 18164
rect 51423 18124 51440 18164
rect 51480 18124 51489 18164
rect 51103 18101 51169 18124
rect 51255 18101 51337 18124
rect 51423 18101 51489 18124
rect 51103 18082 51489 18101
rect 55103 18187 55489 18206
rect 55103 18164 55169 18187
rect 55255 18164 55337 18187
rect 55423 18164 55489 18187
rect 55103 18124 55112 18164
rect 55152 18124 55169 18164
rect 55255 18124 55276 18164
rect 55316 18124 55337 18164
rect 55423 18124 55440 18164
rect 55480 18124 55489 18164
rect 55103 18101 55169 18124
rect 55255 18101 55337 18124
rect 55423 18101 55489 18124
rect 55103 18082 55489 18101
rect 59103 18187 59489 18206
rect 59103 18164 59169 18187
rect 59255 18164 59337 18187
rect 59423 18164 59489 18187
rect 59103 18124 59112 18164
rect 59152 18124 59169 18164
rect 59255 18124 59276 18164
rect 59316 18124 59337 18164
rect 59423 18124 59440 18164
rect 59480 18124 59489 18164
rect 59103 18101 59169 18124
rect 59255 18101 59337 18124
rect 59423 18101 59489 18124
rect 59103 18082 59489 18101
rect 63103 18187 63489 18206
rect 63103 18164 63169 18187
rect 63255 18164 63337 18187
rect 63423 18164 63489 18187
rect 63103 18124 63112 18164
rect 63152 18124 63169 18164
rect 63255 18124 63276 18164
rect 63316 18124 63337 18164
rect 63423 18124 63440 18164
rect 63480 18124 63489 18164
rect 63103 18101 63169 18124
rect 63255 18101 63337 18124
rect 63423 18101 63489 18124
rect 63103 18082 63489 18101
rect 67103 18187 67489 18206
rect 67103 18164 67169 18187
rect 67255 18164 67337 18187
rect 67423 18164 67489 18187
rect 67103 18124 67112 18164
rect 67152 18124 67169 18164
rect 67255 18124 67276 18164
rect 67316 18124 67337 18164
rect 67423 18124 67440 18164
rect 67480 18124 67489 18164
rect 67103 18101 67169 18124
rect 67255 18101 67337 18124
rect 67423 18101 67489 18124
rect 67103 18082 67489 18101
rect 71103 18187 71489 18206
rect 71103 18164 71169 18187
rect 71255 18164 71337 18187
rect 71423 18164 71489 18187
rect 71103 18124 71112 18164
rect 71152 18124 71169 18164
rect 71255 18124 71276 18164
rect 71316 18124 71337 18164
rect 71423 18124 71440 18164
rect 71480 18124 71489 18164
rect 71103 18101 71169 18124
rect 71255 18101 71337 18124
rect 71423 18101 71489 18124
rect 71103 18082 71489 18101
rect 75103 18187 75489 18206
rect 75103 18164 75169 18187
rect 75255 18164 75337 18187
rect 75423 18164 75489 18187
rect 75103 18124 75112 18164
rect 75152 18124 75169 18164
rect 75255 18124 75276 18164
rect 75316 18124 75337 18164
rect 75423 18124 75440 18164
rect 75480 18124 75489 18164
rect 75103 18101 75169 18124
rect 75255 18101 75337 18124
rect 75423 18101 75489 18124
rect 75103 18082 75489 18101
rect 79103 18187 79489 18206
rect 79103 18164 79169 18187
rect 79255 18164 79337 18187
rect 79423 18164 79489 18187
rect 79103 18124 79112 18164
rect 79152 18124 79169 18164
rect 79255 18124 79276 18164
rect 79316 18124 79337 18164
rect 79423 18124 79440 18164
rect 79480 18124 79489 18164
rect 79103 18101 79169 18124
rect 79255 18101 79337 18124
rect 79423 18101 79489 18124
rect 79103 18082 79489 18101
rect 83103 18187 83489 18206
rect 83103 18164 83169 18187
rect 83255 18164 83337 18187
rect 83423 18164 83489 18187
rect 83103 18124 83112 18164
rect 83152 18124 83169 18164
rect 83255 18124 83276 18164
rect 83316 18124 83337 18164
rect 83423 18124 83440 18164
rect 83480 18124 83489 18164
rect 83103 18101 83169 18124
rect 83255 18101 83337 18124
rect 83423 18101 83489 18124
rect 83103 18082 83489 18101
rect 87103 18187 87489 18206
rect 87103 18164 87169 18187
rect 87255 18164 87337 18187
rect 87423 18164 87489 18187
rect 87103 18124 87112 18164
rect 87152 18124 87169 18164
rect 87255 18124 87276 18164
rect 87316 18124 87337 18164
rect 87423 18124 87440 18164
rect 87480 18124 87489 18164
rect 87103 18101 87169 18124
rect 87255 18101 87337 18124
rect 87423 18101 87489 18124
rect 87103 18082 87489 18101
rect 91103 18187 91489 18206
rect 91103 18164 91169 18187
rect 91255 18164 91337 18187
rect 91423 18164 91489 18187
rect 91103 18124 91112 18164
rect 91152 18124 91169 18164
rect 91255 18124 91276 18164
rect 91316 18124 91337 18164
rect 91423 18124 91440 18164
rect 91480 18124 91489 18164
rect 91103 18101 91169 18124
rect 91255 18101 91337 18124
rect 91423 18101 91489 18124
rect 91103 18082 91489 18101
rect 95103 18187 95489 18206
rect 95103 18164 95169 18187
rect 95255 18164 95337 18187
rect 95423 18164 95489 18187
rect 95103 18124 95112 18164
rect 95152 18124 95169 18164
rect 95255 18124 95276 18164
rect 95316 18124 95337 18164
rect 95423 18124 95440 18164
rect 95480 18124 95489 18164
rect 95103 18101 95169 18124
rect 95255 18101 95337 18124
rect 95423 18101 95489 18124
rect 95103 18082 95489 18101
rect 99103 18187 99489 18206
rect 99103 18164 99169 18187
rect 99255 18164 99337 18187
rect 99423 18164 99489 18187
rect 99103 18124 99112 18164
rect 99152 18124 99169 18164
rect 99255 18124 99276 18164
rect 99316 18124 99337 18164
rect 99423 18124 99440 18164
rect 99480 18124 99489 18164
rect 99103 18101 99169 18124
rect 99255 18101 99337 18124
rect 99423 18101 99489 18124
rect 99103 18082 99489 18101
rect 4343 17431 4729 17450
rect 4343 17408 4409 17431
rect 4495 17408 4577 17431
rect 4663 17408 4729 17431
rect 4343 17368 4352 17408
rect 4392 17368 4409 17408
rect 4495 17368 4516 17408
rect 4556 17368 4577 17408
rect 4663 17368 4680 17408
rect 4720 17368 4729 17408
rect 4343 17345 4409 17368
rect 4495 17345 4577 17368
rect 4663 17345 4729 17368
rect 4343 17326 4729 17345
rect 8343 17431 8729 17450
rect 8343 17408 8409 17431
rect 8495 17408 8577 17431
rect 8663 17408 8729 17431
rect 8343 17368 8352 17408
rect 8392 17368 8409 17408
rect 8495 17368 8516 17408
rect 8556 17368 8577 17408
rect 8663 17368 8680 17408
rect 8720 17368 8729 17408
rect 8343 17345 8409 17368
rect 8495 17345 8577 17368
rect 8663 17345 8729 17368
rect 8343 17326 8729 17345
rect 12343 17431 12729 17450
rect 12343 17408 12409 17431
rect 12495 17408 12577 17431
rect 12663 17408 12729 17431
rect 12343 17368 12352 17408
rect 12392 17368 12409 17408
rect 12495 17368 12516 17408
rect 12556 17368 12577 17408
rect 12663 17368 12680 17408
rect 12720 17368 12729 17408
rect 12343 17345 12409 17368
rect 12495 17345 12577 17368
rect 12663 17345 12729 17368
rect 12343 17326 12729 17345
rect 16343 17431 16729 17450
rect 16343 17408 16409 17431
rect 16495 17408 16577 17431
rect 16663 17408 16729 17431
rect 16343 17368 16352 17408
rect 16392 17368 16409 17408
rect 16495 17368 16516 17408
rect 16556 17368 16577 17408
rect 16663 17368 16680 17408
rect 16720 17368 16729 17408
rect 16343 17345 16409 17368
rect 16495 17345 16577 17368
rect 16663 17345 16729 17368
rect 16343 17326 16729 17345
rect 20343 17431 20729 17450
rect 20343 17408 20409 17431
rect 20495 17408 20577 17431
rect 20663 17408 20729 17431
rect 20343 17368 20352 17408
rect 20392 17368 20409 17408
rect 20495 17368 20516 17408
rect 20556 17368 20577 17408
rect 20663 17368 20680 17408
rect 20720 17368 20729 17408
rect 20343 17345 20409 17368
rect 20495 17345 20577 17368
rect 20663 17345 20729 17368
rect 20343 17326 20729 17345
rect 24343 17431 24729 17450
rect 24343 17408 24409 17431
rect 24495 17408 24577 17431
rect 24663 17408 24729 17431
rect 24343 17368 24352 17408
rect 24392 17368 24409 17408
rect 24495 17368 24516 17408
rect 24556 17368 24577 17408
rect 24663 17368 24680 17408
rect 24720 17368 24729 17408
rect 24343 17345 24409 17368
rect 24495 17345 24577 17368
rect 24663 17345 24729 17368
rect 24343 17326 24729 17345
rect 28343 17431 28729 17450
rect 28343 17408 28409 17431
rect 28495 17408 28577 17431
rect 28663 17408 28729 17431
rect 28343 17368 28352 17408
rect 28392 17368 28409 17408
rect 28495 17368 28516 17408
rect 28556 17368 28577 17408
rect 28663 17368 28680 17408
rect 28720 17368 28729 17408
rect 28343 17345 28409 17368
rect 28495 17345 28577 17368
rect 28663 17345 28729 17368
rect 28343 17326 28729 17345
rect 32343 17431 32729 17450
rect 32343 17408 32409 17431
rect 32495 17408 32577 17431
rect 32663 17408 32729 17431
rect 32343 17368 32352 17408
rect 32392 17368 32409 17408
rect 32495 17368 32516 17408
rect 32556 17368 32577 17408
rect 32663 17368 32680 17408
rect 32720 17368 32729 17408
rect 32343 17345 32409 17368
rect 32495 17345 32577 17368
rect 32663 17345 32729 17368
rect 32343 17326 32729 17345
rect 36343 17431 36729 17450
rect 36343 17408 36409 17431
rect 36495 17408 36577 17431
rect 36663 17408 36729 17431
rect 36343 17368 36352 17408
rect 36392 17368 36409 17408
rect 36495 17368 36516 17408
rect 36556 17368 36577 17408
rect 36663 17368 36680 17408
rect 36720 17368 36729 17408
rect 36343 17345 36409 17368
rect 36495 17345 36577 17368
rect 36663 17345 36729 17368
rect 36343 17326 36729 17345
rect 40343 17431 40729 17450
rect 40343 17408 40409 17431
rect 40495 17408 40577 17431
rect 40663 17408 40729 17431
rect 40343 17368 40352 17408
rect 40392 17368 40409 17408
rect 40495 17368 40516 17408
rect 40556 17368 40577 17408
rect 40663 17368 40680 17408
rect 40720 17368 40729 17408
rect 40343 17345 40409 17368
rect 40495 17345 40577 17368
rect 40663 17345 40729 17368
rect 40343 17326 40729 17345
rect 44343 17431 44729 17450
rect 44343 17408 44409 17431
rect 44495 17408 44577 17431
rect 44663 17408 44729 17431
rect 44343 17368 44352 17408
rect 44392 17368 44409 17408
rect 44495 17368 44516 17408
rect 44556 17368 44577 17408
rect 44663 17368 44680 17408
rect 44720 17368 44729 17408
rect 44343 17345 44409 17368
rect 44495 17345 44577 17368
rect 44663 17345 44729 17368
rect 44343 17326 44729 17345
rect 48343 17431 48729 17450
rect 48343 17408 48409 17431
rect 48495 17408 48577 17431
rect 48663 17408 48729 17431
rect 48343 17368 48352 17408
rect 48392 17368 48409 17408
rect 48495 17368 48516 17408
rect 48556 17368 48577 17408
rect 48663 17368 48680 17408
rect 48720 17368 48729 17408
rect 48343 17345 48409 17368
rect 48495 17345 48577 17368
rect 48663 17345 48729 17368
rect 48343 17326 48729 17345
rect 52343 17431 52729 17450
rect 52343 17408 52409 17431
rect 52495 17408 52577 17431
rect 52663 17408 52729 17431
rect 52343 17368 52352 17408
rect 52392 17368 52409 17408
rect 52495 17368 52516 17408
rect 52556 17368 52577 17408
rect 52663 17368 52680 17408
rect 52720 17368 52729 17408
rect 52343 17345 52409 17368
rect 52495 17345 52577 17368
rect 52663 17345 52729 17368
rect 52343 17326 52729 17345
rect 56343 17431 56729 17450
rect 56343 17408 56409 17431
rect 56495 17408 56577 17431
rect 56663 17408 56729 17431
rect 56343 17368 56352 17408
rect 56392 17368 56409 17408
rect 56495 17368 56516 17408
rect 56556 17368 56577 17408
rect 56663 17368 56680 17408
rect 56720 17368 56729 17408
rect 56343 17345 56409 17368
rect 56495 17345 56577 17368
rect 56663 17345 56729 17368
rect 56343 17326 56729 17345
rect 60343 17431 60729 17450
rect 60343 17408 60409 17431
rect 60495 17408 60577 17431
rect 60663 17408 60729 17431
rect 60343 17368 60352 17408
rect 60392 17368 60409 17408
rect 60495 17368 60516 17408
rect 60556 17368 60577 17408
rect 60663 17368 60680 17408
rect 60720 17368 60729 17408
rect 60343 17345 60409 17368
rect 60495 17345 60577 17368
rect 60663 17345 60729 17368
rect 60343 17326 60729 17345
rect 64343 17431 64729 17450
rect 64343 17408 64409 17431
rect 64495 17408 64577 17431
rect 64663 17408 64729 17431
rect 64343 17368 64352 17408
rect 64392 17368 64409 17408
rect 64495 17368 64516 17408
rect 64556 17368 64577 17408
rect 64663 17368 64680 17408
rect 64720 17368 64729 17408
rect 64343 17345 64409 17368
rect 64495 17345 64577 17368
rect 64663 17345 64729 17368
rect 64343 17326 64729 17345
rect 68343 17431 68729 17450
rect 68343 17408 68409 17431
rect 68495 17408 68577 17431
rect 68663 17408 68729 17431
rect 68343 17368 68352 17408
rect 68392 17368 68409 17408
rect 68495 17368 68516 17408
rect 68556 17368 68577 17408
rect 68663 17368 68680 17408
rect 68720 17368 68729 17408
rect 68343 17345 68409 17368
rect 68495 17345 68577 17368
rect 68663 17345 68729 17368
rect 68343 17326 68729 17345
rect 72343 17431 72729 17450
rect 72343 17408 72409 17431
rect 72495 17408 72577 17431
rect 72663 17408 72729 17431
rect 72343 17368 72352 17408
rect 72392 17368 72409 17408
rect 72495 17368 72516 17408
rect 72556 17368 72577 17408
rect 72663 17368 72680 17408
rect 72720 17368 72729 17408
rect 72343 17345 72409 17368
rect 72495 17345 72577 17368
rect 72663 17345 72729 17368
rect 72343 17326 72729 17345
rect 76343 17431 76729 17450
rect 76343 17408 76409 17431
rect 76495 17408 76577 17431
rect 76663 17408 76729 17431
rect 76343 17368 76352 17408
rect 76392 17368 76409 17408
rect 76495 17368 76516 17408
rect 76556 17368 76577 17408
rect 76663 17368 76680 17408
rect 76720 17368 76729 17408
rect 76343 17345 76409 17368
rect 76495 17345 76577 17368
rect 76663 17345 76729 17368
rect 76343 17326 76729 17345
rect 80343 17431 80729 17450
rect 80343 17408 80409 17431
rect 80495 17408 80577 17431
rect 80663 17408 80729 17431
rect 80343 17368 80352 17408
rect 80392 17368 80409 17408
rect 80495 17368 80516 17408
rect 80556 17368 80577 17408
rect 80663 17368 80680 17408
rect 80720 17368 80729 17408
rect 80343 17345 80409 17368
rect 80495 17345 80577 17368
rect 80663 17345 80729 17368
rect 80343 17326 80729 17345
rect 84343 17431 84729 17450
rect 84343 17408 84409 17431
rect 84495 17408 84577 17431
rect 84663 17408 84729 17431
rect 84343 17368 84352 17408
rect 84392 17368 84409 17408
rect 84495 17368 84516 17408
rect 84556 17368 84577 17408
rect 84663 17368 84680 17408
rect 84720 17368 84729 17408
rect 84343 17345 84409 17368
rect 84495 17345 84577 17368
rect 84663 17345 84729 17368
rect 84343 17326 84729 17345
rect 88343 17431 88729 17450
rect 88343 17408 88409 17431
rect 88495 17408 88577 17431
rect 88663 17408 88729 17431
rect 88343 17368 88352 17408
rect 88392 17368 88409 17408
rect 88495 17368 88516 17408
rect 88556 17368 88577 17408
rect 88663 17368 88680 17408
rect 88720 17368 88729 17408
rect 88343 17345 88409 17368
rect 88495 17345 88577 17368
rect 88663 17345 88729 17368
rect 88343 17326 88729 17345
rect 92343 17431 92729 17450
rect 92343 17408 92409 17431
rect 92495 17408 92577 17431
rect 92663 17408 92729 17431
rect 92343 17368 92352 17408
rect 92392 17368 92409 17408
rect 92495 17368 92516 17408
rect 92556 17368 92577 17408
rect 92663 17368 92680 17408
rect 92720 17368 92729 17408
rect 92343 17345 92409 17368
rect 92495 17345 92577 17368
rect 92663 17345 92729 17368
rect 92343 17326 92729 17345
rect 96343 17431 96729 17450
rect 96343 17408 96409 17431
rect 96495 17408 96577 17431
rect 96663 17408 96729 17431
rect 96343 17368 96352 17408
rect 96392 17368 96409 17408
rect 96495 17368 96516 17408
rect 96556 17368 96577 17408
rect 96663 17368 96680 17408
rect 96720 17368 96729 17408
rect 96343 17345 96409 17368
rect 96495 17345 96577 17368
rect 96663 17345 96729 17368
rect 96343 17326 96729 17345
rect 3103 16675 3489 16694
rect 3103 16652 3169 16675
rect 3255 16652 3337 16675
rect 3423 16652 3489 16675
rect 3103 16612 3112 16652
rect 3152 16612 3169 16652
rect 3255 16612 3276 16652
rect 3316 16612 3337 16652
rect 3423 16612 3440 16652
rect 3480 16612 3489 16652
rect 3103 16589 3169 16612
rect 3255 16589 3337 16612
rect 3423 16589 3489 16612
rect 3103 16570 3489 16589
rect 7103 16675 7489 16694
rect 7103 16652 7169 16675
rect 7255 16652 7337 16675
rect 7423 16652 7489 16675
rect 7103 16612 7112 16652
rect 7152 16612 7169 16652
rect 7255 16612 7276 16652
rect 7316 16612 7337 16652
rect 7423 16612 7440 16652
rect 7480 16612 7489 16652
rect 7103 16589 7169 16612
rect 7255 16589 7337 16612
rect 7423 16589 7489 16612
rect 7103 16570 7489 16589
rect 11103 16675 11489 16694
rect 11103 16652 11169 16675
rect 11255 16652 11337 16675
rect 11423 16652 11489 16675
rect 11103 16612 11112 16652
rect 11152 16612 11169 16652
rect 11255 16612 11276 16652
rect 11316 16612 11337 16652
rect 11423 16612 11440 16652
rect 11480 16612 11489 16652
rect 11103 16589 11169 16612
rect 11255 16589 11337 16612
rect 11423 16589 11489 16612
rect 11103 16570 11489 16589
rect 15103 16675 15489 16694
rect 15103 16652 15169 16675
rect 15255 16652 15337 16675
rect 15423 16652 15489 16675
rect 15103 16612 15112 16652
rect 15152 16612 15169 16652
rect 15255 16612 15276 16652
rect 15316 16612 15337 16652
rect 15423 16612 15440 16652
rect 15480 16612 15489 16652
rect 15103 16589 15169 16612
rect 15255 16589 15337 16612
rect 15423 16589 15489 16612
rect 15103 16570 15489 16589
rect 19103 16675 19489 16694
rect 19103 16652 19169 16675
rect 19255 16652 19337 16675
rect 19423 16652 19489 16675
rect 19103 16612 19112 16652
rect 19152 16612 19169 16652
rect 19255 16612 19276 16652
rect 19316 16612 19337 16652
rect 19423 16612 19440 16652
rect 19480 16612 19489 16652
rect 19103 16589 19169 16612
rect 19255 16589 19337 16612
rect 19423 16589 19489 16612
rect 19103 16570 19489 16589
rect 23103 16675 23489 16694
rect 23103 16652 23169 16675
rect 23255 16652 23337 16675
rect 23423 16652 23489 16675
rect 23103 16612 23112 16652
rect 23152 16612 23169 16652
rect 23255 16612 23276 16652
rect 23316 16612 23337 16652
rect 23423 16612 23440 16652
rect 23480 16612 23489 16652
rect 23103 16589 23169 16612
rect 23255 16589 23337 16612
rect 23423 16589 23489 16612
rect 23103 16570 23489 16589
rect 27103 16675 27489 16694
rect 27103 16652 27169 16675
rect 27255 16652 27337 16675
rect 27423 16652 27489 16675
rect 27103 16612 27112 16652
rect 27152 16612 27169 16652
rect 27255 16612 27276 16652
rect 27316 16612 27337 16652
rect 27423 16612 27440 16652
rect 27480 16612 27489 16652
rect 27103 16589 27169 16612
rect 27255 16589 27337 16612
rect 27423 16589 27489 16612
rect 27103 16570 27489 16589
rect 31103 16675 31489 16694
rect 31103 16652 31169 16675
rect 31255 16652 31337 16675
rect 31423 16652 31489 16675
rect 31103 16612 31112 16652
rect 31152 16612 31169 16652
rect 31255 16612 31276 16652
rect 31316 16612 31337 16652
rect 31423 16612 31440 16652
rect 31480 16612 31489 16652
rect 31103 16589 31169 16612
rect 31255 16589 31337 16612
rect 31423 16589 31489 16612
rect 31103 16570 31489 16589
rect 35103 16675 35489 16694
rect 35103 16652 35169 16675
rect 35255 16652 35337 16675
rect 35423 16652 35489 16675
rect 35103 16612 35112 16652
rect 35152 16612 35169 16652
rect 35255 16612 35276 16652
rect 35316 16612 35337 16652
rect 35423 16612 35440 16652
rect 35480 16612 35489 16652
rect 35103 16589 35169 16612
rect 35255 16589 35337 16612
rect 35423 16589 35489 16612
rect 35103 16570 35489 16589
rect 39103 16675 39489 16694
rect 39103 16652 39169 16675
rect 39255 16652 39337 16675
rect 39423 16652 39489 16675
rect 39103 16612 39112 16652
rect 39152 16612 39169 16652
rect 39255 16612 39276 16652
rect 39316 16612 39337 16652
rect 39423 16612 39440 16652
rect 39480 16612 39489 16652
rect 39103 16589 39169 16612
rect 39255 16589 39337 16612
rect 39423 16589 39489 16612
rect 39103 16570 39489 16589
rect 43103 16675 43489 16694
rect 43103 16652 43169 16675
rect 43255 16652 43337 16675
rect 43423 16652 43489 16675
rect 43103 16612 43112 16652
rect 43152 16612 43169 16652
rect 43255 16612 43276 16652
rect 43316 16612 43337 16652
rect 43423 16612 43440 16652
rect 43480 16612 43489 16652
rect 43103 16589 43169 16612
rect 43255 16589 43337 16612
rect 43423 16589 43489 16612
rect 43103 16570 43489 16589
rect 47103 16675 47489 16694
rect 47103 16652 47169 16675
rect 47255 16652 47337 16675
rect 47423 16652 47489 16675
rect 47103 16612 47112 16652
rect 47152 16612 47169 16652
rect 47255 16612 47276 16652
rect 47316 16612 47337 16652
rect 47423 16612 47440 16652
rect 47480 16612 47489 16652
rect 47103 16589 47169 16612
rect 47255 16589 47337 16612
rect 47423 16589 47489 16612
rect 47103 16570 47489 16589
rect 51103 16675 51489 16694
rect 51103 16652 51169 16675
rect 51255 16652 51337 16675
rect 51423 16652 51489 16675
rect 51103 16612 51112 16652
rect 51152 16612 51169 16652
rect 51255 16612 51276 16652
rect 51316 16612 51337 16652
rect 51423 16612 51440 16652
rect 51480 16612 51489 16652
rect 51103 16589 51169 16612
rect 51255 16589 51337 16612
rect 51423 16589 51489 16612
rect 51103 16570 51489 16589
rect 55103 16675 55489 16694
rect 55103 16652 55169 16675
rect 55255 16652 55337 16675
rect 55423 16652 55489 16675
rect 55103 16612 55112 16652
rect 55152 16612 55169 16652
rect 55255 16612 55276 16652
rect 55316 16612 55337 16652
rect 55423 16612 55440 16652
rect 55480 16612 55489 16652
rect 55103 16589 55169 16612
rect 55255 16589 55337 16612
rect 55423 16589 55489 16612
rect 55103 16570 55489 16589
rect 59103 16675 59489 16694
rect 59103 16652 59169 16675
rect 59255 16652 59337 16675
rect 59423 16652 59489 16675
rect 59103 16612 59112 16652
rect 59152 16612 59169 16652
rect 59255 16612 59276 16652
rect 59316 16612 59337 16652
rect 59423 16612 59440 16652
rect 59480 16612 59489 16652
rect 59103 16589 59169 16612
rect 59255 16589 59337 16612
rect 59423 16589 59489 16612
rect 59103 16570 59489 16589
rect 63103 16675 63489 16694
rect 63103 16652 63169 16675
rect 63255 16652 63337 16675
rect 63423 16652 63489 16675
rect 63103 16612 63112 16652
rect 63152 16612 63169 16652
rect 63255 16612 63276 16652
rect 63316 16612 63337 16652
rect 63423 16612 63440 16652
rect 63480 16612 63489 16652
rect 63103 16589 63169 16612
rect 63255 16589 63337 16612
rect 63423 16589 63489 16612
rect 63103 16570 63489 16589
rect 67103 16675 67489 16694
rect 67103 16652 67169 16675
rect 67255 16652 67337 16675
rect 67423 16652 67489 16675
rect 67103 16612 67112 16652
rect 67152 16612 67169 16652
rect 67255 16612 67276 16652
rect 67316 16612 67337 16652
rect 67423 16612 67440 16652
rect 67480 16612 67489 16652
rect 67103 16589 67169 16612
rect 67255 16589 67337 16612
rect 67423 16589 67489 16612
rect 67103 16570 67489 16589
rect 4343 15919 4729 15938
rect 4343 15896 4409 15919
rect 4495 15896 4577 15919
rect 4663 15896 4729 15919
rect 4343 15856 4352 15896
rect 4392 15856 4409 15896
rect 4495 15856 4516 15896
rect 4556 15856 4577 15896
rect 4663 15856 4680 15896
rect 4720 15856 4729 15896
rect 4343 15833 4409 15856
rect 4495 15833 4577 15856
rect 4663 15833 4729 15856
rect 4343 15814 4729 15833
rect 8343 15919 8729 15938
rect 8343 15896 8409 15919
rect 8495 15896 8577 15919
rect 8663 15896 8729 15919
rect 8343 15856 8352 15896
rect 8392 15856 8409 15896
rect 8495 15856 8516 15896
rect 8556 15856 8577 15896
rect 8663 15856 8680 15896
rect 8720 15856 8729 15896
rect 8343 15833 8409 15856
rect 8495 15833 8577 15856
rect 8663 15833 8729 15856
rect 8343 15814 8729 15833
rect 12343 15919 12729 15938
rect 12343 15896 12409 15919
rect 12495 15896 12577 15919
rect 12663 15896 12729 15919
rect 12343 15856 12352 15896
rect 12392 15856 12409 15896
rect 12495 15856 12516 15896
rect 12556 15856 12577 15896
rect 12663 15856 12680 15896
rect 12720 15856 12729 15896
rect 12343 15833 12409 15856
rect 12495 15833 12577 15856
rect 12663 15833 12729 15856
rect 12343 15814 12729 15833
rect 16343 15919 16729 15938
rect 16343 15896 16409 15919
rect 16495 15896 16577 15919
rect 16663 15896 16729 15919
rect 16343 15856 16352 15896
rect 16392 15856 16409 15896
rect 16495 15856 16516 15896
rect 16556 15856 16577 15896
rect 16663 15856 16680 15896
rect 16720 15856 16729 15896
rect 16343 15833 16409 15856
rect 16495 15833 16577 15856
rect 16663 15833 16729 15856
rect 16343 15814 16729 15833
rect 20343 15919 20729 15938
rect 20343 15896 20409 15919
rect 20495 15896 20577 15919
rect 20663 15896 20729 15919
rect 20343 15856 20352 15896
rect 20392 15856 20409 15896
rect 20495 15856 20516 15896
rect 20556 15856 20577 15896
rect 20663 15856 20680 15896
rect 20720 15856 20729 15896
rect 20343 15833 20409 15856
rect 20495 15833 20577 15856
rect 20663 15833 20729 15856
rect 20343 15814 20729 15833
rect 24343 15919 24729 15938
rect 24343 15896 24409 15919
rect 24495 15896 24577 15919
rect 24663 15896 24729 15919
rect 24343 15856 24352 15896
rect 24392 15856 24409 15896
rect 24495 15856 24516 15896
rect 24556 15856 24577 15896
rect 24663 15856 24680 15896
rect 24720 15856 24729 15896
rect 24343 15833 24409 15856
rect 24495 15833 24577 15856
rect 24663 15833 24729 15856
rect 24343 15814 24729 15833
rect 28343 15919 28729 15938
rect 28343 15896 28409 15919
rect 28495 15896 28577 15919
rect 28663 15896 28729 15919
rect 28343 15856 28352 15896
rect 28392 15856 28409 15896
rect 28495 15856 28516 15896
rect 28556 15856 28577 15896
rect 28663 15856 28680 15896
rect 28720 15856 28729 15896
rect 28343 15833 28409 15856
rect 28495 15833 28577 15856
rect 28663 15833 28729 15856
rect 28343 15814 28729 15833
rect 32343 15919 32729 15938
rect 32343 15896 32409 15919
rect 32495 15896 32577 15919
rect 32663 15896 32729 15919
rect 32343 15856 32352 15896
rect 32392 15856 32409 15896
rect 32495 15856 32516 15896
rect 32556 15856 32577 15896
rect 32663 15856 32680 15896
rect 32720 15856 32729 15896
rect 32343 15833 32409 15856
rect 32495 15833 32577 15856
rect 32663 15833 32729 15856
rect 32343 15814 32729 15833
rect 36343 15919 36729 15938
rect 36343 15896 36409 15919
rect 36495 15896 36577 15919
rect 36663 15896 36729 15919
rect 36343 15856 36352 15896
rect 36392 15856 36409 15896
rect 36495 15856 36516 15896
rect 36556 15856 36577 15896
rect 36663 15856 36680 15896
rect 36720 15856 36729 15896
rect 36343 15833 36409 15856
rect 36495 15833 36577 15856
rect 36663 15833 36729 15856
rect 36343 15814 36729 15833
rect 40343 15919 40729 15938
rect 40343 15896 40409 15919
rect 40495 15896 40577 15919
rect 40663 15896 40729 15919
rect 40343 15856 40352 15896
rect 40392 15856 40409 15896
rect 40495 15856 40516 15896
rect 40556 15856 40577 15896
rect 40663 15856 40680 15896
rect 40720 15856 40729 15896
rect 40343 15833 40409 15856
rect 40495 15833 40577 15856
rect 40663 15833 40729 15856
rect 40343 15814 40729 15833
rect 44343 15919 44729 15938
rect 44343 15896 44409 15919
rect 44495 15896 44577 15919
rect 44663 15896 44729 15919
rect 44343 15856 44352 15896
rect 44392 15856 44409 15896
rect 44495 15856 44516 15896
rect 44556 15856 44577 15896
rect 44663 15856 44680 15896
rect 44720 15856 44729 15896
rect 44343 15833 44409 15856
rect 44495 15833 44577 15856
rect 44663 15833 44729 15856
rect 44343 15814 44729 15833
rect 48343 15919 48729 15938
rect 48343 15896 48409 15919
rect 48495 15896 48577 15919
rect 48663 15896 48729 15919
rect 48343 15856 48352 15896
rect 48392 15856 48409 15896
rect 48495 15856 48516 15896
rect 48556 15856 48577 15896
rect 48663 15856 48680 15896
rect 48720 15856 48729 15896
rect 48343 15833 48409 15856
rect 48495 15833 48577 15856
rect 48663 15833 48729 15856
rect 48343 15814 48729 15833
rect 52343 15919 52729 15938
rect 52343 15896 52409 15919
rect 52495 15896 52577 15919
rect 52663 15896 52729 15919
rect 52343 15856 52352 15896
rect 52392 15856 52409 15896
rect 52495 15856 52516 15896
rect 52556 15856 52577 15896
rect 52663 15856 52680 15896
rect 52720 15856 52729 15896
rect 52343 15833 52409 15856
rect 52495 15833 52577 15856
rect 52663 15833 52729 15856
rect 52343 15814 52729 15833
rect 56343 15919 56729 15938
rect 56343 15896 56409 15919
rect 56495 15896 56577 15919
rect 56663 15896 56729 15919
rect 56343 15856 56352 15896
rect 56392 15856 56409 15896
rect 56495 15856 56516 15896
rect 56556 15856 56577 15896
rect 56663 15856 56680 15896
rect 56720 15856 56729 15896
rect 56343 15833 56409 15856
rect 56495 15833 56577 15856
rect 56663 15833 56729 15856
rect 56343 15814 56729 15833
rect 60343 15919 60729 15938
rect 60343 15896 60409 15919
rect 60495 15896 60577 15919
rect 60663 15896 60729 15919
rect 60343 15856 60352 15896
rect 60392 15856 60409 15896
rect 60495 15856 60516 15896
rect 60556 15856 60577 15896
rect 60663 15856 60680 15896
rect 60720 15856 60729 15896
rect 60343 15833 60409 15856
rect 60495 15833 60577 15856
rect 60663 15833 60729 15856
rect 60343 15814 60729 15833
rect 64343 15919 64729 15938
rect 64343 15896 64409 15919
rect 64495 15896 64577 15919
rect 64663 15896 64729 15919
rect 64343 15856 64352 15896
rect 64392 15856 64409 15896
rect 64495 15856 64516 15896
rect 64556 15856 64577 15896
rect 64663 15856 64680 15896
rect 64720 15856 64729 15896
rect 64343 15833 64409 15856
rect 64495 15833 64577 15856
rect 64663 15833 64729 15856
rect 64343 15814 64729 15833
rect 68343 15919 68729 15938
rect 68343 15896 68409 15919
rect 68495 15896 68577 15919
rect 68663 15896 68729 15919
rect 68343 15856 68352 15896
rect 68392 15856 68409 15896
rect 68495 15856 68516 15896
rect 68556 15856 68577 15896
rect 68663 15856 68680 15896
rect 68720 15856 68729 15896
rect 68343 15833 68409 15856
rect 68495 15833 68577 15856
rect 68663 15833 68729 15856
rect 68343 15814 68729 15833
rect 3103 15163 3489 15182
rect 3103 15140 3169 15163
rect 3255 15140 3337 15163
rect 3423 15140 3489 15163
rect 3103 15100 3112 15140
rect 3152 15100 3169 15140
rect 3255 15100 3276 15140
rect 3316 15100 3337 15140
rect 3423 15100 3440 15140
rect 3480 15100 3489 15140
rect 3103 15077 3169 15100
rect 3255 15077 3337 15100
rect 3423 15077 3489 15100
rect 3103 15058 3489 15077
rect 7103 15163 7489 15182
rect 7103 15140 7169 15163
rect 7255 15140 7337 15163
rect 7423 15140 7489 15163
rect 7103 15100 7112 15140
rect 7152 15100 7169 15140
rect 7255 15100 7276 15140
rect 7316 15100 7337 15140
rect 7423 15100 7440 15140
rect 7480 15100 7489 15140
rect 7103 15077 7169 15100
rect 7255 15077 7337 15100
rect 7423 15077 7489 15100
rect 7103 15058 7489 15077
rect 11103 15163 11489 15182
rect 11103 15140 11169 15163
rect 11255 15140 11337 15163
rect 11423 15140 11489 15163
rect 11103 15100 11112 15140
rect 11152 15100 11169 15140
rect 11255 15100 11276 15140
rect 11316 15100 11337 15140
rect 11423 15100 11440 15140
rect 11480 15100 11489 15140
rect 11103 15077 11169 15100
rect 11255 15077 11337 15100
rect 11423 15077 11489 15100
rect 11103 15058 11489 15077
rect 15103 15163 15489 15182
rect 15103 15140 15169 15163
rect 15255 15140 15337 15163
rect 15423 15140 15489 15163
rect 15103 15100 15112 15140
rect 15152 15100 15169 15140
rect 15255 15100 15276 15140
rect 15316 15100 15337 15140
rect 15423 15100 15440 15140
rect 15480 15100 15489 15140
rect 15103 15077 15169 15100
rect 15255 15077 15337 15100
rect 15423 15077 15489 15100
rect 15103 15058 15489 15077
rect 19103 15163 19489 15182
rect 19103 15140 19169 15163
rect 19255 15140 19337 15163
rect 19423 15140 19489 15163
rect 19103 15100 19112 15140
rect 19152 15100 19169 15140
rect 19255 15100 19276 15140
rect 19316 15100 19337 15140
rect 19423 15100 19440 15140
rect 19480 15100 19489 15140
rect 19103 15077 19169 15100
rect 19255 15077 19337 15100
rect 19423 15077 19489 15100
rect 19103 15058 19489 15077
rect 23103 15163 23489 15182
rect 23103 15140 23169 15163
rect 23255 15140 23337 15163
rect 23423 15140 23489 15163
rect 23103 15100 23112 15140
rect 23152 15100 23169 15140
rect 23255 15100 23276 15140
rect 23316 15100 23337 15140
rect 23423 15100 23440 15140
rect 23480 15100 23489 15140
rect 23103 15077 23169 15100
rect 23255 15077 23337 15100
rect 23423 15077 23489 15100
rect 23103 15058 23489 15077
rect 27103 15163 27489 15182
rect 27103 15140 27169 15163
rect 27255 15140 27337 15163
rect 27423 15140 27489 15163
rect 27103 15100 27112 15140
rect 27152 15100 27169 15140
rect 27255 15100 27276 15140
rect 27316 15100 27337 15140
rect 27423 15100 27440 15140
rect 27480 15100 27489 15140
rect 27103 15077 27169 15100
rect 27255 15077 27337 15100
rect 27423 15077 27489 15100
rect 27103 15058 27489 15077
rect 31103 15163 31489 15182
rect 31103 15140 31169 15163
rect 31255 15140 31337 15163
rect 31423 15140 31489 15163
rect 31103 15100 31112 15140
rect 31152 15100 31169 15140
rect 31255 15100 31276 15140
rect 31316 15100 31337 15140
rect 31423 15100 31440 15140
rect 31480 15100 31489 15140
rect 31103 15077 31169 15100
rect 31255 15077 31337 15100
rect 31423 15077 31489 15100
rect 31103 15058 31489 15077
rect 35103 15163 35489 15182
rect 35103 15140 35169 15163
rect 35255 15140 35337 15163
rect 35423 15140 35489 15163
rect 35103 15100 35112 15140
rect 35152 15100 35169 15140
rect 35255 15100 35276 15140
rect 35316 15100 35337 15140
rect 35423 15100 35440 15140
rect 35480 15100 35489 15140
rect 35103 15077 35169 15100
rect 35255 15077 35337 15100
rect 35423 15077 35489 15100
rect 35103 15058 35489 15077
rect 39103 15163 39489 15182
rect 39103 15140 39169 15163
rect 39255 15140 39337 15163
rect 39423 15140 39489 15163
rect 39103 15100 39112 15140
rect 39152 15100 39169 15140
rect 39255 15100 39276 15140
rect 39316 15100 39337 15140
rect 39423 15100 39440 15140
rect 39480 15100 39489 15140
rect 39103 15077 39169 15100
rect 39255 15077 39337 15100
rect 39423 15077 39489 15100
rect 39103 15058 39489 15077
rect 43103 15163 43489 15182
rect 43103 15140 43169 15163
rect 43255 15140 43337 15163
rect 43423 15140 43489 15163
rect 43103 15100 43112 15140
rect 43152 15100 43169 15140
rect 43255 15100 43276 15140
rect 43316 15100 43337 15140
rect 43423 15100 43440 15140
rect 43480 15100 43489 15140
rect 43103 15077 43169 15100
rect 43255 15077 43337 15100
rect 43423 15077 43489 15100
rect 43103 15058 43489 15077
rect 47103 15163 47489 15182
rect 47103 15140 47169 15163
rect 47255 15140 47337 15163
rect 47423 15140 47489 15163
rect 47103 15100 47112 15140
rect 47152 15100 47169 15140
rect 47255 15100 47276 15140
rect 47316 15100 47337 15140
rect 47423 15100 47440 15140
rect 47480 15100 47489 15140
rect 47103 15077 47169 15100
rect 47255 15077 47337 15100
rect 47423 15077 47489 15100
rect 47103 15058 47489 15077
rect 51103 15163 51489 15182
rect 51103 15140 51169 15163
rect 51255 15140 51337 15163
rect 51423 15140 51489 15163
rect 51103 15100 51112 15140
rect 51152 15100 51169 15140
rect 51255 15100 51276 15140
rect 51316 15100 51337 15140
rect 51423 15100 51440 15140
rect 51480 15100 51489 15140
rect 51103 15077 51169 15100
rect 51255 15077 51337 15100
rect 51423 15077 51489 15100
rect 51103 15058 51489 15077
rect 55103 15163 55489 15182
rect 55103 15140 55169 15163
rect 55255 15140 55337 15163
rect 55423 15140 55489 15163
rect 55103 15100 55112 15140
rect 55152 15100 55169 15140
rect 55255 15100 55276 15140
rect 55316 15100 55337 15140
rect 55423 15100 55440 15140
rect 55480 15100 55489 15140
rect 55103 15077 55169 15100
rect 55255 15077 55337 15100
rect 55423 15077 55489 15100
rect 55103 15058 55489 15077
rect 59103 15163 59489 15182
rect 59103 15140 59169 15163
rect 59255 15140 59337 15163
rect 59423 15140 59489 15163
rect 59103 15100 59112 15140
rect 59152 15100 59169 15140
rect 59255 15100 59276 15140
rect 59316 15100 59337 15140
rect 59423 15100 59440 15140
rect 59480 15100 59489 15140
rect 59103 15077 59169 15100
rect 59255 15077 59337 15100
rect 59423 15077 59489 15100
rect 59103 15058 59489 15077
rect 63103 15163 63489 15182
rect 63103 15140 63169 15163
rect 63255 15140 63337 15163
rect 63423 15140 63489 15163
rect 63103 15100 63112 15140
rect 63152 15100 63169 15140
rect 63255 15100 63276 15140
rect 63316 15100 63337 15140
rect 63423 15100 63440 15140
rect 63480 15100 63489 15140
rect 63103 15077 63169 15100
rect 63255 15077 63337 15100
rect 63423 15077 63489 15100
rect 63103 15058 63489 15077
rect 67103 15163 67489 15182
rect 67103 15140 67169 15163
rect 67255 15140 67337 15163
rect 67423 15140 67489 15163
rect 67103 15100 67112 15140
rect 67152 15100 67169 15140
rect 67255 15100 67276 15140
rect 67316 15100 67337 15140
rect 67423 15100 67440 15140
rect 67480 15100 67489 15140
rect 67103 15077 67169 15100
rect 67255 15077 67337 15100
rect 67423 15077 67489 15100
rect 67103 15058 67489 15077
rect 72316 15122 72756 15252
rect 72316 15036 72409 15122
rect 72495 15036 72577 15122
rect 72663 15036 72756 15122
rect 72316 14954 72756 15036
rect 72316 14868 72409 14954
rect 72495 14868 72577 14954
rect 72663 14868 72756 14954
rect 72316 14786 72756 14868
rect 72316 14700 72409 14786
rect 72495 14700 72577 14786
rect 72663 14700 72756 14786
rect 72316 14618 72756 14700
rect 72316 14532 72409 14618
rect 72495 14532 72577 14618
rect 72663 14532 72756 14618
rect 72316 14450 72756 14532
rect 4343 14407 4729 14426
rect 4343 14384 4409 14407
rect 4495 14384 4577 14407
rect 4663 14384 4729 14407
rect 4343 14344 4352 14384
rect 4392 14344 4409 14384
rect 4495 14344 4516 14384
rect 4556 14344 4577 14384
rect 4663 14344 4680 14384
rect 4720 14344 4729 14384
rect 4343 14321 4409 14344
rect 4495 14321 4577 14344
rect 4663 14321 4729 14344
rect 4343 14302 4729 14321
rect 8343 14407 8729 14426
rect 8343 14384 8409 14407
rect 8495 14384 8577 14407
rect 8663 14384 8729 14407
rect 8343 14344 8352 14384
rect 8392 14344 8409 14384
rect 8495 14344 8516 14384
rect 8556 14344 8577 14384
rect 8663 14344 8680 14384
rect 8720 14344 8729 14384
rect 8343 14321 8409 14344
rect 8495 14321 8577 14344
rect 8663 14321 8729 14344
rect 8343 14302 8729 14321
rect 12343 14407 12729 14426
rect 12343 14384 12409 14407
rect 12495 14384 12577 14407
rect 12663 14384 12729 14407
rect 12343 14344 12352 14384
rect 12392 14344 12409 14384
rect 12495 14344 12516 14384
rect 12556 14344 12577 14384
rect 12663 14344 12680 14384
rect 12720 14344 12729 14384
rect 12343 14321 12409 14344
rect 12495 14321 12577 14344
rect 12663 14321 12729 14344
rect 12343 14302 12729 14321
rect 16343 14407 16729 14426
rect 16343 14384 16409 14407
rect 16495 14384 16577 14407
rect 16663 14384 16729 14407
rect 16343 14344 16352 14384
rect 16392 14344 16409 14384
rect 16495 14344 16516 14384
rect 16556 14344 16577 14384
rect 16663 14344 16680 14384
rect 16720 14344 16729 14384
rect 16343 14321 16409 14344
rect 16495 14321 16577 14344
rect 16663 14321 16729 14344
rect 16343 14302 16729 14321
rect 20343 14407 20729 14426
rect 20343 14384 20409 14407
rect 20495 14384 20577 14407
rect 20663 14384 20729 14407
rect 20343 14344 20352 14384
rect 20392 14344 20409 14384
rect 20495 14344 20516 14384
rect 20556 14344 20577 14384
rect 20663 14344 20680 14384
rect 20720 14344 20729 14384
rect 20343 14321 20409 14344
rect 20495 14321 20577 14344
rect 20663 14321 20729 14344
rect 20343 14302 20729 14321
rect 24343 14407 24729 14426
rect 24343 14384 24409 14407
rect 24495 14384 24577 14407
rect 24663 14384 24729 14407
rect 24343 14344 24352 14384
rect 24392 14344 24409 14384
rect 24495 14344 24516 14384
rect 24556 14344 24577 14384
rect 24663 14344 24680 14384
rect 24720 14344 24729 14384
rect 24343 14321 24409 14344
rect 24495 14321 24577 14344
rect 24663 14321 24729 14344
rect 24343 14302 24729 14321
rect 28343 14407 28729 14426
rect 28343 14384 28409 14407
rect 28495 14384 28577 14407
rect 28663 14384 28729 14407
rect 28343 14344 28352 14384
rect 28392 14344 28409 14384
rect 28495 14344 28516 14384
rect 28556 14344 28577 14384
rect 28663 14344 28680 14384
rect 28720 14344 28729 14384
rect 28343 14321 28409 14344
rect 28495 14321 28577 14344
rect 28663 14321 28729 14344
rect 28343 14302 28729 14321
rect 32343 14407 32729 14426
rect 32343 14384 32409 14407
rect 32495 14384 32577 14407
rect 32663 14384 32729 14407
rect 32343 14344 32352 14384
rect 32392 14344 32409 14384
rect 32495 14344 32516 14384
rect 32556 14344 32577 14384
rect 32663 14344 32680 14384
rect 32720 14344 32729 14384
rect 32343 14321 32409 14344
rect 32495 14321 32577 14344
rect 32663 14321 32729 14344
rect 32343 14302 32729 14321
rect 36343 14407 36729 14426
rect 36343 14384 36409 14407
rect 36495 14384 36577 14407
rect 36663 14384 36729 14407
rect 36343 14344 36352 14384
rect 36392 14344 36409 14384
rect 36495 14344 36516 14384
rect 36556 14344 36577 14384
rect 36663 14344 36680 14384
rect 36720 14344 36729 14384
rect 36343 14321 36409 14344
rect 36495 14321 36577 14344
rect 36663 14321 36729 14344
rect 36343 14302 36729 14321
rect 40343 14407 40729 14426
rect 40343 14384 40409 14407
rect 40495 14384 40577 14407
rect 40663 14384 40729 14407
rect 40343 14344 40352 14384
rect 40392 14344 40409 14384
rect 40495 14344 40516 14384
rect 40556 14344 40577 14384
rect 40663 14344 40680 14384
rect 40720 14344 40729 14384
rect 40343 14321 40409 14344
rect 40495 14321 40577 14344
rect 40663 14321 40729 14344
rect 40343 14302 40729 14321
rect 44343 14407 44729 14426
rect 44343 14384 44409 14407
rect 44495 14384 44577 14407
rect 44663 14384 44729 14407
rect 44343 14344 44352 14384
rect 44392 14344 44409 14384
rect 44495 14344 44516 14384
rect 44556 14344 44577 14384
rect 44663 14344 44680 14384
rect 44720 14344 44729 14384
rect 44343 14321 44409 14344
rect 44495 14321 44577 14344
rect 44663 14321 44729 14344
rect 44343 14302 44729 14321
rect 48343 14407 48729 14426
rect 48343 14384 48409 14407
rect 48495 14384 48577 14407
rect 48663 14384 48729 14407
rect 48343 14344 48352 14384
rect 48392 14344 48409 14384
rect 48495 14344 48516 14384
rect 48556 14344 48577 14384
rect 48663 14344 48680 14384
rect 48720 14344 48729 14384
rect 48343 14321 48409 14344
rect 48495 14321 48577 14344
rect 48663 14321 48729 14344
rect 48343 14302 48729 14321
rect 52343 14407 52729 14426
rect 52343 14384 52409 14407
rect 52495 14384 52577 14407
rect 52663 14384 52729 14407
rect 52343 14344 52352 14384
rect 52392 14344 52409 14384
rect 52495 14344 52516 14384
rect 52556 14344 52577 14384
rect 52663 14344 52680 14384
rect 52720 14344 52729 14384
rect 52343 14321 52409 14344
rect 52495 14321 52577 14344
rect 52663 14321 52729 14344
rect 52343 14302 52729 14321
rect 56343 14407 56729 14426
rect 56343 14384 56409 14407
rect 56495 14384 56577 14407
rect 56663 14384 56729 14407
rect 56343 14344 56352 14384
rect 56392 14344 56409 14384
rect 56495 14344 56516 14384
rect 56556 14344 56577 14384
rect 56663 14344 56680 14384
rect 56720 14344 56729 14384
rect 56343 14321 56409 14344
rect 56495 14321 56577 14344
rect 56663 14321 56729 14344
rect 56343 14302 56729 14321
rect 60343 14407 60729 14426
rect 60343 14384 60409 14407
rect 60495 14384 60577 14407
rect 60663 14384 60729 14407
rect 60343 14344 60352 14384
rect 60392 14344 60409 14384
rect 60495 14344 60516 14384
rect 60556 14344 60577 14384
rect 60663 14344 60680 14384
rect 60720 14344 60729 14384
rect 60343 14321 60409 14344
rect 60495 14321 60577 14344
rect 60663 14321 60729 14344
rect 60343 14302 60729 14321
rect 64343 14407 64729 14426
rect 64343 14384 64409 14407
rect 64495 14384 64577 14407
rect 64663 14384 64729 14407
rect 64343 14344 64352 14384
rect 64392 14344 64409 14384
rect 64495 14344 64516 14384
rect 64556 14344 64577 14384
rect 64663 14344 64680 14384
rect 64720 14344 64729 14384
rect 64343 14321 64409 14344
rect 64495 14321 64577 14344
rect 64663 14321 64729 14344
rect 64343 14302 64729 14321
rect 68343 14407 68729 14426
rect 68343 14384 68409 14407
rect 68495 14384 68577 14407
rect 68663 14384 68729 14407
rect 68343 14344 68352 14384
rect 68392 14344 68409 14384
rect 68495 14344 68516 14384
rect 68556 14344 68577 14384
rect 68663 14344 68680 14384
rect 68720 14344 68729 14384
rect 68343 14321 68409 14344
rect 68495 14321 68577 14344
rect 68663 14321 68729 14344
rect 68343 14302 68729 14321
rect 72316 14364 72409 14450
rect 72495 14364 72577 14450
rect 72663 14364 72756 14450
rect 72316 14282 72756 14364
rect 72316 14196 72409 14282
rect 72495 14196 72577 14282
rect 72663 14196 72756 14282
rect 72316 14114 72756 14196
rect 72316 14028 72409 14114
rect 72495 14028 72577 14114
rect 72663 14028 72756 14114
rect 72316 13946 72756 14028
rect 72316 13860 72409 13946
rect 72495 13860 72577 13946
rect 72663 13860 72756 13946
rect 72316 13778 72756 13860
rect 72316 13692 72409 13778
rect 72495 13692 72577 13778
rect 72663 13692 72756 13778
rect 3103 13651 3489 13670
rect 3103 13628 3169 13651
rect 3255 13628 3337 13651
rect 3423 13628 3489 13651
rect 3103 13588 3112 13628
rect 3152 13588 3169 13628
rect 3255 13588 3276 13628
rect 3316 13588 3337 13628
rect 3423 13588 3440 13628
rect 3480 13588 3489 13628
rect 3103 13565 3169 13588
rect 3255 13565 3337 13588
rect 3423 13565 3489 13588
rect 3103 13546 3489 13565
rect 7103 13651 7489 13670
rect 7103 13628 7169 13651
rect 7255 13628 7337 13651
rect 7423 13628 7489 13651
rect 7103 13588 7112 13628
rect 7152 13588 7169 13628
rect 7255 13588 7276 13628
rect 7316 13588 7337 13628
rect 7423 13588 7440 13628
rect 7480 13588 7489 13628
rect 7103 13565 7169 13588
rect 7255 13565 7337 13588
rect 7423 13565 7489 13588
rect 7103 13546 7489 13565
rect 11103 13651 11489 13670
rect 11103 13628 11169 13651
rect 11255 13628 11337 13651
rect 11423 13628 11489 13651
rect 11103 13588 11112 13628
rect 11152 13588 11169 13628
rect 11255 13588 11276 13628
rect 11316 13588 11337 13628
rect 11423 13588 11440 13628
rect 11480 13588 11489 13628
rect 11103 13565 11169 13588
rect 11255 13565 11337 13588
rect 11423 13565 11489 13588
rect 11103 13546 11489 13565
rect 15103 13651 15489 13670
rect 15103 13628 15169 13651
rect 15255 13628 15337 13651
rect 15423 13628 15489 13651
rect 15103 13588 15112 13628
rect 15152 13588 15169 13628
rect 15255 13588 15276 13628
rect 15316 13588 15337 13628
rect 15423 13588 15440 13628
rect 15480 13588 15489 13628
rect 15103 13565 15169 13588
rect 15255 13565 15337 13588
rect 15423 13565 15489 13588
rect 15103 13546 15489 13565
rect 19103 13651 19489 13670
rect 19103 13628 19169 13651
rect 19255 13628 19337 13651
rect 19423 13628 19489 13651
rect 19103 13588 19112 13628
rect 19152 13588 19169 13628
rect 19255 13588 19276 13628
rect 19316 13588 19337 13628
rect 19423 13588 19440 13628
rect 19480 13588 19489 13628
rect 19103 13565 19169 13588
rect 19255 13565 19337 13588
rect 19423 13565 19489 13588
rect 19103 13546 19489 13565
rect 23103 13651 23489 13670
rect 23103 13628 23169 13651
rect 23255 13628 23337 13651
rect 23423 13628 23489 13651
rect 23103 13588 23112 13628
rect 23152 13588 23169 13628
rect 23255 13588 23276 13628
rect 23316 13588 23337 13628
rect 23423 13588 23440 13628
rect 23480 13588 23489 13628
rect 23103 13565 23169 13588
rect 23255 13565 23337 13588
rect 23423 13565 23489 13588
rect 23103 13546 23489 13565
rect 27103 13651 27489 13670
rect 27103 13628 27169 13651
rect 27255 13628 27337 13651
rect 27423 13628 27489 13651
rect 27103 13588 27112 13628
rect 27152 13588 27169 13628
rect 27255 13588 27276 13628
rect 27316 13588 27337 13628
rect 27423 13588 27440 13628
rect 27480 13588 27489 13628
rect 27103 13565 27169 13588
rect 27255 13565 27337 13588
rect 27423 13565 27489 13588
rect 27103 13546 27489 13565
rect 31103 13651 31489 13670
rect 31103 13628 31169 13651
rect 31255 13628 31337 13651
rect 31423 13628 31489 13651
rect 31103 13588 31112 13628
rect 31152 13588 31169 13628
rect 31255 13588 31276 13628
rect 31316 13588 31337 13628
rect 31423 13588 31440 13628
rect 31480 13588 31489 13628
rect 31103 13565 31169 13588
rect 31255 13565 31337 13588
rect 31423 13565 31489 13588
rect 31103 13546 31489 13565
rect 35103 13651 35489 13670
rect 35103 13628 35169 13651
rect 35255 13628 35337 13651
rect 35423 13628 35489 13651
rect 35103 13588 35112 13628
rect 35152 13588 35169 13628
rect 35255 13588 35276 13628
rect 35316 13588 35337 13628
rect 35423 13588 35440 13628
rect 35480 13588 35489 13628
rect 35103 13565 35169 13588
rect 35255 13565 35337 13588
rect 35423 13565 35489 13588
rect 35103 13546 35489 13565
rect 39103 13651 39489 13670
rect 39103 13628 39169 13651
rect 39255 13628 39337 13651
rect 39423 13628 39489 13651
rect 39103 13588 39112 13628
rect 39152 13588 39169 13628
rect 39255 13588 39276 13628
rect 39316 13588 39337 13628
rect 39423 13588 39440 13628
rect 39480 13588 39489 13628
rect 39103 13565 39169 13588
rect 39255 13565 39337 13588
rect 39423 13565 39489 13588
rect 39103 13546 39489 13565
rect 43103 13651 43489 13670
rect 43103 13628 43169 13651
rect 43255 13628 43337 13651
rect 43423 13628 43489 13651
rect 43103 13588 43112 13628
rect 43152 13588 43169 13628
rect 43255 13588 43276 13628
rect 43316 13588 43337 13628
rect 43423 13588 43440 13628
rect 43480 13588 43489 13628
rect 43103 13565 43169 13588
rect 43255 13565 43337 13588
rect 43423 13565 43489 13588
rect 43103 13546 43489 13565
rect 47103 13651 47489 13670
rect 47103 13628 47169 13651
rect 47255 13628 47337 13651
rect 47423 13628 47489 13651
rect 47103 13588 47112 13628
rect 47152 13588 47169 13628
rect 47255 13588 47276 13628
rect 47316 13588 47337 13628
rect 47423 13588 47440 13628
rect 47480 13588 47489 13628
rect 47103 13565 47169 13588
rect 47255 13565 47337 13588
rect 47423 13565 47489 13588
rect 47103 13546 47489 13565
rect 51103 13651 51489 13670
rect 51103 13628 51169 13651
rect 51255 13628 51337 13651
rect 51423 13628 51489 13651
rect 51103 13588 51112 13628
rect 51152 13588 51169 13628
rect 51255 13588 51276 13628
rect 51316 13588 51337 13628
rect 51423 13588 51440 13628
rect 51480 13588 51489 13628
rect 51103 13565 51169 13588
rect 51255 13565 51337 13588
rect 51423 13565 51489 13588
rect 51103 13546 51489 13565
rect 55103 13651 55489 13670
rect 55103 13628 55169 13651
rect 55255 13628 55337 13651
rect 55423 13628 55489 13651
rect 55103 13588 55112 13628
rect 55152 13588 55169 13628
rect 55255 13588 55276 13628
rect 55316 13588 55337 13628
rect 55423 13588 55440 13628
rect 55480 13588 55489 13628
rect 55103 13565 55169 13588
rect 55255 13565 55337 13588
rect 55423 13565 55489 13588
rect 55103 13546 55489 13565
rect 59103 13651 59489 13670
rect 59103 13628 59169 13651
rect 59255 13628 59337 13651
rect 59423 13628 59489 13651
rect 59103 13588 59112 13628
rect 59152 13588 59169 13628
rect 59255 13588 59276 13628
rect 59316 13588 59337 13628
rect 59423 13588 59440 13628
rect 59480 13588 59489 13628
rect 59103 13565 59169 13588
rect 59255 13565 59337 13588
rect 59423 13565 59489 13588
rect 59103 13546 59489 13565
rect 63103 13651 63489 13670
rect 63103 13628 63169 13651
rect 63255 13628 63337 13651
rect 63423 13628 63489 13651
rect 63103 13588 63112 13628
rect 63152 13588 63169 13628
rect 63255 13588 63276 13628
rect 63316 13588 63337 13628
rect 63423 13588 63440 13628
rect 63480 13588 63489 13628
rect 63103 13565 63169 13588
rect 63255 13565 63337 13588
rect 63423 13565 63489 13588
rect 63103 13546 63489 13565
rect 67103 13651 67489 13670
rect 67103 13628 67169 13651
rect 67255 13628 67337 13651
rect 67423 13628 67489 13651
rect 67103 13588 67112 13628
rect 67152 13588 67169 13628
rect 67255 13588 67276 13628
rect 67316 13588 67337 13628
rect 67423 13588 67440 13628
rect 67480 13588 67489 13628
rect 67103 13565 67169 13588
rect 67255 13565 67337 13588
rect 67423 13565 67489 13588
rect 67103 13546 67489 13565
rect 72316 13610 72756 13692
rect 72316 13524 72409 13610
rect 72495 13524 72577 13610
rect 72663 13524 72756 13610
rect 72316 13442 72756 13524
rect 72316 13356 72409 13442
rect 72495 13356 72577 13442
rect 72663 13356 72756 13442
rect 72316 13274 72756 13356
rect 72316 13188 72409 13274
rect 72495 13188 72577 13274
rect 72663 13188 72756 13274
rect 72316 13106 72756 13188
rect 72316 13020 72409 13106
rect 72495 13020 72577 13106
rect 72663 13020 72756 13106
rect 4343 12895 4729 12914
rect 4343 12872 4409 12895
rect 4495 12872 4577 12895
rect 4663 12872 4729 12895
rect 4343 12832 4352 12872
rect 4392 12832 4409 12872
rect 4495 12832 4516 12872
rect 4556 12832 4577 12872
rect 4663 12832 4680 12872
rect 4720 12832 4729 12872
rect 4343 12809 4409 12832
rect 4495 12809 4577 12832
rect 4663 12809 4729 12832
rect 4343 12790 4729 12809
rect 8343 12895 8729 12914
rect 8343 12872 8409 12895
rect 8495 12872 8577 12895
rect 8663 12872 8729 12895
rect 8343 12832 8352 12872
rect 8392 12832 8409 12872
rect 8495 12832 8516 12872
rect 8556 12832 8577 12872
rect 8663 12832 8680 12872
rect 8720 12832 8729 12872
rect 8343 12809 8409 12832
rect 8495 12809 8577 12832
rect 8663 12809 8729 12832
rect 8343 12790 8729 12809
rect 12343 12895 12729 12914
rect 12343 12872 12409 12895
rect 12495 12872 12577 12895
rect 12663 12872 12729 12895
rect 12343 12832 12352 12872
rect 12392 12832 12409 12872
rect 12495 12832 12516 12872
rect 12556 12832 12577 12872
rect 12663 12832 12680 12872
rect 12720 12832 12729 12872
rect 12343 12809 12409 12832
rect 12495 12809 12577 12832
rect 12663 12809 12729 12832
rect 12343 12790 12729 12809
rect 16343 12895 16729 12914
rect 16343 12872 16409 12895
rect 16495 12872 16577 12895
rect 16663 12872 16729 12895
rect 16343 12832 16352 12872
rect 16392 12832 16409 12872
rect 16495 12832 16516 12872
rect 16556 12832 16577 12872
rect 16663 12832 16680 12872
rect 16720 12832 16729 12872
rect 16343 12809 16409 12832
rect 16495 12809 16577 12832
rect 16663 12809 16729 12832
rect 16343 12790 16729 12809
rect 20343 12895 20729 12914
rect 20343 12872 20409 12895
rect 20495 12872 20577 12895
rect 20663 12872 20729 12895
rect 20343 12832 20352 12872
rect 20392 12832 20409 12872
rect 20495 12832 20516 12872
rect 20556 12832 20577 12872
rect 20663 12832 20680 12872
rect 20720 12832 20729 12872
rect 20343 12809 20409 12832
rect 20495 12809 20577 12832
rect 20663 12809 20729 12832
rect 20343 12790 20729 12809
rect 24343 12895 24729 12914
rect 24343 12872 24409 12895
rect 24495 12872 24577 12895
rect 24663 12872 24729 12895
rect 24343 12832 24352 12872
rect 24392 12832 24409 12872
rect 24495 12832 24516 12872
rect 24556 12832 24577 12872
rect 24663 12832 24680 12872
rect 24720 12832 24729 12872
rect 24343 12809 24409 12832
rect 24495 12809 24577 12832
rect 24663 12809 24729 12832
rect 24343 12790 24729 12809
rect 28343 12895 28729 12914
rect 28343 12872 28409 12895
rect 28495 12872 28577 12895
rect 28663 12872 28729 12895
rect 28343 12832 28352 12872
rect 28392 12832 28409 12872
rect 28495 12832 28516 12872
rect 28556 12832 28577 12872
rect 28663 12832 28680 12872
rect 28720 12832 28729 12872
rect 28343 12809 28409 12832
rect 28495 12809 28577 12832
rect 28663 12809 28729 12832
rect 28343 12790 28729 12809
rect 32343 12895 32729 12914
rect 32343 12872 32409 12895
rect 32495 12872 32577 12895
rect 32663 12872 32729 12895
rect 32343 12832 32352 12872
rect 32392 12832 32409 12872
rect 32495 12832 32516 12872
rect 32556 12832 32577 12872
rect 32663 12832 32680 12872
rect 32720 12832 32729 12872
rect 32343 12809 32409 12832
rect 32495 12809 32577 12832
rect 32663 12809 32729 12832
rect 32343 12790 32729 12809
rect 36343 12895 36729 12914
rect 36343 12872 36409 12895
rect 36495 12872 36577 12895
rect 36663 12872 36729 12895
rect 36343 12832 36352 12872
rect 36392 12832 36409 12872
rect 36495 12832 36516 12872
rect 36556 12832 36577 12872
rect 36663 12832 36680 12872
rect 36720 12832 36729 12872
rect 36343 12809 36409 12832
rect 36495 12809 36577 12832
rect 36663 12809 36729 12832
rect 36343 12790 36729 12809
rect 40343 12895 40729 12914
rect 40343 12872 40409 12895
rect 40495 12872 40577 12895
rect 40663 12872 40729 12895
rect 40343 12832 40352 12872
rect 40392 12832 40409 12872
rect 40495 12832 40516 12872
rect 40556 12832 40577 12872
rect 40663 12832 40680 12872
rect 40720 12832 40729 12872
rect 40343 12809 40409 12832
rect 40495 12809 40577 12832
rect 40663 12809 40729 12832
rect 40343 12790 40729 12809
rect 44343 12895 44729 12914
rect 44343 12872 44409 12895
rect 44495 12872 44577 12895
rect 44663 12872 44729 12895
rect 44343 12832 44352 12872
rect 44392 12832 44409 12872
rect 44495 12832 44516 12872
rect 44556 12832 44577 12872
rect 44663 12832 44680 12872
rect 44720 12832 44729 12872
rect 44343 12809 44409 12832
rect 44495 12809 44577 12832
rect 44663 12809 44729 12832
rect 44343 12790 44729 12809
rect 48343 12895 48729 12914
rect 48343 12872 48409 12895
rect 48495 12872 48577 12895
rect 48663 12872 48729 12895
rect 48343 12832 48352 12872
rect 48392 12832 48409 12872
rect 48495 12832 48516 12872
rect 48556 12832 48577 12872
rect 48663 12832 48680 12872
rect 48720 12832 48729 12872
rect 48343 12809 48409 12832
rect 48495 12809 48577 12832
rect 48663 12809 48729 12832
rect 48343 12790 48729 12809
rect 52343 12895 52729 12914
rect 52343 12872 52409 12895
rect 52495 12872 52577 12895
rect 52663 12872 52729 12895
rect 52343 12832 52352 12872
rect 52392 12832 52409 12872
rect 52495 12832 52516 12872
rect 52556 12832 52577 12872
rect 52663 12832 52680 12872
rect 52720 12832 52729 12872
rect 52343 12809 52409 12832
rect 52495 12809 52577 12832
rect 52663 12809 52729 12832
rect 52343 12790 52729 12809
rect 56343 12895 56729 12914
rect 56343 12872 56409 12895
rect 56495 12872 56577 12895
rect 56663 12872 56729 12895
rect 56343 12832 56352 12872
rect 56392 12832 56409 12872
rect 56495 12832 56516 12872
rect 56556 12832 56577 12872
rect 56663 12832 56680 12872
rect 56720 12832 56729 12872
rect 56343 12809 56409 12832
rect 56495 12809 56577 12832
rect 56663 12809 56729 12832
rect 56343 12790 56729 12809
rect 60343 12895 60729 12914
rect 60343 12872 60409 12895
rect 60495 12872 60577 12895
rect 60663 12872 60729 12895
rect 60343 12832 60352 12872
rect 60392 12832 60409 12872
rect 60495 12832 60516 12872
rect 60556 12832 60577 12872
rect 60663 12832 60680 12872
rect 60720 12832 60729 12872
rect 60343 12809 60409 12832
rect 60495 12809 60577 12832
rect 60663 12809 60729 12832
rect 60343 12790 60729 12809
rect 64343 12895 64729 12914
rect 64343 12872 64409 12895
rect 64495 12872 64577 12895
rect 64663 12872 64729 12895
rect 64343 12832 64352 12872
rect 64392 12832 64409 12872
rect 64495 12832 64516 12872
rect 64556 12832 64577 12872
rect 64663 12832 64680 12872
rect 64720 12832 64729 12872
rect 64343 12809 64409 12832
rect 64495 12809 64577 12832
rect 64663 12809 64729 12832
rect 64343 12790 64729 12809
rect 68343 12895 68729 12914
rect 68343 12872 68409 12895
rect 68495 12872 68577 12895
rect 68663 12872 68729 12895
rect 72316 12890 72756 13020
rect 76316 15122 76756 15252
rect 76316 15036 76409 15122
rect 76495 15036 76577 15122
rect 76663 15036 76756 15122
rect 76316 14954 76756 15036
rect 76316 14868 76409 14954
rect 76495 14868 76577 14954
rect 76663 14868 76756 14954
rect 76316 14786 76756 14868
rect 76316 14700 76409 14786
rect 76495 14700 76577 14786
rect 76663 14700 76756 14786
rect 76316 14618 76756 14700
rect 76316 14532 76409 14618
rect 76495 14532 76577 14618
rect 76663 14532 76756 14618
rect 76316 14450 76756 14532
rect 76316 14364 76409 14450
rect 76495 14364 76577 14450
rect 76663 14364 76756 14450
rect 76316 14282 76756 14364
rect 76316 14196 76409 14282
rect 76495 14196 76577 14282
rect 76663 14196 76756 14282
rect 76316 14114 76756 14196
rect 76316 14028 76409 14114
rect 76495 14028 76577 14114
rect 76663 14028 76756 14114
rect 76316 13946 76756 14028
rect 76316 13860 76409 13946
rect 76495 13860 76577 13946
rect 76663 13860 76756 13946
rect 76316 13778 76756 13860
rect 76316 13692 76409 13778
rect 76495 13692 76577 13778
rect 76663 13692 76756 13778
rect 76316 13610 76756 13692
rect 76316 13524 76409 13610
rect 76495 13524 76577 13610
rect 76663 13524 76756 13610
rect 76316 13442 76756 13524
rect 76316 13356 76409 13442
rect 76495 13356 76577 13442
rect 76663 13356 76756 13442
rect 76316 13274 76756 13356
rect 76316 13188 76409 13274
rect 76495 13188 76577 13274
rect 76663 13188 76756 13274
rect 76316 13106 76756 13188
rect 76316 13020 76409 13106
rect 76495 13020 76577 13106
rect 76663 13020 76756 13106
rect 76316 12890 76756 13020
rect 80316 15122 80756 15252
rect 80316 15036 80409 15122
rect 80495 15036 80577 15122
rect 80663 15036 80756 15122
rect 80316 14954 80756 15036
rect 80316 14868 80409 14954
rect 80495 14868 80577 14954
rect 80663 14868 80756 14954
rect 80316 14786 80756 14868
rect 80316 14700 80409 14786
rect 80495 14700 80577 14786
rect 80663 14700 80756 14786
rect 80316 14618 80756 14700
rect 80316 14532 80409 14618
rect 80495 14532 80577 14618
rect 80663 14532 80756 14618
rect 80316 14450 80756 14532
rect 80316 14364 80409 14450
rect 80495 14364 80577 14450
rect 80663 14364 80756 14450
rect 80316 14282 80756 14364
rect 80316 14196 80409 14282
rect 80495 14196 80577 14282
rect 80663 14196 80756 14282
rect 80316 14114 80756 14196
rect 80316 14028 80409 14114
rect 80495 14028 80577 14114
rect 80663 14028 80756 14114
rect 80316 13946 80756 14028
rect 80316 13860 80409 13946
rect 80495 13860 80577 13946
rect 80663 13860 80756 13946
rect 80316 13778 80756 13860
rect 80316 13692 80409 13778
rect 80495 13692 80577 13778
rect 80663 13692 80756 13778
rect 80316 13610 80756 13692
rect 80316 13524 80409 13610
rect 80495 13524 80577 13610
rect 80663 13524 80756 13610
rect 80316 13442 80756 13524
rect 80316 13356 80409 13442
rect 80495 13356 80577 13442
rect 80663 13356 80756 13442
rect 80316 13274 80756 13356
rect 80316 13188 80409 13274
rect 80495 13188 80577 13274
rect 80663 13188 80756 13274
rect 80316 13106 80756 13188
rect 80316 13020 80409 13106
rect 80495 13020 80577 13106
rect 80663 13020 80756 13106
rect 80316 12890 80756 13020
rect 84316 15122 84756 15252
rect 84316 15036 84409 15122
rect 84495 15036 84577 15122
rect 84663 15036 84756 15122
rect 84316 14954 84756 15036
rect 84316 14868 84409 14954
rect 84495 14868 84577 14954
rect 84663 14868 84756 14954
rect 84316 14786 84756 14868
rect 84316 14700 84409 14786
rect 84495 14700 84577 14786
rect 84663 14700 84756 14786
rect 84316 14618 84756 14700
rect 84316 14532 84409 14618
rect 84495 14532 84577 14618
rect 84663 14532 84756 14618
rect 84316 14450 84756 14532
rect 84316 14364 84409 14450
rect 84495 14364 84577 14450
rect 84663 14364 84756 14450
rect 84316 14282 84756 14364
rect 84316 14196 84409 14282
rect 84495 14196 84577 14282
rect 84663 14196 84756 14282
rect 84316 14114 84756 14196
rect 84316 14028 84409 14114
rect 84495 14028 84577 14114
rect 84663 14028 84756 14114
rect 84316 13946 84756 14028
rect 84316 13860 84409 13946
rect 84495 13860 84577 13946
rect 84663 13860 84756 13946
rect 84316 13778 84756 13860
rect 84316 13692 84409 13778
rect 84495 13692 84577 13778
rect 84663 13692 84756 13778
rect 84316 13610 84756 13692
rect 84316 13524 84409 13610
rect 84495 13524 84577 13610
rect 84663 13524 84756 13610
rect 84316 13442 84756 13524
rect 84316 13356 84409 13442
rect 84495 13356 84577 13442
rect 84663 13356 84756 13442
rect 84316 13274 84756 13356
rect 84316 13188 84409 13274
rect 84495 13188 84577 13274
rect 84663 13188 84756 13274
rect 84316 13106 84756 13188
rect 84316 13020 84409 13106
rect 84495 13020 84577 13106
rect 84663 13020 84756 13106
rect 84316 12890 84756 13020
rect 88316 15122 88756 15252
rect 88316 15036 88409 15122
rect 88495 15036 88577 15122
rect 88663 15036 88756 15122
rect 88316 14954 88756 15036
rect 88316 14868 88409 14954
rect 88495 14868 88577 14954
rect 88663 14868 88756 14954
rect 88316 14786 88756 14868
rect 88316 14700 88409 14786
rect 88495 14700 88577 14786
rect 88663 14700 88756 14786
rect 88316 14618 88756 14700
rect 88316 14532 88409 14618
rect 88495 14532 88577 14618
rect 88663 14532 88756 14618
rect 88316 14450 88756 14532
rect 88316 14364 88409 14450
rect 88495 14364 88577 14450
rect 88663 14364 88756 14450
rect 88316 14282 88756 14364
rect 88316 14196 88409 14282
rect 88495 14196 88577 14282
rect 88663 14196 88756 14282
rect 88316 14114 88756 14196
rect 88316 14028 88409 14114
rect 88495 14028 88577 14114
rect 88663 14028 88756 14114
rect 88316 13946 88756 14028
rect 88316 13860 88409 13946
rect 88495 13860 88577 13946
rect 88663 13860 88756 13946
rect 88316 13778 88756 13860
rect 88316 13692 88409 13778
rect 88495 13692 88577 13778
rect 88663 13692 88756 13778
rect 88316 13610 88756 13692
rect 88316 13524 88409 13610
rect 88495 13524 88577 13610
rect 88663 13524 88756 13610
rect 88316 13442 88756 13524
rect 88316 13356 88409 13442
rect 88495 13356 88577 13442
rect 88663 13356 88756 13442
rect 88316 13274 88756 13356
rect 88316 13188 88409 13274
rect 88495 13188 88577 13274
rect 88663 13188 88756 13274
rect 88316 13106 88756 13188
rect 88316 13020 88409 13106
rect 88495 13020 88577 13106
rect 88663 13020 88756 13106
rect 88316 12890 88756 13020
rect 92316 15122 92756 15252
rect 92316 15036 92409 15122
rect 92495 15036 92577 15122
rect 92663 15036 92756 15122
rect 92316 14954 92756 15036
rect 92316 14868 92409 14954
rect 92495 14868 92577 14954
rect 92663 14868 92756 14954
rect 92316 14786 92756 14868
rect 92316 14700 92409 14786
rect 92495 14700 92577 14786
rect 92663 14700 92756 14786
rect 92316 14618 92756 14700
rect 92316 14532 92409 14618
rect 92495 14532 92577 14618
rect 92663 14532 92756 14618
rect 92316 14450 92756 14532
rect 92316 14364 92409 14450
rect 92495 14364 92577 14450
rect 92663 14364 92756 14450
rect 92316 14282 92756 14364
rect 92316 14196 92409 14282
rect 92495 14196 92577 14282
rect 92663 14196 92756 14282
rect 92316 14114 92756 14196
rect 92316 14028 92409 14114
rect 92495 14028 92577 14114
rect 92663 14028 92756 14114
rect 92316 13946 92756 14028
rect 92316 13860 92409 13946
rect 92495 13860 92577 13946
rect 92663 13860 92756 13946
rect 92316 13778 92756 13860
rect 92316 13692 92409 13778
rect 92495 13692 92577 13778
rect 92663 13692 92756 13778
rect 92316 13610 92756 13692
rect 92316 13524 92409 13610
rect 92495 13524 92577 13610
rect 92663 13524 92756 13610
rect 92316 13442 92756 13524
rect 92316 13356 92409 13442
rect 92495 13356 92577 13442
rect 92663 13356 92756 13442
rect 92316 13274 92756 13356
rect 92316 13188 92409 13274
rect 92495 13188 92577 13274
rect 92663 13188 92756 13274
rect 92316 13106 92756 13188
rect 92316 13020 92409 13106
rect 92495 13020 92577 13106
rect 92663 13020 92756 13106
rect 92316 12890 92756 13020
rect 96316 15122 96756 15252
rect 96316 15036 96409 15122
rect 96495 15036 96577 15122
rect 96663 15036 96756 15122
rect 96316 14954 96756 15036
rect 96316 14868 96409 14954
rect 96495 14868 96577 14954
rect 96663 14868 96756 14954
rect 96316 14786 96756 14868
rect 96316 14700 96409 14786
rect 96495 14700 96577 14786
rect 96663 14700 96756 14786
rect 96316 14618 96756 14700
rect 96316 14532 96409 14618
rect 96495 14532 96577 14618
rect 96663 14532 96756 14618
rect 96316 14450 96756 14532
rect 96316 14364 96409 14450
rect 96495 14364 96577 14450
rect 96663 14364 96756 14450
rect 96316 14282 96756 14364
rect 96316 14196 96409 14282
rect 96495 14196 96577 14282
rect 96663 14196 96756 14282
rect 96316 14114 96756 14196
rect 96316 14028 96409 14114
rect 96495 14028 96577 14114
rect 96663 14028 96756 14114
rect 96316 13946 96756 14028
rect 96316 13860 96409 13946
rect 96495 13860 96577 13946
rect 96663 13860 96756 13946
rect 96316 13778 96756 13860
rect 96316 13692 96409 13778
rect 96495 13692 96577 13778
rect 96663 13692 96756 13778
rect 96316 13610 96756 13692
rect 96316 13524 96409 13610
rect 96495 13524 96577 13610
rect 96663 13524 96756 13610
rect 96316 13442 96756 13524
rect 96316 13356 96409 13442
rect 96495 13356 96577 13442
rect 96663 13356 96756 13442
rect 96316 13274 96756 13356
rect 96316 13188 96409 13274
rect 96495 13188 96577 13274
rect 96663 13188 96756 13274
rect 96316 13106 96756 13188
rect 96316 13020 96409 13106
rect 96495 13020 96577 13106
rect 96663 13020 96756 13106
rect 96316 12890 96756 13020
rect 68343 12832 68352 12872
rect 68392 12832 68409 12872
rect 68495 12832 68516 12872
rect 68556 12832 68577 12872
rect 68663 12832 68680 12872
rect 68720 12832 68729 12872
rect 68343 12809 68409 12832
rect 68495 12809 68577 12832
rect 68663 12809 68729 12832
rect 68343 12790 68729 12809
rect 75076 12246 75516 12376
rect 75076 12160 75169 12246
rect 75255 12160 75337 12246
rect 75423 12160 75516 12246
rect 3103 12139 3489 12158
rect 3103 12116 3169 12139
rect 3255 12116 3337 12139
rect 3423 12116 3489 12139
rect 3103 12076 3112 12116
rect 3152 12076 3169 12116
rect 3255 12076 3276 12116
rect 3316 12076 3337 12116
rect 3423 12076 3440 12116
rect 3480 12076 3489 12116
rect 3103 12053 3169 12076
rect 3255 12053 3337 12076
rect 3423 12053 3489 12076
rect 3103 12034 3489 12053
rect 7103 12139 7489 12158
rect 7103 12116 7169 12139
rect 7255 12116 7337 12139
rect 7423 12116 7489 12139
rect 7103 12076 7112 12116
rect 7152 12076 7169 12116
rect 7255 12076 7276 12116
rect 7316 12076 7337 12116
rect 7423 12076 7440 12116
rect 7480 12076 7489 12116
rect 7103 12053 7169 12076
rect 7255 12053 7337 12076
rect 7423 12053 7489 12076
rect 7103 12034 7489 12053
rect 11103 12139 11489 12158
rect 11103 12116 11169 12139
rect 11255 12116 11337 12139
rect 11423 12116 11489 12139
rect 11103 12076 11112 12116
rect 11152 12076 11169 12116
rect 11255 12076 11276 12116
rect 11316 12076 11337 12116
rect 11423 12076 11440 12116
rect 11480 12076 11489 12116
rect 11103 12053 11169 12076
rect 11255 12053 11337 12076
rect 11423 12053 11489 12076
rect 11103 12034 11489 12053
rect 15103 12139 15489 12158
rect 15103 12116 15169 12139
rect 15255 12116 15337 12139
rect 15423 12116 15489 12139
rect 15103 12076 15112 12116
rect 15152 12076 15169 12116
rect 15255 12076 15276 12116
rect 15316 12076 15337 12116
rect 15423 12076 15440 12116
rect 15480 12076 15489 12116
rect 15103 12053 15169 12076
rect 15255 12053 15337 12076
rect 15423 12053 15489 12076
rect 15103 12034 15489 12053
rect 19103 12139 19489 12158
rect 19103 12116 19169 12139
rect 19255 12116 19337 12139
rect 19423 12116 19489 12139
rect 19103 12076 19112 12116
rect 19152 12076 19169 12116
rect 19255 12076 19276 12116
rect 19316 12076 19337 12116
rect 19423 12076 19440 12116
rect 19480 12076 19489 12116
rect 19103 12053 19169 12076
rect 19255 12053 19337 12076
rect 19423 12053 19489 12076
rect 19103 12034 19489 12053
rect 23103 12139 23489 12158
rect 23103 12116 23169 12139
rect 23255 12116 23337 12139
rect 23423 12116 23489 12139
rect 23103 12076 23112 12116
rect 23152 12076 23169 12116
rect 23255 12076 23276 12116
rect 23316 12076 23337 12116
rect 23423 12076 23440 12116
rect 23480 12076 23489 12116
rect 23103 12053 23169 12076
rect 23255 12053 23337 12076
rect 23423 12053 23489 12076
rect 23103 12034 23489 12053
rect 27103 12139 27489 12158
rect 27103 12116 27169 12139
rect 27255 12116 27337 12139
rect 27423 12116 27489 12139
rect 27103 12076 27112 12116
rect 27152 12076 27169 12116
rect 27255 12076 27276 12116
rect 27316 12076 27337 12116
rect 27423 12076 27440 12116
rect 27480 12076 27489 12116
rect 27103 12053 27169 12076
rect 27255 12053 27337 12076
rect 27423 12053 27489 12076
rect 27103 12034 27489 12053
rect 31103 12139 31489 12158
rect 31103 12116 31169 12139
rect 31255 12116 31337 12139
rect 31423 12116 31489 12139
rect 31103 12076 31112 12116
rect 31152 12076 31169 12116
rect 31255 12076 31276 12116
rect 31316 12076 31337 12116
rect 31423 12076 31440 12116
rect 31480 12076 31489 12116
rect 31103 12053 31169 12076
rect 31255 12053 31337 12076
rect 31423 12053 31489 12076
rect 31103 12034 31489 12053
rect 35103 12139 35489 12158
rect 35103 12116 35169 12139
rect 35255 12116 35337 12139
rect 35423 12116 35489 12139
rect 35103 12076 35112 12116
rect 35152 12076 35169 12116
rect 35255 12076 35276 12116
rect 35316 12076 35337 12116
rect 35423 12076 35440 12116
rect 35480 12076 35489 12116
rect 35103 12053 35169 12076
rect 35255 12053 35337 12076
rect 35423 12053 35489 12076
rect 35103 12034 35489 12053
rect 39103 12139 39489 12158
rect 39103 12116 39169 12139
rect 39255 12116 39337 12139
rect 39423 12116 39489 12139
rect 39103 12076 39112 12116
rect 39152 12076 39169 12116
rect 39255 12076 39276 12116
rect 39316 12076 39337 12116
rect 39423 12076 39440 12116
rect 39480 12076 39489 12116
rect 39103 12053 39169 12076
rect 39255 12053 39337 12076
rect 39423 12053 39489 12076
rect 39103 12034 39489 12053
rect 43103 12139 43489 12158
rect 43103 12116 43169 12139
rect 43255 12116 43337 12139
rect 43423 12116 43489 12139
rect 43103 12076 43112 12116
rect 43152 12076 43169 12116
rect 43255 12076 43276 12116
rect 43316 12076 43337 12116
rect 43423 12076 43440 12116
rect 43480 12076 43489 12116
rect 43103 12053 43169 12076
rect 43255 12053 43337 12076
rect 43423 12053 43489 12076
rect 43103 12034 43489 12053
rect 47103 12139 47489 12158
rect 47103 12116 47169 12139
rect 47255 12116 47337 12139
rect 47423 12116 47489 12139
rect 47103 12076 47112 12116
rect 47152 12076 47169 12116
rect 47255 12076 47276 12116
rect 47316 12076 47337 12116
rect 47423 12076 47440 12116
rect 47480 12076 47489 12116
rect 47103 12053 47169 12076
rect 47255 12053 47337 12076
rect 47423 12053 47489 12076
rect 47103 12034 47489 12053
rect 51103 12139 51489 12158
rect 51103 12116 51169 12139
rect 51255 12116 51337 12139
rect 51423 12116 51489 12139
rect 51103 12076 51112 12116
rect 51152 12076 51169 12116
rect 51255 12076 51276 12116
rect 51316 12076 51337 12116
rect 51423 12076 51440 12116
rect 51480 12076 51489 12116
rect 51103 12053 51169 12076
rect 51255 12053 51337 12076
rect 51423 12053 51489 12076
rect 51103 12034 51489 12053
rect 55103 12139 55489 12158
rect 55103 12116 55169 12139
rect 55255 12116 55337 12139
rect 55423 12116 55489 12139
rect 55103 12076 55112 12116
rect 55152 12076 55169 12116
rect 55255 12076 55276 12116
rect 55316 12076 55337 12116
rect 55423 12076 55440 12116
rect 55480 12076 55489 12116
rect 55103 12053 55169 12076
rect 55255 12053 55337 12076
rect 55423 12053 55489 12076
rect 55103 12034 55489 12053
rect 59103 12139 59489 12158
rect 59103 12116 59169 12139
rect 59255 12116 59337 12139
rect 59423 12116 59489 12139
rect 59103 12076 59112 12116
rect 59152 12076 59169 12116
rect 59255 12076 59276 12116
rect 59316 12076 59337 12116
rect 59423 12076 59440 12116
rect 59480 12076 59489 12116
rect 59103 12053 59169 12076
rect 59255 12053 59337 12076
rect 59423 12053 59489 12076
rect 59103 12034 59489 12053
rect 63103 12139 63489 12158
rect 63103 12116 63169 12139
rect 63255 12116 63337 12139
rect 63423 12116 63489 12139
rect 63103 12076 63112 12116
rect 63152 12076 63169 12116
rect 63255 12076 63276 12116
rect 63316 12076 63337 12116
rect 63423 12076 63440 12116
rect 63480 12076 63489 12116
rect 63103 12053 63169 12076
rect 63255 12053 63337 12076
rect 63423 12053 63489 12076
rect 63103 12034 63489 12053
rect 67103 12139 67489 12158
rect 67103 12116 67169 12139
rect 67255 12116 67337 12139
rect 67423 12116 67489 12139
rect 67103 12076 67112 12116
rect 67152 12076 67169 12116
rect 67255 12076 67276 12116
rect 67316 12076 67337 12116
rect 67423 12076 67440 12116
rect 67480 12076 67489 12116
rect 67103 12053 67169 12076
rect 67255 12053 67337 12076
rect 67423 12053 67489 12076
rect 67103 12034 67489 12053
rect 75076 12078 75516 12160
rect 75076 11992 75169 12078
rect 75255 11992 75337 12078
rect 75423 11992 75516 12078
rect 75076 11910 75516 11992
rect 75076 11824 75169 11910
rect 75255 11824 75337 11910
rect 75423 11824 75516 11910
rect 75076 11742 75516 11824
rect 75076 11656 75169 11742
rect 75255 11656 75337 11742
rect 75423 11656 75516 11742
rect 75076 11574 75516 11656
rect 75076 11488 75169 11574
rect 75255 11488 75337 11574
rect 75423 11488 75516 11574
rect 75076 11406 75516 11488
rect 4343 11383 4729 11402
rect 4343 11360 4409 11383
rect 4495 11360 4577 11383
rect 4663 11360 4729 11383
rect 4343 11320 4352 11360
rect 4392 11320 4409 11360
rect 4495 11320 4516 11360
rect 4556 11320 4577 11360
rect 4663 11320 4680 11360
rect 4720 11320 4729 11360
rect 4343 11297 4409 11320
rect 4495 11297 4577 11320
rect 4663 11297 4729 11320
rect 4343 11278 4729 11297
rect 8343 11383 8729 11402
rect 8343 11360 8409 11383
rect 8495 11360 8577 11383
rect 8663 11360 8729 11383
rect 8343 11320 8352 11360
rect 8392 11320 8409 11360
rect 8495 11320 8516 11360
rect 8556 11320 8577 11360
rect 8663 11320 8680 11360
rect 8720 11320 8729 11360
rect 8343 11297 8409 11320
rect 8495 11297 8577 11320
rect 8663 11297 8729 11320
rect 8343 11278 8729 11297
rect 12343 11383 12729 11402
rect 12343 11360 12409 11383
rect 12495 11360 12577 11383
rect 12663 11360 12729 11383
rect 12343 11320 12352 11360
rect 12392 11320 12409 11360
rect 12495 11320 12516 11360
rect 12556 11320 12577 11360
rect 12663 11320 12680 11360
rect 12720 11320 12729 11360
rect 12343 11297 12409 11320
rect 12495 11297 12577 11320
rect 12663 11297 12729 11320
rect 12343 11278 12729 11297
rect 16343 11383 16729 11402
rect 16343 11360 16409 11383
rect 16495 11360 16577 11383
rect 16663 11360 16729 11383
rect 16343 11320 16352 11360
rect 16392 11320 16409 11360
rect 16495 11320 16516 11360
rect 16556 11320 16577 11360
rect 16663 11320 16680 11360
rect 16720 11320 16729 11360
rect 16343 11297 16409 11320
rect 16495 11297 16577 11320
rect 16663 11297 16729 11320
rect 16343 11278 16729 11297
rect 20343 11383 20729 11402
rect 20343 11360 20409 11383
rect 20495 11360 20577 11383
rect 20663 11360 20729 11383
rect 20343 11320 20352 11360
rect 20392 11320 20409 11360
rect 20495 11320 20516 11360
rect 20556 11320 20577 11360
rect 20663 11320 20680 11360
rect 20720 11320 20729 11360
rect 20343 11297 20409 11320
rect 20495 11297 20577 11320
rect 20663 11297 20729 11320
rect 20343 11278 20729 11297
rect 24343 11383 24729 11402
rect 24343 11360 24409 11383
rect 24495 11360 24577 11383
rect 24663 11360 24729 11383
rect 24343 11320 24352 11360
rect 24392 11320 24409 11360
rect 24495 11320 24516 11360
rect 24556 11320 24577 11360
rect 24663 11320 24680 11360
rect 24720 11320 24729 11360
rect 24343 11297 24409 11320
rect 24495 11297 24577 11320
rect 24663 11297 24729 11320
rect 24343 11278 24729 11297
rect 28343 11383 28729 11402
rect 28343 11360 28409 11383
rect 28495 11360 28577 11383
rect 28663 11360 28729 11383
rect 28343 11320 28352 11360
rect 28392 11320 28409 11360
rect 28495 11320 28516 11360
rect 28556 11320 28577 11360
rect 28663 11320 28680 11360
rect 28720 11320 28729 11360
rect 28343 11297 28409 11320
rect 28495 11297 28577 11320
rect 28663 11297 28729 11320
rect 28343 11278 28729 11297
rect 32343 11383 32729 11402
rect 32343 11360 32409 11383
rect 32495 11360 32577 11383
rect 32663 11360 32729 11383
rect 32343 11320 32352 11360
rect 32392 11320 32409 11360
rect 32495 11320 32516 11360
rect 32556 11320 32577 11360
rect 32663 11320 32680 11360
rect 32720 11320 32729 11360
rect 32343 11297 32409 11320
rect 32495 11297 32577 11320
rect 32663 11297 32729 11320
rect 32343 11278 32729 11297
rect 36343 11383 36729 11402
rect 36343 11360 36409 11383
rect 36495 11360 36577 11383
rect 36663 11360 36729 11383
rect 36343 11320 36352 11360
rect 36392 11320 36409 11360
rect 36495 11320 36516 11360
rect 36556 11320 36577 11360
rect 36663 11320 36680 11360
rect 36720 11320 36729 11360
rect 36343 11297 36409 11320
rect 36495 11297 36577 11320
rect 36663 11297 36729 11320
rect 36343 11278 36729 11297
rect 40343 11383 40729 11402
rect 40343 11360 40409 11383
rect 40495 11360 40577 11383
rect 40663 11360 40729 11383
rect 40343 11320 40352 11360
rect 40392 11320 40409 11360
rect 40495 11320 40516 11360
rect 40556 11320 40577 11360
rect 40663 11320 40680 11360
rect 40720 11320 40729 11360
rect 40343 11297 40409 11320
rect 40495 11297 40577 11320
rect 40663 11297 40729 11320
rect 40343 11278 40729 11297
rect 44343 11383 44729 11402
rect 44343 11360 44409 11383
rect 44495 11360 44577 11383
rect 44663 11360 44729 11383
rect 44343 11320 44352 11360
rect 44392 11320 44409 11360
rect 44495 11320 44516 11360
rect 44556 11320 44577 11360
rect 44663 11320 44680 11360
rect 44720 11320 44729 11360
rect 44343 11297 44409 11320
rect 44495 11297 44577 11320
rect 44663 11297 44729 11320
rect 44343 11278 44729 11297
rect 48343 11383 48729 11402
rect 48343 11360 48409 11383
rect 48495 11360 48577 11383
rect 48663 11360 48729 11383
rect 48343 11320 48352 11360
rect 48392 11320 48409 11360
rect 48495 11320 48516 11360
rect 48556 11320 48577 11360
rect 48663 11320 48680 11360
rect 48720 11320 48729 11360
rect 48343 11297 48409 11320
rect 48495 11297 48577 11320
rect 48663 11297 48729 11320
rect 48343 11278 48729 11297
rect 52343 11383 52729 11402
rect 52343 11360 52409 11383
rect 52495 11360 52577 11383
rect 52663 11360 52729 11383
rect 52343 11320 52352 11360
rect 52392 11320 52409 11360
rect 52495 11320 52516 11360
rect 52556 11320 52577 11360
rect 52663 11320 52680 11360
rect 52720 11320 52729 11360
rect 52343 11297 52409 11320
rect 52495 11297 52577 11320
rect 52663 11297 52729 11320
rect 52343 11278 52729 11297
rect 56343 11383 56729 11402
rect 56343 11360 56409 11383
rect 56495 11360 56577 11383
rect 56663 11360 56729 11383
rect 56343 11320 56352 11360
rect 56392 11320 56409 11360
rect 56495 11320 56516 11360
rect 56556 11320 56577 11360
rect 56663 11320 56680 11360
rect 56720 11320 56729 11360
rect 56343 11297 56409 11320
rect 56495 11297 56577 11320
rect 56663 11297 56729 11320
rect 56343 11278 56729 11297
rect 60343 11383 60729 11402
rect 60343 11360 60409 11383
rect 60495 11360 60577 11383
rect 60663 11360 60729 11383
rect 60343 11320 60352 11360
rect 60392 11320 60409 11360
rect 60495 11320 60516 11360
rect 60556 11320 60577 11360
rect 60663 11320 60680 11360
rect 60720 11320 60729 11360
rect 60343 11297 60409 11320
rect 60495 11297 60577 11320
rect 60663 11297 60729 11320
rect 60343 11278 60729 11297
rect 64343 11383 64729 11402
rect 64343 11360 64409 11383
rect 64495 11360 64577 11383
rect 64663 11360 64729 11383
rect 64343 11320 64352 11360
rect 64392 11320 64409 11360
rect 64495 11320 64516 11360
rect 64556 11320 64577 11360
rect 64663 11320 64680 11360
rect 64720 11320 64729 11360
rect 64343 11297 64409 11320
rect 64495 11297 64577 11320
rect 64663 11297 64729 11320
rect 64343 11278 64729 11297
rect 68343 11383 68729 11402
rect 68343 11360 68409 11383
rect 68495 11360 68577 11383
rect 68663 11360 68729 11383
rect 68343 11320 68352 11360
rect 68392 11320 68409 11360
rect 68495 11320 68516 11360
rect 68556 11320 68577 11360
rect 68663 11320 68680 11360
rect 68720 11320 68729 11360
rect 68343 11297 68409 11320
rect 68495 11297 68577 11320
rect 68663 11297 68729 11320
rect 68343 11278 68729 11297
rect 75076 11320 75169 11406
rect 75255 11320 75337 11406
rect 75423 11320 75516 11406
rect 75076 11238 75516 11320
rect 75076 11152 75169 11238
rect 75255 11152 75337 11238
rect 75423 11152 75516 11238
rect 75076 11070 75516 11152
rect 75076 10984 75169 11070
rect 75255 10984 75337 11070
rect 75423 10984 75516 11070
rect 75076 10902 75516 10984
rect 75076 10816 75169 10902
rect 75255 10816 75337 10902
rect 75423 10816 75516 10902
rect 75076 10734 75516 10816
rect 75076 10648 75169 10734
rect 75255 10648 75337 10734
rect 75423 10648 75516 10734
rect 3103 10627 3489 10646
rect 3103 10604 3169 10627
rect 3255 10604 3337 10627
rect 3423 10604 3489 10627
rect 3103 10564 3112 10604
rect 3152 10564 3169 10604
rect 3255 10564 3276 10604
rect 3316 10564 3337 10604
rect 3423 10564 3440 10604
rect 3480 10564 3489 10604
rect 3103 10541 3169 10564
rect 3255 10541 3337 10564
rect 3423 10541 3489 10564
rect 3103 10522 3489 10541
rect 7103 10627 7489 10646
rect 7103 10604 7169 10627
rect 7255 10604 7337 10627
rect 7423 10604 7489 10627
rect 7103 10564 7112 10604
rect 7152 10564 7169 10604
rect 7255 10564 7276 10604
rect 7316 10564 7337 10604
rect 7423 10564 7440 10604
rect 7480 10564 7489 10604
rect 7103 10541 7169 10564
rect 7255 10541 7337 10564
rect 7423 10541 7489 10564
rect 7103 10522 7489 10541
rect 11103 10627 11489 10646
rect 11103 10604 11169 10627
rect 11255 10604 11337 10627
rect 11423 10604 11489 10627
rect 11103 10564 11112 10604
rect 11152 10564 11169 10604
rect 11255 10564 11276 10604
rect 11316 10564 11337 10604
rect 11423 10564 11440 10604
rect 11480 10564 11489 10604
rect 11103 10541 11169 10564
rect 11255 10541 11337 10564
rect 11423 10541 11489 10564
rect 11103 10522 11489 10541
rect 15103 10627 15489 10646
rect 15103 10604 15169 10627
rect 15255 10604 15337 10627
rect 15423 10604 15489 10627
rect 15103 10564 15112 10604
rect 15152 10564 15169 10604
rect 15255 10564 15276 10604
rect 15316 10564 15337 10604
rect 15423 10564 15440 10604
rect 15480 10564 15489 10604
rect 15103 10541 15169 10564
rect 15255 10541 15337 10564
rect 15423 10541 15489 10564
rect 15103 10522 15489 10541
rect 19103 10627 19489 10646
rect 19103 10604 19169 10627
rect 19255 10604 19337 10627
rect 19423 10604 19489 10627
rect 19103 10564 19112 10604
rect 19152 10564 19169 10604
rect 19255 10564 19276 10604
rect 19316 10564 19337 10604
rect 19423 10564 19440 10604
rect 19480 10564 19489 10604
rect 19103 10541 19169 10564
rect 19255 10541 19337 10564
rect 19423 10541 19489 10564
rect 19103 10522 19489 10541
rect 23103 10627 23489 10646
rect 23103 10604 23169 10627
rect 23255 10604 23337 10627
rect 23423 10604 23489 10627
rect 23103 10564 23112 10604
rect 23152 10564 23169 10604
rect 23255 10564 23276 10604
rect 23316 10564 23337 10604
rect 23423 10564 23440 10604
rect 23480 10564 23489 10604
rect 23103 10541 23169 10564
rect 23255 10541 23337 10564
rect 23423 10541 23489 10564
rect 23103 10522 23489 10541
rect 27103 10627 27489 10646
rect 27103 10604 27169 10627
rect 27255 10604 27337 10627
rect 27423 10604 27489 10627
rect 27103 10564 27112 10604
rect 27152 10564 27169 10604
rect 27255 10564 27276 10604
rect 27316 10564 27337 10604
rect 27423 10564 27440 10604
rect 27480 10564 27489 10604
rect 27103 10541 27169 10564
rect 27255 10541 27337 10564
rect 27423 10541 27489 10564
rect 27103 10522 27489 10541
rect 31103 10627 31489 10646
rect 31103 10604 31169 10627
rect 31255 10604 31337 10627
rect 31423 10604 31489 10627
rect 31103 10564 31112 10604
rect 31152 10564 31169 10604
rect 31255 10564 31276 10604
rect 31316 10564 31337 10604
rect 31423 10564 31440 10604
rect 31480 10564 31489 10604
rect 31103 10541 31169 10564
rect 31255 10541 31337 10564
rect 31423 10541 31489 10564
rect 31103 10522 31489 10541
rect 35103 10627 35489 10646
rect 35103 10604 35169 10627
rect 35255 10604 35337 10627
rect 35423 10604 35489 10627
rect 35103 10564 35112 10604
rect 35152 10564 35169 10604
rect 35255 10564 35276 10604
rect 35316 10564 35337 10604
rect 35423 10564 35440 10604
rect 35480 10564 35489 10604
rect 35103 10541 35169 10564
rect 35255 10541 35337 10564
rect 35423 10541 35489 10564
rect 35103 10522 35489 10541
rect 39103 10627 39489 10646
rect 39103 10604 39169 10627
rect 39255 10604 39337 10627
rect 39423 10604 39489 10627
rect 39103 10564 39112 10604
rect 39152 10564 39169 10604
rect 39255 10564 39276 10604
rect 39316 10564 39337 10604
rect 39423 10564 39440 10604
rect 39480 10564 39489 10604
rect 39103 10541 39169 10564
rect 39255 10541 39337 10564
rect 39423 10541 39489 10564
rect 39103 10522 39489 10541
rect 43103 10627 43489 10646
rect 43103 10604 43169 10627
rect 43255 10604 43337 10627
rect 43423 10604 43489 10627
rect 43103 10564 43112 10604
rect 43152 10564 43169 10604
rect 43255 10564 43276 10604
rect 43316 10564 43337 10604
rect 43423 10564 43440 10604
rect 43480 10564 43489 10604
rect 43103 10541 43169 10564
rect 43255 10541 43337 10564
rect 43423 10541 43489 10564
rect 43103 10522 43489 10541
rect 47103 10627 47489 10646
rect 47103 10604 47169 10627
rect 47255 10604 47337 10627
rect 47423 10604 47489 10627
rect 47103 10564 47112 10604
rect 47152 10564 47169 10604
rect 47255 10564 47276 10604
rect 47316 10564 47337 10604
rect 47423 10564 47440 10604
rect 47480 10564 47489 10604
rect 47103 10541 47169 10564
rect 47255 10541 47337 10564
rect 47423 10541 47489 10564
rect 47103 10522 47489 10541
rect 51103 10627 51489 10646
rect 51103 10604 51169 10627
rect 51255 10604 51337 10627
rect 51423 10604 51489 10627
rect 51103 10564 51112 10604
rect 51152 10564 51169 10604
rect 51255 10564 51276 10604
rect 51316 10564 51337 10604
rect 51423 10564 51440 10604
rect 51480 10564 51489 10604
rect 51103 10541 51169 10564
rect 51255 10541 51337 10564
rect 51423 10541 51489 10564
rect 51103 10522 51489 10541
rect 55103 10627 55489 10646
rect 55103 10604 55169 10627
rect 55255 10604 55337 10627
rect 55423 10604 55489 10627
rect 55103 10564 55112 10604
rect 55152 10564 55169 10604
rect 55255 10564 55276 10604
rect 55316 10564 55337 10604
rect 55423 10564 55440 10604
rect 55480 10564 55489 10604
rect 55103 10541 55169 10564
rect 55255 10541 55337 10564
rect 55423 10541 55489 10564
rect 55103 10522 55489 10541
rect 59103 10627 59489 10646
rect 59103 10604 59169 10627
rect 59255 10604 59337 10627
rect 59423 10604 59489 10627
rect 59103 10564 59112 10604
rect 59152 10564 59169 10604
rect 59255 10564 59276 10604
rect 59316 10564 59337 10604
rect 59423 10564 59440 10604
rect 59480 10564 59489 10604
rect 59103 10541 59169 10564
rect 59255 10541 59337 10564
rect 59423 10541 59489 10564
rect 59103 10522 59489 10541
rect 63103 10627 63489 10646
rect 63103 10604 63169 10627
rect 63255 10604 63337 10627
rect 63423 10604 63489 10627
rect 63103 10564 63112 10604
rect 63152 10564 63169 10604
rect 63255 10564 63276 10604
rect 63316 10564 63337 10604
rect 63423 10564 63440 10604
rect 63480 10564 63489 10604
rect 63103 10541 63169 10564
rect 63255 10541 63337 10564
rect 63423 10541 63489 10564
rect 63103 10522 63489 10541
rect 67103 10627 67489 10646
rect 67103 10604 67169 10627
rect 67255 10604 67337 10627
rect 67423 10604 67489 10627
rect 67103 10564 67112 10604
rect 67152 10564 67169 10604
rect 67255 10564 67276 10604
rect 67316 10564 67337 10604
rect 67423 10564 67440 10604
rect 67480 10564 67489 10604
rect 67103 10541 67169 10564
rect 67255 10541 67337 10564
rect 67423 10541 67489 10564
rect 67103 10522 67489 10541
rect 75076 10566 75516 10648
rect 75076 10480 75169 10566
rect 75255 10480 75337 10566
rect 75423 10480 75516 10566
rect 75076 10398 75516 10480
rect 75076 10312 75169 10398
rect 75255 10312 75337 10398
rect 75423 10312 75516 10398
rect 75076 10230 75516 10312
rect 75076 10144 75169 10230
rect 75255 10144 75337 10230
rect 75423 10144 75516 10230
rect 75076 10014 75516 10144
rect 79076 12246 79516 12376
rect 79076 12160 79169 12246
rect 79255 12160 79337 12246
rect 79423 12160 79516 12246
rect 79076 12078 79516 12160
rect 79076 11992 79169 12078
rect 79255 11992 79337 12078
rect 79423 11992 79516 12078
rect 79076 11910 79516 11992
rect 79076 11824 79169 11910
rect 79255 11824 79337 11910
rect 79423 11824 79516 11910
rect 79076 11742 79516 11824
rect 79076 11656 79169 11742
rect 79255 11656 79337 11742
rect 79423 11656 79516 11742
rect 79076 11574 79516 11656
rect 79076 11488 79169 11574
rect 79255 11488 79337 11574
rect 79423 11488 79516 11574
rect 79076 11406 79516 11488
rect 79076 11320 79169 11406
rect 79255 11320 79337 11406
rect 79423 11320 79516 11406
rect 79076 11238 79516 11320
rect 79076 11152 79169 11238
rect 79255 11152 79337 11238
rect 79423 11152 79516 11238
rect 79076 11070 79516 11152
rect 79076 10984 79169 11070
rect 79255 10984 79337 11070
rect 79423 10984 79516 11070
rect 79076 10902 79516 10984
rect 79076 10816 79169 10902
rect 79255 10816 79337 10902
rect 79423 10816 79516 10902
rect 79076 10734 79516 10816
rect 79076 10648 79169 10734
rect 79255 10648 79337 10734
rect 79423 10648 79516 10734
rect 79076 10566 79516 10648
rect 79076 10480 79169 10566
rect 79255 10480 79337 10566
rect 79423 10480 79516 10566
rect 79076 10398 79516 10480
rect 79076 10312 79169 10398
rect 79255 10312 79337 10398
rect 79423 10312 79516 10398
rect 79076 10230 79516 10312
rect 79076 10144 79169 10230
rect 79255 10144 79337 10230
rect 79423 10144 79516 10230
rect 79076 10014 79516 10144
rect 83076 12246 83516 12376
rect 83076 12160 83169 12246
rect 83255 12160 83337 12246
rect 83423 12160 83516 12246
rect 83076 12078 83516 12160
rect 83076 11992 83169 12078
rect 83255 11992 83337 12078
rect 83423 11992 83516 12078
rect 83076 11910 83516 11992
rect 83076 11824 83169 11910
rect 83255 11824 83337 11910
rect 83423 11824 83516 11910
rect 83076 11742 83516 11824
rect 83076 11656 83169 11742
rect 83255 11656 83337 11742
rect 83423 11656 83516 11742
rect 83076 11574 83516 11656
rect 83076 11488 83169 11574
rect 83255 11488 83337 11574
rect 83423 11488 83516 11574
rect 83076 11406 83516 11488
rect 83076 11320 83169 11406
rect 83255 11320 83337 11406
rect 83423 11320 83516 11406
rect 83076 11238 83516 11320
rect 83076 11152 83169 11238
rect 83255 11152 83337 11238
rect 83423 11152 83516 11238
rect 83076 11070 83516 11152
rect 83076 10984 83169 11070
rect 83255 10984 83337 11070
rect 83423 10984 83516 11070
rect 83076 10902 83516 10984
rect 83076 10816 83169 10902
rect 83255 10816 83337 10902
rect 83423 10816 83516 10902
rect 83076 10734 83516 10816
rect 83076 10648 83169 10734
rect 83255 10648 83337 10734
rect 83423 10648 83516 10734
rect 83076 10566 83516 10648
rect 83076 10480 83169 10566
rect 83255 10480 83337 10566
rect 83423 10480 83516 10566
rect 83076 10398 83516 10480
rect 83076 10312 83169 10398
rect 83255 10312 83337 10398
rect 83423 10312 83516 10398
rect 83076 10230 83516 10312
rect 83076 10144 83169 10230
rect 83255 10144 83337 10230
rect 83423 10144 83516 10230
rect 83076 10014 83516 10144
rect 87076 12246 87516 12376
rect 87076 12160 87169 12246
rect 87255 12160 87337 12246
rect 87423 12160 87516 12246
rect 87076 12078 87516 12160
rect 87076 11992 87169 12078
rect 87255 11992 87337 12078
rect 87423 11992 87516 12078
rect 87076 11910 87516 11992
rect 87076 11824 87169 11910
rect 87255 11824 87337 11910
rect 87423 11824 87516 11910
rect 87076 11742 87516 11824
rect 87076 11656 87169 11742
rect 87255 11656 87337 11742
rect 87423 11656 87516 11742
rect 87076 11574 87516 11656
rect 87076 11488 87169 11574
rect 87255 11488 87337 11574
rect 87423 11488 87516 11574
rect 87076 11406 87516 11488
rect 87076 11320 87169 11406
rect 87255 11320 87337 11406
rect 87423 11320 87516 11406
rect 87076 11238 87516 11320
rect 87076 11152 87169 11238
rect 87255 11152 87337 11238
rect 87423 11152 87516 11238
rect 87076 11070 87516 11152
rect 87076 10984 87169 11070
rect 87255 10984 87337 11070
rect 87423 10984 87516 11070
rect 87076 10902 87516 10984
rect 87076 10816 87169 10902
rect 87255 10816 87337 10902
rect 87423 10816 87516 10902
rect 87076 10734 87516 10816
rect 87076 10648 87169 10734
rect 87255 10648 87337 10734
rect 87423 10648 87516 10734
rect 87076 10566 87516 10648
rect 87076 10480 87169 10566
rect 87255 10480 87337 10566
rect 87423 10480 87516 10566
rect 87076 10398 87516 10480
rect 87076 10312 87169 10398
rect 87255 10312 87337 10398
rect 87423 10312 87516 10398
rect 87076 10230 87516 10312
rect 87076 10144 87169 10230
rect 87255 10144 87337 10230
rect 87423 10144 87516 10230
rect 87076 10014 87516 10144
rect 91076 12246 91516 12376
rect 91076 12160 91169 12246
rect 91255 12160 91337 12246
rect 91423 12160 91516 12246
rect 91076 12078 91516 12160
rect 91076 11992 91169 12078
rect 91255 11992 91337 12078
rect 91423 11992 91516 12078
rect 91076 11910 91516 11992
rect 91076 11824 91169 11910
rect 91255 11824 91337 11910
rect 91423 11824 91516 11910
rect 91076 11742 91516 11824
rect 91076 11656 91169 11742
rect 91255 11656 91337 11742
rect 91423 11656 91516 11742
rect 91076 11574 91516 11656
rect 91076 11488 91169 11574
rect 91255 11488 91337 11574
rect 91423 11488 91516 11574
rect 91076 11406 91516 11488
rect 91076 11320 91169 11406
rect 91255 11320 91337 11406
rect 91423 11320 91516 11406
rect 91076 11238 91516 11320
rect 91076 11152 91169 11238
rect 91255 11152 91337 11238
rect 91423 11152 91516 11238
rect 91076 11070 91516 11152
rect 91076 10984 91169 11070
rect 91255 10984 91337 11070
rect 91423 10984 91516 11070
rect 91076 10902 91516 10984
rect 91076 10816 91169 10902
rect 91255 10816 91337 10902
rect 91423 10816 91516 10902
rect 91076 10734 91516 10816
rect 91076 10648 91169 10734
rect 91255 10648 91337 10734
rect 91423 10648 91516 10734
rect 91076 10566 91516 10648
rect 91076 10480 91169 10566
rect 91255 10480 91337 10566
rect 91423 10480 91516 10566
rect 91076 10398 91516 10480
rect 91076 10312 91169 10398
rect 91255 10312 91337 10398
rect 91423 10312 91516 10398
rect 91076 10230 91516 10312
rect 91076 10144 91169 10230
rect 91255 10144 91337 10230
rect 91423 10144 91516 10230
rect 91076 10014 91516 10144
rect 95076 12246 95516 12376
rect 95076 12160 95169 12246
rect 95255 12160 95337 12246
rect 95423 12160 95516 12246
rect 95076 12078 95516 12160
rect 95076 11992 95169 12078
rect 95255 11992 95337 12078
rect 95423 11992 95516 12078
rect 95076 11910 95516 11992
rect 95076 11824 95169 11910
rect 95255 11824 95337 11910
rect 95423 11824 95516 11910
rect 95076 11742 95516 11824
rect 95076 11656 95169 11742
rect 95255 11656 95337 11742
rect 95423 11656 95516 11742
rect 95076 11574 95516 11656
rect 95076 11488 95169 11574
rect 95255 11488 95337 11574
rect 95423 11488 95516 11574
rect 95076 11406 95516 11488
rect 95076 11320 95169 11406
rect 95255 11320 95337 11406
rect 95423 11320 95516 11406
rect 95076 11238 95516 11320
rect 95076 11152 95169 11238
rect 95255 11152 95337 11238
rect 95423 11152 95516 11238
rect 95076 11070 95516 11152
rect 95076 10984 95169 11070
rect 95255 10984 95337 11070
rect 95423 10984 95516 11070
rect 95076 10902 95516 10984
rect 95076 10816 95169 10902
rect 95255 10816 95337 10902
rect 95423 10816 95516 10902
rect 95076 10734 95516 10816
rect 95076 10648 95169 10734
rect 95255 10648 95337 10734
rect 95423 10648 95516 10734
rect 95076 10566 95516 10648
rect 95076 10480 95169 10566
rect 95255 10480 95337 10566
rect 95423 10480 95516 10566
rect 95076 10398 95516 10480
rect 95076 10312 95169 10398
rect 95255 10312 95337 10398
rect 95423 10312 95516 10398
rect 95076 10230 95516 10312
rect 95076 10144 95169 10230
rect 95255 10144 95337 10230
rect 95423 10144 95516 10230
rect 95076 10014 95516 10144
rect 4343 9871 4729 9890
rect 4343 9848 4409 9871
rect 4495 9848 4577 9871
rect 4663 9848 4729 9871
rect 4343 9808 4352 9848
rect 4392 9808 4409 9848
rect 4495 9808 4516 9848
rect 4556 9808 4577 9848
rect 4663 9808 4680 9848
rect 4720 9808 4729 9848
rect 4343 9785 4409 9808
rect 4495 9785 4577 9808
rect 4663 9785 4729 9808
rect 4343 9766 4729 9785
rect 8343 9871 8729 9890
rect 8343 9848 8409 9871
rect 8495 9848 8577 9871
rect 8663 9848 8729 9871
rect 8343 9808 8352 9848
rect 8392 9808 8409 9848
rect 8495 9808 8516 9848
rect 8556 9808 8577 9848
rect 8663 9808 8680 9848
rect 8720 9808 8729 9848
rect 8343 9785 8409 9808
rect 8495 9785 8577 9808
rect 8663 9785 8729 9808
rect 8343 9766 8729 9785
rect 12343 9871 12729 9890
rect 12343 9848 12409 9871
rect 12495 9848 12577 9871
rect 12663 9848 12729 9871
rect 12343 9808 12352 9848
rect 12392 9808 12409 9848
rect 12495 9808 12516 9848
rect 12556 9808 12577 9848
rect 12663 9808 12680 9848
rect 12720 9808 12729 9848
rect 12343 9785 12409 9808
rect 12495 9785 12577 9808
rect 12663 9785 12729 9808
rect 12343 9766 12729 9785
rect 16343 9871 16729 9890
rect 16343 9848 16409 9871
rect 16495 9848 16577 9871
rect 16663 9848 16729 9871
rect 16343 9808 16352 9848
rect 16392 9808 16409 9848
rect 16495 9808 16516 9848
rect 16556 9808 16577 9848
rect 16663 9808 16680 9848
rect 16720 9808 16729 9848
rect 16343 9785 16409 9808
rect 16495 9785 16577 9808
rect 16663 9785 16729 9808
rect 16343 9766 16729 9785
rect 20343 9871 20729 9890
rect 20343 9848 20409 9871
rect 20495 9848 20577 9871
rect 20663 9848 20729 9871
rect 20343 9808 20352 9848
rect 20392 9808 20409 9848
rect 20495 9808 20516 9848
rect 20556 9808 20577 9848
rect 20663 9808 20680 9848
rect 20720 9808 20729 9848
rect 20343 9785 20409 9808
rect 20495 9785 20577 9808
rect 20663 9785 20729 9808
rect 20343 9766 20729 9785
rect 24343 9871 24729 9890
rect 24343 9848 24409 9871
rect 24495 9848 24577 9871
rect 24663 9848 24729 9871
rect 24343 9808 24352 9848
rect 24392 9808 24409 9848
rect 24495 9808 24516 9848
rect 24556 9808 24577 9848
rect 24663 9808 24680 9848
rect 24720 9808 24729 9848
rect 24343 9785 24409 9808
rect 24495 9785 24577 9808
rect 24663 9785 24729 9808
rect 24343 9766 24729 9785
rect 28343 9871 28729 9890
rect 28343 9848 28409 9871
rect 28495 9848 28577 9871
rect 28663 9848 28729 9871
rect 28343 9808 28352 9848
rect 28392 9808 28409 9848
rect 28495 9808 28516 9848
rect 28556 9808 28577 9848
rect 28663 9808 28680 9848
rect 28720 9808 28729 9848
rect 28343 9785 28409 9808
rect 28495 9785 28577 9808
rect 28663 9785 28729 9808
rect 28343 9766 28729 9785
rect 32343 9871 32729 9890
rect 32343 9848 32409 9871
rect 32495 9848 32577 9871
rect 32663 9848 32729 9871
rect 32343 9808 32352 9848
rect 32392 9808 32409 9848
rect 32495 9808 32516 9848
rect 32556 9808 32577 9848
rect 32663 9808 32680 9848
rect 32720 9808 32729 9848
rect 32343 9785 32409 9808
rect 32495 9785 32577 9808
rect 32663 9785 32729 9808
rect 32343 9766 32729 9785
rect 36343 9871 36729 9890
rect 36343 9848 36409 9871
rect 36495 9848 36577 9871
rect 36663 9848 36729 9871
rect 36343 9808 36352 9848
rect 36392 9808 36409 9848
rect 36495 9808 36516 9848
rect 36556 9808 36577 9848
rect 36663 9808 36680 9848
rect 36720 9808 36729 9848
rect 36343 9785 36409 9808
rect 36495 9785 36577 9808
rect 36663 9785 36729 9808
rect 36343 9766 36729 9785
rect 40343 9871 40729 9890
rect 40343 9848 40409 9871
rect 40495 9848 40577 9871
rect 40663 9848 40729 9871
rect 40343 9808 40352 9848
rect 40392 9808 40409 9848
rect 40495 9808 40516 9848
rect 40556 9808 40577 9848
rect 40663 9808 40680 9848
rect 40720 9808 40729 9848
rect 40343 9785 40409 9808
rect 40495 9785 40577 9808
rect 40663 9785 40729 9808
rect 40343 9766 40729 9785
rect 44343 9871 44729 9890
rect 44343 9848 44409 9871
rect 44495 9848 44577 9871
rect 44663 9848 44729 9871
rect 44343 9808 44352 9848
rect 44392 9808 44409 9848
rect 44495 9808 44516 9848
rect 44556 9808 44577 9848
rect 44663 9808 44680 9848
rect 44720 9808 44729 9848
rect 44343 9785 44409 9808
rect 44495 9785 44577 9808
rect 44663 9785 44729 9808
rect 44343 9766 44729 9785
rect 48343 9871 48729 9890
rect 48343 9848 48409 9871
rect 48495 9848 48577 9871
rect 48663 9848 48729 9871
rect 48343 9808 48352 9848
rect 48392 9808 48409 9848
rect 48495 9808 48516 9848
rect 48556 9808 48577 9848
rect 48663 9808 48680 9848
rect 48720 9808 48729 9848
rect 48343 9785 48409 9808
rect 48495 9785 48577 9808
rect 48663 9785 48729 9808
rect 48343 9766 48729 9785
rect 52343 9871 52729 9890
rect 52343 9848 52409 9871
rect 52495 9848 52577 9871
rect 52663 9848 52729 9871
rect 52343 9808 52352 9848
rect 52392 9808 52409 9848
rect 52495 9808 52516 9848
rect 52556 9808 52577 9848
rect 52663 9808 52680 9848
rect 52720 9808 52729 9848
rect 52343 9785 52409 9808
rect 52495 9785 52577 9808
rect 52663 9785 52729 9808
rect 52343 9766 52729 9785
rect 56343 9871 56729 9890
rect 56343 9848 56409 9871
rect 56495 9848 56577 9871
rect 56663 9848 56729 9871
rect 56343 9808 56352 9848
rect 56392 9808 56409 9848
rect 56495 9808 56516 9848
rect 56556 9808 56577 9848
rect 56663 9808 56680 9848
rect 56720 9808 56729 9848
rect 56343 9785 56409 9808
rect 56495 9785 56577 9808
rect 56663 9785 56729 9808
rect 56343 9766 56729 9785
rect 60343 9871 60729 9890
rect 60343 9848 60409 9871
rect 60495 9848 60577 9871
rect 60663 9848 60729 9871
rect 60343 9808 60352 9848
rect 60392 9808 60409 9848
rect 60495 9808 60516 9848
rect 60556 9808 60577 9848
rect 60663 9808 60680 9848
rect 60720 9808 60729 9848
rect 60343 9785 60409 9808
rect 60495 9785 60577 9808
rect 60663 9785 60729 9808
rect 60343 9766 60729 9785
rect 64343 9871 64729 9890
rect 64343 9848 64409 9871
rect 64495 9848 64577 9871
rect 64663 9848 64729 9871
rect 64343 9808 64352 9848
rect 64392 9808 64409 9848
rect 64495 9808 64516 9848
rect 64556 9808 64577 9848
rect 64663 9808 64680 9848
rect 64720 9808 64729 9848
rect 64343 9785 64409 9808
rect 64495 9785 64577 9808
rect 64663 9785 64729 9808
rect 64343 9766 64729 9785
rect 68343 9871 68729 9890
rect 68343 9848 68409 9871
rect 68495 9848 68577 9871
rect 68663 9848 68729 9871
rect 68343 9808 68352 9848
rect 68392 9808 68409 9848
rect 68495 9808 68516 9848
rect 68556 9808 68577 9848
rect 68663 9808 68680 9848
rect 68720 9808 68729 9848
rect 68343 9785 68409 9808
rect 68495 9785 68577 9808
rect 68663 9785 68729 9808
rect 68343 9766 68729 9785
rect 3103 9115 3489 9134
rect 3103 9092 3169 9115
rect 3255 9092 3337 9115
rect 3423 9092 3489 9115
rect 3103 9052 3112 9092
rect 3152 9052 3169 9092
rect 3255 9052 3276 9092
rect 3316 9052 3337 9092
rect 3423 9052 3440 9092
rect 3480 9052 3489 9092
rect 3103 9029 3169 9052
rect 3255 9029 3337 9052
rect 3423 9029 3489 9052
rect 3103 9010 3489 9029
rect 7103 9115 7489 9134
rect 7103 9092 7169 9115
rect 7255 9092 7337 9115
rect 7423 9092 7489 9115
rect 7103 9052 7112 9092
rect 7152 9052 7169 9092
rect 7255 9052 7276 9092
rect 7316 9052 7337 9092
rect 7423 9052 7440 9092
rect 7480 9052 7489 9092
rect 7103 9029 7169 9052
rect 7255 9029 7337 9052
rect 7423 9029 7489 9052
rect 7103 9010 7489 9029
rect 11103 9115 11489 9134
rect 11103 9092 11169 9115
rect 11255 9092 11337 9115
rect 11423 9092 11489 9115
rect 11103 9052 11112 9092
rect 11152 9052 11169 9092
rect 11255 9052 11276 9092
rect 11316 9052 11337 9092
rect 11423 9052 11440 9092
rect 11480 9052 11489 9092
rect 11103 9029 11169 9052
rect 11255 9029 11337 9052
rect 11423 9029 11489 9052
rect 11103 9010 11489 9029
rect 15103 9115 15489 9134
rect 15103 9092 15169 9115
rect 15255 9092 15337 9115
rect 15423 9092 15489 9115
rect 15103 9052 15112 9092
rect 15152 9052 15169 9092
rect 15255 9052 15276 9092
rect 15316 9052 15337 9092
rect 15423 9052 15440 9092
rect 15480 9052 15489 9092
rect 15103 9029 15169 9052
rect 15255 9029 15337 9052
rect 15423 9029 15489 9052
rect 15103 9010 15489 9029
rect 19103 9115 19489 9134
rect 19103 9092 19169 9115
rect 19255 9092 19337 9115
rect 19423 9092 19489 9115
rect 19103 9052 19112 9092
rect 19152 9052 19169 9092
rect 19255 9052 19276 9092
rect 19316 9052 19337 9092
rect 19423 9052 19440 9092
rect 19480 9052 19489 9092
rect 19103 9029 19169 9052
rect 19255 9029 19337 9052
rect 19423 9029 19489 9052
rect 19103 9010 19489 9029
rect 23103 9115 23489 9134
rect 23103 9092 23169 9115
rect 23255 9092 23337 9115
rect 23423 9092 23489 9115
rect 23103 9052 23112 9092
rect 23152 9052 23169 9092
rect 23255 9052 23276 9092
rect 23316 9052 23337 9092
rect 23423 9052 23440 9092
rect 23480 9052 23489 9092
rect 23103 9029 23169 9052
rect 23255 9029 23337 9052
rect 23423 9029 23489 9052
rect 23103 9010 23489 9029
rect 27103 9115 27489 9134
rect 27103 9092 27169 9115
rect 27255 9092 27337 9115
rect 27423 9092 27489 9115
rect 27103 9052 27112 9092
rect 27152 9052 27169 9092
rect 27255 9052 27276 9092
rect 27316 9052 27337 9092
rect 27423 9052 27440 9092
rect 27480 9052 27489 9092
rect 27103 9029 27169 9052
rect 27255 9029 27337 9052
rect 27423 9029 27489 9052
rect 27103 9010 27489 9029
rect 31103 9115 31489 9134
rect 31103 9092 31169 9115
rect 31255 9092 31337 9115
rect 31423 9092 31489 9115
rect 31103 9052 31112 9092
rect 31152 9052 31169 9092
rect 31255 9052 31276 9092
rect 31316 9052 31337 9092
rect 31423 9052 31440 9092
rect 31480 9052 31489 9092
rect 31103 9029 31169 9052
rect 31255 9029 31337 9052
rect 31423 9029 31489 9052
rect 31103 9010 31489 9029
rect 35103 9115 35489 9134
rect 35103 9092 35169 9115
rect 35255 9092 35337 9115
rect 35423 9092 35489 9115
rect 35103 9052 35112 9092
rect 35152 9052 35169 9092
rect 35255 9052 35276 9092
rect 35316 9052 35337 9092
rect 35423 9052 35440 9092
rect 35480 9052 35489 9092
rect 35103 9029 35169 9052
rect 35255 9029 35337 9052
rect 35423 9029 35489 9052
rect 35103 9010 35489 9029
rect 39103 9115 39489 9134
rect 39103 9092 39169 9115
rect 39255 9092 39337 9115
rect 39423 9092 39489 9115
rect 39103 9052 39112 9092
rect 39152 9052 39169 9092
rect 39255 9052 39276 9092
rect 39316 9052 39337 9092
rect 39423 9052 39440 9092
rect 39480 9052 39489 9092
rect 39103 9029 39169 9052
rect 39255 9029 39337 9052
rect 39423 9029 39489 9052
rect 39103 9010 39489 9029
rect 43103 9115 43489 9134
rect 43103 9092 43169 9115
rect 43255 9092 43337 9115
rect 43423 9092 43489 9115
rect 43103 9052 43112 9092
rect 43152 9052 43169 9092
rect 43255 9052 43276 9092
rect 43316 9052 43337 9092
rect 43423 9052 43440 9092
rect 43480 9052 43489 9092
rect 43103 9029 43169 9052
rect 43255 9029 43337 9052
rect 43423 9029 43489 9052
rect 43103 9010 43489 9029
rect 47103 9115 47489 9134
rect 47103 9092 47169 9115
rect 47255 9092 47337 9115
rect 47423 9092 47489 9115
rect 47103 9052 47112 9092
rect 47152 9052 47169 9092
rect 47255 9052 47276 9092
rect 47316 9052 47337 9092
rect 47423 9052 47440 9092
rect 47480 9052 47489 9092
rect 47103 9029 47169 9052
rect 47255 9029 47337 9052
rect 47423 9029 47489 9052
rect 47103 9010 47489 9029
rect 51103 9115 51489 9134
rect 51103 9092 51169 9115
rect 51255 9092 51337 9115
rect 51423 9092 51489 9115
rect 51103 9052 51112 9092
rect 51152 9052 51169 9092
rect 51255 9052 51276 9092
rect 51316 9052 51337 9092
rect 51423 9052 51440 9092
rect 51480 9052 51489 9092
rect 51103 9029 51169 9052
rect 51255 9029 51337 9052
rect 51423 9029 51489 9052
rect 51103 9010 51489 9029
rect 55103 9115 55489 9134
rect 55103 9092 55169 9115
rect 55255 9092 55337 9115
rect 55423 9092 55489 9115
rect 55103 9052 55112 9092
rect 55152 9052 55169 9092
rect 55255 9052 55276 9092
rect 55316 9052 55337 9092
rect 55423 9052 55440 9092
rect 55480 9052 55489 9092
rect 55103 9029 55169 9052
rect 55255 9029 55337 9052
rect 55423 9029 55489 9052
rect 55103 9010 55489 9029
rect 59103 9115 59489 9134
rect 59103 9092 59169 9115
rect 59255 9092 59337 9115
rect 59423 9092 59489 9115
rect 59103 9052 59112 9092
rect 59152 9052 59169 9092
rect 59255 9052 59276 9092
rect 59316 9052 59337 9092
rect 59423 9052 59440 9092
rect 59480 9052 59489 9092
rect 59103 9029 59169 9052
rect 59255 9029 59337 9052
rect 59423 9029 59489 9052
rect 59103 9010 59489 9029
rect 63103 9115 63489 9134
rect 63103 9092 63169 9115
rect 63255 9092 63337 9115
rect 63423 9092 63489 9115
rect 63103 9052 63112 9092
rect 63152 9052 63169 9092
rect 63255 9052 63276 9092
rect 63316 9052 63337 9092
rect 63423 9052 63440 9092
rect 63480 9052 63489 9092
rect 63103 9029 63169 9052
rect 63255 9029 63337 9052
rect 63423 9029 63489 9052
rect 63103 9010 63489 9029
rect 67103 9115 67489 9134
rect 67103 9092 67169 9115
rect 67255 9092 67337 9115
rect 67423 9092 67489 9115
rect 67103 9052 67112 9092
rect 67152 9052 67169 9092
rect 67255 9052 67276 9092
rect 67316 9052 67337 9092
rect 67423 9052 67440 9092
rect 67480 9052 67489 9092
rect 67103 9029 67169 9052
rect 67255 9029 67337 9052
rect 67423 9029 67489 9052
rect 67103 9010 67489 9029
rect 4343 8359 4729 8378
rect 4343 8336 4409 8359
rect 4495 8336 4577 8359
rect 4663 8336 4729 8359
rect 4343 8296 4352 8336
rect 4392 8296 4409 8336
rect 4495 8296 4516 8336
rect 4556 8296 4577 8336
rect 4663 8296 4680 8336
rect 4720 8296 4729 8336
rect 4343 8273 4409 8296
rect 4495 8273 4577 8296
rect 4663 8273 4729 8296
rect 4343 8254 4729 8273
rect 8343 8359 8729 8378
rect 8343 8336 8409 8359
rect 8495 8336 8577 8359
rect 8663 8336 8729 8359
rect 8343 8296 8352 8336
rect 8392 8296 8409 8336
rect 8495 8296 8516 8336
rect 8556 8296 8577 8336
rect 8663 8296 8680 8336
rect 8720 8296 8729 8336
rect 8343 8273 8409 8296
rect 8495 8273 8577 8296
rect 8663 8273 8729 8296
rect 8343 8254 8729 8273
rect 12343 8359 12729 8378
rect 12343 8336 12409 8359
rect 12495 8336 12577 8359
rect 12663 8336 12729 8359
rect 12343 8296 12352 8336
rect 12392 8296 12409 8336
rect 12495 8296 12516 8336
rect 12556 8296 12577 8336
rect 12663 8296 12680 8336
rect 12720 8296 12729 8336
rect 12343 8273 12409 8296
rect 12495 8273 12577 8296
rect 12663 8273 12729 8296
rect 12343 8254 12729 8273
rect 16343 8359 16729 8378
rect 16343 8336 16409 8359
rect 16495 8336 16577 8359
rect 16663 8336 16729 8359
rect 16343 8296 16352 8336
rect 16392 8296 16409 8336
rect 16495 8296 16516 8336
rect 16556 8296 16577 8336
rect 16663 8296 16680 8336
rect 16720 8296 16729 8336
rect 16343 8273 16409 8296
rect 16495 8273 16577 8296
rect 16663 8273 16729 8296
rect 16343 8254 16729 8273
rect 20343 8359 20729 8378
rect 20343 8336 20409 8359
rect 20495 8336 20577 8359
rect 20663 8336 20729 8359
rect 20343 8296 20352 8336
rect 20392 8296 20409 8336
rect 20495 8296 20516 8336
rect 20556 8296 20577 8336
rect 20663 8296 20680 8336
rect 20720 8296 20729 8336
rect 20343 8273 20409 8296
rect 20495 8273 20577 8296
rect 20663 8273 20729 8296
rect 20343 8254 20729 8273
rect 24343 8359 24729 8378
rect 24343 8336 24409 8359
rect 24495 8336 24577 8359
rect 24663 8336 24729 8359
rect 24343 8296 24352 8336
rect 24392 8296 24409 8336
rect 24495 8296 24516 8336
rect 24556 8296 24577 8336
rect 24663 8296 24680 8336
rect 24720 8296 24729 8336
rect 24343 8273 24409 8296
rect 24495 8273 24577 8296
rect 24663 8273 24729 8296
rect 24343 8254 24729 8273
rect 28343 8359 28729 8378
rect 28343 8336 28409 8359
rect 28495 8336 28577 8359
rect 28663 8336 28729 8359
rect 28343 8296 28352 8336
rect 28392 8296 28409 8336
rect 28495 8296 28516 8336
rect 28556 8296 28577 8336
rect 28663 8296 28680 8336
rect 28720 8296 28729 8336
rect 28343 8273 28409 8296
rect 28495 8273 28577 8296
rect 28663 8273 28729 8296
rect 28343 8254 28729 8273
rect 32343 8359 32729 8378
rect 32343 8336 32409 8359
rect 32495 8336 32577 8359
rect 32663 8336 32729 8359
rect 32343 8296 32352 8336
rect 32392 8296 32409 8336
rect 32495 8296 32516 8336
rect 32556 8296 32577 8336
rect 32663 8296 32680 8336
rect 32720 8296 32729 8336
rect 32343 8273 32409 8296
rect 32495 8273 32577 8296
rect 32663 8273 32729 8296
rect 32343 8254 32729 8273
rect 36343 8359 36729 8378
rect 36343 8336 36409 8359
rect 36495 8336 36577 8359
rect 36663 8336 36729 8359
rect 36343 8296 36352 8336
rect 36392 8296 36409 8336
rect 36495 8296 36516 8336
rect 36556 8296 36577 8336
rect 36663 8296 36680 8336
rect 36720 8296 36729 8336
rect 36343 8273 36409 8296
rect 36495 8273 36577 8296
rect 36663 8273 36729 8296
rect 36343 8254 36729 8273
rect 40343 8359 40729 8378
rect 40343 8336 40409 8359
rect 40495 8336 40577 8359
rect 40663 8336 40729 8359
rect 40343 8296 40352 8336
rect 40392 8296 40409 8336
rect 40495 8296 40516 8336
rect 40556 8296 40577 8336
rect 40663 8296 40680 8336
rect 40720 8296 40729 8336
rect 40343 8273 40409 8296
rect 40495 8273 40577 8296
rect 40663 8273 40729 8296
rect 40343 8254 40729 8273
rect 44343 8359 44729 8378
rect 44343 8336 44409 8359
rect 44495 8336 44577 8359
rect 44663 8336 44729 8359
rect 44343 8296 44352 8336
rect 44392 8296 44409 8336
rect 44495 8296 44516 8336
rect 44556 8296 44577 8336
rect 44663 8296 44680 8336
rect 44720 8296 44729 8336
rect 44343 8273 44409 8296
rect 44495 8273 44577 8296
rect 44663 8273 44729 8296
rect 44343 8254 44729 8273
rect 48343 8359 48729 8378
rect 48343 8336 48409 8359
rect 48495 8336 48577 8359
rect 48663 8336 48729 8359
rect 48343 8296 48352 8336
rect 48392 8296 48409 8336
rect 48495 8296 48516 8336
rect 48556 8296 48577 8336
rect 48663 8296 48680 8336
rect 48720 8296 48729 8336
rect 48343 8273 48409 8296
rect 48495 8273 48577 8296
rect 48663 8273 48729 8296
rect 48343 8254 48729 8273
rect 52343 8359 52729 8378
rect 52343 8336 52409 8359
rect 52495 8336 52577 8359
rect 52663 8336 52729 8359
rect 52343 8296 52352 8336
rect 52392 8296 52409 8336
rect 52495 8296 52516 8336
rect 52556 8296 52577 8336
rect 52663 8296 52680 8336
rect 52720 8296 52729 8336
rect 52343 8273 52409 8296
rect 52495 8273 52577 8296
rect 52663 8273 52729 8296
rect 52343 8254 52729 8273
rect 56343 8359 56729 8378
rect 56343 8336 56409 8359
rect 56495 8336 56577 8359
rect 56663 8336 56729 8359
rect 56343 8296 56352 8336
rect 56392 8296 56409 8336
rect 56495 8296 56516 8336
rect 56556 8296 56577 8336
rect 56663 8296 56680 8336
rect 56720 8296 56729 8336
rect 56343 8273 56409 8296
rect 56495 8273 56577 8296
rect 56663 8273 56729 8296
rect 56343 8254 56729 8273
rect 60343 8359 60729 8378
rect 60343 8336 60409 8359
rect 60495 8336 60577 8359
rect 60663 8336 60729 8359
rect 60343 8296 60352 8336
rect 60392 8296 60409 8336
rect 60495 8296 60516 8336
rect 60556 8296 60577 8336
rect 60663 8296 60680 8336
rect 60720 8296 60729 8336
rect 60343 8273 60409 8296
rect 60495 8273 60577 8296
rect 60663 8273 60729 8296
rect 60343 8254 60729 8273
rect 64343 8359 64729 8378
rect 64343 8336 64409 8359
rect 64495 8336 64577 8359
rect 64663 8336 64729 8359
rect 64343 8296 64352 8336
rect 64392 8296 64409 8336
rect 64495 8296 64516 8336
rect 64556 8296 64577 8336
rect 64663 8296 64680 8336
rect 64720 8296 64729 8336
rect 64343 8273 64409 8296
rect 64495 8273 64577 8296
rect 64663 8273 64729 8296
rect 64343 8254 64729 8273
rect 68343 8359 68729 8378
rect 68343 8336 68409 8359
rect 68495 8336 68577 8359
rect 68663 8336 68729 8359
rect 68343 8296 68352 8336
rect 68392 8296 68409 8336
rect 68495 8296 68516 8336
rect 68556 8296 68577 8336
rect 68663 8296 68680 8336
rect 68720 8296 68729 8336
rect 68343 8273 68409 8296
rect 68495 8273 68577 8296
rect 68663 8273 68729 8296
rect 68343 8254 68729 8273
rect 3103 7603 3489 7622
rect 3103 7580 3169 7603
rect 3255 7580 3337 7603
rect 3423 7580 3489 7603
rect 3103 7540 3112 7580
rect 3152 7540 3169 7580
rect 3255 7540 3276 7580
rect 3316 7540 3337 7580
rect 3423 7540 3440 7580
rect 3480 7540 3489 7580
rect 3103 7517 3169 7540
rect 3255 7517 3337 7540
rect 3423 7517 3489 7540
rect 3103 7498 3489 7517
rect 7103 7603 7489 7622
rect 7103 7580 7169 7603
rect 7255 7580 7337 7603
rect 7423 7580 7489 7603
rect 7103 7540 7112 7580
rect 7152 7540 7169 7580
rect 7255 7540 7276 7580
rect 7316 7540 7337 7580
rect 7423 7540 7440 7580
rect 7480 7540 7489 7580
rect 7103 7517 7169 7540
rect 7255 7517 7337 7540
rect 7423 7517 7489 7540
rect 7103 7498 7489 7517
rect 11103 7603 11489 7622
rect 11103 7580 11169 7603
rect 11255 7580 11337 7603
rect 11423 7580 11489 7603
rect 11103 7540 11112 7580
rect 11152 7540 11169 7580
rect 11255 7540 11276 7580
rect 11316 7540 11337 7580
rect 11423 7540 11440 7580
rect 11480 7540 11489 7580
rect 11103 7517 11169 7540
rect 11255 7517 11337 7540
rect 11423 7517 11489 7540
rect 11103 7498 11489 7517
rect 15103 7603 15489 7622
rect 15103 7580 15169 7603
rect 15255 7580 15337 7603
rect 15423 7580 15489 7603
rect 15103 7540 15112 7580
rect 15152 7540 15169 7580
rect 15255 7540 15276 7580
rect 15316 7540 15337 7580
rect 15423 7540 15440 7580
rect 15480 7540 15489 7580
rect 15103 7517 15169 7540
rect 15255 7517 15337 7540
rect 15423 7517 15489 7540
rect 15103 7498 15489 7517
rect 19103 7603 19489 7622
rect 19103 7580 19169 7603
rect 19255 7580 19337 7603
rect 19423 7580 19489 7603
rect 19103 7540 19112 7580
rect 19152 7540 19169 7580
rect 19255 7540 19276 7580
rect 19316 7540 19337 7580
rect 19423 7540 19440 7580
rect 19480 7540 19489 7580
rect 19103 7517 19169 7540
rect 19255 7517 19337 7540
rect 19423 7517 19489 7540
rect 19103 7498 19489 7517
rect 23103 7603 23489 7622
rect 23103 7580 23169 7603
rect 23255 7580 23337 7603
rect 23423 7580 23489 7603
rect 23103 7540 23112 7580
rect 23152 7540 23169 7580
rect 23255 7540 23276 7580
rect 23316 7540 23337 7580
rect 23423 7540 23440 7580
rect 23480 7540 23489 7580
rect 23103 7517 23169 7540
rect 23255 7517 23337 7540
rect 23423 7517 23489 7540
rect 23103 7498 23489 7517
rect 27103 7603 27489 7622
rect 27103 7580 27169 7603
rect 27255 7580 27337 7603
rect 27423 7580 27489 7603
rect 27103 7540 27112 7580
rect 27152 7540 27169 7580
rect 27255 7540 27276 7580
rect 27316 7540 27337 7580
rect 27423 7540 27440 7580
rect 27480 7540 27489 7580
rect 27103 7517 27169 7540
rect 27255 7517 27337 7540
rect 27423 7517 27489 7540
rect 27103 7498 27489 7517
rect 31103 7603 31489 7622
rect 31103 7580 31169 7603
rect 31255 7580 31337 7603
rect 31423 7580 31489 7603
rect 31103 7540 31112 7580
rect 31152 7540 31169 7580
rect 31255 7540 31276 7580
rect 31316 7540 31337 7580
rect 31423 7540 31440 7580
rect 31480 7540 31489 7580
rect 31103 7517 31169 7540
rect 31255 7517 31337 7540
rect 31423 7517 31489 7540
rect 31103 7498 31489 7517
rect 35103 7603 35489 7622
rect 35103 7580 35169 7603
rect 35255 7580 35337 7603
rect 35423 7580 35489 7603
rect 35103 7540 35112 7580
rect 35152 7540 35169 7580
rect 35255 7540 35276 7580
rect 35316 7540 35337 7580
rect 35423 7540 35440 7580
rect 35480 7540 35489 7580
rect 35103 7517 35169 7540
rect 35255 7517 35337 7540
rect 35423 7517 35489 7540
rect 35103 7498 35489 7517
rect 39103 7603 39489 7622
rect 39103 7580 39169 7603
rect 39255 7580 39337 7603
rect 39423 7580 39489 7603
rect 39103 7540 39112 7580
rect 39152 7540 39169 7580
rect 39255 7540 39276 7580
rect 39316 7540 39337 7580
rect 39423 7540 39440 7580
rect 39480 7540 39489 7580
rect 39103 7517 39169 7540
rect 39255 7517 39337 7540
rect 39423 7517 39489 7540
rect 39103 7498 39489 7517
rect 43103 7603 43489 7622
rect 43103 7580 43169 7603
rect 43255 7580 43337 7603
rect 43423 7580 43489 7603
rect 43103 7540 43112 7580
rect 43152 7540 43169 7580
rect 43255 7540 43276 7580
rect 43316 7540 43337 7580
rect 43423 7540 43440 7580
rect 43480 7540 43489 7580
rect 43103 7517 43169 7540
rect 43255 7517 43337 7540
rect 43423 7517 43489 7540
rect 43103 7498 43489 7517
rect 47103 7603 47489 7622
rect 47103 7580 47169 7603
rect 47255 7580 47337 7603
rect 47423 7580 47489 7603
rect 47103 7540 47112 7580
rect 47152 7540 47169 7580
rect 47255 7540 47276 7580
rect 47316 7540 47337 7580
rect 47423 7540 47440 7580
rect 47480 7540 47489 7580
rect 47103 7517 47169 7540
rect 47255 7517 47337 7540
rect 47423 7517 47489 7540
rect 47103 7498 47489 7517
rect 51103 7603 51489 7622
rect 51103 7580 51169 7603
rect 51255 7580 51337 7603
rect 51423 7580 51489 7603
rect 51103 7540 51112 7580
rect 51152 7540 51169 7580
rect 51255 7540 51276 7580
rect 51316 7540 51337 7580
rect 51423 7540 51440 7580
rect 51480 7540 51489 7580
rect 51103 7517 51169 7540
rect 51255 7517 51337 7540
rect 51423 7517 51489 7540
rect 51103 7498 51489 7517
rect 55103 7603 55489 7622
rect 55103 7580 55169 7603
rect 55255 7580 55337 7603
rect 55423 7580 55489 7603
rect 55103 7540 55112 7580
rect 55152 7540 55169 7580
rect 55255 7540 55276 7580
rect 55316 7540 55337 7580
rect 55423 7540 55440 7580
rect 55480 7540 55489 7580
rect 55103 7517 55169 7540
rect 55255 7517 55337 7540
rect 55423 7517 55489 7540
rect 55103 7498 55489 7517
rect 59103 7603 59489 7622
rect 59103 7580 59169 7603
rect 59255 7580 59337 7603
rect 59423 7580 59489 7603
rect 59103 7540 59112 7580
rect 59152 7540 59169 7580
rect 59255 7540 59276 7580
rect 59316 7540 59337 7580
rect 59423 7540 59440 7580
rect 59480 7540 59489 7580
rect 59103 7517 59169 7540
rect 59255 7517 59337 7540
rect 59423 7517 59489 7540
rect 59103 7498 59489 7517
rect 63103 7603 63489 7622
rect 63103 7580 63169 7603
rect 63255 7580 63337 7603
rect 63423 7580 63489 7603
rect 63103 7540 63112 7580
rect 63152 7540 63169 7580
rect 63255 7540 63276 7580
rect 63316 7540 63337 7580
rect 63423 7540 63440 7580
rect 63480 7540 63489 7580
rect 63103 7517 63169 7540
rect 63255 7517 63337 7540
rect 63423 7517 63489 7540
rect 63103 7498 63489 7517
rect 67103 7603 67489 7622
rect 67103 7580 67169 7603
rect 67255 7580 67337 7603
rect 67423 7580 67489 7603
rect 67103 7540 67112 7580
rect 67152 7540 67169 7580
rect 67255 7540 67276 7580
rect 67316 7540 67337 7580
rect 67423 7540 67440 7580
rect 67480 7540 67489 7580
rect 67103 7517 67169 7540
rect 67255 7517 67337 7540
rect 67423 7517 67489 7540
rect 67103 7498 67489 7517
rect 71103 7603 71489 7622
rect 71103 7580 71169 7603
rect 71255 7580 71337 7603
rect 71423 7580 71489 7603
rect 71103 7540 71112 7580
rect 71152 7540 71169 7580
rect 71255 7540 71276 7580
rect 71316 7540 71337 7580
rect 71423 7540 71440 7580
rect 71480 7540 71489 7580
rect 71103 7517 71169 7540
rect 71255 7517 71337 7540
rect 71423 7517 71489 7540
rect 71103 7498 71489 7517
rect 75103 7603 75489 7622
rect 75103 7580 75169 7603
rect 75255 7580 75337 7603
rect 75423 7580 75489 7603
rect 75103 7540 75112 7580
rect 75152 7540 75169 7580
rect 75255 7540 75276 7580
rect 75316 7540 75337 7580
rect 75423 7540 75440 7580
rect 75480 7540 75489 7580
rect 75103 7517 75169 7540
rect 75255 7517 75337 7540
rect 75423 7517 75489 7540
rect 75103 7498 75489 7517
rect 79103 7603 79489 7622
rect 79103 7580 79169 7603
rect 79255 7580 79337 7603
rect 79423 7580 79489 7603
rect 79103 7540 79112 7580
rect 79152 7540 79169 7580
rect 79255 7540 79276 7580
rect 79316 7540 79337 7580
rect 79423 7540 79440 7580
rect 79480 7540 79489 7580
rect 79103 7517 79169 7540
rect 79255 7517 79337 7540
rect 79423 7517 79489 7540
rect 79103 7498 79489 7517
rect 83103 7603 83489 7622
rect 83103 7580 83169 7603
rect 83255 7580 83337 7603
rect 83423 7580 83489 7603
rect 83103 7540 83112 7580
rect 83152 7540 83169 7580
rect 83255 7540 83276 7580
rect 83316 7540 83337 7580
rect 83423 7540 83440 7580
rect 83480 7540 83489 7580
rect 83103 7517 83169 7540
rect 83255 7517 83337 7540
rect 83423 7517 83489 7540
rect 83103 7498 83489 7517
rect 87103 7603 87489 7622
rect 87103 7580 87169 7603
rect 87255 7580 87337 7603
rect 87423 7580 87489 7603
rect 87103 7540 87112 7580
rect 87152 7540 87169 7580
rect 87255 7540 87276 7580
rect 87316 7540 87337 7580
rect 87423 7540 87440 7580
rect 87480 7540 87489 7580
rect 87103 7517 87169 7540
rect 87255 7517 87337 7540
rect 87423 7517 87489 7540
rect 87103 7498 87489 7517
rect 91103 7603 91489 7622
rect 91103 7580 91169 7603
rect 91255 7580 91337 7603
rect 91423 7580 91489 7603
rect 91103 7540 91112 7580
rect 91152 7540 91169 7580
rect 91255 7540 91276 7580
rect 91316 7540 91337 7580
rect 91423 7540 91440 7580
rect 91480 7540 91489 7580
rect 91103 7517 91169 7540
rect 91255 7517 91337 7540
rect 91423 7517 91489 7540
rect 91103 7498 91489 7517
rect 95103 7603 95489 7622
rect 95103 7580 95169 7603
rect 95255 7580 95337 7603
rect 95423 7580 95489 7603
rect 95103 7540 95112 7580
rect 95152 7540 95169 7580
rect 95255 7540 95276 7580
rect 95316 7540 95337 7580
rect 95423 7540 95440 7580
rect 95480 7540 95489 7580
rect 95103 7517 95169 7540
rect 95255 7517 95337 7540
rect 95423 7517 95489 7540
rect 95103 7498 95489 7517
rect 99103 7603 99489 7622
rect 99103 7580 99169 7603
rect 99255 7580 99337 7603
rect 99423 7580 99489 7603
rect 99103 7540 99112 7580
rect 99152 7540 99169 7580
rect 99255 7540 99276 7580
rect 99316 7540 99337 7580
rect 99423 7540 99440 7580
rect 99480 7540 99489 7580
rect 99103 7517 99169 7540
rect 99255 7517 99337 7540
rect 99423 7517 99489 7540
rect 99103 7498 99489 7517
rect 86450 7435 86574 7454
rect 86450 7349 86469 7435
rect 86555 7412 86574 7435
rect 86555 7372 86668 7412
rect 86708 7372 86717 7412
rect 86555 7349 86574 7372
rect 86450 7330 86574 7349
rect 4343 6847 4729 6866
rect 4343 6824 4409 6847
rect 4495 6824 4577 6847
rect 4663 6824 4729 6847
rect 4343 6784 4352 6824
rect 4392 6784 4409 6824
rect 4495 6784 4516 6824
rect 4556 6784 4577 6824
rect 4663 6784 4680 6824
rect 4720 6784 4729 6824
rect 4343 6761 4409 6784
rect 4495 6761 4577 6784
rect 4663 6761 4729 6784
rect 4343 6742 4729 6761
rect 8343 6847 8729 6866
rect 8343 6824 8409 6847
rect 8495 6824 8577 6847
rect 8663 6824 8729 6847
rect 8343 6784 8352 6824
rect 8392 6784 8409 6824
rect 8495 6784 8516 6824
rect 8556 6784 8577 6824
rect 8663 6784 8680 6824
rect 8720 6784 8729 6824
rect 8343 6761 8409 6784
rect 8495 6761 8577 6784
rect 8663 6761 8729 6784
rect 8343 6742 8729 6761
rect 12343 6847 12729 6866
rect 12343 6824 12409 6847
rect 12495 6824 12577 6847
rect 12663 6824 12729 6847
rect 12343 6784 12352 6824
rect 12392 6784 12409 6824
rect 12495 6784 12516 6824
rect 12556 6784 12577 6824
rect 12663 6784 12680 6824
rect 12720 6784 12729 6824
rect 12343 6761 12409 6784
rect 12495 6761 12577 6784
rect 12663 6761 12729 6784
rect 12343 6742 12729 6761
rect 16343 6847 16729 6866
rect 16343 6824 16409 6847
rect 16495 6824 16577 6847
rect 16663 6824 16729 6847
rect 16343 6784 16352 6824
rect 16392 6784 16409 6824
rect 16495 6784 16516 6824
rect 16556 6784 16577 6824
rect 16663 6784 16680 6824
rect 16720 6784 16729 6824
rect 16343 6761 16409 6784
rect 16495 6761 16577 6784
rect 16663 6761 16729 6784
rect 16343 6742 16729 6761
rect 20343 6847 20729 6866
rect 20343 6824 20409 6847
rect 20495 6824 20577 6847
rect 20663 6824 20729 6847
rect 20343 6784 20352 6824
rect 20392 6784 20409 6824
rect 20495 6784 20516 6824
rect 20556 6784 20577 6824
rect 20663 6784 20680 6824
rect 20720 6784 20729 6824
rect 20343 6761 20409 6784
rect 20495 6761 20577 6784
rect 20663 6761 20729 6784
rect 20343 6742 20729 6761
rect 24343 6847 24729 6866
rect 24343 6824 24409 6847
rect 24495 6824 24577 6847
rect 24663 6824 24729 6847
rect 24343 6784 24352 6824
rect 24392 6784 24409 6824
rect 24495 6784 24516 6824
rect 24556 6784 24577 6824
rect 24663 6784 24680 6824
rect 24720 6784 24729 6824
rect 24343 6761 24409 6784
rect 24495 6761 24577 6784
rect 24663 6761 24729 6784
rect 24343 6742 24729 6761
rect 28343 6847 28729 6866
rect 28343 6824 28409 6847
rect 28495 6824 28577 6847
rect 28663 6824 28729 6847
rect 28343 6784 28352 6824
rect 28392 6784 28409 6824
rect 28495 6784 28516 6824
rect 28556 6784 28577 6824
rect 28663 6784 28680 6824
rect 28720 6784 28729 6824
rect 28343 6761 28409 6784
rect 28495 6761 28577 6784
rect 28663 6761 28729 6784
rect 28343 6742 28729 6761
rect 32343 6847 32729 6866
rect 32343 6824 32409 6847
rect 32495 6824 32577 6847
rect 32663 6824 32729 6847
rect 32343 6784 32352 6824
rect 32392 6784 32409 6824
rect 32495 6784 32516 6824
rect 32556 6784 32577 6824
rect 32663 6784 32680 6824
rect 32720 6784 32729 6824
rect 32343 6761 32409 6784
rect 32495 6761 32577 6784
rect 32663 6761 32729 6784
rect 32343 6742 32729 6761
rect 36343 6847 36729 6866
rect 36343 6824 36409 6847
rect 36495 6824 36577 6847
rect 36663 6824 36729 6847
rect 36343 6784 36352 6824
rect 36392 6784 36409 6824
rect 36495 6784 36516 6824
rect 36556 6784 36577 6824
rect 36663 6784 36680 6824
rect 36720 6784 36729 6824
rect 36343 6761 36409 6784
rect 36495 6761 36577 6784
rect 36663 6761 36729 6784
rect 36343 6742 36729 6761
rect 40343 6847 40729 6866
rect 40343 6824 40409 6847
rect 40495 6824 40577 6847
rect 40663 6824 40729 6847
rect 40343 6784 40352 6824
rect 40392 6784 40409 6824
rect 40495 6784 40516 6824
rect 40556 6784 40577 6824
rect 40663 6784 40680 6824
rect 40720 6784 40729 6824
rect 40343 6761 40409 6784
rect 40495 6761 40577 6784
rect 40663 6761 40729 6784
rect 40343 6742 40729 6761
rect 44343 6847 44729 6866
rect 44343 6824 44409 6847
rect 44495 6824 44577 6847
rect 44663 6824 44729 6847
rect 44343 6784 44352 6824
rect 44392 6784 44409 6824
rect 44495 6784 44516 6824
rect 44556 6784 44577 6824
rect 44663 6784 44680 6824
rect 44720 6784 44729 6824
rect 44343 6761 44409 6784
rect 44495 6761 44577 6784
rect 44663 6761 44729 6784
rect 44343 6742 44729 6761
rect 48343 6847 48729 6866
rect 48343 6824 48409 6847
rect 48495 6824 48577 6847
rect 48663 6824 48729 6847
rect 48343 6784 48352 6824
rect 48392 6784 48409 6824
rect 48495 6784 48516 6824
rect 48556 6784 48577 6824
rect 48663 6784 48680 6824
rect 48720 6784 48729 6824
rect 48343 6761 48409 6784
rect 48495 6761 48577 6784
rect 48663 6761 48729 6784
rect 48343 6742 48729 6761
rect 52343 6847 52729 6866
rect 52343 6824 52409 6847
rect 52495 6824 52577 6847
rect 52663 6824 52729 6847
rect 52343 6784 52352 6824
rect 52392 6784 52409 6824
rect 52495 6784 52516 6824
rect 52556 6784 52577 6824
rect 52663 6784 52680 6824
rect 52720 6784 52729 6824
rect 52343 6761 52409 6784
rect 52495 6761 52577 6784
rect 52663 6761 52729 6784
rect 52343 6742 52729 6761
rect 56343 6847 56729 6866
rect 56343 6824 56409 6847
rect 56495 6824 56577 6847
rect 56663 6824 56729 6847
rect 56343 6784 56352 6824
rect 56392 6784 56409 6824
rect 56495 6784 56516 6824
rect 56556 6784 56577 6824
rect 56663 6784 56680 6824
rect 56720 6784 56729 6824
rect 56343 6761 56409 6784
rect 56495 6761 56577 6784
rect 56663 6761 56729 6784
rect 56343 6742 56729 6761
rect 60343 6847 60729 6866
rect 60343 6824 60409 6847
rect 60495 6824 60577 6847
rect 60663 6824 60729 6847
rect 60343 6784 60352 6824
rect 60392 6784 60409 6824
rect 60495 6784 60516 6824
rect 60556 6784 60577 6824
rect 60663 6784 60680 6824
rect 60720 6784 60729 6824
rect 60343 6761 60409 6784
rect 60495 6761 60577 6784
rect 60663 6761 60729 6784
rect 60343 6742 60729 6761
rect 64343 6847 64729 6866
rect 64343 6824 64409 6847
rect 64495 6824 64577 6847
rect 64663 6824 64729 6847
rect 64343 6784 64352 6824
rect 64392 6784 64409 6824
rect 64495 6784 64516 6824
rect 64556 6784 64577 6824
rect 64663 6784 64680 6824
rect 64720 6784 64729 6824
rect 64343 6761 64409 6784
rect 64495 6761 64577 6784
rect 64663 6761 64729 6784
rect 64343 6742 64729 6761
rect 68343 6847 68729 6866
rect 68343 6824 68409 6847
rect 68495 6824 68577 6847
rect 68663 6824 68729 6847
rect 68343 6784 68352 6824
rect 68392 6784 68409 6824
rect 68495 6784 68516 6824
rect 68556 6784 68577 6824
rect 68663 6784 68680 6824
rect 68720 6784 68729 6824
rect 68343 6761 68409 6784
rect 68495 6761 68577 6784
rect 68663 6761 68729 6784
rect 68343 6742 68729 6761
rect 72343 6847 72729 6866
rect 72343 6824 72409 6847
rect 72495 6824 72577 6847
rect 72663 6824 72729 6847
rect 72343 6784 72352 6824
rect 72392 6784 72409 6824
rect 72495 6784 72516 6824
rect 72556 6784 72577 6824
rect 72663 6784 72680 6824
rect 72720 6784 72729 6824
rect 72343 6761 72409 6784
rect 72495 6761 72577 6784
rect 72663 6761 72729 6784
rect 72343 6742 72729 6761
rect 76343 6847 76729 6866
rect 76343 6824 76409 6847
rect 76495 6824 76577 6847
rect 76663 6824 76729 6847
rect 76343 6784 76352 6824
rect 76392 6784 76409 6824
rect 76495 6784 76516 6824
rect 76556 6784 76577 6824
rect 76663 6784 76680 6824
rect 76720 6784 76729 6824
rect 76343 6761 76409 6784
rect 76495 6761 76577 6784
rect 76663 6761 76729 6784
rect 76343 6742 76729 6761
rect 80343 6847 80729 6866
rect 80343 6824 80409 6847
rect 80495 6824 80577 6847
rect 80663 6824 80729 6847
rect 80343 6784 80352 6824
rect 80392 6784 80409 6824
rect 80495 6784 80516 6824
rect 80556 6784 80577 6824
rect 80663 6784 80680 6824
rect 80720 6784 80729 6824
rect 80343 6761 80409 6784
rect 80495 6761 80577 6784
rect 80663 6761 80729 6784
rect 80343 6742 80729 6761
rect 84343 6847 84729 6866
rect 84343 6824 84409 6847
rect 84495 6824 84577 6847
rect 84663 6824 84729 6847
rect 84343 6784 84352 6824
rect 84392 6784 84409 6824
rect 84495 6784 84516 6824
rect 84556 6784 84577 6824
rect 84663 6784 84680 6824
rect 84720 6784 84729 6824
rect 84343 6761 84409 6784
rect 84495 6761 84577 6784
rect 84663 6761 84729 6784
rect 84343 6742 84729 6761
rect 88343 6847 88729 6866
rect 88343 6824 88409 6847
rect 88495 6824 88577 6847
rect 88663 6824 88729 6847
rect 88343 6784 88352 6824
rect 88392 6784 88409 6824
rect 88495 6784 88516 6824
rect 88556 6784 88577 6824
rect 88663 6784 88680 6824
rect 88720 6784 88729 6824
rect 88343 6761 88409 6784
rect 88495 6761 88577 6784
rect 88663 6761 88729 6784
rect 88343 6742 88729 6761
rect 92343 6847 92729 6866
rect 92343 6824 92409 6847
rect 92495 6824 92577 6847
rect 92663 6824 92729 6847
rect 92343 6784 92352 6824
rect 92392 6784 92409 6824
rect 92495 6784 92516 6824
rect 92556 6784 92577 6824
rect 92663 6784 92680 6824
rect 92720 6784 92729 6824
rect 92343 6761 92409 6784
rect 92495 6761 92577 6784
rect 92663 6761 92729 6784
rect 92343 6742 92729 6761
rect 96343 6847 96729 6866
rect 96343 6824 96409 6847
rect 96495 6824 96577 6847
rect 96663 6824 96729 6847
rect 96343 6784 96352 6824
rect 96392 6784 96409 6824
rect 96495 6784 96516 6824
rect 96556 6784 96577 6824
rect 96663 6784 96680 6824
rect 96720 6784 96729 6824
rect 96343 6761 96409 6784
rect 96495 6761 96577 6784
rect 96663 6761 96729 6784
rect 96343 6742 96729 6761
rect 3103 6091 3489 6110
rect 3103 6068 3169 6091
rect 3255 6068 3337 6091
rect 3423 6068 3489 6091
rect 3103 6028 3112 6068
rect 3152 6028 3169 6068
rect 3255 6028 3276 6068
rect 3316 6028 3337 6068
rect 3423 6028 3440 6068
rect 3480 6028 3489 6068
rect 3103 6005 3169 6028
rect 3255 6005 3337 6028
rect 3423 6005 3489 6028
rect 3103 5986 3489 6005
rect 7103 6091 7489 6110
rect 7103 6068 7169 6091
rect 7255 6068 7337 6091
rect 7423 6068 7489 6091
rect 7103 6028 7112 6068
rect 7152 6028 7169 6068
rect 7255 6028 7276 6068
rect 7316 6028 7337 6068
rect 7423 6028 7440 6068
rect 7480 6028 7489 6068
rect 7103 6005 7169 6028
rect 7255 6005 7337 6028
rect 7423 6005 7489 6028
rect 7103 5986 7489 6005
rect 11103 6091 11489 6110
rect 11103 6068 11169 6091
rect 11255 6068 11337 6091
rect 11423 6068 11489 6091
rect 11103 6028 11112 6068
rect 11152 6028 11169 6068
rect 11255 6028 11276 6068
rect 11316 6028 11337 6068
rect 11423 6028 11440 6068
rect 11480 6028 11489 6068
rect 11103 6005 11169 6028
rect 11255 6005 11337 6028
rect 11423 6005 11489 6028
rect 11103 5986 11489 6005
rect 15103 6091 15489 6110
rect 15103 6068 15169 6091
rect 15255 6068 15337 6091
rect 15423 6068 15489 6091
rect 15103 6028 15112 6068
rect 15152 6028 15169 6068
rect 15255 6028 15276 6068
rect 15316 6028 15337 6068
rect 15423 6028 15440 6068
rect 15480 6028 15489 6068
rect 15103 6005 15169 6028
rect 15255 6005 15337 6028
rect 15423 6005 15489 6028
rect 15103 5986 15489 6005
rect 19103 6091 19489 6110
rect 19103 6068 19169 6091
rect 19255 6068 19337 6091
rect 19423 6068 19489 6091
rect 19103 6028 19112 6068
rect 19152 6028 19169 6068
rect 19255 6028 19276 6068
rect 19316 6028 19337 6068
rect 19423 6028 19440 6068
rect 19480 6028 19489 6068
rect 19103 6005 19169 6028
rect 19255 6005 19337 6028
rect 19423 6005 19489 6028
rect 19103 5986 19489 6005
rect 23103 6091 23489 6110
rect 23103 6068 23169 6091
rect 23255 6068 23337 6091
rect 23423 6068 23489 6091
rect 23103 6028 23112 6068
rect 23152 6028 23169 6068
rect 23255 6028 23276 6068
rect 23316 6028 23337 6068
rect 23423 6028 23440 6068
rect 23480 6028 23489 6068
rect 23103 6005 23169 6028
rect 23255 6005 23337 6028
rect 23423 6005 23489 6028
rect 23103 5986 23489 6005
rect 27103 6091 27489 6110
rect 27103 6068 27169 6091
rect 27255 6068 27337 6091
rect 27423 6068 27489 6091
rect 27103 6028 27112 6068
rect 27152 6028 27169 6068
rect 27255 6028 27276 6068
rect 27316 6028 27337 6068
rect 27423 6028 27440 6068
rect 27480 6028 27489 6068
rect 27103 6005 27169 6028
rect 27255 6005 27337 6028
rect 27423 6005 27489 6028
rect 27103 5986 27489 6005
rect 31103 6091 31489 6110
rect 31103 6068 31169 6091
rect 31255 6068 31337 6091
rect 31423 6068 31489 6091
rect 31103 6028 31112 6068
rect 31152 6028 31169 6068
rect 31255 6028 31276 6068
rect 31316 6028 31337 6068
rect 31423 6028 31440 6068
rect 31480 6028 31489 6068
rect 31103 6005 31169 6028
rect 31255 6005 31337 6028
rect 31423 6005 31489 6028
rect 31103 5986 31489 6005
rect 35103 6091 35489 6110
rect 35103 6068 35169 6091
rect 35255 6068 35337 6091
rect 35423 6068 35489 6091
rect 35103 6028 35112 6068
rect 35152 6028 35169 6068
rect 35255 6028 35276 6068
rect 35316 6028 35337 6068
rect 35423 6028 35440 6068
rect 35480 6028 35489 6068
rect 35103 6005 35169 6028
rect 35255 6005 35337 6028
rect 35423 6005 35489 6028
rect 35103 5986 35489 6005
rect 39103 6091 39489 6110
rect 39103 6068 39169 6091
rect 39255 6068 39337 6091
rect 39423 6068 39489 6091
rect 39103 6028 39112 6068
rect 39152 6028 39169 6068
rect 39255 6028 39276 6068
rect 39316 6028 39337 6068
rect 39423 6028 39440 6068
rect 39480 6028 39489 6068
rect 39103 6005 39169 6028
rect 39255 6005 39337 6028
rect 39423 6005 39489 6028
rect 39103 5986 39489 6005
rect 43103 6091 43489 6110
rect 43103 6068 43169 6091
rect 43255 6068 43337 6091
rect 43423 6068 43489 6091
rect 43103 6028 43112 6068
rect 43152 6028 43169 6068
rect 43255 6028 43276 6068
rect 43316 6028 43337 6068
rect 43423 6028 43440 6068
rect 43480 6028 43489 6068
rect 43103 6005 43169 6028
rect 43255 6005 43337 6028
rect 43423 6005 43489 6028
rect 43103 5986 43489 6005
rect 47103 6091 47489 6110
rect 47103 6068 47169 6091
rect 47255 6068 47337 6091
rect 47423 6068 47489 6091
rect 47103 6028 47112 6068
rect 47152 6028 47169 6068
rect 47255 6028 47276 6068
rect 47316 6028 47337 6068
rect 47423 6028 47440 6068
rect 47480 6028 47489 6068
rect 47103 6005 47169 6028
rect 47255 6005 47337 6028
rect 47423 6005 47489 6028
rect 47103 5986 47489 6005
rect 51103 6091 51489 6110
rect 51103 6068 51169 6091
rect 51255 6068 51337 6091
rect 51423 6068 51489 6091
rect 51103 6028 51112 6068
rect 51152 6028 51169 6068
rect 51255 6028 51276 6068
rect 51316 6028 51337 6068
rect 51423 6028 51440 6068
rect 51480 6028 51489 6068
rect 51103 6005 51169 6028
rect 51255 6005 51337 6028
rect 51423 6005 51489 6028
rect 51103 5986 51489 6005
rect 55103 6091 55489 6110
rect 55103 6068 55169 6091
rect 55255 6068 55337 6091
rect 55423 6068 55489 6091
rect 55103 6028 55112 6068
rect 55152 6028 55169 6068
rect 55255 6028 55276 6068
rect 55316 6028 55337 6068
rect 55423 6028 55440 6068
rect 55480 6028 55489 6068
rect 55103 6005 55169 6028
rect 55255 6005 55337 6028
rect 55423 6005 55489 6028
rect 55103 5986 55489 6005
rect 59103 6091 59489 6110
rect 59103 6068 59169 6091
rect 59255 6068 59337 6091
rect 59423 6068 59489 6091
rect 59103 6028 59112 6068
rect 59152 6028 59169 6068
rect 59255 6028 59276 6068
rect 59316 6028 59337 6068
rect 59423 6028 59440 6068
rect 59480 6028 59489 6068
rect 59103 6005 59169 6028
rect 59255 6005 59337 6028
rect 59423 6005 59489 6028
rect 59103 5986 59489 6005
rect 63103 6091 63489 6110
rect 63103 6068 63169 6091
rect 63255 6068 63337 6091
rect 63423 6068 63489 6091
rect 63103 6028 63112 6068
rect 63152 6028 63169 6068
rect 63255 6028 63276 6068
rect 63316 6028 63337 6068
rect 63423 6028 63440 6068
rect 63480 6028 63489 6068
rect 63103 6005 63169 6028
rect 63255 6005 63337 6028
rect 63423 6005 63489 6028
rect 63103 5986 63489 6005
rect 67103 6091 67489 6110
rect 67103 6068 67169 6091
rect 67255 6068 67337 6091
rect 67423 6068 67489 6091
rect 67103 6028 67112 6068
rect 67152 6028 67169 6068
rect 67255 6028 67276 6068
rect 67316 6028 67337 6068
rect 67423 6028 67440 6068
rect 67480 6028 67489 6068
rect 67103 6005 67169 6028
rect 67255 6005 67337 6028
rect 67423 6005 67489 6028
rect 67103 5986 67489 6005
rect 71103 6091 71489 6110
rect 71103 6068 71169 6091
rect 71255 6068 71337 6091
rect 71423 6068 71489 6091
rect 71103 6028 71112 6068
rect 71152 6028 71169 6068
rect 71255 6028 71276 6068
rect 71316 6028 71337 6068
rect 71423 6028 71440 6068
rect 71480 6028 71489 6068
rect 71103 6005 71169 6028
rect 71255 6005 71337 6028
rect 71423 6005 71489 6028
rect 71103 5986 71489 6005
rect 75103 6091 75489 6110
rect 75103 6068 75169 6091
rect 75255 6068 75337 6091
rect 75423 6068 75489 6091
rect 75103 6028 75112 6068
rect 75152 6028 75169 6068
rect 75255 6028 75276 6068
rect 75316 6028 75337 6068
rect 75423 6028 75440 6068
rect 75480 6028 75489 6068
rect 75103 6005 75169 6028
rect 75255 6005 75337 6028
rect 75423 6005 75489 6028
rect 75103 5986 75489 6005
rect 79103 6091 79489 6110
rect 79103 6068 79169 6091
rect 79255 6068 79337 6091
rect 79423 6068 79489 6091
rect 79103 6028 79112 6068
rect 79152 6028 79169 6068
rect 79255 6028 79276 6068
rect 79316 6028 79337 6068
rect 79423 6028 79440 6068
rect 79480 6028 79489 6068
rect 79103 6005 79169 6028
rect 79255 6005 79337 6028
rect 79423 6005 79489 6028
rect 79103 5986 79489 6005
rect 83103 6091 83489 6110
rect 83103 6068 83169 6091
rect 83255 6068 83337 6091
rect 83423 6068 83489 6091
rect 83103 6028 83112 6068
rect 83152 6028 83169 6068
rect 83255 6028 83276 6068
rect 83316 6028 83337 6068
rect 83423 6028 83440 6068
rect 83480 6028 83489 6068
rect 83103 6005 83169 6028
rect 83255 6005 83337 6028
rect 83423 6005 83489 6028
rect 83103 5986 83489 6005
rect 87103 6091 87489 6110
rect 87103 6068 87169 6091
rect 87255 6068 87337 6091
rect 87423 6068 87489 6091
rect 87103 6028 87112 6068
rect 87152 6028 87169 6068
rect 87255 6028 87276 6068
rect 87316 6028 87337 6068
rect 87423 6028 87440 6068
rect 87480 6028 87489 6068
rect 87103 6005 87169 6028
rect 87255 6005 87337 6028
rect 87423 6005 87489 6028
rect 87103 5986 87489 6005
rect 91103 6091 91489 6110
rect 91103 6068 91169 6091
rect 91255 6068 91337 6091
rect 91423 6068 91489 6091
rect 91103 6028 91112 6068
rect 91152 6028 91169 6068
rect 91255 6028 91276 6068
rect 91316 6028 91337 6068
rect 91423 6028 91440 6068
rect 91480 6028 91489 6068
rect 91103 6005 91169 6028
rect 91255 6005 91337 6028
rect 91423 6005 91489 6028
rect 91103 5986 91489 6005
rect 95103 6091 95489 6110
rect 95103 6068 95169 6091
rect 95255 6068 95337 6091
rect 95423 6068 95489 6091
rect 95103 6028 95112 6068
rect 95152 6028 95169 6068
rect 95255 6028 95276 6068
rect 95316 6028 95337 6068
rect 95423 6028 95440 6068
rect 95480 6028 95489 6068
rect 95103 6005 95169 6028
rect 95255 6005 95337 6028
rect 95423 6005 95489 6028
rect 95103 5986 95489 6005
rect 99103 6091 99489 6110
rect 99103 6068 99169 6091
rect 99255 6068 99337 6091
rect 99423 6068 99489 6091
rect 99103 6028 99112 6068
rect 99152 6028 99169 6068
rect 99255 6028 99276 6068
rect 99316 6028 99337 6068
rect 99423 6028 99440 6068
rect 99480 6028 99489 6068
rect 99103 6005 99169 6028
rect 99255 6005 99337 6028
rect 99423 6005 99489 6028
rect 99103 5986 99489 6005
rect 4343 5335 4729 5354
rect 4343 5312 4409 5335
rect 4495 5312 4577 5335
rect 4663 5312 4729 5335
rect 4343 5272 4352 5312
rect 4392 5272 4409 5312
rect 4495 5272 4516 5312
rect 4556 5272 4577 5312
rect 4663 5272 4680 5312
rect 4720 5272 4729 5312
rect 4343 5249 4409 5272
rect 4495 5249 4577 5272
rect 4663 5249 4729 5272
rect 4343 5230 4729 5249
rect 8343 5335 8729 5354
rect 8343 5312 8409 5335
rect 8495 5312 8577 5335
rect 8663 5312 8729 5335
rect 8343 5272 8352 5312
rect 8392 5272 8409 5312
rect 8495 5272 8516 5312
rect 8556 5272 8577 5312
rect 8663 5272 8680 5312
rect 8720 5272 8729 5312
rect 8343 5249 8409 5272
rect 8495 5249 8577 5272
rect 8663 5249 8729 5272
rect 8343 5230 8729 5249
rect 12343 5335 12729 5354
rect 12343 5312 12409 5335
rect 12495 5312 12577 5335
rect 12663 5312 12729 5335
rect 12343 5272 12352 5312
rect 12392 5272 12409 5312
rect 12495 5272 12516 5312
rect 12556 5272 12577 5312
rect 12663 5272 12680 5312
rect 12720 5272 12729 5312
rect 12343 5249 12409 5272
rect 12495 5249 12577 5272
rect 12663 5249 12729 5272
rect 12343 5230 12729 5249
rect 16343 5335 16729 5354
rect 16343 5312 16409 5335
rect 16495 5312 16577 5335
rect 16663 5312 16729 5335
rect 16343 5272 16352 5312
rect 16392 5272 16409 5312
rect 16495 5272 16516 5312
rect 16556 5272 16577 5312
rect 16663 5272 16680 5312
rect 16720 5272 16729 5312
rect 16343 5249 16409 5272
rect 16495 5249 16577 5272
rect 16663 5249 16729 5272
rect 16343 5230 16729 5249
rect 20343 5335 20729 5354
rect 20343 5312 20409 5335
rect 20495 5312 20577 5335
rect 20663 5312 20729 5335
rect 20343 5272 20352 5312
rect 20392 5272 20409 5312
rect 20495 5272 20516 5312
rect 20556 5272 20577 5312
rect 20663 5272 20680 5312
rect 20720 5272 20729 5312
rect 20343 5249 20409 5272
rect 20495 5249 20577 5272
rect 20663 5249 20729 5272
rect 20343 5230 20729 5249
rect 24343 5335 24729 5354
rect 24343 5312 24409 5335
rect 24495 5312 24577 5335
rect 24663 5312 24729 5335
rect 24343 5272 24352 5312
rect 24392 5272 24409 5312
rect 24495 5272 24516 5312
rect 24556 5272 24577 5312
rect 24663 5272 24680 5312
rect 24720 5272 24729 5312
rect 24343 5249 24409 5272
rect 24495 5249 24577 5272
rect 24663 5249 24729 5272
rect 24343 5230 24729 5249
rect 28343 5335 28729 5354
rect 28343 5312 28409 5335
rect 28495 5312 28577 5335
rect 28663 5312 28729 5335
rect 28343 5272 28352 5312
rect 28392 5272 28409 5312
rect 28495 5272 28516 5312
rect 28556 5272 28577 5312
rect 28663 5272 28680 5312
rect 28720 5272 28729 5312
rect 28343 5249 28409 5272
rect 28495 5249 28577 5272
rect 28663 5249 28729 5272
rect 28343 5230 28729 5249
rect 32343 5335 32729 5354
rect 32343 5312 32409 5335
rect 32495 5312 32577 5335
rect 32663 5312 32729 5335
rect 32343 5272 32352 5312
rect 32392 5272 32409 5312
rect 32495 5272 32516 5312
rect 32556 5272 32577 5312
rect 32663 5272 32680 5312
rect 32720 5272 32729 5312
rect 32343 5249 32409 5272
rect 32495 5249 32577 5272
rect 32663 5249 32729 5272
rect 32343 5230 32729 5249
rect 36343 5335 36729 5354
rect 36343 5312 36409 5335
rect 36495 5312 36577 5335
rect 36663 5312 36729 5335
rect 36343 5272 36352 5312
rect 36392 5272 36409 5312
rect 36495 5272 36516 5312
rect 36556 5272 36577 5312
rect 36663 5272 36680 5312
rect 36720 5272 36729 5312
rect 36343 5249 36409 5272
rect 36495 5249 36577 5272
rect 36663 5249 36729 5272
rect 36343 5230 36729 5249
rect 40343 5335 40729 5354
rect 40343 5312 40409 5335
rect 40495 5312 40577 5335
rect 40663 5312 40729 5335
rect 40343 5272 40352 5312
rect 40392 5272 40409 5312
rect 40495 5272 40516 5312
rect 40556 5272 40577 5312
rect 40663 5272 40680 5312
rect 40720 5272 40729 5312
rect 40343 5249 40409 5272
rect 40495 5249 40577 5272
rect 40663 5249 40729 5272
rect 40343 5230 40729 5249
rect 44343 5335 44729 5354
rect 44343 5312 44409 5335
rect 44495 5312 44577 5335
rect 44663 5312 44729 5335
rect 44343 5272 44352 5312
rect 44392 5272 44409 5312
rect 44495 5272 44516 5312
rect 44556 5272 44577 5312
rect 44663 5272 44680 5312
rect 44720 5272 44729 5312
rect 44343 5249 44409 5272
rect 44495 5249 44577 5272
rect 44663 5249 44729 5272
rect 44343 5230 44729 5249
rect 48343 5335 48729 5354
rect 48343 5312 48409 5335
rect 48495 5312 48577 5335
rect 48663 5312 48729 5335
rect 48343 5272 48352 5312
rect 48392 5272 48409 5312
rect 48495 5272 48516 5312
rect 48556 5272 48577 5312
rect 48663 5272 48680 5312
rect 48720 5272 48729 5312
rect 48343 5249 48409 5272
rect 48495 5249 48577 5272
rect 48663 5249 48729 5272
rect 48343 5230 48729 5249
rect 52343 5335 52729 5354
rect 52343 5312 52409 5335
rect 52495 5312 52577 5335
rect 52663 5312 52729 5335
rect 52343 5272 52352 5312
rect 52392 5272 52409 5312
rect 52495 5272 52516 5312
rect 52556 5272 52577 5312
rect 52663 5272 52680 5312
rect 52720 5272 52729 5312
rect 52343 5249 52409 5272
rect 52495 5249 52577 5272
rect 52663 5249 52729 5272
rect 52343 5230 52729 5249
rect 56343 5335 56729 5354
rect 56343 5312 56409 5335
rect 56495 5312 56577 5335
rect 56663 5312 56729 5335
rect 56343 5272 56352 5312
rect 56392 5272 56409 5312
rect 56495 5272 56516 5312
rect 56556 5272 56577 5312
rect 56663 5272 56680 5312
rect 56720 5272 56729 5312
rect 56343 5249 56409 5272
rect 56495 5249 56577 5272
rect 56663 5249 56729 5272
rect 56343 5230 56729 5249
rect 60343 5335 60729 5354
rect 60343 5312 60409 5335
rect 60495 5312 60577 5335
rect 60663 5312 60729 5335
rect 60343 5272 60352 5312
rect 60392 5272 60409 5312
rect 60495 5272 60516 5312
rect 60556 5272 60577 5312
rect 60663 5272 60680 5312
rect 60720 5272 60729 5312
rect 60343 5249 60409 5272
rect 60495 5249 60577 5272
rect 60663 5249 60729 5272
rect 60343 5230 60729 5249
rect 64343 5335 64729 5354
rect 64343 5312 64409 5335
rect 64495 5312 64577 5335
rect 64663 5312 64729 5335
rect 64343 5272 64352 5312
rect 64392 5272 64409 5312
rect 64495 5272 64516 5312
rect 64556 5272 64577 5312
rect 64663 5272 64680 5312
rect 64720 5272 64729 5312
rect 64343 5249 64409 5272
rect 64495 5249 64577 5272
rect 64663 5249 64729 5272
rect 64343 5230 64729 5249
rect 68343 5335 68729 5354
rect 68343 5312 68409 5335
rect 68495 5312 68577 5335
rect 68663 5312 68729 5335
rect 68343 5272 68352 5312
rect 68392 5272 68409 5312
rect 68495 5272 68516 5312
rect 68556 5272 68577 5312
rect 68663 5272 68680 5312
rect 68720 5272 68729 5312
rect 68343 5249 68409 5272
rect 68495 5249 68577 5272
rect 68663 5249 68729 5272
rect 68343 5230 68729 5249
rect 72343 5335 72729 5354
rect 72343 5312 72409 5335
rect 72495 5312 72577 5335
rect 72663 5312 72729 5335
rect 72343 5272 72352 5312
rect 72392 5272 72409 5312
rect 72495 5272 72516 5312
rect 72556 5272 72577 5312
rect 72663 5272 72680 5312
rect 72720 5272 72729 5312
rect 72343 5249 72409 5272
rect 72495 5249 72577 5272
rect 72663 5249 72729 5272
rect 72343 5230 72729 5249
rect 76343 5335 76729 5354
rect 76343 5312 76409 5335
rect 76495 5312 76577 5335
rect 76663 5312 76729 5335
rect 76343 5272 76352 5312
rect 76392 5272 76409 5312
rect 76495 5272 76516 5312
rect 76556 5272 76577 5312
rect 76663 5272 76680 5312
rect 76720 5272 76729 5312
rect 76343 5249 76409 5272
rect 76495 5249 76577 5272
rect 76663 5249 76729 5272
rect 76343 5230 76729 5249
rect 80343 5335 80729 5354
rect 80343 5312 80409 5335
rect 80495 5312 80577 5335
rect 80663 5312 80729 5335
rect 80343 5272 80352 5312
rect 80392 5272 80409 5312
rect 80495 5272 80516 5312
rect 80556 5272 80577 5312
rect 80663 5272 80680 5312
rect 80720 5272 80729 5312
rect 80343 5249 80409 5272
rect 80495 5249 80577 5272
rect 80663 5249 80729 5272
rect 80343 5230 80729 5249
rect 84343 5335 84729 5354
rect 84343 5312 84409 5335
rect 84495 5312 84577 5335
rect 84663 5312 84729 5335
rect 84343 5272 84352 5312
rect 84392 5272 84409 5312
rect 84495 5272 84516 5312
rect 84556 5272 84577 5312
rect 84663 5272 84680 5312
rect 84720 5272 84729 5312
rect 84343 5249 84409 5272
rect 84495 5249 84577 5272
rect 84663 5249 84729 5272
rect 84343 5230 84729 5249
rect 88343 5335 88729 5354
rect 88343 5312 88409 5335
rect 88495 5312 88577 5335
rect 88663 5312 88729 5335
rect 88343 5272 88352 5312
rect 88392 5272 88409 5312
rect 88495 5272 88516 5312
rect 88556 5272 88577 5312
rect 88663 5272 88680 5312
rect 88720 5272 88729 5312
rect 88343 5249 88409 5272
rect 88495 5249 88577 5272
rect 88663 5249 88729 5272
rect 88343 5230 88729 5249
rect 92343 5335 92729 5354
rect 92343 5312 92409 5335
rect 92495 5312 92577 5335
rect 92663 5312 92729 5335
rect 92343 5272 92352 5312
rect 92392 5272 92409 5312
rect 92495 5272 92516 5312
rect 92556 5272 92577 5312
rect 92663 5272 92680 5312
rect 92720 5272 92729 5312
rect 92343 5249 92409 5272
rect 92495 5249 92577 5272
rect 92663 5249 92729 5272
rect 92343 5230 92729 5249
rect 96343 5335 96729 5354
rect 96343 5312 96409 5335
rect 96495 5312 96577 5335
rect 96663 5312 96729 5335
rect 96343 5272 96352 5312
rect 96392 5272 96409 5312
rect 96495 5272 96516 5312
rect 96556 5272 96577 5312
rect 96663 5272 96680 5312
rect 96720 5272 96729 5312
rect 96343 5249 96409 5272
rect 96495 5249 96577 5272
rect 96663 5249 96729 5272
rect 96343 5230 96729 5249
rect 3103 4579 3489 4598
rect 3103 4556 3169 4579
rect 3255 4556 3337 4579
rect 3423 4556 3489 4579
rect 3103 4516 3112 4556
rect 3152 4516 3169 4556
rect 3255 4516 3276 4556
rect 3316 4516 3337 4556
rect 3423 4516 3440 4556
rect 3480 4516 3489 4556
rect 3103 4493 3169 4516
rect 3255 4493 3337 4516
rect 3423 4493 3489 4516
rect 3103 4474 3489 4493
rect 7103 4579 7489 4598
rect 7103 4556 7169 4579
rect 7255 4556 7337 4579
rect 7423 4556 7489 4579
rect 7103 4516 7112 4556
rect 7152 4516 7169 4556
rect 7255 4516 7276 4556
rect 7316 4516 7337 4556
rect 7423 4516 7440 4556
rect 7480 4516 7489 4556
rect 7103 4493 7169 4516
rect 7255 4493 7337 4516
rect 7423 4493 7489 4516
rect 7103 4474 7489 4493
rect 11103 4579 11489 4598
rect 11103 4556 11169 4579
rect 11255 4556 11337 4579
rect 11423 4556 11489 4579
rect 11103 4516 11112 4556
rect 11152 4516 11169 4556
rect 11255 4516 11276 4556
rect 11316 4516 11337 4556
rect 11423 4516 11440 4556
rect 11480 4516 11489 4556
rect 11103 4493 11169 4516
rect 11255 4493 11337 4516
rect 11423 4493 11489 4516
rect 11103 4474 11489 4493
rect 15103 4579 15489 4598
rect 15103 4556 15169 4579
rect 15255 4556 15337 4579
rect 15423 4556 15489 4579
rect 15103 4516 15112 4556
rect 15152 4516 15169 4556
rect 15255 4516 15276 4556
rect 15316 4516 15337 4556
rect 15423 4516 15440 4556
rect 15480 4516 15489 4556
rect 15103 4493 15169 4516
rect 15255 4493 15337 4516
rect 15423 4493 15489 4516
rect 15103 4474 15489 4493
rect 19103 4579 19489 4598
rect 19103 4556 19169 4579
rect 19255 4556 19337 4579
rect 19423 4556 19489 4579
rect 19103 4516 19112 4556
rect 19152 4516 19169 4556
rect 19255 4516 19276 4556
rect 19316 4516 19337 4556
rect 19423 4516 19440 4556
rect 19480 4516 19489 4556
rect 19103 4493 19169 4516
rect 19255 4493 19337 4516
rect 19423 4493 19489 4516
rect 19103 4474 19489 4493
rect 23103 4579 23489 4598
rect 23103 4556 23169 4579
rect 23255 4556 23337 4579
rect 23423 4556 23489 4579
rect 23103 4516 23112 4556
rect 23152 4516 23169 4556
rect 23255 4516 23276 4556
rect 23316 4516 23337 4556
rect 23423 4516 23440 4556
rect 23480 4516 23489 4556
rect 23103 4493 23169 4516
rect 23255 4493 23337 4516
rect 23423 4493 23489 4516
rect 23103 4474 23489 4493
rect 27103 4579 27489 4598
rect 27103 4556 27169 4579
rect 27255 4556 27337 4579
rect 27423 4556 27489 4579
rect 27103 4516 27112 4556
rect 27152 4516 27169 4556
rect 27255 4516 27276 4556
rect 27316 4516 27337 4556
rect 27423 4516 27440 4556
rect 27480 4516 27489 4556
rect 27103 4493 27169 4516
rect 27255 4493 27337 4516
rect 27423 4493 27489 4516
rect 27103 4474 27489 4493
rect 31103 4579 31489 4598
rect 31103 4556 31169 4579
rect 31255 4556 31337 4579
rect 31423 4556 31489 4579
rect 31103 4516 31112 4556
rect 31152 4516 31169 4556
rect 31255 4516 31276 4556
rect 31316 4516 31337 4556
rect 31423 4516 31440 4556
rect 31480 4516 31489 4556
rect 31103 4493 31169 4516
rect 31255 4493 31337 4516
rect 31423 4493 31489 4516
rect 31103 4474 31489 4493
rect 35103 4579 35489 4598
rect 35103 4556 35169 4579
rect 35255 4556 35337 4579
rect 35423 4556 35489 4579
rect 35103 4516 35112 4556
rect 35152 4516 35169 4556
rect 35255 4516 35276 4556
rect 35316 4516 35337 4556
rect 35423 4516 35440 4556
rect 35480 4516 35489 4556
rect 35103 4493 35169 4516
rect 35255 4493 35337 4516
rect 35423 4493 35489 4516
rect 35103 4474 35489 4493
rect 39103 4579 39489 4598
rect 39103 4556 39169 4579
rect 39255 4556 39337 4579
rect 39423 4556 39489 4579
rect 39103 4516 39112 4556
rect 39152 4516 39169 4556
rect 39255 4516 39276 4556
rect 39316 4516 39337 4556
rect 39423 4516 39440 4556
rect 39480 4516 39489 4556
rect 39103 4493 39169 4516
rect 39255 4493 39337 4516
rect 39423 4493 39489 4516
rect 39103 4474 39489 4493
rect 43103 4579 43489 4598
rect 43103 4556 43169 4579
rect 43255 4556 43337 4579
rect 43423 4556 43489 4579
rect 43103 4516 43112 4556
rect 43152 4516 43169 4556
rect 43255 4516 43276 4556
rect 43316 4516 43337 4556
rect 43423 4516 43440 4556
rect 43480 4516 43489 4556
rect 43103 4493 43169 4516
rect 43255 4493 43337 4516
rect 43423 4493 43489 4516
rect 43103 4474 43489 4493
rect 47103 4579 47489 4598
rect 47103 4556 47169 4579
rect 47255 4556 47337 4579
rect 47423 4556 47489 4579
rect 47103 4516 47112 4556
rect 47152 4516 47169 4556
rect 47255 4516 47276 4556
rect 47316 4516 47337 4556
rect 47423 4516 47440 4556
rect 47480 4516 47489 4556
rect 47103 4493 47169 4516
rect 47255 4493 47337 4516
rect 47423 4493 47489 4516
rect 47103 4474 47489 4493
rect 51103 4579 51489 4598
rect 51103 4556 51169 4579
rect 51255 4556 51337 4579
rect 51423 4556 51489 4579
rect 51103 4516 51112 4556
rect 51152 4516 51169 4556
rect 51255 4516 51276 4556
rect 51316 4516 51337 4556
rect 51423 4516 51440 4556
rect 51480 4516 51489 4556
rect 51103 4493 51169 4516
rect 51255 4493 51337 4516
rect 51423 4493 51489 4516
rect 51103 4474 51489 4493
rect 55103 4579 55489 4598
rect 55103 4556 55169 4579
rect 55255 4556 55337 4579
rect 55423 4556 55489 4579
rect 55103 4516 55112 4556
rect 55152 4516 55169 4556
rect 55255 4516 55276 4556
rect 55316 4516 55337 4556
rect 55423 4516 55440 4556
rect 55480 4516 55489 4556
rect 55103 4493 55169 4516
rect 55255 4493 55337 4516
rect 55423 4493 55489 4516
rect 55103 4474 55489 4493
rect 59103 4579 59489 4598
rect 59103 4556 59169 4579
rect 59255 4556 59337 4579
rect 59423 4556 59489 4579
rect 59103 4516 59112 4556
rect 59152 4516 59169 4556
rect 59255 4516 59276 4556
rect 59316 4516 59337 4556
rect 59423 4516 59440 4556
rect 59480 4516 59489 4556
rect 59103 4493 59169 4516
rect 59255 4493 59337 4516
rect 59423 4493 59489 4516
rect 59103 4474 59489 4493
rect 63103 4579 63489 4598
rect 63103 4556 63169 4579
rect 63255 4556 63337 4579
rect 63423 4556 63489 4579
rect 63103 4516 63112 4556
rect 63152 4516 63169 4556
rect 63255 4516 63276 4556
rect 63316 4516 63337 4556
rect 63423 4516 63440 4556
rect 63480 4516 63489 4556
rect 63103 4493 63169 4516
rect 63255 4493 63337 4516
rect 63423 4493 63489 4516
rect 63103 4474 63489 4493
rect 67103 4579 67489 4598
rect 67103 4556 67169 4579
rect 67255 4556 67337 4579
rect 67423 4556 67489 4579
rect 67103 4516 67112 4556
rect 67152 4516 67169 4556
rect 67255 4516 67276 4556
rect 67316 4516 67337 4556
rect 67423 4516 67440 4556
rect 67480 4516 67489 4556
rect 67103 4493 67169 4516
rect 67255 4493 67337 4516
rect 67423 4493 67489 4516
rect 67103 4474 67489 4493
rect 71103 4579 71489 4598
rect 71103 4556 71169 4579
rect 71255 4556 71337 4579
rect 71423 4556 71489 4579
rect 71103 4516 71112 4556
rect 71152 4516 71169 4556
rect 71255 4516 71276 4556
rect 71316 4516 71337 4556
rect 71423 4516 71440 4556
rect 71480 4516 71489 4556
rect 71103 4493 71169 4516
rect 71255 4493 71337 4516
rect 71423 4493 71489 4516
rect 71103 4474 71489 4493
rect 75103 4579 75489 4598
rect 75103 4556 75169 4579
rect 75255 4556 75337 4579
rect 75423 4556 75489 4579
rect 75103 4516 75112 4556
rect 75152 4516 75169 4556
rect 75255 4516 75276 4556
rect 75316 4516 75337 4556
rect 75423 4516 75440 4556
rect 75480 4516 75489 4556
rect 75103 4493 75169 4516
rect 75255 4493 75337 4516
rect 75423 4493 75489 4516
rect 75103 4474 75489 4493
rect 79103 4579 79489 4598
rect 79103 4556 79169 4579
rect 79255 4556 79337 4579
rect 79423 4556 79489 4579
rect 79103 4516 79112 4556
rect 79152 4516 79169 4556
rect 79255 4516 79276 4556
rect 79316 4516 79337 4556
rect 79423 4516 79440 4556
rect 79480 4516 79489 4556
rect 79103 4493 79169 4516
rect 79255 4493 79337 4516
rect 79423 4493 79489 4516
rect 79103 4474 79489 4493
rect 83103 4579 83489 4598
rect 83103 4556 83169 4579
rect 83255 4556 83337 4579
rect 83423 4556 83489 4579
rect 83103 4516 83112 4556
rect 83152 4516 83169 4556
rect 83255 4516 83276 4556
rect 83316 4516 83337 4556
rect 83423 4516 83440 4556
rect 83480 4516 83489 4556
rect 83103 4493 83169 4516
rect 83255 4493 83337 4516
rect 83423 4493 83489 4516
rect 83103 4474 83489 4493
rect 87103 4579 87489 4598
rect 87103 4556 87169 4579
rect 87255 4556 87337 4579
rect 87423 4556 87489 4579
rect 87103 4516 87112 4556
rect 87152 4516 87169 4556
rect 87255 4516 87276 4556
rect 87316 4516 87337 4556
rect 87423 4516 87440 4556
rect 87480 4516 87489 4556
rect 87103 4493 87169 4516
rect 87255 4493 87337 4516
rect 87423 4493 87489 4516
rect 87103 4474 87489 4493
rect 91103 4579 91489 4598
rect 91103 4556 91169 4579
rect 91255 4556 91337 4579
rect 91423 4556 91489 4579
rect 91103 4516 91112 4556
rect 91152 4516 91169 4556
rect 91255 4516 91276 4556
rect 91316 4516 91337 4556
rect 91423 4516 91440 4556
rect 91480 4516 91489 4556
rect 91103 4493 91169 4516
rect 91255 4493 91337 4516
rect 91423 4493 91489 4516
rect 91103 4474 91489 4493
rect 95103 4579 95489 4598
rect 95103 4556 95169 4579
rect 95255 4556 95337 4579
rect 95423 4556 95489 4579
rect 95103 4516 95112 4556
rect 95152 4516 95169 4556
rect 95255 4516 95276 4556
rect 95316 4516 95337 4556
rect 95423 4516 95440 4556
rect 95480 4516 95489 4556
rect 95103 4493 95169 4516
rect 95255 4493 95337 4516
rect 95423 4493 95489 4516
rect 95103 4474 95489 4493
rect 99103 4579 99489 4598
rect 99103 4556 99169 4579
rect 99255 4556 99337 4579
rect 99423 4556 99489 4579
rect 99103 4516 99112 4556
rect 99152 4516 99169 4556
rect 99255 4516 99276 4556
rect 99316 4516 99337 4556
rect 99423 4516 99440 4556
rect 99480 4516 99489 4556
rect 99103 4493 99169 4516
rect 99255 4493 99337 4516
rect 99423 4493 99489 4516
rect 99103 4474 99489 4493
rect 4343 3823 4729 3842
rect 4343 3800 4409 3823
rect 4495 3800 4577 3823
rect 4663 3800 4729 3823
rect 4343 3760 4352 3800
rect 4392 3760 4409 3800
rect 4495 3760 4516 3800
rect 4556 3760 4577 3800
rect 4663 3760 4680 3800
rect 4720 3760 4729 3800
rect 4343 3737 4409 3760
rect 4495 3737 4577 3760
rect 4663 3737 4729 3760
rect 4343 3718 4729 3737
rect 8343 3823 8729 3842
rect 8343 3800 8409 3823
rect 8495 3800 8577 3823
rect 8663 3800 8729 3823
rect 8343 3760 8352 3800
rect 8392 3760 8409 3800
rect 8495 3760 8516 3800
rect 8556 3760 8577 3800
rect 8663 3760 8680 3800
rect 8720 3760 8729 3800
rect 8343 3737 8409 3760
rect 8495 3737 8577 3760
rect 8663 3737 8729 3760
rect 8343 3718 8729 3737
rect 12343 3823 12729 3842
rect 12343 3800 12409 3823
rect 12495 3800 12577 3823
rect 12663 3800 12729 3823
rect 12343 3760 12352 3800
rect 12392 3760 12409 3800
rect 12495 3760 12516 3800
rect 12556 3760 12577 3800
rect 12663 3760 12680 3800
rect 12720 3760 12729 3800
rect 12343 3737 12409 3760
rect 12495 3737 12577 3760
rect 12663 3737 12729 3760
rect 12343 3718 12729 3737
rect 16343 3823 16729 3842
rect 16343 3800 16409 3823
rect 16495 3800 16577 3823
rect 16663 3800 16729 3823
rect 16343 3760 16352 3800
rect 16392 3760 16409 3800
rect 16495 3760 16516 3800
rect 16556 3760 16577 3800
rect 16663 3760 16680 3800
rect 16720 3760 16729 3800
rect 16343 3737 16409 3760
rect 16495 3737 16577 3760
rect 16663 3737 16729 3760
rect 16343 3718 16729 3737
rect 20343 3823 20729 3842
rect 20343 3800 20409 3823
rect 20495 3800 20577 3823
rect 20663 3800 20729 3823
rect 20343 3760 20352 3800
rect 20392 3760 20409 3800
rect 20495 3760 20516 3800
rect 20556 3760 20577 3800
rect 20663 3760 20680 3800
rect 20720 3760 20729 3800
rect 20343 3737 20409 3760
rect 20495 3737 20577 3760
rect 20663 3737 20729 3760
rect 20343 3718 20729 3737
rect 24343 3823 24729 3842
rect 24343 3800 24409 3823
rect 24495 3800 24577 3823
rect 24663 3800 24729 3823
rect 24343 3760 24352 3800
rect 24392 3760 24409 3800
rect 24495 3760 24516 3800
rect 24556 3760 24577 3800
rect 24663 3760 24680 3800
rect 24720 3760 24729 3800
rect 24343 3737 24409 3760
rect 24495 3737 24577 3760
rect 24663 3737 24729 3760
rect 24343 3718 24729 3737
rect 28343 3823 28729 3842
rect 28343 3800 28409 3823
rect 28495 3800 28577 3823
rect 28663 3800 28729 3823
rect 28343 3760 28352 3800
rect 28392 3760 28409 3800
rect 28495 3760 28516 3800
rect 28556 3760 28577 3800
rect 28663 3760 28680 3800
rect 28720 3760 28729 3800
rect 28343 3737 28409 3760
rect 28495 3737 28577 3760
rect 28663 3737 28729 3760
rect 28343 3718 28729 3737
rect 32343 3823 32729 3842
rect 32343 3800 32409 3823
rect 32495 3800 32577 3823
rect 32663 3800 32729 3823
rect 32343 3760 32352 3800
rect 32392 3760 32409 3800
rect 32495 3760 32516 3800
rect 32556 3760 32577 3800
rect 32663 3760 32680 3800
rect 32720 3760 32729 3800
rect 32343 3737 32409 3760
rect 32495 3737 32577 3760
rect 32663 3737 32729 3760
rect 32343 3718 32729 3737
rect 36343 3823 36729 3842
rect 36343 3800 36409 3823
rect 36495 3800 36577 3823
rect 36663 3800 36729 3823
rect 36343 3760 36352 3800
rect 36392 3760 36409 3800
rect 36495 3760 36516 3800
rect 36556 3760 36577 3800
rect 36663 3760 36680 3800
rect 36720 3760 36729 3800
rect 36343 3737 36409 3760
rect 36495 3737 36577 3760
rect 36663 3737 36729 3760
rect 36343 3718 36729 3737
rect 40343 3823 40729 3842
rect 40343 3800 40409 3823
rect 40495 3800 40577 3823
rect 40663 3800 40729 3823
rect 40343 3760 40352 3800
rect 40392 3760 40409 3800
rect 40495 3760 40516 3800
rect 40556 3760 40577 3800
rect 40663 3760 40680 3800
rect 40720 3760 40729 3800
rect 40343 3737 40409 3760
rect 40495 3737 40577 3760
rect 40663 3737 40729 3760
rect 40343 3718 40729 3737
rect 44343 3823 44729 3842
rect 44343 3800 44409 3823
rect 44495 3800 44577 3823
rect 44663 3800 44729 3823
rect 44343 3760 44352 3800
rect 44392 3760 44409 3800
rect 44495 3760 44516 3800
rect 44556 3760 44577 3800
rect 44663 3760 44680 3800
rect 44720 3760 44729 3800
rect 44343 3737 44409 3760
rect 44495 3737 44577 3760
rect 44663 3737 44729 3760
rect 44343 3718 44729 3737
rect 48343 3823 48729 3842
rect 48343 3800 48409 3823
rect 48495 3800 48577 3823
rect 48663 3800 48729 3823
rect 48343 3760 48352 3800
rect 48392 3760 48409 3800
rect 48495 3760 48516 3800
rect 48556 3760 48577 3800
rect 48663 3760 48680 3800
rect 48720 3760 48729 3800
rect 48343 3737 48409 3760
rect 48495 3737 48577 3760
rect 48663 3737 48729 3760
rect 48343 3718 48729 3737
rect 52343 3823 52729 3842
rect 52343 3800 52409 3823
rect 52495 3800 52577 3823
rect 52663 3800 52729 3823
rect 52343 3760 52352 3800
rect 52392 3760 52409 3800
rect 52495 3760 52516 3800
rect 52556 3760 52577 3800
rect 52663 3760 52680 3800
rect 52720 3760 52729 3800
rect 52343 3737 52409 3760
rect 52495 3737 52577 3760
rect 52663 3737 52729 3760
rect 52343 3718 52729 3737
rect 56343 3823 56729 3842
rect 56343 3800 56409 3823
rect 56495 3800 56577 3823
rect 56663 3800 56729 3823
rect 56343 3760 56352 3800
rect 56392 3760 56409 3800
rect 56495 3760 56516 3800
rect 56556 3760 56577 3800
rect 56663 3760 56680 3800
rect 56720 3760 56729 3800
rect 56343 3737 56409 3760
rect 56495 3737 56577 3760
rect 56663 3737 56729 3760
rect 56343 3718 56729 3737
rect 60343 3823 60729 3842
rect 60343 3800 60409 3823
rect 60495 3800 60577 3823
rect 60663 3800 60729 3823
rect 60343 3760 60352 3800
rect 60392 3760 60409 3800
rect 60495 3760 60516 3800
rect 60556 3760 60577 3800
rect 60663 3760 60680 3800
rect 60720 3760 60729 3800
rect 60343 3737 60409 3760
rect 60495 3737 60577 3760
rect 60663 3737 60729 3760
rect 60343 3718 60729 3737
rect 64343 3823 64729 3842
rect 64343 3800 64409 3823
rect 64495 3800 64577 3823
rect 64663 3800 64729 3823
rect 64343 3760 64352 3800
rect 64392 3760 64409 3800
rect 64495 3760 64516 3800
rect 64556 3760 64577 3800
rect 64663 3760 64680 3800
rect 64720 3760 64729 3800
rect 64343 3737 64409 3760
rect 64495 3737 64577 3760
rect 64663 3737 64729 3760
rect 64343 3718 64729 3737
rect 68343 3823 68729 3842
rect 68343 3800 68409 3823
rect 68495 3800 68577 3823
rect 68663 3800 68729 3823
rect 68343 3760 68352 3800
rect 68392 3760 68409 3800
rect 68495 3760 68516 3800
rect 68556 3760 68577 3800
rect 68663 3760 68680 3800
rect 68720 3760 68729 3800
rect 68343 3737 68409 3760
rect 68495 3737 68577 3760
rect 68663 3737 68729 3760
rect 68343 3718 68729 3737
rect 72343 3823 72729 3842
rect 72343 3800 72409 3823
rect 72495 3800 72577 3823
rect 72663 3800 72729 3823
rect 72343 3760 72352 3800
rect 72392 3760 72409 3800
rect 72495 3760 72516 3800
rect 72556 3760 72577 3800
rect 72663 3760 72680 3800
rect 72720 3760 72729 3800
rect 72343 3737 72409 3760
rect 72495 3737 72577 3760
rect 72663 3737 72729 3760
rect 72343 3718 72729 3737
rect 76343 3823 76729 3842
rect 76343 3800 76409 3823
rect 76495 3800 76577 3823
rect 76663 3800 76729 3823
rect 76343 3760 76352 3800
rect 76392 3760 76409 3800
rect 76495 3760 76516 3800
rect 76556 3760 76577 3800
rect 76663 3760 76680 3800
rect 76720 3760 76729 3800
rect 76343 3737 76409 3760
rect 76495 3737 76577 3760
rect 76663 3737 76729 3760
rect 76343 3718 76729 3737
rect 80343 3823 80729 3842
rect 80343 3800 80409 3823
rect 80495 3800 80577 3823
rect 80663 3800 80729 3823
rect 80343 3760 80352 3800
rect 80392 3760 80409 3800
rect 80495 3760 80516 3800
rect 80556 3760 80577 3800
rect 80663 3760 80680 3800
rect 80720 3760 80729 3800
rect 80343 3737 80409 3760
rect 80495 3737 80577 3760
rect 80663 3737 80729 3760
rect 80343 3718 80729 3737
rect 84343 3823 84729 3842
rect 84343 3800 84409 3823
rect 84495 3800 84577 3823
rect 84663 3800 84729 3823
rect 84343 3760 84352 3800
rect 84392 3760 84409 3800
rect 84495 3760 84516 3800
rect 84556 3760 84577 3800
rect 84663 3760 84680 3800
rect 84720 3760 84729 3800
rect 84343 3737 84409 3760
rect 84495 3737 84577 3760
rect 84663 3737 84729 3760
rect 84343 3718 84729 3737
rect 88343 3823 88729 3842
rect 88343 3800 88409 3823
rect 88495 3800 88577 3823
rect 88663 3800 88729 3823
rect 88343 3760 88352 3800
rect 88392 3760 88409 3800
rect 88495 3760 88516 3800
rect 88556 3760 88577 3800
rect 88663 3760 88680 3800
rect 88720 3760 88729 3800
rect 88343 3737 88409 3760
rect 88495 3737 88577 3760
rect 88663 3737 88729 3760
rect 88343 3718 88729 3737
rect 92343 3823 92729 3842
rect 92343 3800 92409 3823
rect 92495 3800 92577 3823
rect 92663 3800 92729 3823
rect 92343 3760 92352 3800
rect 92392 3760 92409 3800
rect 92495 3760 92516 3800
rect 92556 3760 92577 3800
rect 92663 3760 92680 3800
rect 92720 3760 92729 3800
rect 92343 3737 92409 3760
rect 92495 3737 92577 3760
rect 92663 3737 92729 3760
rect 92343 3718 92729 3737
rect 96343 3823 96729 3842
rect 96343 3800 96409 3823
rect 96495 3800 96577 3823
rect 96663 3800 96729 3823
rect 96343 3760 96352 3800
rect 96392 3760 96409 3800
rect 96495 3760 96516 3800
rect 96556 3760 96577 3800
rect 96663 3760 96680 3800
rect 96720 3760 96729 3800
rect 96343 3737 96409 3760
rect 96495 3737 96577 3760
rect 96663 3737 96729 3760
rect 96343 3718 96729 3737
rect 3103 3067 3489 3086
rect 3103 3044 3169 3067
rect 3255 3044 3337 3067
rect 3423 3044 3489 3067
rect 3103 3004 3112 3044
rect 3152 3004 3169 3044
rect 3255 3004 3276 3044
rect 3316 3004 3337 3044
rect 3423 3004 3440 3044
rect 3480 3004 3489 3044
rect 3103 2981 3169 3004
rect 3255 2981 3337 3004
rect 3423 2981 3489 3004
rect 3103 2962 3489 2981
rect 7103 3067 7489 3086
rect 7103 3044 7169 3067
rect 7255 3044 7337 3067
rect 7423 3044 7489 3067
rect 7103 3004 7112 3044
rect 7152 3004 7169 3044
rect 7255 3004 7276 3044
rect 7316 3004 7337 3044
rect 7423 3004 7440 3044
rect 7480 3004 7489 3044
rect 7103 2981 7169 3004
rect 7255 2981 7337 3004
rect 7423 2981 7489 3004
rect 7103 2962 7489 2981
rect 11103 3067 11489 3086
rect 11103 3044 11169 3067
rect 11255 3044 11337 3067
rect 11423 3044 11489 3067
rect 11103 3004 11112 3044
rect 11152 3004 11169 3044
rect 11255 3004 11276 3044
rect 11316 3004 11337 3044
rect 11423 3004 11440 3044
rect 11480 3004 11489 3044
rect 11103 2981 11169 3004
rect 11255 2981 11337 3004
rect 11423 2981 11489 3004
rect 11103 2962 11489 2981
rect 15103 3067 15489 3086
rect 15103 3044 15169 3067
rect 15255 3044 15337 3067
rect 15423 3044 15489 3067
rect 15103 3004 15112 3044
rect 15152 3004 15169 3044
rect 15255 3004 15276 3044
rect 15316 3004 15337 3044
rect 15423 3004 15440 3044
rect 15480 3004 15489 3044
rect 15103 2981 15169 3004
rect 15255 2981 15337 3004
rect 15423 2981 15489 3004
rect 15103 2962 15489 2981
rect 19103 3067 19489 3086
rect 19103 3044 19169 3067
rect 19255 3044 19337 3067
rect 19423 3044 19489 3067
rect 19103 3004 19112 3044
rect 19152 3004 19169 3044
rect 19255 3004 19276 3044
rect 19316 3004 19337 3044
rect 19423 3004 19440 3044
rect 19480 3004 19489 3044
rect 19103 2981 19169 3004
rect 19255 2981 19337 3004
rect 19423 2981 19489 3004
rect 19103 2962 19489 2981
rect 23103 3067 23489 3086
rect 23103 3044 23169 3067
rect 23255 3044 23337 3067
rect 23423 3044 23489 3067
rect 23103 3004 23112 3044
rect 23152 3004 23169 3044
rect 23255 3004 23276 3044
rect 23316 3004 23337 3044
rect 23423 3004 23440 3044
rect 23480 3004 23489 3044
rect 23103 2981 23169 3004
rect 23255 2981 23337 3004
rect 23423 2981 23489 3004
rect 23103 2962 23489 2981
rect 27103 3067 27489 3086
rect 27103 3044 27169 3067
rect 27255 3044 27337 3067
rect 27423 3044 27489 3067
rect 27103 3004 27112 3044
rect 27152 3004 27169 3044
rect 27255 3004 27276 3044
rect 27316 3004 27337 3044
rect 27423 3004 27440 3044
rect 27480 3004 27489 3044
rect 27103 2981 27169 3004
rect 27255 2981 27337 3004
rect 27423 2981 27489 3004
rect 27103 2962 27489 2981
rect 31103 3067 31489 3086
rect 31103 3044 31169 3067
rect 31255 3044 31337 3067
rect 31423 3044 31489 3067
rect 31103 3004 31112 3044
rect 31152 3004 31169 3044
rect 31255 3004 31276 3044
rect 31316 3004 31337 3044
rect 31423 3004 31440 3044
rect 31480 3004 31489 3044
rect 31103 2981 31169 3004
rect 31255 2981 31337 3004
rect 31423 2981 31489 3004
rect 31103 2962 31489 2981
rect 35103 3067 35489 3086
rect 35103 3044 35169 3067
rect 35255 3044 35337 3067
rect 35423 3044 35489 3067
rect 35103 3004 35112 3044
rect 35152 3004 35169 3044
rect 35255 3004 35276 3044
rect 35316 3004 35337 3044
rect 35423 3004 35440 3044
rect 35480 3004 35489 3044
rect 35103 2981 35169 3004
rect 35255 2981 35337 3004
rect 35423 2981 35489 3004
rect 35103 2962 35489 2981
rect 39103 3067 39489 3086
rect 39103 3044 39169 3067
rect 39255 3044 39337 3067
rect 39423 3044 39489 3067
rect 39103 3004 39112 3044
rect 39152 3004 39169 3044
rect 39255 3004 39276 3044
rect 39316 3004 39337 3044
rect 39423 3004 39440 3044
rect 39480 3004 39489 3044
rect 39103 2981 39169 3004
rect 39255 2981 39337 3004
rect 39423 2981 39489 3004
rect 39103 2962 39489 2981
rect 43103 3067 43489 3086
rect 43103 3044 43169 3067
rect 43255 3044 43337 3067
rect 43423 3044 43489 3067
rect 43103 3004 43112 3044
rect 43152 3004 43169 3044
rect 43255 3004 43276 3044
rect 43316 3004 43337 3044
rect 43423 3004 43440 3044
rect 43480 3004 43489 3044
rect 43103 2981 43169 3004
rect 43255 2981 43337 3004
rect 43423 2981 43489 3004
rect 43103 2962 43489 2981
rect 47103 3067 47489 3086
rect 47103 3044 47169 3067
rect 47255 3044 47337 3067
rect 47423 3044 47489 3067
rect 47103 3004 47112 3044
rect 47152 3004 47169 3044
rect 47255 3004 47276 3044
rect 47316 3004 47337 3044
rect 47423 3004 47440 3044
rect 47480 3004 47489 3044
rect 47103 2981 47169 3004
rect 47255 2981 47337 3004
rect 47423 2981 47489 3004
rect 47103 2962 47489 2981
rect 51103 3067 51489 3086
rect 51103 3044 51169 3067
rect 51255 3044 51337 3067
rect 51423 3044 51489 3067
rect 51103 3004 51112 3044
rect 51152 3004 51169 3044
rect 51255 3004 51276 3044
rect 51316 3004 51337 3044
rect 51423 3004 51440 3044
rect 51480 3004 51489 3044
rect 51103 2981 51169 3004
rect 51255 2981 51337 3004
rect 51423 2981 51489 3004
rect 51103 2962 51489 2981
rect 55103 3067 55489 3086
rect 55103 3044 55169 3067
rect 55255 3044 55337 3067
rect 55423 3044 55489 3067
rect 55103 3004 55112 3044
rect 55152 3004 55169 3044
rect 55255 3004 55276 3044
rect 55316 3004 55337 3044
rect 55423 3004 55440 3044
rect 55480 3004 55489 3044
rect 55103 2981 55169 3004
rect 55255 2981 55337 3004
rect 55423 2981 55489 3004
rect 55103 2962 55489 2981
rect 59103 3067 59489 3086
rect 59103 3044 59169 3067
rect 59255 3044 59337 3067
rect 59423 3044 59489 3067
rect 59103 3004 59112 3044
rect 59152 3004 59169 3044
rect 59255 3004 59276 3044
rect 59316 3004 59337 3044
rect 59423 3004 59440 3044
rect 59480 3004 59489 3044
rect 59103 2981 59169 3004
rect 59255 2981 59337 3004
rect 59423 2981 59489 3004
rect 59103 2962 59489 2981
rect 63103 3067 63489 3086
rect 63103 3044 63169 3067
rect 63255 3044 63337 3067
rect 63423 3044 63489 3067
rect 63103 3004 63112 3044
rect 63152 3004 63169 3044
rect 63255 3004 63276 3044
rect 63316 3004 63337 3044
rect 63423 3004 63440 3044
rect 63480 3004 63489 3044
rect 63103 2981 63169 3004
rect 63255 2981 63337 3004
rect 63423 2981 63489 3004
rect 63103 2962 63489 2981
rect 67103 3067 67489 3086
rect 67103 3044 67169 3067
rect 67255 3044 67337 3067
rect 67423 3044 67489 3067
rect 67103 3004 67112 3044
rect 67152 3004 67169 3044
rect 67255 3004 67276 3044
rect 67316 3004 67337 3044
rect 67423 3004 67440 3044
rect 67480 3004 67489 3044
rect 67103 2981 67169 3004
rect 67255 2981 67337 3004
rect 67423 2981 67489 3004
rect 67103 2962 67489 2981
rect 71103 3067 71489 3086
rect 71103 3044 71169 3067
rect 71255 3044 71337 3067
rect 71423 3044 71489 3067
rect 71103 3004 71112 3044
rect 71152 3004 71169 3044
rect 71255 3004 71276 3044
rect 71316 3004 71337 3044
rect 71423 3004 71440 3044
rect 71480 3004 71489 3044
rect 71103 2981 71169 3004
rect 71255 2981 71337 3004
rect 71423 2981 71489 3004
rect 71103 2962 71489 2981
rect 75103 3067 75489 3086
rect 75103 3044 75169 3067
rect 75255 3044 75337 3067
rect 75423 3044 75489 3067
rect 75103 3004 75112 3044
rect 75152 3004 75169 3044
rect 75255 3004 75276 3044
rect 75316 3004 75337 3044
rect 75423 3004 75440 3044
rect 75480 3004 75489 3044
rect 75103 2981 75169 3004
rect 75255 2981 75337 3004
rect 75423 2981 75489 3004
rect 75103 2962 75489 2981
rect 79103 3067 79489 3086
rect 79103 3044 79169 3067
rect 79255 3044 79337 3067
rect 79423 3044 79489 3067
rect 79103 3004 79112 3044
rect 79152 3004 79169 3044
rect 79255 3004 79276 3044
rect 79316 3004 79337 3044
rect 79423 3004 79440 3044
rect 79480 3004 79489 3044
rect 79103 2981 79169 3004
rect 79255 2981 79337 3004
rect 79423 2981 79489 3004
rect 79103 2962 79489 2981
rect 83103 3067 83489 3086
rect 83103 3044 83169 3067
rect 83255 3044 83337 3067
rect 83423 3044 83489 3067
rect 83103 3004 83112 3044
rect 83152 3004 83169 3044
rect 83255 3004 83276 3044
rect 83316 3004 83337 3044
rect 83423 3004 83440 3044
rect 83480 3004 83489 3044
rect 83103 2981 83169 3004
rect 83255 2981 83337 3004
rect 83423 2981 83489 3004
rect 83103 2962 83489 2981
rect 87103 3067 87489 3086
rect 87103 3044 87169 3067
rect 87255 3044 87337 3067
rect 87423 3044 87489 3067
rect 87103 3004 87112 3044
rect 87152 3004 87169 3044
rect 87255 3004 87276 3044
rect 87316 3004 87337 3044
rect 87423 3004 87440 3044
rect 87480 3004 87489 3044
rect 87103 2981 87169 3004
rect 87255 2981 87337 3004
rect 87423 2981 87489 3004
rect 87103 2962 87489 2981
rect 91103 3067 91489 3086
rect 91103 3044 91169 3067
rect 91255 3044 91337 3067
rect 91423 3044 91489 3067
rect 91103 3004 91112 3044
rect 91152 3004 91169 3044
rect 91255 3004 91276 3044
rect 91316 3004 91337 3044
rect 91423 3004 91440 3044
rect 91480 3004 91489 3044
rect 91103 2981 91169 3004
rect 91255 2981 91337 3004
rect 91423 2981 91489 3004
rect 91103 2962 91489 2981
rect 95103 3067 95489 3086
rect 95103 3044 95169 3067
rect 95255 3044 95337 3067
rect 95423 3044 95489 3067
rect 95103 3004 95112 3044
rect 95152 3004 95169 3044
rect 95255 3004 95276 3044
rect 95316 3004 95337 3044
rect 95423 3004 95440 3044
rect 95480 3004 95489 3044
rect 95103 2981 95169 3004
rect 95255 2981 95337 3004
rect 95423 2981 95489 3004
rect 95103 2962 95489 2981
rect 99103 3067 99489 3086
rect 99103 3044 99169 3067
rect 99255 3044 99337 3067
rect 99423 3044 99489 3067
rect 99103 3004 99112 3044
rect 99152 3004 99169 3044
rect 99255 3004 99276 3044
rect 99316 3004 99337 3044
rect 99423 3004 99440 3044
rect 99480 3004 99489 3044
rect 99103 2981 99169 3004
rect 99255 2981 99337 3004
rect 99423 2981 99489 3004
rect 99103 2962 99489 2981
rect 4343 2311 4729 2330
rect 4343 2288 4409 2311
rect 4495 2288 4577 2311
rect 4663 2288 4729 2311
rect 4343 2248 4352 2288
rect 4392 2248 4409 2288
rect 4495 2248 4516 2288
rect 4556 2248 4577 2288
rect 4663 2248 4680 2288
rect 4720 2248 4729 2288
rect 4343 2225 4409 2248
rect 4495 2225 4577 2248
rect 4663 2225 4729 2248
rect 4343 2206 4729 2225
rect 8343 2311 8729 2330
rect 8343 2288 8409 2311
rect 8495 2288 8577 2311
rect 8663 2288 8729 2311
rect 8343 2248 8352 2288
rect 8392 2248 8409 2288
rect 8495 2248 8516 2288
rect 8556 2248 8577 2288
rect 8663 2248 8680 2288
rect 8720 2248 8729 2288
rect 8343 2225 8409 2248
rect 8495 2225 8577 2248
rect 8663 2225 8729 2248
rect 8343 2206 8729 2225
rect 12343 2311 12729 2330
rect 12343 2288 12409 2311
rect 12495 2288 12577 2311
rect 12663 2288 12729 2311
rect 12343 2248 12352 2288
rect 12392 2248 12409 2288
rect 12495 2248 12516 2288
rect 12556 2248 12577 2288
rect 12663 2248 12680 2288
rect 12720 2248 12729 2288
rect 12343 2225 12409 2248
rect 12495 2225 12577 2248
rect 12663 2225 12729 2248
rect 12343 2206 12729 2225
rect 16343 2311 16729 2330
rect 16343 2288 16409 2311
rect 16495 2288 16577 2311
rect 16663 2288 16729 2311
rect 16343 2248 16352 2288
rect 16392 2248 16409 2288
rect 16495 2248 16516 2288
rect 16556 2248 16577 2288
rect 16663 2248 16680 2288
rect 16720 2248 16729 2288
rect 16343 2225 16409 2248
rect 16495 2225 16577 2248
rect 16663 2225 16729 2248
rect 16343 2206 16729 2225
rect 20343 2311 20729 2330
rect 20343 2288 20409 2311
rect 20495 2288 20577 2311
rect 20663 2288 20729 2311
rect 20343 2248 20352 2288
rect 20392 2248 20409 2288
rect 20495 2248 20516 2288
rect 20556 2248 20577 2288
rect 20663 2248 20680 2288
rect 20720 2248 20729 2288
rect 20343 2225 20409 2248
rect 20495 2225 20577 2248
rect 20663 2225 20729 2248
rect 20343 2206 20729 2225
rect 24343 2311 24729 2330
rect 24343 2288 24409 2311
rect 24495 2288 24577 2311
rect 24663 2288 24729 2311
rect 24343 2248 24352 2288
rect 24392 2248 24409 2288
rect 24495 2248 24516 2288
rect 24556 2248 24577 2288
rect 24663 2248 24680 2288
rect 24720 2248 24729 2288
rect 24343 2225 24409 2248
rect 24495 2225 24577 2248
rect 24663 2225 24729 2248
rect 24343 2206 24729 2225
rect 28343 2311 28729 2330
rect 28343 2288 28409 2311
rect 28495 2288 28577 2311
rect 28663 2288 28729 2311
rect 28343 2248 28352 2288
rect 28392 2248 28409 2288
rect 28495 2248 28516 2288
rect 28556 2248 28577 2288
rect 28663 2248 28680 2288
rect 28720 2248 28729 2288
rect 28343 2225 28409 2248
rect 28495 2225 28577 2248
rect 28663 2225 28729 2248
rect 28343 2206 28729 2225
rect 32343 2311 32729 2330
rect 32343 2288 32409 2311
rect 32495 2288 32577 2311
rect 32663 2288 32729 2311
rect 32343 2248 32352 2288
rect 32392 2248 32409 2288
rect 32495 2248 32516 2288
rect 32556 2248 32577 2288
rect 32663 2248 32680 2288
rect 32720 2248 32729 2288
rect 32343 2225 32409 2248
rect 32495 2225 32577 2248
rect 32663 2225 32729 2248
rect 32343 2206 32729 2225
rect 36343 2311 36729 2330
rect 36343 2288 36409 2311
rect 36495 2288 36577 2311
rect 36663 2288 36729 2311
rect 36343 2248 36352 2288
rect 36392 2248 36409 2288
rect 36495 2248 36516 2288
rect 36556 2248 36577 2288
rect 36663 2248 36680 2288
rect 36720 2248 36729 2288
rect 36343 2225 36409 2248
rect 36495 2225 36577 2248
rect 36663 2225 36729 2248
rect 36343 2206 36729 2225
rect 40343 2311 40729 2330
rect 40343 2288 40409 2311
rect 40495 2288 40577 2311
rect 40663 2288 40729 2311
rect 40343 2248 40352 2288
rect 40392 2248 40409 2288
rect 40495 2248 40516 2288
rect 40556 2248 40577 2288
rect 40663 2248 40680 2288
rect 40720 2248 40729 2288
rect 40343 2225 40409 2248
rect 40495 2225 40577 2248
rect 40663 2225 40729 2248
rect 40343 2206 40729 2225
rect 44343 2311 44729 2330
rect 44343 2288 44409 2311
rect 44495 2288 44577 2311
rect 44663 2288 44729 2311
rect 44343 2248 44352 2288
rect 44392 2248 44409 2288
rect 44495 2248 44516 2288
rect 44556 2248 44577 2288
rect 44663 2248 44680 2288
rect 44720 2248 44729 2288
rect 44343 2225 44409 2248
rect 44495 2225 44577 2248
rect 44663 2225 44729 2248
rect 44343 2206 44729 2225
rect 48343 2311 48729 2330
rect 48343 2288 48409 2311
rect 48495 2288 48577 2311
rect 48663 2288 48729 2311
rect 48343 2248 48352 2288
rect 48392 2248 48409 2288
rect 48495 2248 48516 2288
rect 48556 2248 48577 2288
rect 48663 2248 48680 2288
rect 48720 2248 48729 2288
rect 48343 2225 48409 2248
rect 48495 2225 48577 2248
rect 48663 2225 48729 2248
rect 48343 2206 48729 2225
rect 52343 2311 52729 2330
rect 52343 2288 52409 2311
rect 52495 2288 52577 2311
rect 52663 2288 52729 2311
rect 52343 2248 52352 2288
rect 52392 2248 52409 2288
rect 52495 2248 52516 2288
rect 52556 2248 52577 2288
rect 52663 2248 52680 2288
rect 52720 2248 52729 2288
rect 52343 2225 52409 2248
rect 52495 2225 52577 2248
rect 52663 2225 52729 2248
rect 52343 2206 52729 2225
rect 56343 2311 56729 2330
rect 56343 2288 56409 2311
rect 56495 2288 56577 2311
rect 56663 2288 56729 2311
rect 56343 2248 56352 2288
rect 56392 2248 56409 2288
rect 56495 2248 56516 2288
rect 56556 2248 56577 2288
rect 56663 2248 56680 2288
rect 56720 2248 56729 2288
rect 56343 2225 56409 2248
rect 56495 2225 56577 2248
rect 56663 2225 56729 2248
rect 56343 2206 56729 2225
rect 60343 2311 60729 2330
rect 60343 2288 60409 2311
rect 60495 2288 60577 2311
rect 60663 2288 60729 2311
rect 60343 2248 60352 2288
rect 60392 2248 60409 2288
rect 60495 2248 60516 2288
rect 60556 2248 60577 2288
rect 60663 2248 60680 2288
rect 60720 2248 60729 2288
rect 60343 2225 60409 2248
rect 60495 2225 60577 2248
rect 60663 2225 60729 2248
rect 60343 2206 60729 2225
rect 64343 2311 64729 2330
rect 64343 2288 64409 2311
rect 64495 2288 64577 2311
rect 64663 2288 64729 2311
rect 64343 2248 64352 2288
rect 64392 2248 64409 2288
rect 64495 2248 64516 2288
rect 64556 2248 64577 2288
rect 64663 2248 64680 2288
rect 64720 2248 64729 2288
rect 64343 2225 64409 2248
rect 64495 2225 64577 2248
rect 64663 2225 64729 2248
rect 64343 2206 64729 2225
rect 68343 2311 68729 2330
rect 68343 2288 68409 2311
rect 68495 2288 68577 2311
rect 68663 2288 68729 2311
rect 68343 2248 68352 2288
rect 68392 2248 68409 2288
rect 68495 2248 68516 2288
rect 68556 2248 68577 2288
rect 68663 2248 68680 2288
rect 68720 2248 68729 2288
rect 68343 2225 68409 2248
rect 68495 2225 68577 2248
rect 68663 2225 68729 2248
rect 68343 2206 68729 2225
rect 72343 2311 72729 2330
rect 72343 2288 72409 2311
rect 72495 2288 72577 2311
rect 72663 2288 72729 2311
rect 72343 2248 72352 2288
rect 72392 2248 72409 2288
rect 72495 2248 72516 2288
rect 72556 2248 72577 2288
rect 72663 2248 72680 2288
rect 72720 2248 72729 2288
rect 72343 2225 72409 2248
rect 72495 2225 72577 2248
rect 72663 2225 72729 2248
rect 72343 2206 72729 2225
rect 76343 2311 76729 2330
rect 76343 2288 76409 2311
rect 76495 2288 76577 2311
rect 76663 2288 76729 2311
rect 76343 2248 76352 2288
rect 76392 2248 76409 2288
rect 76495 2248 76516 2288
rect 76556 2248 76577 2288
rect 76663 2248 76680 2288
rect 76720 2248 76729 2288
rect 76343 2225 76409 2248
rect 76495 2225 76577 2248
rect 76663 2225 76729 2248
rect 76343 2206 76729 2225
rect 80343 2311 80729 2330
rect 80343 2288 80409 2311
rect 80495 2288 80577 2311
rect 80663 2288 80729 2311
rect 80343 2248 80352 2288
rect 80392 2248 80409 2288
rect 80495 2248 80516 2288
rect 80556 2248 80577 2288
rect 80663 2248 80680 2288
rect 80720 2248 80729 2288
rect 80343 2225 80409 2248
rect 80495 2225 80577 2248
rect 80663 2225 80729 2248
rect 80343 2206 80729 2225
rect 84343 2311 84729 2330
rect 84343 2288 84409 2311
rect 84495 2288 84577 2311
rect 84663 2288 84729 2311
rect 84343 2248 84352 2288
rect 84392 2248 84409 2288
rect 84495 2248 84516 2288
rect 84556 2248 84577 2288
rect 84663 2248 84680 2288
rect 84720 2248 84729 2288
rect 84343 2225 84409 2248
rect 84495 2225 84577 2248
rect 84663 2225 84729 2248
rect 84343 2206 84729 2225
rect 88343 2311 88729 2330
rect 88343 2288 88409 2311
rect 88495 2288 88577 2311
rect 88663 2288 88729 2311
rect 88343 2248 88352 2288
rect 88392 2248 88409 2288
rect 88495 2248 88516 2288
rect 88556 2248 88577 2288
rect 88663 2248 88680 2288
rect 88720 2248 88729 2288
rect 88343 2225 88409 2248
rect 88495 2225 88577 2248
rect 88663 2225 88729 2248
rect 88343 2206 88729 2225
rect 92343 2311 92729 2330
rect 92343 2288 92409 2311
rect 92495 2288 92577 2311
rect 92663 2288 92729 2311
rect 92343 2248 92352 2288
rect 92392 2248 92409 2288
rect 92495 2248 92516 2288
rect 92556 2248 92577 2288
rect 92663 2248 92680 2288
rect 92720 2248 92729 2288
rect 92343 2225 92409 2248
rect 92495 2225 92577 2248
rect 92663 2225 92729 2248
rect 92343 2206 92729 2225
rect 96343 2311 96729 2330
rect 96343 2288 96409 2311
rect 96495 2288 96577 2311
rect 96663 2288 96729 2311
rect 96343 2248 96352 2288
rect 96392 2248 96409 2288
rect 96495 2248 96516 2288
rect 96556 2248 96577 2288
rect 96663 2248 96680 2288
rect 96720 2248 96729 2288
rect 96343 2225 96409 2248
rect 96495 2225 96577 2248
rect 96663 2225 96729 2248
rect 96343 2206 96729 2225
rect 3103 1555 3489 1574
rect 3103 1532 3169 1555
rect 3255 1532 3337 1555
rect 3423 1532 3489 1555
rect 3103 1492 3112 1532
rect 3152 1492 3169 1532
rect 3255 1492 3276 1532
rect 3316 1492 3337 1532
rect 3423 1492 3440 1532
rect 3480 1492 3489 1532
rect 3103 1469 3169 1492
rect 3255 1469 3337 1492
rect 3423 1469 3489 1492
rect 3103 1450 3489 1469
rect 7103 1555 7489 1574
rect 7103 1532 7169 1555
rect 7255 1532 7337 1555
rect 7423 1532 7489 1555
rect 7103 1492 7112 1532
rect 7152 1492 7169 1532
rect 7255 1492 7276 1532
rect 7316 1492 7337 1532
rect 7423 1492 7440 1532
rect 7480 1492 7489 1532
rect 7103 1469 7169 1492
rect 7255 1469 7337 1492
rect 7423 1469 7489 1492
rect 7103 1450 7489 1469
rect 11103 1555 11489 1574
rect 11103 1532 11169 1555
rect 11255 1532 11337 1555
rect 11423 1532 11489 1555
rect 11103 1492 11112 1532
rect 11152 1492 11169 1532
rect 11255 1492 11276 1532
rect 11316 1492 11337 1532
rect 11423 1492 11440 1532
rect 11480 1492 11489 1532
rect 11103 1469 11169 1492
rect 11255 1469 11337 1492
rect 11423 1469 11489 1492
rect 11103 1450 11489 1469
rect 15103 1555 15489 1574
rect 15103 1532 15169 1555
rect 15255 1532 15337 1555
rect 15423 1532 15489 1555
rect 15103 1492 15112 1532
rect 15152 1492 15169 1532
rect 15255 1492 15276 1532
rect 15316 1492 15337 1532
rect 15423 1492 15440 1532
rect 15480 1492 15489 1532
rect 15103 1469 15169 1492
rect 15255 1469 15337 1492
rect 15423 1469 15489 1492
rect 15103 1450 15489 1469
rect 19103 1555 19489 1574
rect 19103 1532 19169 1555
rect 19255 1532 19337 1555
rect 19423 1532 19489 1555
rect 19103 1492 19112 1532
rect 19152 1492 19169 1532
rect 19255 1492 19276 1532
rect 19316 1492 19337 1532
rect 19423 1492 19440 1532
rect 19480 1492 19489 1532
rect 19103 1469 19169 1492
rect 19255 1469 19337 1492
rect 19423 1469 19489 1492
rect 19103 1450 19489 1469
rect 23103 1555 23489 1574
rect 23103 1532 23169 1555
rect 23255 1532 23337 1555
rect 23423 1532 23489 1555
rect 23103 1492 23112 1532
rect 23152 1492 23169 1532
rect 23255 1492 23276 1532
rect 23316 1492 23337 1532
rect 23423 1492 23440 1532
rect 23480 1492 23489 1532
rect 23103 1469 23169 1492
rect 23255 1469 23337 1492
rect 23423 1469 23489 1492
rect 23103 1450 23489 1469
rect 27103 1555 27489 1574
rect 27103 1532 27169 1555
rect 27255 1532 27337 1555
rect 27423 1532 27489 1555
rect 27103 1492 27112 1532
rect 27152 1492 27169 1532
rect 27255 1492 27276 1532
rect 27316 1492 27337 1532
rect 27423 1492 27440 1532
rect 27480 1492 27489 1532
rect 27103 1469 27169 1492
rect 27255 1469 27337 1492
rect 27423 1469 27489 1492
rect 27103 1450 27489 1469
rect 31103 1555 31489 1574
rect 31103 1532 31169 1555
rect 31255 1532 31337 1555
rect 31423 1532 31489 1555
rect 31103 1492 31112 1532
rect 31152 1492 31169 1532
rect 31255 1492 31276 1532
rect 31316 1492 31337 1532
rect 31423 1492 31440 1532
rect 31480 1492 31489 1532
rect 31103 1469 31169 1492
rect 31255 1469 31337 1492
rect 31423 1469 31489 1492
rect 31103 1450 31489 1469
rect 35103 1555 35489 1574
rect 35103 1532 35169 1555
rect 35255 1532 35337 1555
rect 35423 1532 35489 1555
rect 35103 1492 35112 1532
rect 35152 1492 35169 1532
rect 35255 1492 35276 1532
rect 35316 1492 35337 1532
rect 35423 1492 35440 1532
rect 35480 1492 35489 1532
rect 35103 1469 35169 1492
rect 35255 1469 35337 1492
rect 35423 1469 35489 1492
rect 35103 1450 35489 1469
rect 39103 1555 39489 1574
rect 39103 1532 39169 1555
rect 39255 1532 39337 1555
rect 39423 1532 39489 1555
rect 39103 1492 39112 1532
rect 39152 1492 39169 1532
rect 39255 1492 39276 1532
rect 39316 1492 39337 1532
rect 39423 1492 39440 1532
rect 39480 1492 39489 1532
rect 39103 1469 39169 1492
rect 39255 1469 39337 1492
rect 39423 1469 39489 1492
rect 39103 1450 39489 1469
rect 43103 1555 43489 1574
rect 43103 1532 43169 1555
rect 43255 1532 43337 1555
rect 43423 1532 43489 1555
rect 43103 1492 43112 1532
rect 43152 1492 43169 1532
rect 43255 1492 43276 1532
rect 43316 1492 43337 1532
rect 43423 1492 43440 1532
rect 43480 1492 43489 1532
rect 43103 1469 43169 1492
rect 43255 1469 43337 1492
rect 43423 1469 43489 1492
rect 43103 1450 43489 1469
rect 47103 1555 47489 1574
rect 47103 1532 47169 1555
rect 47255 1532 47337 1555
rect 47423 1532 47489 1555
rect 47103 1492 47112 1532
rect 47152 1492 47169 1532
rect 47255 1492 47276 1532
rect 47316 1492 47337 1532
rect 47423 1492 47440 1532
rect 47480 1492 47489 1532
rect 47103 1469 47169 1492
rect 47255 1469 47337 1492
rect 47423 1469 47489 1492
rect 47103 1450 47489 1469
rect 51103 1555 51489 1574
rect 51103 1532 51169 1555
rect 51255 1532 51337 1555
rect 51423 1532 51489 1555
rect 51103 1492 51112 1532
rect 51152 1492 51169 1532
rect 51255 1492 51276 1532
rect 51316 1492 51337 1532
rect 51423 1492 51440 1532
rect 51480 1492 51489 1532
rect 51103 1469 51169 1492
rect 51255 1469 51337 1492
rect 51423 1469 51489 1492
rect 51103 1450 51489 1469
rect 55103 1555 55489 1574
rect 55103 1532 55169 1555
rect 55255 1532 55337 1555
rect 55423 1532 55489 1555
rect 55103 1492 55112 1532
rect 55152 1492 55169 1532
rect 55255 1492 55276 1532
rect 55316 1492 55337 1532
rect 55423 1492 55440 1532
rect 55480 1492 55489 1532
rect 55103 1469 55169 1492
rect 55255 1469 55337 1492
rect 55423 1469 55489 1492
rect 55103 1450 55489 1469
rect 59103 1555 59489 1574
rect 59103 1532 59169 1555
rect 59255 1532 59337 1555
rect 59423 1532 59489 1555
rect 59103 1492 59112 1532
rect 59152 1492 59169 1532
rect 59255 1492 59276 1532
rect 59316 1492 59337 1532
rect 59423 1492 59440 1532
rect 59480 1492 59489 1532
rect 59103 1469 59169 1492
rect 59255 1469 59337 1492
rect 59423 1469 59489 1492
rect 59103 1450 59489 1469
rect 63103 1555 63489 1574
rect 63103 1532 63169 1555
rect 63255 1532 63337 1555
rect 63423 1532 63489 1555
rect 63103 1492 63112 1532
rect 63152 1492 63169 1532
rect 63255 1492 63276 1532
rect 63316 1492 63337 1532
rect 63423 1492 63440 1532
rect 63480 1492 63489 1532
rect 63103 1469 63169 1492
rect 63255 1469 63337 1492
rect 63423 1469 63489 1492
rect 63103 1450 63489 1469
rect 67103 1555 67489 1574
rect 67103 1532 67169 1555
rect 67255 1532 67337 1555
rect 67423 1532 67489 1555
rect 67103 1492 67112 1532
rect 67152 1492 67169 1532
rect 67255 1492 67276 1532
rect 67316 1492 67337 1532
rect 67423 1492 67440 1532
rect 67480 1492 67489 1532
rect 67103 1469 67169 1492
rect 67255 1469 67337 1492
rect 67423 1469 67489 1492
rect 67103 1450 67489 1469
rect 71103 1555 71489 1574
rect 71103 1532 71169 1555
rect 71255 1532 71337 1555
rect 71423 1532 71489 1555
rect 71103 1492 71112 1532
rect 71152 1492 71169 1532
rect 71255 1492 71276 1532
rect 71316 1492 71337 1532
rect 71423 1492 71440 1532
rect 71480 1492 71489 1532
rect 71103 1469 71169 1492
rect 71255 1469 71337 1492
rect 71423 1469 71489 1492
rect 71103 1450 71489 1469
rect 75103 1555 75489 1574
rect 75103 1532 75169 1555
rect 75255 1532 75337 1555
rect 75423 1532 75489 1555
rect 75103 1492 75112 1532
rect 75152 1492 75169 1532
rect 75255 1492 75276 1532
rect 75316 1492 75337 1532
rect 75423 1492 75440 1532
rect 75480 1492 75489 1532
rect 75103 1469 75169 1492
rect 75255 1469 75337 1492
rect 75423 1469 75489 1492
rect 75103 1450 75489 1469
rect 79103 1555 79489 1574
rect 79103 1532 79169 1555
rect 79255 1532 79337 1555
rect 79423 1532 79489 1555
rect 79103 1492 79112 1532
rect 79152 1492 79169 1532
rect 79255 1492 79276 1532
rect 79316 1492 79337 1532
rect 79423 1492 79440 1532
rect 79480 1492 79489 1532
rect 79103 1469 79169 1492
rect 79255 1469 79337 1492
rect 79423 1469 79489 1492
rect 79103 1450 79489 1469
rect 83103 1555 83489 1574
rect 83103 1532 83169 1555
rect 83255 1532 83337 1555
rect 83423 1532 83489 1555
rect 83103 1492 83112 1532
rect 83152 1492 83169 1532
rect 83255 1492 83276 1532
rect 83316 1492 83337 1532
rect 83423 1492 83440 1532
rect 83480 1492 83489 1532
rect 83103 1469 83169 1492
rect 83255 1469 83337 1492
rect 83423 1469 83489 1492
rect 83103 1450 83489 1469
rect 87103 1555 87489 1574
rect 87103 1532 87169 1555
rect 87255 1532 87337 1555
rect 87423 1532 87489 1555
rect 87103 1492 87112 1532
rect 87152 1492 87169 1532
rect 87255 1492 87276 1532
rect 87316 1492 87337 1532
rect 87423 1492 87440 1532
rect 87480 1492 87489 1532
rect 87103 1469 87169 1492
rect 87255 1469 87337 1492
rect 87423 1469 87489 1492
rect 87103 1450 87489 1469
rect 91103 1555 91489 1574
rect 91103 1532 91169 1555
rect 91255 1532 91337 1555
rect 91423 1532 91489 1555
rect 91103 1492 91112 1532
rect 91152 1492 91169 1532
rect 91255 1492 91276 1532
rect 91316 1492 91337 1532
rect 91423 1492 91440 1532
rect 91480 1492 91489 1532
rect 91103 1469 91169 1492
rect 91255 1469 91337 1492
rect 91423 1469 91489 1492
rect 91103 1450 91489 1469
rect 95103 1555 95489 1574
rect 95103 1532 95169 1555
rect 95255 1532 95337 1555
rect 95423 1532 95489 1555
rect 95103 1492 95112 1532
rect 95152 1492 95169 1532
rect 95255 1492 95276 1532
rect 95316 1492 95337 1532
rect 95423 1492 95440 1532
rect 95480 1492 95489 1532
rect 95103 1469 95169 1492
rect 95255 1469 95337 1492
rect 95423 1469 95489 1492
rect 95103 1450 95489 1469
rect 99103 1555 99489 1574
rect 99103 1532 99169 1555
rect 99255 1532 99337 1555
rect 99423 1532 99489 1555
rect 99103 1492 99112 1532
rect 99152 1492 99169 1532
rect 99255 1492 99276 1532
rect 99316 1492 99337 1532
rect 99423 1492 99440 1532
rect 99480 1492 99489 1532
rect 99103 1469 99169 1492
rect 99255 1469 99337 1492
rect 99423 1469 99489 1492
rect 99103 1450 99489 1469
rect 4343 799 4729 818
rect 4343 776 4409 799
rect 4495 776 4577 799
rect 4663 776 4729 799
rect 4343 736 4352 776
rect 4392 736 4409 776
rect 4495 736 4516 776
rect 4556 736 4577 776
rect 4663 736 4680 776
rect 4720 736 4729 776
rect 4343 713 4409 736
rect 4495 713 4577 736
rect 4663 713 4729 736
rect 4343 694 4729 713
rect 8343 799 8729 818
rect 8343 776 8409 799
rect 8495 776 8577 799
rect 8663 776 8729 799
rect 8343 736 8352 776
rect 8392 736 8409 776
rect 8495 736 8516 776
rect 8556 736 8577 776
rect 8663 736 8680 776
rect 8720 736 8729 776
rect 8343 713 8409 736
rect 8495 713 8577 736
rect 8663 713 8729 736
rect 8343 694 8729 713
rect 12343 799 12729 818
rect 12343 776 12409 799
rect 12495 776 12577 799
rect 12663 776 12729 799
rect 12343 736 12352 776
rect 12392 736 12409 776
rect 12495 736 12516 776
rect 12556 736 12577 776
rect 12663 736 12680 776
rect 12720 736 12729 776
rect 12343 713 12409 736
rect 12495 713 12577 736
rect 12663 713 12729 736
rect 12343 694 12729 713
rect 16343 799 16729 818
rect 16343 776 16409 799
rect 16495 776 16577 799
rect 16663 776 16729 799
rect 16343 736 16352 776
rect 16392 736 16409 776
rect 16495 736 16516 776
rect 16556 736 16577 776
rect 16663 736 16680 776
rect 16720 736 16729 776
rect 16343 713 16409 736
rect 16495 713 16577 736
rect 16663 713 16729 736
rect 16343 694 16729 713
rect 20343 799 20729 818
rect 20343 776 20409 799
rect 20495 776 20577 799
rect 20663 776 20729 799
rect 20343 736 20352 776
rect 20392 736 20409 776
rect 20495 736 20516 776
rect 20556 736 20577 776
rect 20663 736 20680 776
rect 20720 736 20729 776
rect 20343 713 20409 736
rect 20495 713 20577 736
rect 20663 713 20729 736
rect 20343 694 20729 713
rect 24343 799 24729 818
rect 24343 776 24409 799
rect 24495 776 24577 799
rect 24663 776 24729 799
rect 24343 736 24352 776
rect 24392 736 24409 776
rect 24495 736 24516 776
rect 24556 736 24577 776
rect 24663 736 24680 776
rect 24720 736 24729 776
rect 24343 713 24409 736
rect 24495 713 24577 736
rect 24663 713 24729 736
rect 24343 694 24729 713
rect 28343 799 28729 818
rect 28343 776 28409 799
rect 28495 776 28577 799
rect 28663 776 28729 799
rect 28343 736 28352 776
rect 28392 736 28409 776
rect 28495 736 28516 776
rect 28556 736 28577 776
rect 28663 736 28680 776
rect 28720 736 28729 776
rect 28343 713 28409 736
rect 28495 713 28577 736
rect 28663 713 28729 736
rect 28343 694 28729 713
rect 32343 799 32729 818
rect 32343 776 32409 799
rect 32495 776 32577 799
rect 32663 776 32729 799
rect 32343 736 32352 776
rect 32392 736 32409 776
rect 32495 736 32516 776
rect 32556 736 32577 776
rect 32663 736 32680 776
rect 32720 736 32729 776
rect 32343 713 32409 736
rect 32495 713 32577 736
rect 32663 713 32729 736
rect 32343 694 32729 713
rect 36343 799 36729 818
rect 36343 776 36409 799
rect 36495 776 36577 799
rect 36663 776 36729 799
rect 36343 736 36352 776
rect 36392 736 36409 776
rect 36495 736 36516 776
rect 36556 736 36577 776
rect 36663 736 36680 776
rect 36720 736 36729 776
rect 36343 713 36409 736
rect 36495 713 36577 736
rect 36663 713 36729 736
rect 36343 694 36729 713
rect 40343 799 40729 818
rect 40343 776 40409 799
rect 40495 776 40577 799
rect 40663 776 40729 799
rect 40343 736 40352 776
rect 40392 736 40409 776
rect 40495 736 40516 776
rect 40556 736 40577 776
rect 40663 736 40680 776
rect 40720 736 40729 776
rect 40343 713 40409 736
rect 40495 713 40577 736
rect 40663 713 40729 736
rect 40343 694 40729 713
rect 44343 799 44729 818
rect 44343 776 44409 799
rect 44495 776 44577 799
rect 44663 776 44729 799
rect 44343 736 44352 776
rect 44392 736 44409 776
rect 44495 736 44516 776
rect 44556 736 44577 776
rect 44663 736 44680 776
rect 44720 736 44729 776
rect 44343 713 44409 736
rect 44495 713 44577 736
rect 44663 713 44729 736
rect 44343 694 44729 713
rect 48343 799 48729 818
rect 48343 776 48409 799
rect 48495 776 48577 799
rect 48663 776 48729 799
rect 48343 736 48352 776
rect 48392 736 48409 776
rect 48495 736 48516 776
rect 48556 736 48577 776
rect 48663 736 48680 776
rect 48720 736 48729 776
rect 48343 713 48409 736
rect 48495 713 48577 736
rect 48663 713 48729 736
rect 48343 694 48729 713
rect 52343 799 52729 818
rect 52343 776 52409 799
rect 52495 776 52577 799
rect 52663 776 52729 799
rect 52343 736 52352 776
rect 52392 736 52409 776
rect 52495 736 52516 776
rect 52556 736 52577 776
rect 52663 736 52680 776
rect 52720 736 52729 776
rect 52343 713 52409 736
rect 52495 713 52577 736
rect 52663 713 52729 736
rect 52343 694 52729 713
rect 56343 799 56729 818
rect 56343 776 56409 799
rect 56495 776 56577 799
rect 56663 776 56729 799
rect 56343 736 56352 776
rect 56392 736 56409 776
rect 56495 736 56516 776
rect 56556 736 56577 776
rect 56663 736 56680 776
rect 56720 736 56729 776
rect 56343 713 56409 736
rect 56495 713 56577 736
rect 56663 713 56729 736
rect 56343 694 56729 713
rect 60343 799 60729 818
rect 60343 776 60409 799
rect 60495 776 60577 799
rect 60663 776 60729 799
rect 60343 736 60352 776
rect 60392 736 60409 776
rect 60495 736 60516 776
rect 60556 736 60577 776
rect 60663 736 60680 776
rect 60720 736 60729 776
rect 60343 713 60409 736
rect 60495 713 60577 736
rect 60663 713 60729 736
rect 60343 694 60729 713
rect 64343 799 64729 818
rect 64343 776 64409 799
rect 64495 776 64577 799
rect 64663 776 64729 799
rect 64343 736 64352 776
rect 64392 736 64409 776
rect 64495 736 64516 776
rect 64556 736 64577 776
rect 64663 736 64680 776
rect 64720 736 64729 776
rect 64343 713 64409 736
rect 64495 713 64577 736
rect 64663 713 64729 736
rect 64343 694 64729 713
rect 68343 799 68729 818
rect 68343 776 68409 799
rect 68495 776 68577 799
rect 68663 776 68729 799
rect 68343 736 68352 776
rect 68392 736 68409 776
rect 68495 736 68516 776
rect 68556 736 68577 776
rect 68663 736 68680 776
rect 68720 736 68729 776
rect 68343 713 68409 736
rect 68495 713 68577 736
rect 68663 713 68729 736
rect 68343 694 68729 713
rect 72343 799 72729 818
rect 72343 776 72409 799
rect 72495 776 72577 799
rect 72663 776 72729 799
rect 72343 736 72352 776
rect 72392 736 72409 776
rect 72495 736 72516 776
rect 72556 736 72577 776
rect 72663 736 72680 776
rect 72720 736 72729 776
rect 72343 713 72409 736
rect 72495 713 72577 736
rect 72663 713 72729 736
rect 72343 694 72729 713
rect 76343 799 76729 818
rect 76343 776 76409 799
rect 76495 776 76577 799
rect 76663 776 76729 799
rect 76343 736 76352 776
rect 76392 736 76409 776
rect 76495 736 76516 776
rect 76556 736 76577 776
rect 76663 736 76680 776
rect 76720 736 76729 776
rect 76343 713 76409 736
rect 76495 713 76577 736
rect 76663 713 76729 736
rect 76343 694 76729 713
rect 80343 799 80729 818
rect 80343 776 80409 799
rect 80495 776 80577 799
rect 80663 776 80729 799
rect 80343 736 80352 776
rect 80392 736 80409 776
rect 80495 736 80516 776
rect 80556 736 80577 776
rect 80663 736 80680 776
rect 80720 736 80729 776
rect 80343 713 80409 736
rect 80495 713 80577 736
rect 80663 713 80729 736
rect 80343 694 80729 713
rect 84343 799 84729 818
rect 84343 776 84409 799
rect 84495 776 84577 799
rect 84663 776 84729 799
rect 84343 736 84352 776
rect 84392 736 84409 776
rect 84495 736 84516 776
rect 84556 736 84577 776
rect 84663 736 84680 776
rect 84720 736 84729 776
rect 84343 713 84409 736
rect 84495 713 84577 736
rect 84663 713 84729 736
rect 84343 694 84729 713
rect 88343 799 88729 818
rect 88343 776 88409 799
rect 88495 776 88577 799
rect 88663 776 88729 799
rect 88343 736 88352 776
rect 88392 736 88409 776
rect 88495 736 88516 776
rect 88556 736 88577 776
rect 88663 736 88680 776
rect 88720 736 88729 776
rect 88343 713 88409 736
rect 88495 713 88577 736
rect 88663 713 88729 736
rect 88343 694 88729 713
rect 92343 799 92729 818
rect 92343 776 92409 799
rect 92495 776 92577 799
rect 92663 776 92729 799
rect 92343 736 92352 776
rect 92392 736 92409 776
rect 92495 736 92516 776
rect 92556 736 92577 776
rect 92663 736 92680 776
rect 92720 736 92729 776
rect 92343 713 92409 736
rect 92495 713 92577 736
rect 92663 713 92729 736
rect 92343 694 92729 713
rect 96343 799 96729 818
rect 96343 776 96409 799
rect 96495 776 96577 799
rect 96663 776 96729 799
rect 96343 736 96352 776
rect 96392 736 96409 776
rect 96495 736 96516 776
rect 96556 736 96577 776
rect 96663 736 96680 776
rect 96720 736 96729 776
rect 96343 713 96409 736
rect 96495 713 96577 736
rect 96663 713 96729 736
rect 96343 694 96729 713
<< via5 >>
rect 4409 38576 4495 38599
rect 4577 38576 4663 38599
rect 4409 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4495 38576
rect 4577 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4663 38576
rect 4409 38513 4495 38536
rect 4577 38513 4663 38536
rect 8409 38576 8495 38599
rect 8577 38576 8663 38599
rect 8409 38536 8434 38576
rect 8434 38536 8474 38576
rect 8474 38536 8495 38576
rect 8577 38536 8598 38576
rect 8598 38536 8638 38576
rect 8638 38536 8663 38576
rect 8409 38513 8495 38536
rect 8577 38513 8663 38536
rect 12409 38576 12495 38599
rect 12577 38576 12663 38599
rect 12409 38536 12434 38576
rect 12434 38536 12474 38576
rect 12474 38536 12495 38576
rect 12577 38536 12598 38576
rect 12598 38536 12638 38576
rect 12638 38536 12663 38576
rect 12409 38513 12495 38536
rect 12577 38513 12663 38536
rect 16409 38576 16495 38599
rect 16577 38576 16663 38599
rect 16409 38536 16434 38576
rect 16434 38536 16474 38576
rect 16474 38536 16495 38576
rect 16577 38536 16598 38576
rect 16598 38536 16638 38576
rect 16638 38536 16663 38576
rect 16409 38513 16495 38536
rect 16577 38513 16663 38536
rect 20409 38576 20495 38599
rect 20577 38576 20663 38599
rect 20409 38536 20434 38576
rect 20434 38536 20474 38576
rect 20474 38536 20495 38576
rect 20577 38536 20598 38576
rect 20598 38536 20638 38576
rect 20638 38536 20663 38576
rect 20409 38513 20495 38536
rect 20577 38513 20663 38536
rect 24409 38576 24495 38599
rect 24577 38576 24663 38599
rect 24409 38536 24434 38576
rect 24434 38536 24474 38576
rect 24474 38536 24495 38576
rect 24577 38536 24598 38576
rect 24598 38536 24638 38576
rect 24638 38536 24663 38576
rect 24409 38513 24495 38536
rect 24577 38513 24663 38536
rect 28409 38576 28495 38599
rect 28577 38576 28663 38599
rect 28409 38536 28434 38576
rect 28434 38536 28474 38576
rect 28474 38536 28495 38576
rect 28577 38536 28598 38576
rect 28598 38536 28638 38576
rect 28638 38536 28663 38576
rect 28409 38513 28495 38536
rect 28577 38513 28663 38536
rect 32409 38576 32495 38599
rect 32577 38576 32663 38599
rect 32409 38536 32434 38576
rect 32434 38536 32474 38576
rect 32474 38536 32495 38576
rect 32577 38536 32598 38576
rect 32598 38536 32638 38576
rect 32638 38536 32663 38576
rect 32409 38513 32495 38536
rect 32577 38513 32663 38536
rect 36409 38576 36495 38599
rect 36577 38576 36663 38599
rect 36409 38536 36434 38576
rect 36434 38536 36474 38576
rect 36474 38536 36495 38576
rect 36577 38536 36598 38576
rect 36598 38536 36638 38576
rect 36638 38536 36663 38576
rect 36409 38513 36495 38536
rect 36577 38513 36663 38536
rect 40409 38576 40495 38599
rect 40577 38576 40663 38599
rect 40409 38536 40434 38576
rect 40434 38536 40474 38576
rect 40474 38536 40495 38576
rect 40577 38536 40598 38576
rect 40598 38536 40638 38576
rect 40638 38536 40663 38576
rect 40409 38513 40495 38536
rect 40577 38513 40663 38536
rect 44409 38576 44495 38599
rect 44577 38576 44663 38599
rect 44409 38536 44434 38576
rect 44434 38536 44474 38576
rect 44474 38536 44495 38576
rect 44577 38536 44598 38576
rect 44598 38536 44638 38576
rect 44638 38536 44663 38576
rect 44409 38513 44495 38536
rect 44577 38513 44663 38536
rect 48409 38576 48495 38599
rect 48577 38576 48663 38599
rect 48409 38536 48434 38576
rect 48434 38536 48474 38576
rect 48474 38536 48495 38576
rect 48577 38536 48598 38576
rect 48598 38536 48638 38576
rect 48638 38536 48663 38576
rect 48409 38513 48495 38536
rect 48577 38513 48663 38536
rect 52409 38576 52495 38599
rect 52577 38576 52663 38599
rect 52409 38536 52434 38576
rect 52434 38536 52474 38576
rect 52474 38536 52495 38576
rect 52577 38536 52598 38576
rect 52598 38536 52638 38576
rect 52638 38536 52663 38576
rect 52409 38513 52495 38536
rect 52577 38513 52663 38536
rect 56409 38576 56495 38599
rect 56577 38576 56663 38599
rect 56409 38536 56434 38576
rect 56434 38536 56474 38576
rect 56474 38536 56495 38576
rect 56577 38536 56598 38576
rect 56598 38536 56638 38576
rect 56638 38536 56663 38576
rect 56409 38513 56495 38536
rect 56577 38513 56663 38536
rect 60409 38576 60495 38599
rect 60577 38576 60663 38599
rect 60409 38536 60434 38576
rect 60434 38536 60474 38576
rect 60474 38536 60495 38576
rect 60577 38536 60598 38576
rect 60598 38536 60638 38576
rect 60638 38536 60663 38576
rect 60409 38513 60495 38536
rect 60577 38513 60663 38536
rect 64409 38576 64495 38599
rect 64577 38576 64663 38599
rect 64409 38536 64434 38576
rect 64434 38536 64474 38576
rect 64474 38536 64495 38576
rect 64577 38536 64598 38576
rect 64598 38536 64638 38576
rect 64638 38536 64663 38576
rect 64409 38513 64495 38536
rect 64577 38513 64663 38536
rect 68409 38576 68495 38599
rect 68577 38576 68663 38599
rect 68409 38536 68434 38576
rect 68434 38536 68474 38576
rect 68474 38536 68495 38576
rect 68577 38536 68598 38576
rect 68598 38536 68638 38576
rect 68638 38536 68663 38576
rect 68409 38513 68495 38536
rect 68577 38513 68663 38536
rect 72409 38576 72495 38599
rect 72577 38576 72663 38599
rect 72409 38536 72434 38576
rect 72434 38536 72474 38576
rect 72474 38536 72495 38576
rect 72577 38536 72598 38576
rect 72598 38536 72638 38576
rect 72638 38536 72663 38576
rect 72409 38513 72495 38536
rect 72577 38513 72663 38536
rect 76409 38576 76495 38599
rect 76577 38576 76663 38599
rect 76409 38536 76434 38576
rect 76434 38536 76474 38576
rect 76474 38536 76495 38576
rect 76577 38536 76598 38576
rect 76598 38536 76638 38576
rect 76638 38536 76663 38576
rect 76409 38513 76495 38536
rect 76577 38513 76663 38536
rect 80409 38576 80495 38599
rect 80577 38576 80663 38599
rect 80409 38536 80434 38576
rect 80434 38536 80474 38576
rect 80474 38536 80495 38576
rect 80577 38536 80598 38576
rect 80598 38536 80638 38576
rect 80638 38536 80663 38576
rect 80409 38513 80495 38536
rect 80577 38513 80663 38536
rect 84409 38576 84495 38599
rect 84577 38576 84663 38599
rect 84409 38536 84434 38576
rect 84434 38536 84474 38576
rect 84474 38536 84495 38576
rect 84577 38536 84598 38576
rect 84598 38536 84638 38576
rect 84638 38536 84663 38576
rect 84409 38513 84495 38536
rect 84577 38513 84663 38536
rect 88409 38576 88495 38599
rect 88577 38576 88663 38599
rect 88409 38536 88434 38576
rect 88434 38536 88474 38576
rect 88474 38536 88495 38576
rect 88577 38536 88598 38576
rect 88598 38536 88638 38576
rect 88638 38536 88663 38576
rect 88409 38513 88495 38536
rect 88577 38513 88663 38536
rect 92409 38576 92495 38599
rect 92577 38576 92663 38599
rect 92409 38536 92434 38576
rect 92434 38536 92474 38576
rect 92474 38536 92495 38576
rect 92577 38536 92598 38576
rect 92598 38536 92638 38576
rect 92638 38536 92663 38576
rect 92409 38513 92495 38536
rect 92577 38513 92663 38536
rect 96409 38576 96495 38599
rect 96577 38576 96663 38599
rect 96409 38536 96434 38576
rect 96434 38536 96474 38576
rect 96474 38536 96495 38576
rect 96577 38536 96598 38576
rect 96598 38536 96638 38576
rect 96638 38536 96663 38576
rect 96409 38513 96495 38536
rect 96577 38513 96663 38536
rect 3169 37820 3255 37843
rect 3337 37820 3423 37843
rect 3169 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3255 37820
rect 3337 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3423 37820
rect 3169 37757 3255 37780
rect 3337 37757 3423 37780
rect 7169 37820 7255 37843
rect 7337 37820 7423 37843
rect 7169 37780 7194 37820
rect 7194 37780 7234 37820
rect 7234 37780 7255 37820
rect 7337 37780 7358 37820
rect 7358 37780 7398 37820
rect 7398 37780 7423 37820
rect 7169 37757 7255 37780
rect 7337 37757 7423 37780
rect 11169 37820 11255 37843
rect 11337 37820 11423 37843
rect 11169 37780 11194 37820
rect 11194 37780 11234 37820
rect 11234 37780 11255 37820
rect 11337 37780 11358 37820
rect 11358 37780 11398 37820
rect 11398 37780 11423 37820
rect 11169 37757 11255 37780
rect 11337 37757 11423 37780
rect 15169 37820 15255 37843
rect 15337 37820 15423 37843
rect 15169 37780 15194 37820
rect 15194 37780 15234 37820
rect 15234 37780 15255 37820
rect 15337 37780 15358 37820
rect 15358 37780 15398 37820
rect 15398 37780 15423 37820
rect 15169 37757 15255 37780
rect 15337 37757 15423 37780
rect 19169 37820 19255 37843
rect 19337 37820 19423 37843
rect 19169 37780 19194 37820
rect 19194 37780 19234 37820
rect 19234 37780 19255 37820
rect 19337 37780 19358 37820
rect 19358 37780 19398 37820
rect 19398 37780 19423 37820
rect 19169 37757 19255 37780
rect 19337 37757 19423 37780
rect 23169 37820 23255 37843
rect 23337 37820 23423 37843
rect 23169 37780 23194 37820
rect 23194 37780 23234 37820
rect 23234 37780 23255 37820
rect 23337 37780 23358 37820
rect 23358 37780 23398 37820
rect 23398 37780 23423 37820
rect 23169 37757 23255 37780
rect 23337 37757 23423 37780
rect 27169 37820 27255 37843
rect 27337 37820 27423 37843
rect 27169 37780 27194 37820
rect 27194 37780 27234 37820
rect 27234 37780 27255 37820
rect 27337 37780 27358 37820
rect 27358 37780 27398 37820
rect 27398 37780 27423 37820
rect 27169 37757 27255 37780
rect 27337 37757 27423 37780
rect 31169 37820 31255 37843
rect 31337 37820 31423 37843
rect 31169 37780 31194 37820
rect 31194 37780 31234 37820
rect 31234 37780 31255 37820
rect 31337 37780 31358 37820
rect 31358 37780 31398 37820
rect 31398 37780 31423 37820
rect 31169 37757 31255 37780
rect 31337 37757 31423 37780
rect 35169 37820 35255 37843
rect 35337 37820 35423 37843
rect 35169 37780 35194 37820
rect 35194 37780 35234 37820
rect 35234 37780 35255 37820
rect 35337 37780 35358 37820
rect 35358 37780 35398 37820
rect 35398 37780 35423 37820
rect 35169 37757 35255 37780
rect 35337 37757 35423 37780
rect 39169 37820 39255 37843
rect 39337 37820 39423 37843
rect 39169 37780 39194 37820
rect 39194 37780 39234 37820
rect 39234 37780 39255 37820
rect 39337 37780 39358 37820
rect 39358 37780 39398 37820
rect 39398 37780 39423 37820
rect 39169 37757 39255 37780
rect 39337 37757 39423 37780
rect 43169 37820 43255 37843
rect 43337 37820 43423 37843
rect 43169 37780 43194 37820
rect 43194 37780 43234 37820
rect 43234 37780 43255 37820
rect 43337 37780 43358 37820
rect 43358 37780 43398 37820
rect 43398 37780 43423 37820
rect 43169 37757 43255 37780
rect 43337 37757 43423 37780
rect 47169 37820 47255 37843
rect 47337 37820 47423 37843
rect 47169 37780 47194 37820
rect 47194 37780 47234 37820
rect 47234 37780 47255 37820
rect 47337 37780 47358 37820
rect 47358 37780 47398 37820
rect 47398 37780 47423 37820
rect 47169 37757 47255 37780
rect 47337 37757 47423 37780
rect 51169 37820 51255 37843
rect 51337 37820 51423 37843
rect 51169 37780 51194 37820
rect 51194 37780 51234 37820
rect 51234 37780 51255 37820
rect 51337 37780 51358 37820
rect 51358 37780 51398 37820
rect 51398 37780 51423 37820
rect 51169 37757 51255 37780
rect 51337 37757 51423 37780
rect 55169 37820 55255 37843
rect 55337 37820 55423 37843
rect 55169 37780 55194 37820
rect 55194 37780 55234 37820
rect 55234 37780 55255 37820
rect 55337 37780 55358 37820
rect 55358 37780 55398 37820
rect 55398 37780 55423 37820
rect 55169 37757 55255 37780
rect 55337 37757 55423 37780
rect 59169 37820 59255 37843
rect 59337 37820 59423 37843
rect 59169 37780 59194 37820
rect 59194 37780 59234 37820
rect 59234 37780 59255 37820
rect 59337 37780 59358 37820
rect 59358 37780 59398 37820
rect 59398 37780 59423 37820
rect 59169 37757 59255 37780
rect 59337 37757 59423 37780
rect 63169 37820 63255 37843
rect 63337 37820 63423 37843
rect 63169 37780 63194 37820
rect 63194 37780 63234 37820
rect 63234 37780 63255 37820
rect 63337 37780 63358 37820
rect 63358 37780 63398 37820
rect 63398 37780 63423 37820
rect 63169 37757 63255 37780
rect 63337 37757 63423 37780
rect 67169 37820 67255 37843
rect 67337 37820 67423 37843
rect 67169 37780 67194 37820
rect 67194 37780 67234 37820
rect 67234 37780 67255 37820
rect 67337 37780 67358 37820
rect 67358 37780 67398 37820
rect 67398 37780 67423 37820
rect 67169 37757 67255 37780
rect 67337 37757 67423 37780
rect 71169 37820 71255 37843
rect 71337 37820 71423 37843
rect 71169 37780 71194 37820
rect 71194 37780 71234 37820
rect 71234 37780 71255 37820
rect 71337 37780 71358 37820
rect 71358 37780 71398 37820
rect 71398 37780 71423 37820
rect 71169 37757 71255 37780
rect 71337 37757 71423 37780
rect 75169 37820 75255 37843
rect 75337 37820 75423 37843
rect 75169 37780 75194 37820
rect 75194 37780 75234 37820
rect 75234 37780 75255 37820
rect 75337 37780 75358 37820
rect 75358 37780 75398 37820
rect 75398 37780 75423 37820
rect 75169 37757 75255 37780
rect 75337 37757 75423 37780
rect 79169 37820 79255 37843
rect 79337 37820 79423 37843
rect 79169 37780 79194 37820
rect 79194 37780 79234 37820
rect 79234 37780 79255 37820
rect 79337 37780 79358 37820
rect 79358 37780 79398 37820
rect 79398 37780 79423 37820
rect 79169 37757 79255 37780
rect 79337 37757 79423 37780
rect 83169 37820 83255 37843
rect 83337 37820 83423 37843
rect 83169 37780 83194 37820
rect 83194 37780 83234 37820
rect 83234 37780 83255 37820
rect 83337 37780 83358 37820
rect 83358 37780 83398 37820
rect 83398 37780 83423 37820
rect 83169 37757 83255 37780
rect 83337 37757 83423 37780
rect 87169 37820 87255 37843
rect 87337 37820 87423 37843
rect 87169 37780 87194 37820
rect 87194 37780 87234 37820
rect 87234 37780 87255 37820
rect 87337 37780 87358 37820
rect 87358 37780 87398 37820
rect 87398 37780 87423 37820
rect 87169 37757 87255 37780
rect 87337 37757 87423 37780
rect 91169 37820 91255 37843
rect 91337 37820 91423 37843
rect 91169 37780 91194 37820
rect 91194 37780 91234 37820
rect 91234 37780 91255 37820
rect 91337 37780 91358 37820
rect 91358 37780 91398 37820
rect 91398 37780 91423 37820
rect 91169 37757 91255 37780
rect 91337 37757 91423 37780
rect 95169 37820 95255 37843
rect 95337 37820 95423 37843
rect 95169 37780 95194 37820
rect 95194 37780 95234 37820
rect 95234 37780 95255 37820
rect 95337 37780 95358 37820
rect 95358 37780 95398 37820
rect 95398 37780 95423 37820
rect 95169 37757 95255 37780
rect 95337 37757 95423 37780
rect 99169 37820 99255 37843
rect 99337 37820 99423 37843
rect 99169 37780 99194 37820
rect 99194 37780 99234 37820
rect 99234 37780 99255 37820
rect 99337 37780 99358 37820
rect 99358 37780 99398 37820
rect 99398 37780 99423 37820
rect 99169 37757 99255 37780
rect 99337 37757 99423 37780
rect 4409 37064 4495 37087
rect 4577 37064 4663 37087
rect 4409 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4495 37064
rect 4577 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4663 37064
rect 4409 37001 4495 37024
rect 4577 37001 4663 37024
rect 8409 37064 8495 37087
rect 8577 37064 8663 37087
rect 8409 37024 8434 37064
rect 8434 37024 8474 37064
rect 8474 37024 8495 37064
rect 8577 37024 8598 37064
rect 8598 37024 8638 37064
rect 8638 37024 8663 37064
rect 8409 37001 8495 37024
rect 8577 37001 8663 37024
rect 12409 37064 12495 37087
rect 12577 37064 12663 37087
rect 12409 37024 12434 37064
rect 12434 37024 12474 37064
rect 12474 37024 12495 37064
rect 12577 37024 12598 37064
rect 12598 37024 12638 37064
rect 12638 37024 12663 37064
rect 12409 37001 12495 37024
rect 12577 37001 12663 37024
rect 16409 37064 16495 37087
rect 16577 37064 16663 37087
rect 16409 37024 16434 37064
rect 16434 37024 16474 37064
rect 16474 37024 16495 37064
rect 16577 37024 16598 37064
rect 16598 37024 16638 37064
rect 16638 37024 16663 37064
rect 16409 37001 16495 37024
rect 16577 37001 16663 37024
rect 20409 37064 20495 37087
rect 20577 37064 20663 37087
rect 20409 37024 20434 37064
rect 20434 37024 20474 37064
rect 20474 37024 20495 37064
rect 20577 37024 20598 37064
rect 20598 37024 20638 37064
rect 20638 37024 20663 37064
rect 20409 37001 20495 37024
rect 20577 37001 20663 37024
rect 24409 37064 24495 37087
rect 24577 37064 24663 37087
rect 24409 37024 24434 37064
rect 24434 37024 24474 37064
rect 24474 37024 24495 37064
rect 24577 37024 24598 37064
rect 24598 37024 24638 37064
rect 24638 37024 24663 37064
rect 24409 37001 24495 37024
rect 24577 37001 24663 37024
rect 28409 37064 28495 37087
rect 28577 37064 28663 37087
rect 28409 37024 28434 37064
rect 28434 37024 28474 37064
rect 28474 37024 28495 37064
rect 28577 37024 28598 37064
rect 28598 37024 28638 37064
rect 28638 37024 28663 37064
rect 28409 37001 28495 37024
rect 28577 37001 28663 37024
rect 32409 37064 32495 37087
rect 32577 37064 32663 37087
rect 32409 37024 32434 37064
rect 32434 37024 32474 37064
rect 32474 37024 32495 37064
rect 32577 37024 32598 37064
rect 32598 37024 32638 37064
rect 32638 37024 32663 37064
rect 32409 37001 32495 37024
rect 32577 37001 32663 37024
rect 36409 37064 36495 37087
rect 36577 37064 36663 37087
rect 36409 37024 36434 37064
rect 36434 37024 36474 37064
rect 36474 37024 36495 37064
rect 36577 37024 36598 37064
rect 36598 37024 36638 37064
rect 36638 37024 36663 37064
rect 36409 37001 36495 37024
rect 36577 37001 36663 37024
rect 40409 37064 40495 37087
rect 40577 37064 40663 37087
rect 40409 37024 40434 37064
rect 40434 37024 40474 37064
rect 40474 37024 40495 37064
rect 40577 37024 40598 37064
rect 40598 37024 40638 37064
rect 40638 37024 40663 37064
rect 40409 37001 40495 37024
rect 40577 37001 40663 37024
rect 44409 37064 44495 37087
rect 44577 37064 44663 37087
rect 44409 37024 44434 37064
rect 44434 37024 44474 37064
rect 44474 37024 44495 37064
rect 44577 37024 44598 37064
rect 44598 37024 44638 37064
rect 44638 37024 44663 37064
rect 44409 37001 44495 37024
rect 44577 37001 44663 37024
rect 48409 37064 48495 37087
rect 48577 37064 48663 37087
rect 48409 37024 48434 37064
rect 48434 37024 48474 37064
rect 48474 37024 48495 37064
rect 48577 37024 48598 37064
rect 48598 37024 48638 37064
rect 48638 37024 48663 37064
rect 48409 37001 48495 37024
rect 48577 37001 48663 37024
rect 52409 37064 52495 37087
rect 52577 37064 52663 37087
rect 52409 37024 52434 37064
rect 52434 37024 52474 37064
rect 52474 37024 52495 37064
rect 52577 37024 52598 37064
rect 52598 37024 52638 37064
rect 52638 37024 52663 37064
rect 52409 37001 52495 37024
rect 52577 37001 52663 37024
rect 56409 37064 56495 37087
rect 56577 37064 56663 37087
rect 56409 37024 56434 37064
rect 56434 37024 56474 37064
rect 56474 37024 56495 37064
rect 56577 37024 56598 37064
rect 56598 37024 56638 37064
rect 56638 37024 56663 37064
rect 56409 37001 56495 37024
rect 56577 37001 56663 37024
rect 60409 37064 60495 37087
rect 60577 37064 60663 37087
rect 60409 37024 60434 37064
rect 60434 37024 60474 37064
rect 60474 37024 60495 37064
rect 60577 37024 60598 37064
rect 60598 37024 60638 37064
rect 60638 37024 60663 37064
rect 60409 37001 60495 37024
rect 60577 37001 60663 37024
rect 64409 37064 64495 37087
rect 64577 37064 64663 37087
rect 64409 37024 64434 37064
rect 64434 37024 64474 37064
rect 64474 37024 64495 37064
rect 64577 37024 64598 37064
rect 64598 37024 64638 37064
rect 64638 37024 64663 37064
rect 64409 37001 64495 37024
rect 64577 37001 64663 37024
rect 68409 37064 68495 37087
rect 68577 37064 68663 37087
rect 68409 37024 68434 37064
rect 68434 37024 68474 37064
rect 68474 37024 68495 37064
rect 68577 37024 68598 37064
rect 68598 37024 68638 37064
rect 68638 37024 68663 37064
rect 68409 37001 68495 37024
rect 68577 37001 68663 37024
rect 72409 37064 72495 37087
rect 72577 37064 72663 37087
rect 72409 37024 72434 37064
rect 72434 37024 72474 37064
rect 72474 37024 72495 37064
rect 72577 37024 72598 37064
rect 72598 37024 72638 37064
rect 72638 37024 72663 37064
rect 72409 37001 72495 37024
rect 72577 37001 72663 37024
rect 76409 37064 76495 37087
rect 76577 37064 76663 37087
rect 76409 37024 76434 37064
rect 76434 37024 76474 37064
rect 76474 37024 76495 37064
rect 76577 37024 76598 37064
rect 76598 37024 76638 37064
rect 76638 37024 76663 37064
rect 76409 37001 76495 37024
rect 76577 37001 76663 37024
rect 80409 37064 80495 37087
rect 80577 37064 80663 37087
rect 80409 37024 80434 37064
rect 80434 37024 80474 37064
rect 80474 37024 80495 37064
rect 80577 37024 80598 37064
rect 80598 37024 80638 37064
rect 80638 37024 80663 37064
rect 80409 37001 80495 37024
rect 80577 37001 80663 37024
rect 84409 37064 84495 37087
rect 84577 37064 84663 37087
rect 84409 37024 84434 37064
rect 84434 37024 84474 37064
rect 84474 37024 84495 37064
rect 84577 37024 84598 37064
rect 84598 37024 84638 37064
rect 84638 37024 84663 37064
rect 84409 37001 84495 37024
rect 84577 37001 84663 37024
rect 88409 37064 88495 37087
rect 88577 37064 88663 37087
rect 88409 37024 88434 37064
rect 88434 37024 88474 37064
rect 88474 37024 88495 37064
rect 88577 37024 88598 37064
rect 88598 37024 88638 37064
rect 88638 37024 88663 37064
rect 88409 37001 88495 37024
rect 88577 37001 88663 37024
rect 92409 37064 92495 37087
rect 92577 37064 92663 37087
rect 92409 37024 92434 37064
rect 92434 37024 92474 37064
rect 92474 37024 92495 37064
rect 92577 37024 92598 37064
rect 92598 37024 92638 37064
rect 92638 37024 92663 37064
rect 92409 37001 92495 37024
rect 92577 37001 92663 37024
rect 96409 37064 96495 37087
rect 96577 37064 96663 37087
rect 96409 37024 96434 37064
rect 96434 37024 96474 37064
rect 96474 37024 96495 37064
rect 96577 37024 96598 37064
rect 96598 37024 96638 37064
rect 96638 37024 96663 37064
rect 96409 37001 96495 37024
rect 96577 37001 96663 37024
rect 3169 36308 3255 36331
rect 3337 36308 3423 36331
rect 3169 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3255 36308
rect 3337 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3423 36308
rect 3169 36245 3255 36268
rect 3337 36245 3423 36268
rect 7169 36308 7255 36331
rect 7337 36308 7423 36331
rect 7169 36268 7194 36308
rect 7194 36268 7234 36308
rect 7234 36268 7255 36308
rect 7337 36268 7358 36308
rect 7358 36268 7398 36308
rect 7398 36268 7423 36308
rect 7169 36245 7255 36268
rect 7337 36245 7423 36268
rect 11169 36308 11255 36331
rect 11337 36308 11423 36331
rect 11169 36268 11194 36308
rect 11194 36268 11234 36308
rect 11234 36268 11255 36308
rect 11337 36268 11358 36308
rect 11358 36268 11398 36308
rect 11398 36268 11423 36308
rect 11169 36245 11255 36268
rect 11337 36245 11423 36268
rect 15169 36308 15255 36331
rect 15337 36308 15423 36331
rect 15169 36268 15194 36308
rect 15194 36268 15234 36308
rect 15234 36268 15255 36308
rect 15337 36268 15358 36308
rect 15358 36268 15398 36308
rect 15398 36268 15423 36308
rect 15169 36245 15255 36268
rect 15337 36245 15423 36268
rect 19169 36308 19255 36331
rect 19337 36308 19423 36331
rect 19169 36268 19194 36308
rect 19194 36268 19234 36308
rect 19234 36268 19255 36308
rect 19337 36268 19358 36308
rect 19358 36268 19398 36308
rect 19398 36268 19423 36308
rect 19169 36245 19255 36268
rect 19337 36245 19423 36268
rect 23169 36308 23255 36331
rect 23337 36308 23423 36331
rect 23169 36268 23194 36308
rect 23194 36268 23234 36308
rect 23234 36268 23255 36308
rect 23337 36268 23358 36308
rect 23358 36268 23398 36308
rect 23398 36268 23423 36308
rect 23169 36245 23255 36268
rect 23337 36245 23423 36268
rect 27169 36308 27255 36331
rect 27337 36308 27423 36331
rect 27169 36268 27194 36308
rect 27194 36268 27234 36308
rect 27234 36268 27255 36308
rect 27337 36268 27358 36308
rect 27358 36268 27398 36308
rect 27398 36268 27423 36308
rect 27169 36245 27255 36268
rect 27337 36245 27423 36268
rect 31169 36308 31255 36331
rect 31337 36308 31423 36331
rect 31169 36268 31194 36308
rect 31194 36268 31234 36308
rect 31234 36268 31255 36308
rect 31337 36268 31358 36308
rect 31358 36268 31398 36308
rect 31398 36268 31423 36308
rect 31169 36245 31255 36268
rect 31337 36245 31423 36268
rect 35169 36308 35255 36331
rect 35337 36308 35423 36331
rect 35169 36268 35194 36308
rect 35194 36268 35234 36308
rect 35234 36268 35255 36308
rect 35337 36268 35358 36308
rect 35358 36268 35398 36308
rect 35398 36268 35423 36308
rect 35169 36245 35255 36268
rect 35337 36245 35423 36268
rect 39169 36308 39255 36331
rect 39337 36308 39423 36331
rect 39169 36268 39194 36308
rect 39194 36268 39234 36308
rect 39234 36268 39255 36308
rect 39337 36268 39358 36308
rect 39358 36268 39398 36308
rect 39398 36268 39423 36308
rect 39169 36245 39255 36268
rect 39337 36245 39423 36268
rect 43169 36308 43255 36331
rect 43337 36308 43423 36331
rect 43169 36268 43194 36308
rect 43194 36268 43234 36308
rect 43234 36268 43255 36308
rect 43337 36268 43358 36308
rect 43358 36268 43398 36308
rect 43398 36268 43423 36308
rect 43169 36245 43255 36268
rect 43337 36245 43423 36268
rect 47169 36308 47255 36331
rect 47337 36308 47423 36331
rect 47169 36268 47194 36308
rect 47194 36268 47234 36308
rect 47234 36268 47255 36308
rect 47337 36268 47358 36308
rect 47358 36268 47398 36308
rect 47398 36268 47423 36308
rect 47169 36245 47255 36268
rect 47337 36245 47423 36268
rect 51169 36308 51255 36331
rect 51337 36308 51423 36331
rect 51169 36268 51194 36308
rect 51194 36268 51234 36308
rect 51234 36268 51255 36308
rect 51337 36268 51358 36308
rect 51358 36268 51398 36308
rect 51398 36268 51423 36308
rect 51169 36245 51255 36268
rect 51337 36245 51423 36268
rect 55169 36308 55255 36331
rect 55337 36308 55423 36331
rect 55169 36268 55194 36308
rect 55194 36268 55234 36308
rect 55234 36268 55255 36308
rect 55337 36268 55358 36308
rect 55358 36268 55398 36308
rect 55398 36268 55423 36308
rect 55169 36245 55255 36268
rect 55337 36245 55423 36268
rect 59169 36308 59255 36331
rect 59337 36308 59423 36331
rect 59169 36268 59194 36308
rect 59194 36268 59234 36308
rect 59234 36268 59255 36308
rect 59337 36268 59358 36308
rect 59358 36268 59398 36308
rect 59398 36268 59423 36308
rect 59169 36245 59255 36268
rect 59337 36245 59423 36268
rect 63169 36308 63255 36331
rect 63337 36308 63423 36331
rect 63169 36268 63194 36308
rect 63194 36268 63234 36308
rect 63234 36268 63255 36308
rect 63337 36268 63358 36308
rect 63358 36268 63398 36308
rect 63398 36268 63423 36308
rect 63169 36245 63255 36268
rect 63337 36245 63423 36268
rect 67169 36308 67255 36331
rect 67337 36308 67423 36331
rect 67169 36268 67194 36308
rect 67194 36268 67234 36308
rect 67234 36268 67255 36308
rect 67337 36268 67358 36308
rect 67358 36268 67398 36308
rect 67398 36268 67423 36308
rect 67169 36245 67255 36268
rect 67337 36245 67423 36268
rect 71169 36308 71255 36331
rect 71337 36308 71423 36331
rect 71169 36268 71194 36308
rect 71194 36268 71234 36308
rect 71234 36268 71255 36308
rect 71337 36268 71358 36308
rect 71358 36268 71398 36308
rect 71398 36268 71423 36308
rect 71169 36245 71255 36268
rect 71337 36245 71423 36268
rect 75169 36308 75255 36331
rect 75337 36308 75423 36331
rect 75169 36268 75194 36308
rect 75194 36268 75234 36308
rect 75234 36268 75255 36308
rect 75337 36268 75358 36308
rect 75358 36268 75398 36308
rect 75398 36268 75423 36308
rect 75169 36245 75255 36268
rect 75337 36245 75423 36268
rect 79169 36308 79255 36331
rect 79337 36308 79423 36331
rect 79169 36268 79194 36308
rect 79194 36268 79234 36308
rect 79234 36268 79255 36308
rect 79337 36268 79358 36308
rect 79358 36268 79398 36308
rect 79398 36268 79423 36308
rect 79169 36245 79255 36268
rect 79337 36245 79423 36268
rect 83169 36308 83255 36331
rect 83337 36308 83423 36331
rect 83169 36268 83194 36308
rect 83194 36268 83234 36308
rect 83234 36268 83255 36308
rect 83337 36268 83358 36308
rect 83358 36268 83398 36308
rect 83398 36268 83423 36308
rect 83169 36245 83255 36268
rect 83337 36245 83423 36268
rect 87169 36308 87255 36331
rect 87337 36308 87423 36331
rect 87169 36268 87194 36308
rect 87194 36268 87234 36308
rect 87234 36268 87255 36308
rect 87337 36268 87358 36308
rect 87358 36268 87398 36308
rect 87398 36268 87423 36308
rect 87169 36245 87255 36268
rect 87337 36245 87423 36268
rect 91169 36308 91255 36331
rect 91337 36308 91423 36331
rect 91169 36268 91194 36308
rect 91194 36268 91234 36308
rect 91234 36268 91255 36308
rect 91337 36268 91358 36308
rect 91358 36268 91398 36308
rect 91398 36268 91423 36308
rect 91169 36245 91255 36268
rect 91337 36245 91423 36268
rect 95169 36308 95255 36331
rect 95337 36308 95423 36331
rect 95169 36268 95194 36308
rect 95194 36268 95234 36308
rect 95234 36268 95255 36308
rect 95337 36268 95358 36308
rect 95358 36268 95398 36308
rect 95398 36268 95423 36308
rect 95169 36245 95255 36268
rect 95337 36245 95423 36268
rect 99169 36308 99255 36331
rect 99337 36308 99423 36331
rect 99169 36268 99194 36308
rect 99194 36268 99234 36308
rect 99234 36268 99255 36308
rect 99337 36268 99358 36308
rect 99358 36268 99398 36308
rect 99398 36268 99423 36308
rect 99169 36245 99255 36268
rect 99337 36245 99423 36268
rect 4409 35552 4495 35575
rect 4577 35552 4663 35575
rect 4409 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4495 35552
rect 4577 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4663 35552
rect 4409 35489 4495 35512
rect 4577 35489 4663 35512
rect 8409 35552 8495 35575
rect 8577 35552 8663 35575
rect 8409 35512 8434 35552
rect 8434 35512 8474 35552
rect 8474 35512 8495 35552
rect 8577 35512 8598 35552
rect 8598 35512 8638 35552
rect 8638 35512 8663 35552
rect 8409 35489 8495 35512
rect 8577 35489 8663 35512
rect 12409 35552 12495 35575
rect 12577 35552 12663 35575
rect 12409 35512 12434 35552
rect 12434 35512 12474 35552
rect 12474 35512 12495 35552
rect 12577 35512 12598 35552
rect 12598 35512 12638 35552
rect 12638 35512 12663 35552
rect 12409 35489 12495 35512
rect 12577 35489 12663 35512
rect 16409 35552 16495 35575
rect 16577 35552 16663 35575
rect 16409 35512 16434 35552
rect 16434 35512 16474 35552
rect 16474 35512 16495 35552
rect 16577 35512 16598 35552
rect 16598 35512 16638 35552
rect 16638 35512 16663 35552
rect 16409 35489 16495 35512
rect 16577 35489 16663 35512
rect 20409 35552 20495 35575
rect 20577 35552 20663 35575
rect 20409 35512 20434 35552
rect 20434 35512 20474 35552
rect 20474 35512 20495 35552
rect 20577 35512 20598 35552
rect 20598 35512 20638 35552
rect 20638 35512 20663 35552
rect 20409 35489 20495 35512
rect 20577 35489 20663 35512
rect 24409 35552 24495 35575
rect 24577 35552 24663 35575
rect 24409 35512 24434 35552
rect 24434 35512 24474 35552
rect 24474 35512 24495 35552
rect 24577 35512 24598 35552
rect 24598 35512 24638 35552
rect 24638 35512 24663 35552
rect 24409 35489 24495 35512
rect 24577 35489 24663 35512
rect 28409 35552 28495 35575
rect 28577 35552 28663 35575
rect 28409 35512 28434 35552
rect 28434 35512 28474 35552
rect 28474 35512 28495 35552
rect 28577 35512 28598 35552
rect 28598 35512 28638 35552
rect 28638 35512 28663 35552
rect 28409 35489 28495 35512
rect 28577 35489 28663 35512
rect 32409 35552 32495 35575
rect 32577 35552 32663 35575
rect 32409 35512 32434 35552
rect 32434 35512 32474 35552
rect 32474 35512 32495 35552
rect 32577 35512 32598 35552
rect 32598 35512 32638 35552
rect 32638 35512 32663 35552
rect 32409 35489 32495 35512
rect 32577 35489 32663 35512
rect 36409 35552 36495 35575
rect 36577 35552 36663 35575
rect 36409 35512 36434 35552
rect 36434 35512 36474 35552
rect 36474 35512 36495 35552
rect 36577 35512 36598 35552
rect 36598 35512 36638 35552
rect 36638 35512 36663 35552
rect 36409 35489 36495 35512
rect 36577 35489 36663 35512
rect 40409 35552 40495 35575
rect 40577 35552 40663 35575
rect 40409 35512 40434 35552
rect 40434 35512 40474 35552
rect 40474 35512 40495 35552
rect 40577 35512 40598 35552
rect 40598 35512 40638 35552
rect 40638 35512 40663 35552
rect 40409 35489 40495 35512
rect 40577 35489 40663 35512
rect 44409 35552 44495 35575
rect 44577 35552 44663 35575
rect 44409 35512 44434 35552
rect 44434 35512 44474 35552
rect 44474 35512 44495 35552
rect 44577 35512 44598 35552
rect 44598 35512 44638 35552
rect 44638 35512 44663 35552
rect 44409 35489 44495 35512
rect 44577 35489 44663 35512
rect 48409 35552 48495 35575
rect 48577 35552 48663 35575
rect 48409 35512 48434 35552
rect 48434 35512 48474 35552
rect 48474 35512 48495 35552
rect 48577 35512 48598 35552
rect 48598 35512 48638 35552
rect 48638 35512 48663 35552
rect 48409 35489 48495 35512
rect 48577 35489 48663 35512
rect 52409 35552 52495 35575
rect 52577 35552 52663 35575
rect 52409 35512 52434 35552
rect 52434 35512 52474 35552
rect 52474 35512 52495 35552
rect 52577 35512 52598 35552
rect 52598 35512 52638 35552
rect 52638 35512 52663 35552
rect 52409 35489 52495 35512
rect 52577 35489 52663 35512
rect 56409 35552 56495 35575
rect 56577 35552 56663 35575
rect 56409 35512 56434 35552
rect 56434 35512 56474 35552
rect 56474 35512 56495 35552
rect 56577 35512 56598 35552
rect 56598 35512 56638 35552
rect 56638 35512 56663 35552
rect 56409 35489 56495 35512
rect 56577 35489 56663 35512
rect 60409 35552 60495 35575
rect 60577 35552 60663 35575
rect 60409 35512 60434 35552
rect 60434 35512 60474 35552
rect 60474 35512 60495 35552
rect 60577 35512 60598 35552
rect 60598 35512 60638 35552
rect 60638 35512 60663 35552
rect 60409 35489 60495 35512
rect 60577 35489 60663 35512
rect 64409 35552 64495 35575
rect 64577 35552 64663 35575
rect 64409 35512 64434 35552
rect 64434 35512 64474 35552
rect 64474 35512 64495 35552
rect 64577 35512 64598 35552
rect 64598 35512 64638 35552
rect 64638 35512 64663 35552
rect 64409 35489 64495 35512
rect 64577 35489 64663 35512
rect 68409 35552 68495 35575
rect 68577 35552 68663 35575
rect 68409 35512 68434 35552
rect 68434 35512 68474 35552
rect 68474 35512 68495 35552
rect 68577 35512 68598 35552
rect 68598 35512 68638 35552
rect 68638 35512 68663 35552
rect 68409 35489 68495 35512
rect 68577 35489 68663 35512
rect 72409 35552 72495 35575
rect 72577 35552 72663 35575
rect 72409 35512 72434 35552
rect 72434 35512 72474 35552
rect 72474 35512 72495 35552
rect 72577 35512 72598 35552
rect 72598 35512 72638 35552
rect 72638 35512 72663 35552
rect 72409 35489 72495 35512
rect 72577 35489 72663 35512
rect 76409 35552 76495 35575
rect 76577 35552 76663 35575
rect 76409 35512 76434 35552
rect 76434 35512 76474 35552
rect 76474 35512 76495 35552
rect 76577 35512 76598 35552
rect 76598 35512 76638 35552
rect 76638 35512 76663 35552
rect 76409 35489 76495 35512
rect 76577 35489 76663 35512
rect 80409 35552 80495 35575
rect 80577 35552 80663 35575
rect 80409 35512 80434 35552
rect 80434 35512 80474 35552
rect 80474 35512 80495 35552
rect 80577 35512 80598 35552
rect 80598 35512 80638 35552
rect 80638 35512 80663 35552
rect 80409 35489 80495 35512
rect 80577 35489 80663 35512
rect 84409 35552 84495 35575
rect 84577 35552 84663 35575
rect 84409 35512 84434 35552
rect 84434 35512 84474 35552
rect 84474 35512 84495 35552
rect 84577 35512 84598 35552
rect 84598 35512 84638 35552
rect 84638 35512 84663 35552
rect 84409 35489 84495 35512
rect 84577 35489 84663 35512
rect 88409 35552 88495 35575
rect 88577 35552 88663 35575
rect 88409 35512 88434 35552
rect 88434 35512 88474 35552
rect 88474 35512 88495 35552
rect 88577 35512 88598 35552
rect 88598 35512 88638 35552
rect 88638 35512 88663 35552
rect 88409 35489 88495 35512
rect 88577 35489 88663 35512
rect 92409 35552 92495 35575
rect 92577 35552 92663 35575
rect 92409 35512 92434 35552
rect 92434 35512 92474 35552
rect 92474 35512 92495 35552
rect 92577 35512 92598 35552
rect 92598 35512 92638 35552
rect 92638 35512 92663 35552
rect 92409 35489 92495 35512
rect 92577 35489 92663 35512
rect 96409 35552 96495 35575
rect 96577 35552 96663 35575
rect 96409 35512 96434 35552
rect 96434 35512 96474 35552
rect 96474 35512 96495 35552
rect 96577 35512 96598 35552
rect 96598 35512 96638 35552
rect 96638 35512 96663 35552
rect 96409 35489 96495 35512
rect 96577 35489 96663 35512
rect 86469 34901 86555 34987
rect 3169 34796 3255 34819
rect 3337 34796 3423 34819
rect 3169 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3255 34796
rect 3337 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3423 34796
rect 3169 34733 3255 34756
rect 3337 34733 3423 34756
rect 7169 34796 7255 34819
rect 7337 34796 7423 34819
rect 7169 34756 7194 34796
rect 7194 34756 7234 34796
rect 7234 34756 7255 34796
rect 7337 34756 7358 34796
rect 7358 34756 7398 34796
rect 7398 34756 7423 34796
rect 7169 34733 7255 34756
rect 7337 34733 7423 34756
rect 11169 34796 11255 34819
rect 11337 34796 11423 34819
rect 11169 34756 11194 34796
rect 11194 34756 11234 34796
rect 11234 34756 11255 34796
rect 11337 34756 11358 34796
rect 11358 34756 11398 34796
rect 11398 34756 11423 34796
rect 11169 34733 11255 34756
rect 11337 34733 11423 34756
rect 15169 34796 15255 34819
rect 15337 34796 15423 34819
rect 15169 34756 15194 34796
rect 15194 34756 15234 34796
rect 15234 34756 15255 34796
rect 15337 34756 15358 34796
rect 15358 34756 15398 34796
rect 15398 34756 15423 34796
rect 15169 34733 15255 34756
rect 15337 34733 15423 34756
rect 19169 34796 19255 34819
rect 19337 34796 19423 34819
rect 19169 34756 19194 34796
rect 19194 34756 19234 34796
rect 19234 34756 19255 34796
rect 19337 34756 19358 34796
rect 19358 34756 19398 34796
rect 19398 34756 19423 34796
rect 19169 34733 19255 34756
rect 19337 34733 19423 34756
rect 23169 34796 23255 34819
rect 23337 34796 23423 34819
rect 23169 34756 23194 34796
rect 23194 34756 23234 34796
rect 23234 34756 23255 34796
rect 23337 34756 23358 34796
rect 23358 34756 23398 34796
rect 23398 34756 23423 34796
rect 23169 34733 23255 34756
rect 23337 34733 23423 34756
rect 27169 34796 27255 34819
rect 27337 34796 27423 34819
rect 27169 34756 27194 34796
rect 27194 34756 27234 34796
rect 27234 34756 27255 34796
rect 27337 34756 27358 34796
rect 27358 34756 27398 34796
rect 27398 34756 27423 34796
rect 27169 34733 27255 34756
rect 27337 34733 27423 34756
rect 31169 34796 31255 34819
rect 31337 34796 31423 34819
rect 31169 34756 31194 34796
rect 31194 34756 31234 34796
rect 31234 34756 31255 34796
rect 31337 34756 31358 34796
rect 31358 34756 31398 34796
rect 31398 34756 31423 34796
rect 31169 34733 31255 34756
rect 31337 34733 31423 34756
rect 35169 34796 35255 34819
rect 35337 34796 35423 34819
rect 35169 34756 35194 34796
rect 35194 34756 35234 34796
rect 35234 34756 35255 34796
rect 35337 34756 35358 34796
rect 35358 34756 35398 34796
rect 35398 34756 35423 34796
rect 35169 34733 35255 34756
rect 35337 34733 35423 34756
rect 39169 34796 39255 34819
rect 39337 34796 39423 34819
rect 39169 34756 39194 34796
rect 39194 34756 39234 34796
rect 39234 34756 39255 34796
rect 39337 34756 39358 34796
rect 39358 34756 39398 34796
rect 39398 34756 39423 34796
rect 39169 34733 39255 34756
rect 39337 34733 39423 34756
rect 43169 34796 43255 34819
rect 43337 34796 43423 34819
rect 43169 34756 43194 34796
rect 43194 34756 43234 34796
rect 43234 34756 43255 34796
rect 43337 34756 43358 34796
rect 43358 34756 43398 34796
rect 43398 34756 43423 34796
rect 43169 34733 43255 34756
rect 43337 34733 43423 34756
rect 47169 34796 47255 34819
rect 47337 34796 47423 34819
rect 47169 34756 47194 34796
rect 47194 34756 47234 34796
rect 47234 34756 47255 34796
rect 47337 34756 47358 34796
rect 47358 34756 47398 34796
rect 47398 34756 47423 34796
rect 47169 34733 47255 34756
rect 47337 34733 47423 34756
rect 51169 34796 51255 34819
rect 51337 34796 51423 34819
rect 51169 34756 51194 34796
rect 51194 34756 51234 34796
rect 51234 34756 51255 34796
rect 51337 34756 51358 34796
rect 51358 34756 51398 34796
rect 51398 34756 51423 34796
rect 51169 34733 51255 34756
rect 51337 34733 51423 34756
rect 55169 34796 55255 34819
rect 55337 34796 55423 34819
rect 55169 34756 55194 34796
rect 55194 34756 55234 34796
rect 55234 34756 55255 34796
rect 55337 34756 55358 34796
rect 55358 34756 55398 34796
rect 55398 34756 55423 34796
rect 55169 34733 55255 34756
rect 55337 34733 55423 34756
rect 59169 34796 59255 34819
rect 59337 34796 59423 34819
rect 59169 34756 59194 34796
rect 59194 34756 59234 34796
rect 59234 34756 59255 34796
rect 59337 34756 59358 34796
rect 59358 34756 59398 34796
rect 59398 34756 59423 34796
rect 59169 34733 59255 34756
rect 59337 34733 59423 34756
rect 63169 34796 63255 34819
rect 63337 34796 63423 34819
rect 63169 34756 63194 34796
rect 63194 34756 63234 34796
rect 63234 34756 63255 34796
rect 63337 34756 63358 34796
rect 63358 34756 63398 34796
rect 63398 34756 63423 34796
rect 63169 34733 63255 34756
rect 63337 34733 63423 34756
rect 67169 34796 67255 34819
rect 67337 34796 67423 34819
rect 67169 34756 67194 34796
rect 67194 34756 67234 34796
rect 67234 34756 67255 34796
rect 67337 34756 67358 34796
rect 67358 34756 67398 34796
rect 67398 34756 67423 34796
rect 67169 34733 67255 34756
rect 67337 34733 67423 34756
rect 71169 34796 71255 34819
rect 71337 34796 71423 34819
rect 71169 34756 71194 34796
rect 71194 34756 71234 34796
rect 71234 34756 71255 34796
rect 71337 34756 71358 34796
rect 71358 34756 71398 34796
rect 71398 34756 71423 34796
rect 71169 34733 71255 34756
rect 71337 34733 71423 34756
rect 75169 34796 75255 34819
rect 75337 34796 75423 34819
rect 75169 34756 75194 34796
rect 75194 34756 75234 34796
rect 75234 34756 75255 34796
rect 75337 34756 75358 34796
rect 75358 34756 75398 34796
rect 75398 34756 75423 34796
rect 75169 34733 75255 34756
rect 75337 34733 75423 34756
rect 79169 34796 79255 34819
rect 79337 34796 79423 34819
rect 79169 34756 79194 34796
rect 79194 34756 79234 34796
rect 79234 34756 79255 34796
rect 79337 34756 79358 34796
rect 79358 34756 79398 34796
rect 79398 34756 79423 34796
rect 79169 34733 79255 34756
rect 79337 34733 79423 34756
rect 83169 34796 83255 34819
rect 83337 34796 83423 34819
rect 83169 34756 83194 34796
rect 83194 34756 83234 34796
rect 83234 34756 83255 34796
rect 83337 34756 83358 34796
rect 83358 34756 83398 34796
rect 83398 34756 83423 34796
rect 83169 34733 83255 34756
rect 83337 34733 83423 34756
rect 87169 34796 87255 34819
rect 87337 34796 87423 34819
rect 87169 34756 87194 34796
rect 87194 34756 87234 34796
rect 87234 34756 87255 34796
rect 87337 34756 87358 34796
rect 87358 34756 87398 34796
rect 87398 34756 87423 34796
rect 87169 34733 87255 34756
rect 87337 34733 87423 34756
rect 91169 34796 91255 34819
rect 91337 34796 91423 34819
rect 91169 34756 91194 34796
rect 91194 34756 91234 34796
rect 91234 34756 91255 34796
rect 91337 34756 91358 34796
rect 91358 34756 91398 34796
rect 91398 34756 91423 34796
rect 91169 34733 91255 34756
rect 91337 34733 91423 34756
rect 95169 34796 95255 34819
rect 95337 34796 95423 34819
rect 95169 34756 95194 34796
rect 95194 34756 95234 34796
rect 95234 34756 95255 34796
rect 95337 34756 95358 34796
rect 95358 34756 95398 34796
rect 95398 34756 95423 34796
rect 95169 34733 95255 34756
rect 95337 34733 95423 34756
rect 99169 34796 99255 34819
rect 99337 34796 99423 34819
rect 99169 34756 99194 34796
rect 99194 34756 99234 34796
rect 99234 34756 99255 34796
rect 99337 34756 99358 34796
rect 99358 34756 99398 34796
rect 99398 34756 99423 34796
rect 99169 34733 99255 34756
rect 99337 34733 99423 34756
rect 4409 34040 4495 34063
rect 4577 34040 4663 34063
rect 4409 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4495 34040
rect 4577 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4663 34040
rect 4409 33977 4495 34000
rect 4577 33977 4663 34000
rect 8409 34040 8495 34063
rect 8577 34040 8663 34063
rect 8409 34000 8434 34040
rect 8434 34000 8474 34040
rect 8474 34000 8495 34040
rect 8577 34000 8598 34040
rect 8598 34000 8638 34040
rect 8638 34000 8663 34040
rect 8409 33977 8495 34000
rect 8577 33977 8663 34000
rect 12409 34040 12495 34063
rect 12577 34040 12663 34063
rect 12409 34000 12434 34040
rect 12434 34000 12474 34040
rect 12474 34000 12495 34040
rect 12577 34000 12598 34040
rect 12598 34000 12638 34040
rect 12638 34000 12663 34040
rect 12409 33977 12495 34000
rect 12577 33977 12663 34000
rect 16409 34040 16495 34063
rect 16577 34040 16663 34063
rect 16409 34000 16434 34040
rect 16434 34000 16474 34040
rect 16474 34000 16495 34040
rect 16577 34000 16598 34040
rect 16598 34000 16638 34040
rect 16638 34000 16663 34040
rect 16409 33977 16495 34000
rect 16577 33977 16663 34000
rect 20409 34040 20495 34063
rect 20577 34040 20663 34063
rect 20409 34000 20434 34040
rect 20434 34000 20474 34040
rect 20474 34000 20495 34040
rect 20577 34000 20598 34040
rect 20598 34000 20638 34040
rect 20638 34000 20663 34040
rect 20409 33977 20495 34000
rect 20577 33977 20663 34000
rect 24409 34040 24495 34063
rect 24577 34040 24663 34063
rect 24409 34000 24434 34040
rect 24434 34000 24474 34040
rect 24474 34000 24495 34040
rect 24577 34000 24598 34040
rect 24598 34000 24638 34040
rect 24638 34000 24663 34040
rect 24409 33977 24495 34000
rect 24577 33977 24663 34000
rect 28409 34040 28495 34063
rect 28577 34040 28663 34063
rect 28409 34000 28434 34040
rect 28434 34000 28474 34040
rect 28474 34000 28495 34040
rect 28577 34000 28598 34040
rect 28598 34000 28638 34040
rect 28638 34000 28663 34040
rect 28409 33977 28495 34000
rect 28577 33977 28663 34000
rect 32409 34040 32495 34063
rect 32577 34040 32663 34063
rect 32409 34000 32434 34040
rect 32434 34000 32474 34040
rect 32474 34000 32495 34040
rect 32577 34000 32598 34040
rect 32598 34000 32638 34040
rect 32638 34000 32663 34040
rect 32409 33977 32495 34000
rect 32577 33977 32663 34000
rect 36409 34040 36495 34063
rect 36577 34040 36663 34063
rect 36409 34000 36434 34040
rect 36434 34000 36474 34040
rect 36474 34000 36495 34040
rect 36577 34000 36598 34040
rect 36598 34000 36638 34040
rect 36638 34000 36663 34040
rect 36409 33977 36495 34000
rect 36577 33977 36663 34000
rect 40409 34040 40495 34063
rect 40577 34040 40663 34063
rect 40409 34000 40434 34040
rect 40434 34000 40474 34040
rect 40474 34000 40495 34040
rect 40577 34000 40598 34040
rect 40598 34000 40638 34040
rect 40638 34000 40663 34040
rect 40409 33977 40495 34000
rect 40577 33977 40663 34000
rect 44409 34040 44495 34063
rect 44577 34040 44663 34063
rect 44409 34000 44434 34040
rect 44434 34000 44474 34040
rect 44474 34000 44495 34040
rect 44577 34000 44598 34040
rect 44598 34000 44638 34040
rect 44638 34000 44663 34040
rect 44409 33977 44495 34000
rect 44577 33977 44663 34000
rect 48409 34040 48495 34063
rect 48577 34040 48663 34063
rect 48409 34000 48434 34040
rect 48434 34000 48474 34040
rect 48474 34000 48495 34040
rect 48577 34000 48598 34040
rect 48598 34000 48638 34040
rect 48638 34000 48663 34040
rect 48409 33977 48495 34000
rect 48577 33977 48663 34000
rect 52409 34040 52495 34063
rect 52577 34040 52663 34063
rect 52409 34000 52434 34040
rect 52434 34000 52474 34040
rect 52474 34000 52495 34040
rect 52577 34000 52598 34040
rect 52598 34000 52638 34040
rect 52638 34000 52663 34040
rect 52409 33977 52495 34000
rect 52577 33977 52663 34000
rect 56409 34040 56495 34063
rect 56577 34040 56663 34063
rect 56409 34000 56434 34040
rect 56434 34000 56474 34040
rect 56474 34000 56495 34040
rect 56577 34000 56598 34040
rect 56598 34000 56638 34040
rect 56638 34000 56663 34040
rect 56409 33977 56495 34000
rect 56577 33977 56663 34000
rect 60409 34040 60495 34063
rect 60577 34040 60663 34063
rect 60409 34000 60434 34040
rect 60434 34000 60474 34040
rect 60474 34000 60495 34040
rect 60577 34000 60598 34040
rect 60598 34000 60638 34040
rect 60638 34000 60663 34040
rect 60409 33977 60495 34000
rect 60577 33977 60663 34000
rect 64409 34040 64495 34063
rect 64577 34040 64663 34063
rect 64409 34000 64434 34040
rect 64434 34000 64474 34040
rect 64474 34000 64495 34040
rect 64577 34000 64598 34040
rect 64598 34000 64638 34040
rect 64638 34000 64663 34040
rect 64409 33977 64495 34000
rect 64577 33977 64663 34000
rect 68409 34040 68495 34063
rect 68577 34040 68663 34063
rect 68409 34000 68434 34040
rect 68434 34000 68474 34040
rect 68474 34000 68495 34040
rect 68577 34000 68598 34040
rect 68598 34000 68638 34040
rect 68638 34000 68663 34040
rect 68409 33977 68495 34000
rect 68577 33977 68663 34000
rect 72409 34040 72495 34063
rect 72577 34040 72663 34063
rect 72409 34000 72434 34040
rect 72434 34000 72474 34040
rect 72474 34000 72495 34040
rect 72577 34000 72598 34040
rect 72598 34000 72638 34040
rect 72638 34000 72663 34040
rect 72409 33977 72495 34000
rect 72577 33977 72663 34000
rect 76409 34040 76495 34063
rect 76577 34040 76663 34063
rect 76409 34000 76434 34040
rect 76434 34000 76474 34040
rect 76474 34000 76495 34040
rect 76577 34000 76598 34040
rect 76598 34000 76638 34040
rect 76638 34000 76663 34040
rect 76409 33977 76495 34000
rect 76577 33977 76663 34000
rect 80409 34040 80495 34063
rect 80577 34040 80663 34063
rect 80409 34000 80434 34040
rect 80434 34000 80474 34040
rect 80474 34000 80495 34040
rect 80577 34000 80598 34040
rect 80598 34000 80638 34040
rect 80638 34000 80663 34040
rect 80409 33977 80495 34000
rect 80577 33977 80663 34000
rect 84409 34040 84495 34063
rect 84577 34040 84663 34063
rect 84409 34000 84434 34040
rect 84434 34000 84474 34040
rect 84474 34000 84495 34040
rect 84577 34000 84598 34040
rect 84598 34000 84638 34040
rect 84638 34000 84663 34040
rect 84409 33977 84495 34000
rect 84577 33977 84663 34000
rect 88409 34040 88495 34063
rect 88577 34040 88663 34063
rect 88409 34000 88434 34040
rect 88434 34000 88474 34040
rect 88474 34000 88495 34040
rect 88577 34000 88598 34040
rect 88598 34000 88638 34040
rect 88638 34000 88663 34040
rect 88409 33977 88495 34000
rect 88577 33977 88663 34000
rect 92409 34040 92495 34063
rect 92577 34040 92663 34063
rect 92409 34000 92434 34040
rect 92434 34000 92474 34040
rect 92474 34000 92495 34040
rect 92577 34000 92598 34040
rect 92598 34000 92638 34040
rect 92638 34000 92663 34040
rect 92409 33977 92495 34000
rect 92577 33977 92663 34000
rect 96409 34040 96495 34063
rect 96577 34040 96663 34063
rect 96409 34000 96434 34040
rect 96434 34000 96474 34040
rect 96474 34000 96495 34040
rect 96577 34000 96598 34040
rect 96598 34000 96638 34040
rect 96638 34000 96663 34040
rect 96409 33977 96495 34000
rect 96577 33977 96663 34000
rect 3169 33284 3255 33307
rect 3337 33284 3423 33307
rect 3169 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3255 33284
rect 3337 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3423 33284
rect 3169 33221 3255 33244
rect 3337 33221 3423 33244
rect 7169 33284 7255 33307
rect 7337 33284 7423 33307
rect 7169 33244 7194 33284
rect 7194 33244 7234 33284
rect 7234 33244 7255 33284
rect 7337 33244 7358 33284
rect 7358 33244 7398 33284
rect 7398 33244 7423 33284
rect 7169 33221 7255 33244
rect 7337 33221 7423 33244
rect 11169 33284 11255 33307
rect 11337 33284 11423 33307
rect 11169 33244 11194 33284
rect 11194 33244 11234 33284
rect 11234 33244 11255 33284
rect 11337 33244 11358 33284
rect 11358 33244 11398 33284
rect 11398 33244 11423 33284
rect 11169 33221 11255 33244
rect 11337 33221 11423 33244
rect 15169 33284 15255 33307
rect 15337 33284 15423 33307
rect 15169 33244 15194 33284
rect 15194 33244 15234 33284
rect 15234 33244 15255 33284
rect 15337 33244 15358 33284
rect 15358 33244 15398 33284
rect 15398 33244 15423 33284
rect 15169 33221 15255 33244
rect 15337 33221 15423 33244
rect 19169 33284 19255 33307
rect 19337 33284 19423 33307
rect 19169 33244 19194 33284
rect 19194 33244 19234 33284
rect 19234 33244 19255 33284
rect 19337 33244 19358 33284
rect 19358 33244 19398 33284
rect 19398 33244 19423 33284
rect 19169 33221 19255 33244
rect 19337 33221 19423 33244
rect 23169 33284 23255 33307
rect 23337 33284 23423 33307
rect 23169 33244 23194 33284
rect 23194 33244 23234 33284
rect 23234 33244 23255 33284
rect 23337 33244 23358 33284
rect 23358 33244 23398 33284
rect 23398 33244 23423 33284
rect 23169 33221 23255 33244
rect 23337 33221 23423 33244
rect 27169 33284 27255 33307
rect 27337 33284 27423 33307
rect 27169 33244 27194 33284
rect 27194 33244 27234 33284
rect 27234 33244 27255 33284
rect 27337 33244 27358 33284
rect 27358 33244 27398 33284
rect 27398 33244 27423 33284
rect 27169 33221 27255 33244
rect 27337 33221 27423 33244
rect 31169 33284 31255 33307
rect 31337 33284 31423 33307
rect 31169 33244 31194 33284
rect 31194 33244 31234 33284
rect 31234 33244 31255 33284
rect 31337 33244 31358 33284
rect 31358 33244 31398 33284
rect 31398 33244 31423 33284
rect 31169 33221 31255 33244
rect 31337 33221 31423 33244
rect 35169 33284 35255 33307
rect 35337 33284 35423 33307
rect 35169 33244 35194 33284
rect 35194 33244 35234 33284
rect 35234 33244 35255 33284
rect 35337 33244 35358 33284
rect 35358 33244 35398 33284
rect 35398 33244 35423 33284
rect 35169 33221 35255 33244
rect 35337 33221 35423 33244
rect 39169 33284 39255 33307
rect 39337 33284 39423 33307
rect 39169 33244 39194 33284
rect 39194 33244 39234 33284
rect 39234 33244 39255 33284
rect 39337 33244 39358 33284
rect 39358 33244 39398 33284
rect 39398 33244 39423 33284
rect 39169 33221 39255 33244
rect 39337 33221 39423 33244
rect 43169 33284 43255 33307
rect 43337 33284 43423 33307
rect 43169 33244 43194 33284
rect 43194 33244 43234 33284
rect 43234 33244 43255 33284
rect 43337 33244 43358 33284
rect 43358 33244 43398 33284
rect 43398 33244 43423 33284
rect 43169 33221 43255 33244
rect 43337 33221 43423 33244
rect 47169 33284 47255 33307
rect 47337 33284 47423 33307
rect 47169 33244 47194 33284
rect 47194 33244 47234 33284
rect 47234 33244 47255 33284
rect 47337 33244 47358 33284
rect 47358 33244 47398 33284
rect 47398 33244 47423 33284
rect 47169 33221 47255 33244
rect 47337 33221 47423 33244
rect 51169 33284 51255 33307
rect 51337 33284 51423 33307
rect 51169 33244 51194 33284
rect 51194 33244 51234 33284
rect 51234 33244 51255 33284
rect 51337 33244 51358 33284
rect 51358 33244 51398 33284
rect 51398 33244 51423 33284
rect 51169 33221 51255 33244
rect 51337 33221 51423 33244
rect 55169 33284 55255 33307
rect 55337 33284 55423 33307
rect 55169 33244 55194 33284
rect 55194 33244 55234 33284
rect 55234 33244 55255 33284
rect 55337 33244 55358 33284
rect 55358 33244 55398 33284
rect 55398 33244 55423 33284
rect 55169 33221 55255 33244
rect 55337 33221 55423 33244
rect 59169 33284 59255 33307
rect 59337 33284 59423 33307
rect 59169 33244 59194 33284
rect 59194 33244 59234 33284
rect 59234 33244 59255 33284
rect 59337 33244 59358 33284
rect 59358 33244 59398 33284
rect 59398 33244 59423 33284
rect 59169 33221 59255 33244
rect 59337 33221 59423 33244
rect 63169 33284 63255 33307
rect 63337 33284 63423 33307
rect 63169 33244 63194 33284
rect 63194 33244 63234 33284
rect 63234 33244 63255 33284
rect 63337 33244 63358 33284
rect 63358 33244 63398 33284
rect 63398 33244 63423 33284
rect 63169 33221 63255 33244
rect 63337 33221 63423 33244
rect 67169 33284 67255 33307
rect 67337 33284 67423 33307
rect 67169 33244 67194 33284
rect 67194 33244 67234 33284
rect 67234 33244 67255 33284
rect 67337 33244 67358 33284
rect 67358 33244 67398 33284
rect 67398 33244 67423 33284
rect 67169 33221 67255 33244
rect 67337 33221 67423 33244
rect 4409 32528 4495 32551
rect 4577 32528 4663 32551
rect 4409 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4495 32528
rect 4577 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4663 32528
rect 4409 32465 4495 32488
rect 4577 32465 4663 32488
rect 8409 32528 8495 32551
rect 8577 32528 8663 32551
rect 8409 32488 8434 32528
rect 8434 32488 8474 32528
rect 8474 32488 8495 32528
rect 8577 32488 8598 32528
rect 8598 32488 8638 32528
rect 8638 32488 8663 32528
rect 8409 32465 8495 32488
rect 8577 32465 8663 32488
rect 12409 32528 12495 32551
rect 12577 32528 12663 32551
rect 12409 32488 12434 32528
rect 12434 32488 12474 32528
rect 12474 32488 12495 32528
rect 12577 32488 12598 32528
rect 12598 32488 12638 32528
rect 12638 32488 12663 32528
rect 12409 32465 12495 32488
rect 12577 32465 12663 32488
rect 16409 32528 16495 32551
rect 16577 32528 16663 32551
rect 16409 32488 16434 32528
rect 16434 32488 16474 32528
rect 16474 32488 16495 32528
rect 16577 32488 16598 32528
rect 16598 32488 16638 32528
rect 16638 32488 16663 32528
rect 16409 32465 16495 32488
rect 16577 32465 16663 32488
rect 20409 32528 20495 32551
rect 20577 32528 20663 32551
rect 20409 32488 20434 32528
rect 20434 32488 20474 32528
rect 20474 32488 20495 32528
rect 20577 32488 20598 32528
rect 20598 32488 20638 32528
rect 20638 32488 20663 32528
rect 20409 32465 20495 32488
rect 20577 32465 20663 32488
rect 24409 32528 24495 32551
rect 24577 32528 24663 32551
rect 24409 32488 24434 32528
rect 24434 32488 24474 32528
rect 24474 32488 24495 32528
rect 24577 32488 24598 32528
rect 24598 32488 24638 32528
rect 24638 32488 24663 32528
rect 24409 32465 24495 32488
rect 24577 32465 24663 32488
rect 28409 32528 28495 32551
rect 28577 32528 28663 32551
rect 28409 32488 28434 32528
rect 28434 32488 28474 32528
rect 28474 32488 28495 32528
rect 28577 32488 28598 32528
rect 28598 32488 28638 32528
rect 28638 32488 28663 32528
rect 28409 32465 28495 32488
rect 28577 32465 28663 32488
rect 32409 32528 32495 32551
rect 32577 32528 32663 32551
rect 32409 32488 32434 32528
rect 32434 32488 32474 32528
rect 32474 32488 32495 32528
rect 32577 32488 32598 32528
rect 32598 32488 32638 32528
rect 32638 32488 32663 32528
rect 32409 32465 32495 32488
rect 32577 32465 32663 32488
rect 36409 32528 36495 32551
rect 36577 32528 36663 32551
rect 36409 32488 36434 32528
rect 36434 32488 36474 32528
rect 36474 32488 36495 32528
rect 36577 32488 36598 32528
rect 36598 32488 36638 32528
rect 36638 32488 36663 32528
rect 36409 32465 36495 32488
rect 36577 32465 36663 32488
rect 40409 32528 40495 32551
rect 40577 32528 40663 32551
rect 40409 32488 40434 32528
rect 40434 32488 40474 32528
rect 40474 32488 40495 32528
rect 40577 32488 40598 32528
rect 40598 32488 40638 32528
rect 40638 32488 40663 32528
rect 40409 32465 40495 32488
rect 40577 32465 40663 32488
rect 44409 32528 44495 32551
rect 44577 32528 44663 32551
rect 44409 32488 44434 32528
rect 44434 32488 44474 32528
rect 44474 32488 44495 32528
rect 44577 32488 44598 32528
rect 44598 32488 44638 32528
rect 44638 32488 44663 32528
rect 44409 32465 44495 32488
rect 44577 32465 44663 32488
rect 48409 32528 48495 32551
rect 48577 32528 48663 32551
rect 48409 32488 48434 32528
rect 48434 32488 48474 32528
rect 48474 32488 48495 32528
rect 48577 32488 48598 32528
rect 48598 32488 48638 32528
rect 48638 32488 48663 32528
rect 48409 32465 48495 32488
rect 48577 32465 48663 32488
rect 52409 32528 52495 32551
rect 52577 32528 52663 32551
rect 52409 32488 52434 32528
rect 52434 32488 52474 32528
rect 52474 32488 52495 32528
rect 52577 32488 52598 32528
rect 52598 32488 52638 32528
rect 52638 32488 52663 32528
rect 52409 32465 52495 32488
rect 52577 32465 52663 32488
rect 56409 32528 56495 32551
rect 56577 32528 56663 32551
rect 56409 32488 56434 32528
rect 56434 32488 56474 32528
rect 56474 32488 56495 32528
rect 56577 32488 56598 32528
rect 56598 32488 56638 32528
rect 56638 32488 56663 32528
rect 56409 32465 56495 32488
rect 56577 32465 56663 32488
rect 60409 32528 60495 32551
rect 60577 32528 60663 32551
rect 60409 32488 60434 32528
rect 60434 32488 60474 32528
rect 60474 32488 60495 32528
rect 60577 32488 60598 32528
rect 60598 32488 60638 32528
rect 60638 32488 60663 32528
rect 60409 32465 60495 32488
rect 60577 32465 60663 32488
rect 64409 32528 64495 32551
rect 64577 32528 64663 32551
rect 64409 32488 64434 32528
rect 64434 32488 64474 32528
rect 64474 32488 64495 32528
rect 64577 32488 64598 32528
rect 64598 32488 64638 32528
rect 64638 32488 64663 32528
rect 64409 32465 64495 32488
rect 64577 32465 64663 32488
rect 68409 32528 68495 32551
rect 68577 32528 68663 32551
rect 68409 32488 68434 32528
rect 68434 32488 68474 32528
rect 68474 32488 68495 32528
rect 68577 32488 68598 32528
rect 68598 32488 68638 32528
rect 68638 32488 68663 32528
rect 68409 32465 68495 32488
rect 68577 32465 68663 32488
rect 3169 31772 3255 31795
rect 3337 31772 3423 31795
rect 3169 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3255 31772
rect 3337 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3423 31772
rect 3169 31709 3255 31732
rect 3337 31709 3423 31732
rect 7169 31772 7255 31795
rect 7337 31772 7423 31795
rect 7169 31732 7194 31772
rect 7194 31732 7234 31772
rect 7234 31732 7255 31772
rect 7337 31732 7358 31772
rect 7358 31732 7398 31772
rect 7398 31732 7423 31772
rect 7169 31709 7255 31732
rect 7337 31709 7423 31732
rect 11169 31772 11255 31795
rect 11337 31772 11423 31795
rect 11169 31732 11194 31772
rect 11194 31732 11234 31772
rect 11234 31732 11255 31772
rect 11337 31732 11358 31772
rect 11358 31732 11398 31772
rect 11398 31732 11423 31772
rect 11169 31709 11255 31732
rect 11337 31709 11423 31732
rect 15169 31772 15255 31795
rect 15337 31772 15423 31795
rect 15169 31732 15194 31772
rect 15194 31732 15234 31772
rect 15234 31732 15255 31772
rect 15337 31732 15358 31772
rect 15358 31732 15398 31772
rect 15398 31732 15423 31772
rect 15169 31709 15255 31732
rect 15337 31709 15423 31732
rect 19169 31772 19255 31795
rect 19337 31772 19423 31795
rect 19169 31732 19194 31772
rect 19194 31732 19234 31772
rect 19234 31732 19255 31772
rect 19337 31732 19358 31772
rect 19358 31732 19398 31772
rect 19398 31732 19423 31772
rect 19169 31709 19255 31732
rect 19337 31709 19423 31732
rect 23169 31772 23255 31795
rect 23337 31772 23423 31795
rect 23169 31732 23194 31772
rect 23194 31732 23234 31772
rect 23234 31732 23255 31772
rect 23337 31732 23358 31772
rect 23358 31732 23398 31772
rect 23398 31732 23423 31772
rect 23169 31709 23255 31732
rect 23337 31709 23423 31732
rect 27169 31772 27255 31795
rect 27337 31772 27423 31795
rect 27169 31732 27194 31772
rect 27194 31732 27234 31772
rect 27234 31732 27255 31772
rect 27337 31732 27358 31772
rect 27358 31732 27398 31772
rect 27398 31732 27423 31772
rect 27169 31709 27255 31732
rect 27337 31709 27423 31732
rect 31169 31772 31255 31795
rect 31337 31772 31423 31795
rect 31169 31732 31194 31772
rect 31194 31732 31234 31772
rect 31234 31732 31255 31772
rect 31337 31732 31358 31772
rect 31358 31732 31398 31772
rect 31398 31732 31423 31772
rect 31169 31709 31255 31732
rect 31337 31709 31423 31732
rect 35169 31772 35255 31795
rect 35337 31772 35423 31795
rect 35169 31732 35194 31772
rect 35194 31732 35234 31772
rect 35234 31732 35255 31772
rect 35337 31732 35358 31772
rect 35358 31732 35398 31772
rect 35398 31732 35423 31772
rect 35169 31709 35255 31732
rect 35337 31709 35423 31732
rect 39169 31772 39255 31795
rect 39337 31772 39423 31795
rect 39169 31732 39194 31772
rect 39194 31732 39234 31772
rect 39234 31732 39255 31772
rect 39337 31732 39358 31772
rect 39358 31732 39398 31772
rect 39398 31732 39423 31772
rect 39169 31709 39255 31732
rect 39337 31709 39423 31732
rect 43169 31772 43255 31795
rect 43337 31772 43423 31795
rect 43169 31732 43194 31772
rect 43194 31732 43234 31772
rect 43234 31732 43255 31772
rect 43337 31732 43358 31772
rect 43358 31732 43398 31772
rect 43398 31732 43423 31772
rect 43169 31709 43255 31732
rect 43337 31709 43423 31732
rect 47169 31772 47255 31795
rect 47337 31772 47423 31795
rect 47169 31732 47194 31772
rect 47194 31732 47234 31772
rect 47234 31732 47255 31772
rect 47337 31732 47358 31772
rect 47358 31732 47398 31772
rect 47398 31732 47423 31772
rect 47169 31709 47255 31732
rect 47337 31709 47423 31732
rect 51169 31772 51255 31795
rect 51337 31772 51423 31795
rect 51169 31732 51194 31772
rect 51194 31732 51234 31772
rect 51234 31732 51255 31772
rect 51337 31732 51358 31772
rect 51358 31732 51398 31772
rect 51398 31732 51423 31772
rect 51169 31709 51255 31732
rect 51337 31709 51423 31732
rect 55169 31772 55255 31795
rect 55337 31772 55423 31795
rect 55169 31732 55194 31772
rect 55194 31732 55234 31772
rect 55234 31732 55255 31772
rect 55337 31732 55358 31772
rect 55358 31732 55398 31772
rect 55398 31732 55423 31772
rect 55169 31709 55255 31732
rect 55337 31709 55423 31732
rect 59169 31772 59255 31795
rect 59337 31772 59423 31795
rect 59169 31732 59194 31772
rect 59194 31732 59234 31772
rect 59234 31732 59255 31772
rect 59337 31732 59358 31772
rect 59358 31732 59398 31772
rect 59398 31732 59423 31772
rect 59169 31709 59255 31732
rect 59337 31709 59423 31732
rect 63169 31772 63255 31795
rect 63337 31772 63423 31795
rect 63169 31732 63194 31772
rect 63194 31732 63234 31772
rect 63234 31732 63255 31772
rect 63337 31732 63358 31772
rect 63358 31732 63398 31772
rect 63398 31732 63423 31772
rect 63169 31709 63255 31732
rect 63337 31709 63423 31732
rect 67169 31772 67255 31795
rect 67337 31772 67423 31795
rect 67169 31732 67194 31772
rect 67194 31732 67234 31772
rect 67234 31732 67255 31772
rect 67337 31732 67358 31772
rect 67358 31732 67398 31772
rect 67398 31732 67423 31772
rect 67169 31709 67255 31732
rect 67337 31709 67423 31732
rect 4409 31016 4495 31039
rect 4577 31016 4663 31039
rect 4409 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4495 31016
rect 4577 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4663 31016
rect 4409 30953 4495 30976
rect 4577 30953 4663 30976
rect 8409 31016 8495 31039
rect 8577 31016 8663 31039
rect 8409 30976 8434 31016
rect 8434 30976 8474 31016
rect 8474 30976 8495 31016
rect 8577 30976 8598 31016
rect 8598 30976 8638 31016
rect 8638 30976 8663 31016
rect 8409 30953 8495 30976
rect 8577 30953 8663 30976
rect 12409 31016 12495 31039
rect 12577 31016 12663 31039
rect 12409 30976 12434 31016
rect 12434 30976 12474 31016
rect 12474 30976 12495 31016
rect 12577 30976 12598 31016
rect 12598 30976 12638 31016
rect 12638 30976 12663 31016
rect 12409 30953 12495 30976
rect 12577 30953 12663 30976
rect 16409 31016 16495 31039
rect 16577 31016 16663 31039
rect 16409 30976 16434 31016
rect 16434 30976 16474 31016
rect 16474 30976 16495 31016
rect 16577 30976 16598 31016
rect 16598 30976 16638 31016
rect 16638 30976 16663 31016
rect 16409 30953 16495 30976
rect 16577 30953 16663 30976
rect 20409 31016 20495 31039
rect 20577 31016 20663 31039
rect 20409 30976 20434 31016
rect 20434 30976 20474 31016
rect 20474 30976 20495 31016
rect 20577 30976 20598 31016
rect 20598 30976 20638 31016
rect 20638 30976 20663 31016
rect 20409 30953 20495 30976
rect 20577 30953 20663 30976
rect 24409 31016 24495 31039
rect 24577 31016 24663 31039
rect 24409 30976 24434 31016
rect 24434 30976 24474 31016
rect 24474 30976 24495 31016
rect 24577 30976 24598 31016
rect 24598 30976 24638 31016
rect 24638 30976 24663 31016
rect 24409 30953 24495 30976
rect 24577 30953 24663 30976
rect 28409 31016 28495 31039
rect 28577 31016 28663 31039
rect 28409 30976 28434 31016
rect 28434 30976 28474 31016
rect 28474 30976 28495 31016
rect 28577 30976 28598 31016
rect 28598 30976 28638 31016
rect 28638 30976 28663 31016
rect 28409 30953 28495 30976
rect 28577 30953 28663 30976
rect 32409 31016 32495 31039
rect 32577 31016 32663 31039
rect 32409 30976 32434 31016
rect 32434 30976 32474 31016
rect 32474 30976 32495 31016
rect 32577 30976 32598 31016
rect 32598 30976 32638 31016
rect 32638 30976 32663 31016
rect 32409 30953 32495 30976
rect 32577 30953 32663 30976
rect 36409 31016 36495 31039
rect 36577 31016 36663 31039
rect 36409 30976 36434 31016
rect 36434 30976 36474 31016
rect 36474 30976 36495 31016
rect 36577 30976 36598 31016
rect 36598 30976 36638 31016
rect 36638 30976 36663 31016
rect 36409 30953 36495 30976
rect 36577 30953 36663 30976
rect 40409 31016 40495 31039
rect 40577 31016 40663 31039
rect 40409 30976 40434 31016
rect 40434 30976 40474 31016
rect 40474 30976 40495 31016
rect 40577 30976 40598 31016
rect 40598 30976 40638 31016
rect 40638 30976 40663 31016
rect 40409 30953 40495 30976
rect 40577 30953 40663 30976
rect 44409 31016 44495 31039
rect 44577 31016 44663 31039
rect 44409 30976 44434 31016
rect 44434 30976 44474 31016
rect 44474 30976 44495 31016
rect 44577 30976 44598 31016
rect 44598 30976 44638 31016
rect 44638 30976 44663 31016
rect 44409 30953 44495 30976
rect 44577 30953 44663 30976
rect 48409 31016 48495 31039
rect 48577 31016 48663 31039
rect 48409 30976 48434 31016
rect 48434 30976 48474 31016
rect 48474 30976 48495 31016
rect 48577 30976 48598 31016
rect 48598 30976 48638 31016
rect 48638 30976 48663 31016
rect 48409 30953 48495 30976
rect 48577 30953 48663 30976
rect 52409 31016 52495 31039
rect 52577 31016 52663 31039
rect 52409 30976 52434 31016
rect 52434 30976 52474 31016
rect 52474 30976 52495 31016
rect 52577 30976 52598 31016
rect 52598 30976 52638 31016
rect 52638 30976 52663 31016
rect 52409 30953 52495 30976
rect 52577 30953 52663 30976
rect 56409 31016 56495 31039
rect 56577 31016 56663 31039
rect 56409 30976 56434 31016
rect 56434 30976 56474 31016
rect 56474 30976 56495 31016
rect 56577 30976 56598 31016
rect 56598 30976 56638 31016
rect 56638 30976 56663 31016
rect 56409 30953 56495 30976
rect 56577 30953 56663 30976
rect 60409 31016 60495 31039
rect 60577 31016 60663 31039
rect 60409 30976 60434 31016
rect 60434 30976 60474 31016
rect 60474 30976 60495 31016
rect 60577 30976 60598 31016
rect 60598 30976 60638 31016
rect 60638 30976 60663 31016
rect 60409 30953 60495 30976
rect 60577 30953 60663 30976
rect 64409 31016 64495 31039
rect 64577 31016 64663 31039
rect 64409 30976 64434 31016
rect 64434 30976 64474 31016
rect 64474 30976 64495 31016
rect 64577 30976 64598 31016
rect 64598 30976 64638 31016
rect 64638 30976 64663 31016
rect 64409 30953 64495 30976
rect 64577 30953 64663 30976
rect 68409 31016 68495 31039
rect 68577 31016 68663 31039
rect 68409 30976 68434 31016
rect 68434 30976 68474 31016
rect 68474 30976 68495 31016
rect 68577 30976 68598 31016
rect 68598 30976 68638 31016
rect 68638 30976 68663 31016
rect 68409 30953 68495 30976
rect 68577 30953 68663 30976
rect 72409 31036 72495 31122
rect 72577 31036 72663 31122
rect 72409 30868 72495 30954
rect 72577 30868 72663 30954
rect 72409 30700 72495 30786
rect 72577 30700 72663 30786
rect 72409 30532 72495 30618
rect 72577 30532 72663 30618
rect 72409 30364 72495 30450
rect 72577 30364 72663 30450
rect 3169 30260 3255 30283
rect 3337 30260 3423 30283
rect 3169 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3255 30260
rect 3337 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3423 30260
rect 3169 30197 3255 30220
rect 3337 30197 3423 30220
rect 7169 30260 7255 30283
rect 7337 30260 7423 30283
rect 7169 30220 7194 30260
rect 7194 30220 7234 30260
rect 7234 30220 7255 30260
rect 7337 30220 7358 30260
rect 7358 30220 7398 30260
rect 7398 30220 7423 30260
rect 7169 30197 7255 30220
rect 7337 30197 7423 30220
rect 11169 30260 11255 30283
rect 11337 30260 11423 30283
rect 11169 30220 11194 30260
rect 11194 30220 11234 30260
rect 11234 30220 11255 30260
rect 11337 30220 11358 30260
rect 11358 30220 11398 30260
rect 11398 30220 11423 30260
rect 11169 30197 11255 30220
rect 11337 30197 11423 30220
rect 15169 30260 15255 30283
rect 15337 30260 15423 30283
rect 15169 30220 15194 30260
rect 15194 30220 15234 30260
rect 15234 30220 15255 30260
rect 15337 30220 15358 30260
rect 15358 30220 15398 30260
rect 15398 30220 15423 30260
rect 15169 30197 15255 30220
rect 15337 30197 15423 30220
rect 19169 30260 19255 30283
rect 19337 30260 19423 30283
rect 19169 30220 19194 30260
rect 19194 30220 19234 30260
rect 19234 30220 19255 30260
rect 19337 30220 19358 30260
rect 19358 30220 19398 30260
rect 19398 30220 19423 30260
rect 19169 30197 19255 30220
rect 19337 30197 19423 30220
rect 23169 30260 23255 30283
rect 23337 30260 23423 30283
rect 23169 30220 23194 30260
rect 23194 30220 23234 30260
rect 23234 30220 23255 30260
rect 23337 30220 23358 30260
rect 23358 30220 23398 30260
rect 23398 30220 23423 30260
rect 23169 30197 23255 30220
rect 23337 30197 23423 30220
rect 27169 30260 27255 30283
rect 27337 30260 27423 30283
rect 27169 30220 27194 30260
rect 27194 30220 27234 30260
rect 27234 30220 27255 30260
rect 27337 30220 27358 30260
rect 27358 30220 27398 30260
rect 27398 30220 27423 30260
rect 27169 30197 27255 30220
rect 27337 30197 27423 30220
rect 31169 30260 31255 30283
rect 31337 30260 31423 30283
rect 31169 30220 31194 30260
rect 31194 30220 31234 30260
rect 31234 30220 31255 30260
rect 31337 30220 31358 30260
rect 31358 30220 31398 30260
rect 31398 30220 31423 30260
rect 31169 30197 31255 30220
rect 31337 30197 31423 30220
rect 35169 30260 35255 30283
rect 35337 30260 35423 30283
rect 35169 30220 35194 30260
rect 35194 30220 35234 30260
rect 35234 30220 35255 30260
rect 35337 30220 35358 30260
rect 35358 30220 35398 30260
rect 35398 30220 35423 30260
rect 35169 30197 35255 30220
rect 35337 30197 35423 30220
rect 39169 30260 39255 30283
rect 39337 30260 39423 30283
rect 39169 30220 39194 30260
rect 39194 30220 39234 30260
rect 39234 30220 39255 30260
rect 39337 30220 39358 30260
rect 39358 30220 39398 30260
rect 39398 30220 39423 30260
rect 39169 30197 39255 30220
rect 39337 30197 39423 30220
rect 43169 30260 43255 30283
rect 43337 30260 43423 30283
rect 43169 30220 43194 30260
rect 43194 30220 43234 30260
rect 43234 30220 43255 30260
rect 43337 30220 43358 30260
rect 43358 30220 43398 30260
rect 43398 30220 43423 30260
rect 43169 30197 43255 30220
rect 43337 30197 43423 30220
rect 47169 30260 47255 30283
rect 47337 30260 47423 30283
rect 47169 30220 47194 30260
rect 47194 30220 47234 30260
rect 47234 30220 47255 30260
rect 47337 30220 47358 30260
rect 47358 30220 47398 30260
rect 47398 30220 47423 30260
rect 47169 30197 47255 30220
rect 47337 30197 47423 30220
rect 51169 30260 51255 30283
rect 51337 30260 51423 30283
rect 51169 30220 51194 30260
rect 51194 30220 51234 30260
rect 51234 30220 51255 30260
rect 51337 30220 51358 30260
rect 51358 30220 51398 30260
rect 51398 30220 51423 30260
rect 51169 30197 51255 30220
rect 51337 30197 51423 30220
rect 55169 30260 55255 30283
rect 55337 30260 55423 30283
rect 55169 30220 55194 30260
rect 55194 30220 55234 30260
rect 55234 30220 55255 30260
rect 55337 30220 55358 30260
rect 55358 30220 55398 30260
rect 55398 30220 55423 30260
rect 55169 30197 55255 30220
rect 55337 30197 55423 30220
rect 59169 30260 59255 30283
rect 59337 30260 59423 30283
rect 59169 30220 59194 30260
rect 59194 30220 59234 30260
rect 59234 30220 59255 30260
rect 59337 30220 59358 30260
rect 59358 30220 59398 30260
rect 59398 30220 59423 30260
rect 59169 30197 59255 30220
rect 59337 30197 59423 30220
rect 63169 30260 63255 30283
rect 63337 30260 63423 30283
rect 63169 30220 63194 30260
rect 63194 30220 63234 30260
rect 63234 30220 63255 30260
rect 63337 30220 63358 30260
rect 63358 30220 63398 30260
rect 63398 30220 63423 30260
rect 63169 30197 63255 30220
rect 63337 30197 63423 30220
rect 67169 30260 67255 30283
rect 67337 30260 67423 30283
rect 67169 30220 67194 30260
rect 67194 30220 67234 30260
rect 67234 30220 67255 30260
rect 67337 30220 67358 30260
rect 67358 30220 67398 30260
rect 67398 30220 67423 30260
rect 67169 30197 67255 30220
rect 67337 30197 67423 30220
rect 72409 30196 72495 30282
rect 72577 30196 72663 30282
rect 72409 30028 72495 30114
rect 72577 30028 72663 30114
rect 72409 29860 72495 29946
rect 72577 29860 72663 29946
rect 72409 29692 72495 29778
rect 72577 29692 72663 29778
rect 4409 29504 4495 29527
rect 4577 29504 4663 29527
rect 4409 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4495 29504
rect 4577 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4663 29504
rect 4409 29441 4495 29464
rect 4577 29441 4663 29464
rect 8409 29504 8495 29527
rect 8577 29504 8663 29527
rect 8409 29464 8434 29504
rect 8434 29464 8474 29504
rect 8474 29464 8495 29504
rect 8577 29464 8598 29504
rect 8598 29464 8638 29504
rect 8638 29464 8663 29504
rect 8409 29441 8495 29464
rect 8577 29441 8663 29464
rect 12409 29504 12495 29527
rect 12577 29504 12663 29527
rect 12409 29464 12434 29504
rect 12434 29464 12474 29504
rect 12474 29464 12495 29504
rect 12577 29464 12598 29504
rect 12598 29464 12638 29504
rect 12638 29464 12663 29504
rect 12409 29441 12495 29464
rect 12577 29441 12663 29464
rect 16409 29504 16495 29527
rect 16577 29504 16663 29527
rect 16409 29464 16434 29504
rect 16434 29464 16474 29504
rect 16474 29464 16495 29504
rect 16577 29464 16598 29504
rect 16598 29464 16638 29504
rect 16638 29464 16663 29504
rect 16409 29441 16495 29464
rect 16577 29441 16663 29464
rect 20409 29504 20495 29527
rect 20577 29504 20663 29527
rect 20409 29464 20434 29504
rect 20434 29464 20474 29504
rect 20474 29464 20495 29504
rect 20577 29464 20598 29504
rect 20598 29464 20638 29504
rect 20638 29464 20663 29504
rect 20409 29441 20495 29464
rect 20577 29441 20663 29464
rect 24409 29504 24495 29527
rect 24577 29504 24663 29527
rect 24409 29464 24434 29504
rect 24434 29464 24474 29504
rect 24474 29464 24495 29504
rect 24577 29464 24598 29504
rect 24598 29464 24638 29504
rect 24638 29464 24663 29504
rect 24409 29441 24495 29464
rect 24577 29441 24663 29464
rect 28409 29504 28495 29527
rect 28577 29504 28663 29527
rect 28409 29464 28434 29504
rect 28434 29464 28474 29504
rect 28474 29464 28495 29504
rect 28577 29464 28598 29504
rect 28598 29464 28638 29504
rect 28638 29464 28663 29504
rect 28409 29441 28495 29464
rect 28577 29441 28663 29464
rect 32409 29504 32495 29527
rect 32577 29504 32663 29527
rect 32409 29464 32434 29504
rect 32434 29464 32474 29504
rect 32474 29464 32495 29504
rect 32577 29464 32598 29504
rect 32598 29464 32638 29504
rect 32638 29464 32663 29504
rect 32409 29441 32495 29464
rect 32577 29441 32663 29464
rect 36409 29504 36495 29527
rect 36577 29504 36663 29527
rect 36409 29464 36434 29504
rect 36434 29464 36474 29504
rect 36474 29464 36495 29504
rect 36577 29464 36598 29504
rect 36598 29464 36638 29504
rect 36638 29464 36663 29504
rect 36409 29441 36495 29464
rect 36577 29441 36663 29464
rect 40409 29504 40495 29527
rect 40577 29504 40663 29527
rect 40409 29464 40434 29504
rect 40434 29464 40474 29504
rect 40474 29464 40495 29504
rect 40577 29464 40598 29504
rect 40598 29464 40638 29504
rect 40638 29464 40663 29504
rect 40409 29441 40495 29464
rect 40577 29441 40663 29464
rect 44409 29504 44495 29527
rect 44577 29504 44663 29527
rect 44409 29464 44434 29504
rect 44434 29464 44474 29504
rect 44474 29464 44495 29504
rect 44577 29464 44598 29504
rect 44598 29464 44638 29504
rect 44638 29464 44663 29504
rect 44409 29441 44495 29464
rect 44577 29441 44663 29464
rect 48409 29504 48495 29527
rect 48577 29504 48663 29527
rect 48409 29464 48434 29504
rect 48434 29464 48474 29504
rect 48474 29464 48495 29504
rect 48577 29464 48598 29504
rect 48598 29464 48638 29504
rect 48638 29464 48663 29504
rect 48409 29441 48495 29464
rect 48577 29441 48663 29464
rect 52409 29504 52495 29527
rect 52577 29504 52663 29527
rect 52409 29464 52434 29504
rect 52434 29464 52474 29504
rect 52474 29464 52495 29504
rect 52577 29464 52598 29504
rect 52598 29464 52638 29504
rect 52638 29464 52663 29504
rect 52409 29441 52495 29464
rect 52577 29441 52663 29464
rect 56409 29504 56495 29527
rect 56577 29504 56663 29527
rect 56409 29464 56434 29504
rect 56434 29464 56474 29504
rect 56474 29464 56495 29504
rect 56577 29464 56598 29504
rect 56598 29464 56638 29504
rect 56638 29464 56663 29504
rect 56409 29441 56495 29464
rect 56577 29441 56663 29464
rect 60409 29504 60495 29527
rect 60577 29504 60663 29527
rect 60409 29464 60434 29504
rect 60434 29464 60474 29504
rect 60474 29464 60495 29504
rect 60577 29464 60598 29504
rect 60598 29464 60638 29504
rect 60638 29464 60663 29504
rect 60409 29441 60495 29464
rect 60577 29441 60663 29464
rect 64409 29504 64495 29527
rect 64577 29504 64663 29527
rect 64409 29464 64434 29504
rect 64434 29464 64474 29504
rect 64474 29464 64495 29504
rect 64577 29464 64598 29504
rect 64598 29464 64638 29504
rect 64638 29464 64663 29504
rect 64409 29441 64495 29464
rect 64577 29441 64663 29464
rect 68409 29504 68495 29527
rect 68577 29504 68663 29527
rect 68409 29464 68434 29504
rect 68434 29464 68474 29504
rect 68474 29464 68495 29504
rect 68577 29464 68598 29504
rect 68598 29464 68638 29504
rect 68638 29464 68663 29504
rect 68409 29441 68495 29464
rect 68577 29441 68663 29464
rect 72409 29524 72495 29610
rect 72577 29524 72663 29610
rect 72409 29356 72495 29442
rect 72577 29356 72663 29442
rect 72409 29188 72495 29274
rect 72577 29188 72663 29274
rect 72409 29020 72495 29106
rect 72577 29020 72663 29106
rect 76409 31036 76495 31122
rect 76577 31036 76663 31122
rect 76409 30868 76495 30954
rect 76577 30868 76663 30954
rect 76409 30700 76495 30786
rect 76577 30700 76663 30786
rect 76409 30532 76495 30618
rect 76577 30532 76663 30618
rect 76409 30364 76495 30450
rect 76577 30364 76663 30450
rect 76409 30196 76495 30282
rect 76577 30196 76663 30282
rect 76409 30028 76495 30114
rect 76577 30028 76663 30114
rect 76409 29860 76495 29946
rect 76577 29860 76663 29946
rect 76409 29692 76495 29778
rect 76577 29692 76663 29778
rect 76409 29524 76495 29610
rect 76577 29524 76663 29610
rect 76409 29356 76495 29442
rect 76577 29356 76663 29442
rect 76409 29188 76495 29274
rect 76577 29188 76663 29274
rect 76409 29020 76495 29106
rect 76577 29020 76663 29106
rect 80409 31036 80495 31122
rect 80577 31036 80663 31122
rect 80409 30868 80495 30954
rect 80577 30868 80663 30954
rect 80409 30700 80495 30786
rect 80577 30700 80663 30786
rect 80409 30532 80495 30618
rect 80577 30532 80663 30618
rect 80409 30364 80495 30450
rect 80577 30364 80663 30450
rect 80409 30196 80495 30282
rect 80577 30196 80663 30282
rect 80409 30028 80495 30114
rect 80577 30028 80663 30114
rect 80409 29860 80495 29946
rect 80577 29860 80663 29946
rect 80409 29692 80495 29778
rect 80577 29692 80663 29778
rect 80409 29524 80495 29610
rect 80577 29524 80663 29610
rect 80409 29356 80495 29442
rect 80577 29356 80663 29442
rect 80409 29188 80495 29274
rect 80577 29188 80663 29274
rect 80409 29020 80495 29106
rect 80577 29020 80663 29106
rect 84409 31036 84495 31122
rect 84577 31036 84663 31122
rect 84409 30868 84495 30954
rect 84577 30868 84663 30954
rect 84409 30700 84495 30786
rect 84577 30700 84663 30786
rect 84409 30532 84495 30618
rect 84577 30532 84663 30618
rect 84409 30364 84495 30450
rect 84577 30364 84663 30450
rect 84409 30196 84495 30282
rect 84577 30196 84663 30282
rect 84409 30028 84495 30114
rect 84577 30028 84663 30114
rect 84409 29860 84495 29946
rect 84577 29860 84663 29946
rect 84409 29692 84495 29778
rect 84577 29692 84663 29778
rect 84409 29524 84495 29610
rect 84577 29524 84663 29610
rect 84409 29356 84495 29442
rect 84577 29356 84663 29442
rect 84409 29188 84495 29274
rect 84577 29188 84663 29274
rect 84409 29020 84495 29106
rect 84577 29020 84663 29106
rect 88409 31036 88495 31122
rect 88577 31036 88663 31122
rect 88409 30868 88495 30954
rect 88577 30868 88663 30954
rect 88409 30700 88495 30786
rect 88577 30700 88663 30786
rect 88409 30532 88495 30618
rect 88577 30532 88663 30618
rect 88409 30364 88495 30450
rect 88577 30364 88663 30450
rect 88409 30196 88495 30282
rect 88577 30196 88663 30282
rect 88409 30028 88495 30114
rect 88577 30028 88663 30114
rect 88409 29860 88495 29946
rect 88577 29860 88663 29946
rect 88409 29692 88495 29778
rect 88577 29692 88663 29778
rect 88409 29524 88495 29610
rect 88577 29524 88663 29610
rect 88409 29356 88495 29442
rect 88577 29356 88663 29442
rect 88409 29188 88495 29274
rect 88577 29188 88663 29274
rect 88409 29020 88495 29106
rect 88577 29020 88663 29106
rect 92409 31036 92495 31122
rect 92577 31036 92663 31122
rect 92409 30868 92495 30954
rect 92577 30868 92663 30954
rect 92409 30700 92495 30786
rect 92577 30700 92663 30786
rect 92409 30532 92495 30618
rect 92577 30532 92663 30618
rect 92409 30364 92495 30450
rect 92577 30364 92663 30450
rect 92409 30196 92495 30282
rect 92577 30196 92663 30282
rect 92409 30028 92495 30114
rect 92577 30028 92663 30114
rect 92409 29860 92495 29946
rect 92577 29860 92663 29946
rect 92409 29692 92495 29778
rect 92577 29692 92663 29778
rect 92409 29524 92495 29610
rect 92577 29524 92663 29610
rect 92409 29356 92495 29442
rect 92577 29356 92663 29442
rect 92409 29188 92495 29274
rect 92577 29188 92663 29274
rect 92409 29020 92495 29106
rect 92577 29020 92663 29106
rect 96409 31036 96495 31122
rect 96577 31036 96663 31122
rect 96409 30868 96495 30954
rect 96577 30868 96663 30954
rect 96409 30700 96495 30786
rect 96577 30700 96663 30786
rect 96409 30532 96495 30618
rect 96577 30532 96663 30618
rect 96409 30364 96495 30450
rect 96577 30364 96663 30450
rect 96409 30196 96495 30282
rect 96577 30196 96663 30282
rect 96409 30028 96495 30114
rect 96577 30028 96663 30114
rect 96409 29860 96495 29946
rect 96577 29860 96663 29946
rect 96409 29692 96495 29778
rect 96577 29692 96663 29778
rect 96409 29524 96495 29610
rect 96577 29524 96663 29610
rect 96409 29356 96495 29442
rect 96577 29356 96663 29442
rect 96409 29188 96495 29274
rect 96577 29188 96663 29274
rect 96409 29020 96495 29106
rect 96577 29020 96663 29106
rect 3169 28748 3255 28771
rect 3337 28748 3423 28771
rect 3169 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3255 28748
rect 3337 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3423 28748
rect 3169 28685 3255 28708
rect 3337 28685 3423 28708
rect 7169 28748 7255 28771
rect 7337 28748 7423 28771
rect 7169 28708 7194 28748
rect 7194 28708 7234 28748
rect 7234 28708 7255 28748
rect 7337 28708 7358 28748
rect 7358 28708 7398 28748
rect 7398 28708 7423 28748
rect 7169 28685 7255 28708
rect 7337 28685 7423 28708
rect 11169 28748 11255 28771
rect 11337 28748 11423 28771
rect 11169 28708 11194 28748
rect 11194 28708 11234 28748
rect 11234 28708 11255 28748
rect 11337 28708 11358 28748
rect 11358 28708 11398 28748
rect 11398 28708 11423 28748
rect 11169 28685 11255 28708
rect 11337 28685 11423 28708
rect 15169 28748 15255 28771
rect 15337 28748 15423 28771
rect 15169 28708 15194 28748
rect 15194 28708 15234 28748
rect 15234 28708 15255 28748
rect 15337 28708 15358 28748
rect 15358 28708 15398 28748
rect 15398 28708 15423 28748
rect 15169 28685 15255 28708
rect 15337 28685 15423 28708
rect 19169 28748 19255 28771
rect 19337 28748 19423 28771
rect 19169 28708 19194 28748
rect 19194 28708 19234 28748
rect 19234 28708 19255 28748
rect 19337 28708 19358 28748
rect 19358 28708 19398 28748
rect 19398 28708 19423 28748
rect 19169 28685 19255 28708
rect 19337 28685 19423 28708
rect 23169 28748 23255 28771
rect 23337 28748 23423 28771
rect 23169 28708 23194 28748
rect 23194 28708 23234 28748
rect 23234 28708 23255 28748
rect 23337 28708 23358 28748
rect 23358 28708 23398 28748
rect 23398 28708 23423 28748
rect 23169 28685 23255 28708
rect 23337 28685 23423 28708
rect 27169 28748 27255 28771
rect 27337 28748 27423 28771
rect 27169 28708 27194 28748
rect 27194 28708 27234 28748
rect 27234 28708 27255 28748
rect 27337 28708 27358 28748
rect 27358 28708 27398 28748
rect 27398 28708 27423 28748
rect 27169 28685 27255 28708
rect 27337 28685 27423 28708
rect 31169 28748 31255 28771
rect 31337 28748 31423 28771
rect 31169 28708 31194 28748
rect 31194 28708 31234 28748
rect 31234 28708 31255 28748
rect 31337 28708 31358 28748
rect 31358 28708 31398 28748
rect 31398 28708 31423 28748
rect 31169 28685 31255 28708
rect 31337 28685 31423 28708
rect 35169 28748 35255 28771
rect 35337 28748 35423 28771
rect 35169 28708 35194 28748
rect 35194 28708 35234 28748
rect 35234 28708 35255 28748
rect 35337 28708 35358 28748
rect 35358 28708 35398 28748
rect 35398 28708 35423 28748
rect 35169 28685 35255 28708
rect 35337 28685 35423 28708
rect 39169 28748 39255 28771
rect 39337 28748 39423 28771
rect 39169 28708 39194 28748
rect 39194 28708 39234 28748
rect 39234 28708 39255 28748
rect 39337 28708 39358 28748
rect 39358 28708 39398 28748
rect 39398 28708 39423 28748
rect 39169 28685 39255 28708
rect 39337 28685 39423 28708
rect 43169 28748 43255 28771
rect 43337 28748 43423 28771
rect 43169 28708 43194 28748
rect 43194 28708 43234 28748
rect 43234 28708 43255 28748
rect 43337 28708 43358 28748
rect 43358 28708 43398 28748
rect 43398 28708 43423 28748
rect 43169 28685 43255 28708
rect 43337 28685 43423 28708
rect 47169 28748 47255 28771
rect 47337 28748 47423 28771
rect 47169 28708 47194 28748
rect 47194 28708 47234 28748
rect 47234 28708 47255 28748
rect 47337 28708 47358 28748
rect 47358 28708 47398 28748
rect 47398 28708 47423 28748
rect 47169 28685 47255 28708
rect 47337 28685 47423 28708
rect 51169 28748 51255 28771
rect 51337 28748 51423 28771
rect 51169 28708 51194 28748
rect 51194 28708 51234 28748
rect 51234 28708 51255 28748
rect 51337 28708 51358 28748
rect 51358 28708 51398 28748
rect 51398 28708 51423 28748
rect 51169 28685 51255 28708
rect 51337 28685 51423 28708
rect 55169 28748 55255 28771
rect 55337 28748 55423 28771
rect 55169 28708 55194 28748
rect 55194 28708 55234 28748
rect 55234 28708 55255 28748
rect 55337 28708 55358 28748
rect 55358 28708 55398 28748
rect 55398 28708 55423 28748
rect 55169 28685 55255 28708
rect 55337 28685 55423 28708
rect 59169 28748 59255 28771
rect 59337 28748 59423 28771
rect 59169 28708 59194 28748
rect 59194 28708 59234 28748
rect 59234 28708 59255 28748
rect 59337 28708 59358 28748
rect 59358 28708 59398 28748
rect 59398 28708 59423 28748
rect 59169 28685 59255 28708
rect 59337 28685 59423 28708
rect 63169 28748 63255 28771
rect 63337 28748 63423 28771
rect 63169 28708 63194 28748
rect 63194 28708 63234 28748
rect 63234 28708 63255 28748
rect 63337 28708 63358 28748
rect 63358 28708 63398 28748
rect 63398 28708 63423 28748
rect 63169 28685 63255 28708
rect 63337 28685 63423 28708
rect 67169 28748 67255 28771
rect 67337 28748 67423 28771
rect 67169 28708 67194 28748
rect 67194 28708 67234 28748
rect 67234 28708 67255 28748
rect 67337 28708 67358 28748
rect 67358 28708 67398 28748
rect 67398 28708 67423 28748
rect 67169 28685 67255 28708
rect 67337 28685 67423 28708
rect 75169 28160 75255 28246
rect 75337 28160 75423 28246
rect 4409 27992 4495 28015
rect 4577 27992 4663 28015
rect 4409 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4495 27992
rect 4577 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4663 27992
rect 4409 27929 4495 27952
rect 4577 27929 4663 27952
rect 8409 27992 8495 28015
rect 8577 27992 8663 28015
rect 8409 27952 8434 27992
rect 8434 27952 8474 27992
rect 8474 27952 8495 27992
rect 8577 27952 8598 27992
rect 8598 27952 8638 27992
rect 8638 27952 8663 27992
rect 8409 27929 8495 27952
rect 8577 27929 8663 27952
rect 12409 27992 12495 28015
rect 12577 27992 12663 28015
rect 12409 27952 12434 27992
rect 12434 27952 12474 27992
rect 12474 27952 12495 27992
rect 12577 27952 12598 27992
rect 12598 27952 12638 27992
rect 12638 27952 12663 27992
rect 12409 27929 12495 27952
rect 12577 27929 12663 27952
rect 16409 27992 16495 28015
rect 16577 27992 16663 28015
rect 16409 27952 16434 27992
rect 16434 27952 16474 27992
rect 16474 27952 16495 27992
rect 16577 27952 16598 27992
rect 16598 27952 16638 27992
rect 16638 27952 16663 27992
rect 16409 27929 16495 27952
rect 16577 27929 16663 27952
rect 20409 27992 20495 28015
rect 20577 27992 20663 28015
rect 20409 27952 20434 27992
rect 20434 27952 20474 27992
rect 20474 27952 20495 27992
rect 20577 27952 20598 27992
rect 20598 27952 20638 27992
rect 20638 27952 20663 27992
rect 20409 27929 20495 27952
rect 20577 27929 20663 27952
rect 24409 27992 24495 28015
rect 24577 27992 24663 28015
rect 24409 27952 24434 27992
rect 24434 27952 24474 27992
rect 24474 27952 24495 27992
rect 24577 27952 24598 27992
rect 24598 27952 24638 27992
rect 24638 27952 24663 27992
rect 24409 27929 24495 27952
rect 24577 27929 24663 27952
rect 28409 27992 28495 28015
rect 28577 27992 28663 28015
rect 28409 27952 28434 27992
rect 28434 27952 28474 27992
rect 28474 27952 28495 27992
rect 28577 27952 28598 27992
rect 28598 27952 28638 27992
rect 28638 27952 28663 27992
rect 28409 27929 28495 27952
rect 28577 27929 28663 27952
rect 32409 27992 32495 28015
rect 32577 27992 32663 28015
rect 32409 27952 32434 27992
rect 32434 27952 32474 27992
rect 32474 27952 32495 27992
rect 32577 27952 32598 27992
rect 32598 27952 32638 27992
rect 32638 27952 32663 27992
rect 32409 27929 32495 27952
rect 32577 27929 32663 27952
rect 36409 27992 36495 28015
rect 36577 27992 36663 28015
rect 36409 27952 36434 27992
rect 36434 27952 36474 27992
rect 36474 27952 36495 27992
rect 36577 27952 36598 27992
rect 36598 27952 36638 27992
rect 36638 27952 36663 27992
rect 36409 27929 36495 27952
rect 36577 27929 36663 27952
rect 40409 27992 40495 28015
rect 40577 27992 40663 28015
rect 40409 27952 40434 27992
rect 40434 27952 40474 27992
rect 40474 27952 40495 27992
rect 40577 27952 40598 27992
rect 40598 27952 40638 27992
rect 40638 27952 40663 27992
rect 40409 27929 40495 27952
rect 40577 27929 40663 27952
rect 44409 27992 44495 28015
rect 44577 27992 44663 28015
rect 44409 27952 44434 27992
rect 44434 27952 44474 27992
rect 44474 27952 44495 27992
rect 44577 27952 44598 27992
rect 44598 27952 44638 27992
rect 44638 27952 44663 27992
rect 44409 27929 44495 27952
rect 44577 27929 44663 27952
rect 48409 27992 48495 28015
rect 48577 27992 48663 28015
rect 48409 27952 48434 27992
rect 48434 27952 48474 27992
rect 48474 27952 48495 27992
rect 48577 27952 48598 27992
rect 48598 27952 48638 27992
rect 48638 27952 48663 27992
rect 48409 27929 48495 27952
rect 48577 27929 48663 27952
rect 52409 27992 52495 28015
rect 52577 27992 52663 28015
rect 52409 27952 52434 27992
rect 52434 27952 52474 27992
rect 52474 27952 52495 27992
rect 52577 27952 52598 27992
rect 52598 27952 52638 27992
rect 52638 27952 52663 27992
rect 52409 27929 52495 27952
rect 52577 27929 52663 27952
rect 56409 27992 56495 28015
rect 56577 27992 56663 28015
rect 56409 27952 56434 27992
rect 56434 27952 56474 27992
rect 56474 27952 56495 27992
rect 56577 27952 56598 27992
rect 56598 27952 56638 27992
rect 56638 27952 56663 27992
rect 56409 27929 56495 27952
rect 56577 27929 56663 27952
rect 60409 27992 60495 28015
rect 60577 27992 60663 28015
rect 60409 27952 60434 27992
rect 60434 27952 60474 27992
rect 60474 27952 60495 27992
rect 60577 27952 60598 27992
rect 60598 27952 60638 27992
rect 60638 27952 60663 27992
rect 60409 27929 60495 27952
rect 60577 27929 60663 27952
rect 64409 27992 64495 28015
rect 64577 27992 64663 28015
rect 64409 27952 64434 27992
rect 64434 27952 64474 27992
rect 64474 27952 64495 27992
rect 64577 27952 64598 27992
rect 64598 27952 64638 27992
rect 64638 27952 64663 27992
rect 64409 27929 64495 27952
rect 64577 27929 64663 27952
rect 68409 27992 68495 28015
rect 68577 27992 68663 28015
rect 68409 27952 68434 27992
rect 68434 27952 68474 27992
rect 68474 27952 68495 27992
rect 68577 27952 68598 27992
rect 68598 27952 68638 27992
rect 68638 27952 68663 27992
rect 68409 27929 68495 27952
rect 68577 27929 68663 27952
rect 75169 27992 75255 28078
rect 75337 27992 75423 28078
rect 75169 27824 75255 27910
rect 75337 27824 75423 27910
rect 75169 27656 75255 27742
rect 75337 27656 75423 27742
rect 75169 27488 75255 27574
rect 75337 27488 75423 27574
rect 75169 27320 75255 27406
rect 75337 27320 75423 27406
rect 3169 27236 3255 27259
rect 3337 27236 3423 27259
rect 3169 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3255 27236
rect 3337 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3423 27236
rect 3169 27173 3255 27196
rect 3337 27173 3423 27196
rect 7169 27236 7255 27259
rect 7337 27236 7423 27259
rect 7169 27196 7194 27236
rect 7194 27196 7234 27236
rect 7234 27196 7255 27236
rect 7337 27196 7358 27236
rect 7358 27196 7398 27236
rect 7398 27196 7423 27236
rect 7169 27173 7255 27196
rect 7337 27173 7423 27196
rect 11169 27236 11255 27259
rect 11337 27236 11423 27259
rect 11169 27196 11194 27236
rect 11194 27196 11234 27236
rect 11234 27196 11255 27236
rect 11337 27196 11358 27236
rect 11358 27196 11398 27236
rect 11398 27196 11423 27236
rect 11169 27173 11255 27196
rect 11337 27173 11423 27196
rect 15169 27236 15255 27259
rect 15337 27236 15423 27259
rect 15169 27196 15194 27236
rect 15194 27196 15234 27236
rect 15234 27196 15255 27236
rect 15337 27196 15358 27236
rect 15358 27196 15398 27236
rect 15398 27196 15423 27236
rect 15169 27173 15255 27196
rect 15337 27173 15423 27196
rect 19169 27236 19255 27259
rect 19337 27236 19423 27259
rect 19169 27196 19194 27236
rect 19194 27196 19234 27236
rect 19234 27196 19255 27236
rect 19337 27196 19358 27236
rect 19358 27196 19398 27236
rect 19398 27196 19423 27236
rect 19169 27173 19255 27196
rect 19337 27173 19423 27196
rect 23169 27236 23255 27259
rect 23337 27236 23423 27259
rect 23169 27196 23194 27236
rect 23194 27196 23234 27236
rect 23234 27196 23255 27236
rect 23337 27196 23358 27236
rect 23358 27196 23398 27236
rect 23398 27196 23423 27236
rect 23169 27173 23255 27196
rect 23337 27173 23423 27196
rect 27169 27236 27255 27259
rect 27337 27236 27423 27259
rect 27169 27196 27194 27236
rect 27194 27196 27234 27236
rect 27234 27196 27255 27236
rect 27337 27196 27358 27236
rect 27358 27196 27398 27236
rect 27398 27196 27423 27236
rect 27169 27173 27255 27196
rect 27337 27173 27423 27196
rect 31169 27236 31255 27259
rect 31337 27236 31423 27259
rect 31169 27196 31194 27236
rect 31194 27196 31234 27236
rect 31234 27196 31255 27236
rect 31337 27196 31358 27236
rect 31358 27196 31398 27236
rect 31398 27196 31423 27236
rect 31169 27173 31255 27196
rect 31337 27173 31423 27196
rect 35169 27236 35255 27259
rect 35337 27236 35423 27259
rect 35169 27196 35194 27236
rect 35194 27196 35234 27236
rect 35234 27196 35255 27236
rect 35337 27196 35358 27236
rect 35358 27196 35398 27236
rect 35398 27196 35423 27236
rect 35169 27173 35255 27196
rect 35337 27173 35423 27196
rect 39169 27236 39255 27259
rect 39337 27236 39423 27259
rect 39169 27196 39194 27236
rect 39194 27196 39234 27236
rect 39234 27196 39255 27236
rect 39337 27196 39358 27236
rect 39358 27196 39398 27236
rect 39398 27196 39423 27236
rect 39169 27173 39255 27196
rect 39337 27173 39423 27196
rect 43169 27236 43255 27259
rect 43337 27236 43423 27259
rect 43169 27196 43194 27236
rect 43194 27196 43234 27236
rect 43234 27196 43255 27236
rect 43337 27196 43358 27236
rect 43358 27196 43398 27236
rect 43398 27196 43423 27236
rect 43169 27173 43255 27196
rect 43337 27173 43423 27196
rect 47169 27236 47255 27259
rect 47337 27236 47423 27259
rect 47169 27196 47194 27236
rect 47194 27196 47234 27236
rect 47234 27196 47255 27236
rect 47337 27196 47358 27236
rect 47358 27196 47398 27236
rect 47398 27196 47423 27236
rect 47169 27173 47255 27196
rect 47337 27173 47423 27196
rect 51169 27236 51255 27259
rect 51337 27236 51423 27259
rect 51169 27196 51194 27236
rect 51194 27196 51234 27236
rect 51234 27196 51255 27236
rect 51337 27196 51358 27236
rect 51358 27196 51398 27236
rect 51398 27196 51423 27236
rect 51169 27173 51255 27196
rect 51337 27173 51423 27196
rect 55169 27236 55255 27259
rect 55337 27236 55423 27259
rect 55169 27196 55194 27236
rect 55194 27196 55234 27236
rect 55234 27196 55255 27236
rect 55337 27196 55358 27236
rect 55358 27196 55398 27236
rect 55398 27196 55423 27236
rect 55169 27173 55255 27196
rect 55337 27173 55423 27196
rect 59169 27236 59255 27259
rect 59337 27236 59423 27259
rect 59169 27196 59194 27236
rect 59194 27196 59234 27236
rect 59234 27196 59255 27236
rect 59337 27196 59358 27236
rect 59358 27196 59398 27236
rect 59398 27196 59423 27236
rect 59169 27173 59255 27196
rect 59337 27173 59423 27196
rect 63169 27236 63255 27259
rect 63337 27236 63423 27259
rect 63169 27196 63194 27236
rect 63194 27196 63234 27236
rect 63234 27196 63255 27236
rect 63337 27196 63358 27236
rect 63358 27196 63398 27236
rect 63398 27196 63423 27236
rect 63169 27173 63255 27196
rect 63337 27173 63423 27196
rect 67169 27236 67255 27259
rect 67337 27236 67423 27259
rect 67169 27196 67194 27236
rect 67194 27196 67234 27236
rect 67234 27196 67255 27236
rect 67337 27196 67358 27236
rect 67358 27196 67398 27236
rect 67398 27196 67423 27236
rect 67169 27173 67255 27196
rect 67337 27173 67423 27196
rect 75169 27152 75255 27238
rect 75337 27152 75423 27238
rect 75169 26984 75255 27070
rect 75337 26984 75423 27070
rect 75169 26816 75255 26902
rect 75337 26816 75423 26902
rect 75169 26648 75255 26734
rect 75337 26648 75423 26734
rect 4409 26480 4495 26503
rect 4577 26480 4663 26503
rect 4409 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4495 26480
rect 4577 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4663 26480
rect 4409 26417 4495 26440
rect 4577 26417 4663 26440
rect 8409 26480 8495 26503
rect 8577 26480 8663 26503
rect 8409 26440 8434 26480
rect 8434 26440 8474 26480
rect 8474 26440 8495 26480
rect 8577 26440 8598 26480
rect 8598 26440 8638 26480
rect 8638 26440 8663 26480
rect 8409 26417 8495 26440
rect 8577 26417 8663 26440
rect 12409 26480 12495 26503
rect 12577 26480 12663 26503
rect 12409 26440 12434 26480
rect 12434 26440 12474 26480
rect 12474 26440 12495 26480
rect 12577 26440 12598 26480
rect 12598 26440 12638 26480
rect 12638 26440 12663 26480
rect 12409 26417 12495 26440
rect 12577 26417 12663 26440
rect 16409 26480 16495 26503
rect 16577 26480 16663 26503
rect 16409 26440 16434 26480
rect 16434 26440 16474 26480
rect 16474 26440 16495 26480
rect 16577 26440 16598 26480
rect 16598 26440 16638 26480
rect 16638 26440 16663 26480
rect 16409 26417 16495 26440
rect 16577 26417 16663 26440
rect 20409 26480 20495 26503
rect 20577 26480 20663 26503
rect 20409 26440 20434 26480
rect 20434 26440 20474 26480
rect 20474 26440 20495 26480
rect 20577 26440 20598 26480
rect 20598 26440 20638 26480
rect 20638 26440 20663 26480
rect 20409 26417 20495 26440
rect 20577 26417 20663 26440
rect 24409 26480 24495 26503
rect 24577 26480 24663 26503
rect 24409 26440 24434 26480
rect 24434 26440 24474 26480
rect 24474 26440 24495 26480
rect 24577 26440 24598 26480
rect 24598 26440 24638 26480
rect 24638 26440 24663 26480
rect 24409 26417 24495 26440
rect 24577 26417 24663 26440
rect 28409 26480 28495 26503
rect 28577 26480 28663 26503
rect 28409 26440 28434 26480
rect 28434 26440 28474 26480
rect 28474 26440 28495 26480
rect 28577 26440 28598 26480
rect 28598 26440 28638 26480
rect 28638 26440 28663 26480
rect 28409 26417 28495 26440
rect 28577 26417 28663 26440
rect 32409 26480 32495 26503
rect 32577 26480 32663 26503
rect 32409 26440 32434 26480
rect 32434 26440 32474 26480
rect 32474 26440 32495 26480
rect 32577 26440 32598 26480
rect 32598 26440 32638 26480
rect 32638 26440 32663 26480
rect 32409 26417 32495 26440
rect 32577 26417 32663 26440
rect 36409 26480 36495 26503
rect 36577 26480 36663 26503
rect 36409 26440 36434 26480
rect 36434 26440 36474 26480
rect 36474 26440 36495 26480
rect 36577 26440 36598 26480
rect 36598 26440 36638 26480
rect 36638 26440 36663 26480
rect 36409 26417 36495 26440
rect 36577 26417 36663 26440
rect 40409 26480 40495 26503
rect 40577 26480 40663 26503
rect 40409 26440 40434 26480
rect 40434 26440 40474 26480
rect 40474 26440 40495 26480
rect 40577 26440 40598 26480
rect 40598 26440 40638 26480
rect 40638 26440 40663 26480
rect 40409 26417 40495 26440
rect 40577 26417 40663 26440
rect 44409 26480 44495 26503
rect 44577 26480 44663 26503
rect 44409 26440 44434 26480
rect 44434 26440 44474 26480
rect 44474 26440 44495 26480
rect 44577 26440 44598 26480
rect 44598 26440 44638 26480
rect 44638 26440 44663 26480
rect 44409 26417 44495 26440
rect 44577 26417 44663 26440
rect 48409 26480 48495 26503
rect 48577 26480 48663 26503
rect 48409 26440 48434 26480
rect 48434 26440 48474 26480
rect 48474 26440 48495 26480
rect 48577 26440 48598 26480
rect 48598 26440 48638 26480
rect 48638 26440 48663 26480
rect 48409 26417 48495 26440
rect 48577 26417 48663 26440
rect 52409 26480 52495 26503
rect 52577 26480 52663 26503
rect 52409 26440 52434 26480
rect 52434 26440 52474 26480
rect 52474 26440 52495 26480
rect 52577 26440 52598 26480
rect 52598 26440 52638 26480
rect 52638 26440 52663 26480
rect 52409 26417 52495 26440
rect 52577 26417 52663 26440
rect 56409 26480 56495 26503
rect 56577 26480 56663 26503
rect 56409 26440 56434 26480
rect 56434 26440 56474 26480
rect 56474 26440 56495 26480
rect 56577 26440 56598 26480
rect 56598 26440 56638 26480
rect 56638 26440 56663 26480
rect 56409 26417 56495 26440
rect 56577 26417 56663 26440
rect 60409 26480 60495 26503
rect 60577 26480 60663 26503
rect 60409 26440 60434 26480
rect 60434 26440 60474 26480
rect 60474 26440 60495 26480
rect 60577 26440 60598 26480
rect 60598 26440 60638 26480
rect 60638 26440 60663 26480
rect 60409 26417 60495 26440
rect 60577 26417 60663 26440
rect 64409 26480 64495 26503
rect 64577 26480 64663 26503
rect 64409 26440 64434 26480
rect 64434 26440 64474 26480
rect 64474 26440 64495 26480
rect 64577 26440 64598 26480
rect 64598 26440 64638 26480
rect 64638 26440 64663 26480
rect 64409 26417 64495 26440
rect 64577 26417 64663 26440
rect 68409 26480 68495 26503
rect 68577 26480 68663 26503
rect 68409 26440 68434 26480
rect 68434 26440 68474 26480
rect 68474 26440 68495 26480
rect 68577 26440 68598 26480
rect 68598 26440 68638 26480
rect 68638 26440 68663 26480
rect 68409 26417 68495 26440
rect 68577 26417 68663 26440
rect 75169 26480 75255 26566
rect 75337 26480 75423 26566
rect 75169 26312 75255 26398
rect 75337 26312 75423 26398
rect 75169 26144 75255 26230
rect 75337 26144 75423 26230
rect 79169 28160 79255 28246
rect 79337 28160 79423 28246
rect 79169 27992 79255 28078
rect 79337 27992 79423 28078
rect 79169 27824 79255 27910
rect 79337 27824 79423 27910
rect 79169 27656 79255 27742
rect 79337 27656 79423 27742
rect 79169 27488 79255 27574
rect 79337 27488 79423 27574
rect 79169 27320 79255 27406
rect 79337 27320 79423 27406
rect 79169 27152 79255 27238
rect 79337 27152 79423 27238
rect 79169 26984 79255 27070
rect 79337 26984 79423 27070
rect 79169 26816 79255 26902
rect 79337 26816 79423 26902
rect 79169 26648 79255 26734
rect 79337 26648 79423 26734
rect 79169 26480 79255 26566
rect 79337 26480 79423 26566
rect 79169 26312 79255 26398
rect 79337 26312 79423 26398
rect 79169 26144 79255 26230
rect 79337 26144 79423 26230
rect 83169 28160 83255 28246
rect 83337 28160 83423 28246
rect 83169 27992 83255 28078
rect 83337 27992 83423 28078
rect 83169 27824 83255 27910
rect 83337 27824 83423 27910
rect 83169 27656 83255 27742
rect 83337 27656 83423 27742
rect 83169 27488 83255 27574
rect 83337 27488 83423 27574
rect 83169 27320 83255 27406
rect 83337 27320 83423 27406
rect 83169 27152 83255 27238
rect 83337 27152 83423 27238
rect 83169 26984 83255 27070
rect 83337 26984 83423 27070
rect 83169 26816 83255 26902
rect 83337 26816 83423 26902
rect 83169 26648 83255 26734
rect 83337 26648 83423 26734
rect 83169 26480 83255 26566
rect 83337 26480 83423 26566
rect 83169 26312 83255 26398
rect 83337 26312 83423 26398
rect 83169 26144 83255 26230
rect 83337 26144 83423 26230
rect 87169 28160 87255 28246
rect 87337 28160 87423 28246
rect 87169 27992 87255 28078
rect 87337 27992 87423 28078
rect 87169 27824 87255 27910
rect 87337 27824 87423 27910
rect 87169 27656 87255 27742
rect 87337 27656 87423 27742
rect 87169 27488 87255 27574
rect 87337 27488 87423 27574
rect 87169 27320 87255 27406
rect 87337 27320 87423 27406
rect 87169 27152 87255 27238
rect 87337 27152 87423 27238
rect 87169 26984 87255 27070
rect 87337 26984 87423 27070
rect 87169 26816 87255 26902
rect 87337 26816 87423 26902
rect 87169 26648 87255 26734
rect 87337 26648 87423 26734
rect 87169 26480 87255 26566
rect 87337 26480 87423 26566
rect 87169 26312 87255 26398
rect 87337 26312 87423 26398
rect 87169 26144 87255 26230
rect 87337 26144 87423 26230
rect 91169 28160 91255 28246
rect 91337 28160 91423 28246
rect 91169 27992 91255 28078
rect 91337 27992 91423 28078
rect 91169 27824 91255 27910
rect 91337 27824 91423 27910
rect 91169 27656 91255 27742
rect 91337 27656 91423 27742
rect 91169 27488 91255 27574
rect 91337 27488 91423 27574
rect 91169 27320 91255 27406
rect 91337 27320 91423 27406
rect 91169 27152 91255 27238
rect 91337 27152 91423 27238
rect 91169 26984 91255 27070
rect 91337 26984 91423 27070
rect 91169 26816 91255 26902
rect 91337 26816 91423 26902
rect 91169 26648 91255 26734
rect 91337 26648 91423 26734
rect 91169 26480 91255 26566
rect 91337 26480 91423 26566
rect 91169 26312 91255 26398
rect 91337 26312 91423 26398
rect 91169 26144 91255 26230
rect 91337 26144 91423 26230
rect 95169 28160 95255 28246
rect 95337 28160 95423 28246
rect 95169 27992 95255 28078
rect 95337 27992 95423 28078
rect 95169 27824 95255 27910
rect 95337 27824 95423 27910
rect 95169 27656 95255 27742
rect 95337 27656 95423 27742
rect 95169 27488 95255 27574
rect 95337 27488 95423 27574
rect 95169 27320 95255 27406
rect 95337 27320 95423 27406
rect 95169 27152 95255 27238
rect 95337 27152 95423 27238
rect 95169 26984 95255 27070
rect 95337 26984 95423 27070
rect 95169 26816 95255 26902
rect 95337 26816 95423 26902
rect 95169 26648 95255 26734
rect 95337 26648 95423 26734
rect 95169 26480 95255 26566
rect 95337 26480 95423 26566
rect 95169 26312 95255 26398
rect 95337 26312 95423 26398
rect 95169 26144 95255 26230
rect 95337 26144 95423 26230
rect 3169 25724 3255 25747
rect 3337 25724 3423 25747
rect 3169 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3255 25724
rect 3337 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3423 25724
rect 3169 25661 3255 25684
rect 3337 25661 3423 25684
rect 7169 25724 7255 25747
rect 7337 25724 7423 25747
rect 7169 25684 7194 25724
rect 7194 25684 7234 25724
rect 7234 25684 7255 25724
rect 7337 25684 7358 25724
rect 7358 25684 7398 25724
rect 7398 25684 7423 25724
rect 7169 25661 7255 25684
rect 7337 25661 7423 25684
rect 11169 25724 11255 25747
rect 11337 25724 11423 25747
rect 11169 25684 11194 25724
rect 11194 25684 11234 25724
rect 11234 25684 11255 25724
rect 11337 25684 11358 25724
rect 11358 25684 11398 25724
rect 11398 25684 11423 25724
rect 11169 25661 11255 25684
rect 11337 25661 11423 25684
rect 15169 25724 15255 25747
rect 15337 25724 15423 25747
rect 15169 25684 15194 25724
rect 15194 25684 15234 25724
rect 15234 25684 15255 25724
rect 15337 25684 15358 25724
rect 15358 25684 15398 25724
rect 15398 25684 15423 25724
rect 15169 25661 15255 25684
rect 15337 25661 15423 25684
rect 19169 25724 19255 25747
rect 19337 25724 19423 25747
rect 19169 25684 19194 25724
rect 19194 25684 19234 25724
rect 19234 25684 19255 25724
rect 19337 25684 19358 25724
rect 19358 25684 19398 25724
rect 19398 25684 19423 25724
rect 19169 25661 19255 25684
rect 19337 25661 19423 25684
rect 23169 25724 23255 25747
rect 23337 25724 23423 25747
rect 23169 25684 23194 25724
rect 23194 25684 23234 25724
rect 23234 25684 23255 25724
rect 23337 25684 23358 25724
rect 23358 25684 23398 25724
rect 23398 25684 23423 25724
rect 23169 25661 23255 25684
rect 23337 25661 23423 25684
rect 27169 25724 27255 25747
rect 27337 25724 27423 25747
rect 27169 25684 27194 25724
rect 27194 25684 27234 25724
rect 27234 25684 27255 25724
rect 27337 25684 27358 25724
rect 27358 25684 27398 25724
rect 27398 25684 27423 25724
rect 27169 25661 27255 25684
rect 27337 25661 27423 25684
rect 31169 25724 31255 25747
rect 31337 25724 31423 25747
rect 31169 25684 31194 25724
rect 31194 25684 31234 25724
rect 31234 25684 31255 25724
rect 31337 25684 31358 25724
rect 31358 25684 31398 25724
rect 31398 25684 31423 25724
rect 31169 25661 31255 25684
rect 31337 25661 31423 25684
rect 35169 25724 35255 25747
rect 35337 25724 35423 25747
rect 35169 25684 35194 25724
rect 35194 25684 35234 25724
rect 35234 25684 35255 25724
rect 35337 25684 35358 25724
rect 35358 25684 35398 25724
rect 35398 25684 35423 25724
rect 35169 25661 35255 25684
rect 35337 25661 35423 25684
rect 39169 25724 39255 25747
rect 39337 25724 39423 25747
rect 39169 25684 39194 25724
rect 39194 25684 39234 25724
rect 39234 25684 39255 25724
rect 39337 25684 39358 25724
rect 39358 25684 39398 25724
rect 39398 25684 39423 25724
rect 39169 25661 39255 25684
rect 39337 25661 39423 25684
rect 43169 25724 43255 25747
rect 43337 25724 43423 25747
rect 43169 25684 43194 25724
rect 43194 25684 43234 25724
rect 43234 25684 43255 25724
rect 43337 25684 43358 25724
rect 43358 25684 43398 25724
rect 43398 25684 43423 25724
rect 43169 25661 43255 25684
rect 43337 25661 43423 25684
rect 47169 25724 47255 25747
rect 47337 25724 47423 25747
rect 47169 25684 47194 25724
rect 47194 25684 47234 25724
rect 47234 25684 47255 25724
rect 47337 25684 47358 25724
rect 47358 25684 47398 25724
rect 47398 25684 47423 25724
rect 47169 25661 47255 25684
rect 47337 25661 47423 25684
rect 51169 25724 51255 25747
rect 51337 25724 51423 25747
rect 51169 25684 51194 25724
rect 51194 25684 51234 25724
rect 51234 25684 51255 25724
rect 51337 25684 51358 25724
rect 51358 25684 51398 25724
rect 51398 25684 51423 25724
rect 51169 25661 51255 25684
rect 51337 25661 51423 25684
rect 55169 25724 55255 25747
rect 55337 25724 55423 25747
rect 55169 25684 55194 25724
rect 55194 25684 55234 25724
rect 55234 25684 55255 25724
rect 55337 25684 55358 25724
rect 55358 25684 55398 25724
rect 55398 25684 55423 25724
rect 55169 25661 55255 25684
rect 55337 25661 55423 25684
rect 59169 25724 59255 25747
rect 59337 25724 59423 25747
rect 59169 25684 59194 25724
rect 59194 25684 59234 25724
rect 59234 25684 59255 25724
rect 59337 25684 59358 25724
rect 59358 25684 59398 25724
rect 59398 25684 59423 25724
rect 59169 25661 59255 25684
rect 59337 25661 59423 25684
rect 63169 25724 63255 25747
rect 63337 25724 63423 25747
rect 63169 25684 63194 25724
rect 63194 25684 63234 25724
rect 63234 25684 63255 25724
rect 63337 25684 63358 25724
rect 63358 25684 63398 25724
rect 63398 25684 63423 25724
rect 63169 25661 63255 25684
rect 63337 25661 63423 25684
rect 67169 25724 67255 25747
rect 67337 25724 67423 25747
rect 67169 25684 67194 25724
rect 67194 25684 67234 25724
rect 67234 25684 67255 25724
rect 67337 25684 67358 25724
rect 67358 25684 67398 25724
rect 67398 25684 67423 25724
rect 67169 25661 67255 25684
rect 67337 25661 67423 25684
rect 4409 24968 4495 24991
rect 4577 24968 4663 24991
rect 4409 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4495 24968
rect 4577 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4663 24968
rect 4409 24905 4495 24928
rect 4577 24905 4663 24928
rect 8409 24968 8495 24991
rect 8577 24968 8663 24991
rect 8409 24928 8434 24968
rect 8434 24928 8474 24968
rect 8474 24928 8495 24968
rect 8577 24928 8598 24968
rect 8598 24928 8638 24968
rect 8638 24928 8663 24968
rect 8409 24905 8495 24928
rect 8577 24905 8663 24928
rect 12409 24968 12495 24991
rect 12577 24968 12663 24991
rect 12409 24928 12434 24968
rect 12434 24928 12474 24968
rect 12474 24928 12495 24968
rect 12577 24928 12598 24968
rect 12598 24928 12638 24968
rect 12638 24928 12663 24968
rect 12409 24905 12495 24928
rect 12577 24905 12663 24928
rect 16409 24968 16495 24991
rect 16577 24968 16663 24991
rect 16409 24928 16434 24968
rect 16434 24928 16474 24968
rect 16474 24928 16495 24968
rect 16577 24928 16598 24968
rect 16598 24928 16638 24968
rect 16638 24928 16663 24968
rect 16409 24905 16495 24928
rect 16577 24905 16663 24928
rect 20409 24968 20495 24991
rect 20577 24968 20663 24991
rect 20409 24928 20434 24968
rect 20434 24928 20474 24968
rect 20474 24928 20495 24968
rect 20577 24928 20598 24968
rect 20598 24928 20638 24968
rect 20638 24928 20663 24968
rect 20409 24905 20495 24928
rect 20577 24905 20663 24928
rect 24409 24968 24495 24991
rect 24577 24968 24663 24991
rect 24409 24928 24434 24968
rect 24434 24928 24474 24968
rect 24474 24928 24495 24968
rect 24577 24928 24598 24968
rect 24598 24928 24638 24968
rect 24638 24928 24663 24968
rect 24409 24905 24495 24928
rect 24577 24905 24663 24928
rect 28409 24968 28495 24991
rect 28577 24968 28663 24991
rect 28409 24928 28434 24968
rect 28434 24928 28474 24968
rect 28474 24928 28495 24968
rect 28577 24928 28598 24968
rect 28598 24928 28638 24968
rect 28638 24928 28663 24968
rect 28409 24905 28495 24928
rect 28577 24905 28663 24928
rect 32409 24968 32495 24991
rect 32577 24968 32663 24991
rect 32409 24928 32434 24968
rect 32434 24928 32474 24968
rect 32474 24928 32495 24968
rect 32577 24928 32598 24968
rect 32598 24928 32638 24968
rect 32638 24928 32663 24968
rect 32409 24905 32495 24928
rect 32577 24905 32663 24928
rect 36409 24968 36495 24991
rect 36577 24968 36663 24991
rect 36409 24928 36434 24968
rect 36434 24928 36474 24968
rect 36474 24928 36495 24968
rect 36577 24928 36598 24968
rect 36598 24928 36638 24968
rect 36638 24928 36663 24968
rect 36409 24905 36495 24928
rect 36577 24905 36663 24928
rect 40409 24968 40495 24991
rect 40577 24968 40663 24991
rect 40409 24928 40434 24968
rect 40434 24928 40474 24968
rect 40474 24928 40495 24968
rect 40577 24928 40598 24968
rect 40598 24928 40638 24968
rect 40638 24928 40663 24968
rect 40409 24905 40495 24928
rect 40577 24905 40663 24928
rect 44409 24968 44495 24991
rect 44577 24968 44663 24991
rect 44409 24928 44434 24968
rect 44434 24928 44474 24968
rect 44474 24928 44495 24968
rect 44577 24928 44598 24968
rect 44598 24928 44638 24968
rect 44638 24928 44663 24968
rect 44409 24905 44495 24928
rect 44577 24905 44663 24928
rect 48409 24968 48495 24991
rect 48577 24968 48663 24991
rect 48409 24928 48434 24968
rect 48434 24928 48474 24968
rect 48474 24928 48495 24968
rect 48577 24928 48598 24968
rect 48598 24928 48638 24968
rect 48638 24928 48663 24968
rect 48409 24905 48495 24928
rect 48577 24905 48663 24928
rect 52409 24968 52495 24991
rect 52577 24968 52663 24991
rect 52409 24928 52434 24968
rect 52434 24928 52474 24968
rect 52474 24928 52495 24968
rect 52577 24928 52598 24968
rect 52598 24928 52638 24968
rect 52638 24928 52663 24968
rect 52409 24905 52495 24928
rect 52577 24905 52663 24928
rect 56409 24968 56495 24991
rect 56577 24968 56663 24991
rect 56409 24928 56434 24968
rect 56434 24928 56474 24968
rect 56474 24928 56495 24968
rect 56577 24928 56598 24968
rect 56598 24928 56638 24968
rect 56638 24928 56663 24968
rect 56409 24905 56495 24928
rect 56577 24905 56663 24928
rect 60409 24968 60495 24991
rect 60577 24968 60663 24991
rect 60409 24928 60434 24968
rect 60434 24928 60474 24968
rect 60474 24928 60495 24968
rect 60577 24928 60598 24968
rect 60598 24928 60638 24968
rect 60638 24928 60663 24968
rect 60409 24905 60495 24928
rect 60577 24905 60663 24928
rect 64409 24968 64495 24991
rect 64577 24968 64663 24991
rect 64409 24928 64434 24968
rect 64434 24928 64474 24968
rect 64474 24928 64495 24968
rect 64577 24928 64598 24968
rect 64598 24928 64638 24968
rect 64638 24928 64663 24968
rect 64409 24905 64495 24928
rect 64577 24905 64663 24928
rect 68409 24968 68495 24991
rect 68577 24968 68663 24991
rect 68409 24928 68434 24968
rect 68434 24928 68474 24968
rect 68474 24928 68495 24968
rect 68577 24928 68598 24968
rect 68598 24928 68638 24968
rect 68638 24928 68663 24968
rect 68409 24905 68495 24928
rect 68577 24905 68663 24928
rect 3169 24212 3255 24235
rect 3337 24212 3423 24235
rect 3169 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3255 24212
rect 3337 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3423 24212
rect 3169 24149 3255 24172
rect 3337 24149 3423 24172
rect 7169 24212 7255 24235
rect 7337 24212 7423 24235
rect 7169 24172 7194 24212
rect 7194 24172 7234 24212
rect 7234 24172 7255 24212
rect 7337 24172 7358 24212
rect 7358 24172 7398 24212
rect 7398 24172 7423 24212
rect 7169 24149 7255 24172
rect 7337 24149 7423 24172
rect 11169 24212 11255 24235
rect 11337 24212 11423 24235
rect 11169 24172 11194 24212
rect 11194 24172 11234 24212
rect 11234 24172 11255 24212
rect 11337 24172 11358 24212
rect 11358 24172 11398 24212
rect 11398 24172 11423 24212
rect 11169 24149 11255 24172
rect 11337 24149 11423 24172
rect 15169 24212 15255 24235
rect 15337 24212 15423 24235
rect 15169 24172 15194 24212
rect 15194 24172 15234 24212
rect 15234 24172 15255 24212
rect 15337 24172 15358 24212
rect 15358 24172 15398 24212
rect 15398 24172 15423 24212
rect 15169 24149 15255 24172
rect 15337 24149 15423 24172
rect 19169 24212 19255 24235
rect 19337 24212 19423 24235
rect 19169 24172 19194 24212
rect 19194 24172 19234 24212
rect 19234 24172 19255 24212
rect 19337 24172 19358 24212
rect 19358 24172 19398 24212
rect 19398 24172 19423 24212
rect 19169 24149 19255 24172
rect 19337 24149 19423 24172
rect 23169 24212 23255 24235
rect 23337 24212 23423 24235
rect 23169 24172 23194 24212
rect 23194 24172 23234 24212
rect 23234 24172 23255 24212
rect 23337 24172 23358 24212
rect 23358 24172 23398 24212
rect 23398 24172 23423 24212
rect 23169 24149 23255 24172
rect 23337 24149 23423 24172
rect 27169 24212 27255 24235
rect 27337 24212 27423 24235
rect 27169 24172 27194 24212
rect 27194 24172 27234 24212
rect 27234 24172 27255 24212
rect 27337 24172 27358 24212
rect 27358 24172 27398 24212
rect 27398 24172 27423 24212
rect 27169 24149 27255 24172
rect 27337 24149 27423 24172
rect 31169 24212 31255 24235
rect 31337 24212 31423 24235
rect 31169 24172 31194 24212
rect 31194 24172 31234 24212
rect 31234 24172 31255 24212
rect 31337 24172 31358 24212
rect 31358 24172 31398 24212
rect 31398 24172 31423 24212
rect 31169 24149 31255 24172
rect 31337 24149 31423 24172
rect 35169 24212 35255 24235
rect 35337 24212 35423 24235
rect 35169 24172 35194 24212
rect 35194 24172 35234 24212
rect 35234 24172 35255 24212
rect 35337 24172 35358 24212
rect 35358 24172 35398 24212
rect 35398 24172 35423 24212
rect 35169 24149 35255 24172
rect 35337 24149 35423 24172
rect 39169 24212 39255 24235
rect 39337 24212 39423 24235
rect 39169 24172 39194 24212
rect 39194 24172 39234 24212
rect 39234 24172 39255 24212
rect 39337 24172 39358 24212
rect 39358 24172 39398 24212
rect 39398 24172 39423 24212
rect 39169 24149 39255 24172
rect 39337 24149 39423 24172
rect 43169 24212 43255 24235
rect 43337 24212 43423 24235
rect 43169 24172 43194 24212
rect 43194 24172 43234 24212
rect 43234 24172 43255 24212
rect 43337 24172 43358 24212
rect 43358 24172 43398 24212
rect 43398 24172 43423 24212
rect 43169 24149 43255 24172
rect 43337 24149 43423 24172
rect 47169 24212 47255 24235
rect 47337 24212 47423 24235
rect 47169 24172 47194 24212
rect 47194 24172 47234 24212
rect 47234 24172 47255 24212
rect 47337 24172 47358 24212
rect 47358 24172 47398 24212
rect 47398 24172 47423 24212
rect 47169 24149 47255 24172
rect 47337 24149 47423 24172
rect 51169 24212 51255 24235
rect 51337 24212 51423 24235
rect 51169 24172 51194 24212
rect 51194 24172 51234 24212
rect 51234 24172 51255 24212
rect 51337 24172 51358 24212
rect 51358 24172 51398 24212
rect 51398 24172 51423 24212
rect 51169 24149 51255 24172
rect 51337 24149 51423 24172
rect 55169 24212 55255 24235
rect 55337 24212 55423 24235
rect 55169 24172 55194 24212
rect 55194 24172 55234 24212
rect 55234 24172 55255 24212
rect 55337 24172 55358 24212
rect 55358 24172 55398 24212
rect 55398 24172 55423 24212
rect 55169 24149 55255 24172
rect 55337 24149 55423 24172
rect 59169 24212 59255 24235
rect 59337 24212 59423 24235
rect 59169 24172 59194 24212
rect 59194 24172 59234 24212
rect 59234 24172 59255 24212
rect 59337 24172 59358 24212
rect 59358 24172 59398 24212
rect 59398 24172 59423 24212
rect 59169 24149 59255 24172
rect 59337 24149 59423 24172
rect 63169 24212 63255 24235
rect 63337 24212 63423 24235
rect 63169 24172 63194 24212
rect 63194 24172 63234 24212
rect 63234 24172 63255 24212
rect 63337 24172 63358 24212
rect 63358 24172 63398 24212
rect 63398 24172 63423 24212
rect 63169 24149 63255 24172
rect 63337 24149 63423 24172
rect 67169 24212 67255 24235
rect 67337 24212 67423 24235
rect 67169 24172 67194 24212
rect 67194 24172 67234 24212
rect 67234 24172 67255 24212
rect 67337 24172 67358 24212
rect 67358 24172 67398 24212
rect 67398 24172 67423 24212
rect 67169 24149 67255 24172
rect 67337 24149 67423 24172
rect 4409 23456 4495 23479
rect 4577 23456 4663 23479
rect 4409 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4495 23456
rect 4577 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4663 23456
rect 4409 23393 4495 23416
rect 4577 23393 4663 23416
rect 8409 23456 8495 23479
rect 8577 23456 8663 23479
rect 8409 23416 8434 23456
rect 8434 23416 8474 23456
rect 8474 23416 8495 23456
rect 8577 23416 8598 23456
rect 8598 23416 8638 23456
rect 8638 23416 8663 23456
rect 8409 23393 8495 23416
rect 8577 23393 8663 23416
rect 12409 23456 12495 23479
rect 12577 23456 12663 23479
rect 12409 23416 12434 23456
rect 12434 23416 12474 23456
rect 12474 23416 12495 23456
rect 12577 23416 12598 23456
rect 12598 23416 12638 23456
rect 12638 23416 12663 23456
rect 12409 23393 12495 23416
rect 12577 23393 12663 23416
rect 16409 23456 16495 23479
rect 16577 23456 16663 23479
rect 16409 23416 16434 23456
rect 16434 23416 16474 23456
rect 16474 23416 16495 23456
rect 16577 23416 16598 23456
rect 16598 23416 16638 23456
rect 16638 23416 16663 23456
rect 16409 23393 16495 23416
rect 16577 23393 16663 23416
rect 20409 23456 20495 23479
rect 20577 23456 20663 23479
rect 20409 23416 20434 23456
rect 20434 23416 20474 23456
rect 20474 23416 20495 23456
rect 20577 23416 20598 23456
rect 20598 23416 20638 23456
rect 20638 23416 20663 23456
rect 20409 23393 20495 23416
rect 20577 23393 20663 23416
rect 24409 23456 24495 23479
rect 24577 23456 24663 23479
rect 24409 23416 24434 23456
rect 24434 23416 24474 23456
rect 24474 23416 24495 23456
rect 24577 23416 24598 23456
rect 24598 23416 24638 23456
rect 24638 23416 24663 23456
rect 24409 23393 24495 23416
rect 24577 23393 24663 23416
rect 28409 23456 28495 23479
rect 28577 23456 28663 23479
rect 28409 23416 28434 23456
rect 28434 23416 28474 23456
rect 28474 23416 28495 23456
rect 28577 23416 28598 23456
rect 28598 23416 28638 23456
rect 28638 23416 28663 23456
rect 28409 23393 28495 23416
rect 28577 23393 28663 23416
rect 32409 23456 32495 23479
rect 32577 23456 32663 23479
rect 32409 23416 32434 23456
rect 32434 23416 32474 23456
rect 32474 23416 32495 23456
rect 32577 23416 32598 23456
rect 32598 23416 32638 23456
rect 32638 23416 32663 23456
rect 32409 23393 32495 23416
rect 32577 23393 32663 23416
rect 36409 23456 36495 23479
rect 36577 23456 36663 23479
rect 36409 23416 36434 23456
rect 36434 23416 36474 23456
rect 36474 23416 36495 23456
rect 36577 23416 36598 23456
rect 36598 23416 36638 23456
rect 36638 23416 36663 23456
rect 36409 23393 36495 23416
rect 36577 23393 36663 23416
rect 40409 23456 40495 23479
rect 40577 23456 40663 23479
rect 40409 23416 40434 23456
rect 40434 23416 40474 23456
rect 40474 23416 40495 23456
rect 40577 23416 40598 23456
rect 40598 23416 40638 23456
rect 40638 23416 40663 23456
rect 40409 23393 40495 23416
rect 40577 23393 40663 23416
rect 44409 23456 44495 23479
rect 44577 23456 44663 23479
rect 44409 23416 44434 23456
rect 44434 23416 44474 23456
rect 44474 23416 44495 23456
rect 44577 23416 44598 23456
rect 44598 23416 44638 23456
rect 44638 23416 44663 23456
rect 44409 23393 44495 23416
rect 44577 23393 44663 23416
rect 48409 23456 48495 23479
rect 48577 23456 48663 23479
rect 48409 23416 48434 23456
rect 48434 23416 48474 23456
rect 48474 23416 48495 23456
rect 48577 23416 48598 23456
rect 48598 23416 48638 23456
rect 48638 23416 48663 23456
rect 48409 23393 48495 23416
rect 48577 23393 48663 23416
rect 52409 23456 52495 23479
rect 52577 23456 52663 23479
rect 52409 23416 52434 23456
rect 52434 23416 52474 23456
rect 52474 23416 52495 23456
rect 52577 23416 52598 23456
rect 52598 23416 52638 23456
rect 52638 23416 52663 23456
rect 52409 23393 52495 23416
rect 52577 23393 52663 23416
rect 56409 23456 56495 23479
rect 56577 23456 56663 23479
rect 56409 23416 56434 23456
rect 56434 23416 56474 23456
rect 56474 23416 56495 23456
rect 56577 23416 56598 23456
rect 56598 23416 56638 23456
rect 56638 23416 56663 23456
rect 56409 23393 56495 23416
rect 56577 23393 56663 23416
rect 60409 23456 60495 23479
rect 60577 23456 60663 23479
rect 60409 23416 60434 23456
rect 60434 23416 60474 23456
rect 60474 23416 60495 23456
rect 60577 23416 60598 23456
rect 60598 23416 60638 23456
rect 60638 23416 60663 23456
rect 60409 23393 60495 23416
rect 60577 23393 60663 23416
rect 64409 23456 64495 23479
rect 64577 23456 64663 23479
rect 64409 23416 64434 23456
rect 64434 23416 64474 23456
rect 64474 23416 64495 23456
rect 64577 23416 64598 23456
rect 64598 23416 64638 23456
rect 64638 23416 64663 23456
rect 64409 23393 64495 23416
rect 64577 23393 64663 23416
rect 68409 23456 68495 23479
rect 68577 23456 68663 23479
rect 68409 23416 68434 23456
rect 68434 23416 68474 23456
rect 68474 23416 68495 23456
rect 68577 23416 68598 23456
rect 68598 23416 68638 23456
rect 68638 23416 68663 23456
rect 68409 23393 68495 23416
rect 68577 23393 68663 23416
rect 72409 23456 72495 23479
rect 72577 23456 72663 23479
rect 72409 23416 72434 23456
rect 72434 23416 72474 23456
rect 72474 23416 72495 23456
rect 72577 23416 72598 23456
rect 72598 23416 72638 23456
rect 72638 23416 72663 23456
rect 72409 23393 72495 23416
rect 72577 23393 72663 23416
rect 76409 23456 76495 23479
rect 76577 23456 76663 23479
rect 76409 23416 76434 23456
rect 76434 23416 76474 23456
rect 76474 23416 76495 23456
rect 76577 23416 76598 23456
rect 76598 23416 76638 23456
rect 76638 23416 76663 23456
rect 76409 23393 76495 23416
rect 76577 23393 76663 23416
rect 80409 23456 80495 23479
rect 80577 23456 80663 23479
rect 80409 23416 80434 23456
rect 80434 23416 80474 23456
rect 80474 23416 80495 23456
rect 80577 23416 80598 23456
rect 80598 23416 80638 23456
rect 80638 23416 80663 23456
rect 80409 23393 80495 23416
rect 80577 23393 80663 23416
rect 84409 23456 84495 23479
rect 84577 23456 84663 23479
rect 84409 23416 84434 23456
rect 84434 23416 84474 23456
rect 84474 23416 84495 23456
rect 84577 23416 84598 23456
rect 84598 23416 84638 23456
rect 84638 23416 84663 23456
rect 84409 23393 84495 23416
rect 84577 23393 84663 23416
rect 88409 23456 88495 23479
rect 88577 23456 88663 23479
rect 88409 23416 88434 23456
rect 88434 23416 88474 23456
rect 88474 23416 88495 23456
rect 88577 23416 88598 23456
rect 88598 23416 88638 23456
rect 88638 23416 88663 23456
rect 88409 23393 88495 23416
rect 88577 23393 88663 23416
rect 92409 23456 92495 23479
rect 92577 23456 92663 23479
rect 92409 23416 92434 23456
rect 92434 23416 92474 23456
rect 92474 23416 92495 23456
rect 92577 23416 92598 23456
rect 92598 23416 92638 23456
rect 92638 23416 92663 23456
rect 92409 23393 92495 23416
rect 92577 23393 92663 23416
rect 96409 23456 96495 23479
rect 96577 23456 96663 23479
rect 96409 23416 96434 23456
rect 96434 23416 96474 23456
rect 96474 23416 96495 23456
rect 96577 23416 96598 23456
rect 96598 23416 96638 23456
rect 96638 23416 96663 23456
rect 96409 23393 96495 23416
rect 96577 23393 96663 23416
rect 86469 23057 86555 23143
rect 3169 22700 3255 22723
rect 3337 22700 3423 22723
rect 3169 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3255 22700
rect 3337 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3423 22700
rect 3169 22637 3255 22660
rect 3337 22637 3423 22660
rect 7169 22700 7255 22723
rect 7337 22700 7423 22723
rect 7169 22660 7194 22700
rect 7194 22660 7234 22700
rect 7234 22660 7255 22700
rect 7337 22660 7358 22700
rect 7358 22660 7398 22700
rect 7398 22660 7423 22700
rect 7169 22637 7255 22660
rect 7337 22637 7423 22660
rect 11169 22700 11255 22723
rect 11337 22700 11423 22723
rect 11169 22660 11194 22700
rect 11194 22660 11234 22700
rect 11234 22660 11255 22700
rect 11337 22660 11358 22700
rect 11358 22660 11398 22700
rect 11398 22660 11423 22700
rect 11169 22637 11255 22660
rect 11337 22637 11423 22660
rect 15169 22700 15255 22723
rect 15337 22700 15423 22723
rect 15169 22660 15194 22700
rect 15194 22660 15234 22700
rect 15234 22660 15255 22700
rect 15337 22660 15358 22700
rect 15358 22660 15398 22700
rect 15398 22660 15423 22700
rect 15169 22637 15255 22660
rect 15337 22637 15423 22660
rect 19169 22700 19255 22723
rect 19337 22700 19423 22723
rect 19169 22660 19194 22700
rect 19194 22660 19234 22700
rect 19234 22660 19255 22700
rect 19337 22660 19358 22700
rect 19358 22660 19398 22700
rect 19398 22660 19423 22700
rect 19169 22637 19255 22660
rect 19337 22637 19423 22660
rect 23169 22700 23255 22723
rect 23337 22700 23423 22723
rect 23169 22660 23194 22700
rect 23194 22660 23234 22700
rect 23234 22660 23255 22700
rect 23337 22660 23358 22700
rect 23358 22660 23398 22700
rect 23398 22660 23423 22700
rect 23169 22637 23255 22660
rect 23337 22637 23423 22660
rect 27169 22700 27255 22723
rect 27337 22700 27423 22723
rect 27169 22660 27194 22700
rect 27194 22660 27234 22700
rect 27234 22660 27255 22700
rect 27337 22660 27358 22700
rect 27358 22660 27398 22700
rect 27398 22660 27423 22700
rect 27169 22637 27255 22660
rect 27337 22637 27423 22660
rect 31169 22700 31255 22723
rect 31337 22700 31423 22723
rect 31169 22660 31194 22700
rect 31194 22660 31234 22700
rect 31234 22660 31255 22700
rect 31337 22660 31358 22700
rect 31358 22660 31398 22700
rect 31398 22660 31423 22700
rect 31169 22637 31255 22660
rect 31337 22637 31423 22660
rect 35169 22700 35255 22723
rect 35337 22700 35423 22723
rect 35169 22660 35194 22700
rect 35194 22660 35234 22700
rect 35234 22660 35255 22700
rect 35337 22660 35358 22700
rect 35358 22660 35398 22700
rect 35398 22660 35423 22700
rect 35169 22637 35255 22660
rect 35337 22637 35423 22660
rect 39169 22700 39255 22723
rect 39337 22700 39423 22723
rect 39169 22660 39194 22700
rect 39194 22660 39234 22700
rect 39234 22660 39255 22700
rect 39337 22660 39358 22700
rect 39358 22660 39398 22700
rect 39398 22660 39423 22700
rect 39169 22637 39255 22660
rect 39337 22637 39423 22660
rect 43169 22700 43255 22723
rect 43337 22700 43423 22723
rect 43169 22660 43194 22700
rect 43194 22660 43234 22700
rect 43234 22660 43255 22700
rect 43337 22660 43358 22700
rect 43358 22660 43398 22700
rect 43398 22660 43423 22700
rect 43169 22637 43255 22660
rect 43337 22637 43423 22660
rect 47169 22700 47255 22723
rect 47337 22700 47423 22723
rect 47169 22660 47194 22700
rect 47194 22660 47234 22700
rect 47234 22660 47255 22700
rect 47337 22660 47358 22700
rect 47358 22660 47398 22700
rect 47398 22660 47423 22700
rect 47169 22637 47255 22660
rect 47337 22637 47423 22660
rect 51169 22700 51255 22723
rect 51337 22700 51423 22723
rect 51169 22660 51194 22700
rect 51194 22660 51234 22700
rect 51234 22660 51255 22700
rect 51337 22660 51358 22700
rect 51358 22660 51398 22700
rect 51398 22660 51423 22700
rect 51169 22637 51255 22660
rect 51337 22637 51423 22660
rect 55169 22700 55255 22723
rect 55337 22700 55423 22723
rect 55169 22660 55194 22700
rect 55194 22660 55234 22700
rect 55234 22660 55255 22700
rect 55337 22660 55358 22700
rect 55358 22660 55398 22700
rect 55398 22660 55423 22700
rect 55169 22637 55255 22660
rect 55337 22637 55423 22660
rect 59169 22700 59255 22723
rect 59337 22700 59423 22723
rect 59169 22660 59194 22700
rect 59194 22660 59234 22700
rect 59234 22660 59255 22700
rect 59337 22660 59358 22700
rect 59358 22660 59398 22700
rect 59398 22660 59423 22700
rect 59169 22637 59255 22660
rect 59337 22637 59423 22660
rect 63169 22700 63255 22723
rect 63337 22700 63423 22723
rect 63169 22660 63194 22700
rect 63194 22660 63234 22700
rect 63234 22660 63255 22700
rect 63337 22660 63358 22700
rect 63358 22660 63398 22700
rect 63398 22660 63423 22700
rect 63169 22637 63255 22660
rect 63337 22637 63423 22660
rect 67169 22700 67255 22723
rect 67337 22700 67423 22723
rect 67169 22660 67194 22700
rect 67194 22660 67234 22700
rect 67234 22660 67255 22700
rect 67337 22660 67358 22700
rect 67358 22660 67398 22700
rect 67398 22660 67423 22700
rect 67169 22637 67255 22660
rect 67337 22637 67423 22660
rect 71169 22700 71255 22723
rect 71337 22700 71423 22723
rect 71169 22660 71194 22700
rect 71194 22660 71234 22700
rect 71234 22660 71255 22700
rect 71337 22660 71358 22700
rect 71358 22660 71398 22700
rect 71398 22660 71423 22700
rect 71169 22637 71255 22660
rect 71337 22637 71423 22660
rect 75169 22700 75255 22723
rect 75337 22700 75423 22723
rect 75169 22660 75194 22700
rect 75194 22660 75234 22700
rect 75234 22660 75255 22700
rect 75337 22660 75358 22700
rect 75358 22660 75398 22700
rect 75398 22660 75423 22700
rect 75169 22637 75255 22660
rect 75337 22637 75423 22660
rect 79169 22700 79255 22723
rect 79337 22700 79423 22723
rect 79169 22660 79194 22700
rect 79194 22660 79234 22700
rect 79234 22660 79255 22700
rect 79337 22660 79358 22700
rect 79358 22660 79398 22700
rect 79398 22660 79423 22700
rect 79169 22637 79255 22660
rect 79337 22637 79423 22660
rect 83169 22700 83255 22723
rect 83337 22700 83423 22723
rect 83169 22660 83194 22700
rect 83194 22660 83234 22700
rect 83234 22660 83255 22700
rect 83337 22660 83358 22700
rect 83358 22660 83398 22700
rect 83398 22660 83423 22700
rect 83169 22637 83255 22660
rect 83337 22637 83423 22660
rect 87169 22700 87255 22723
rect 87337 22700 87423 22723
rect 87169 22660 87194 22700
rect 87194 22660 87234 22700
rect 87234 22660 87255 22700
rect 87337 22660 87358 22700
rect 87358 22660 87398 22700
rect 87398 22660 87423 22700
rect 87169 22637 87255 22660
rect 87337 22637 87423 22660
rect 91169 22700 91255 22723
rect 91337 22700 91423 22723
rect 91169 22660 91194 22700
rect 91194 22660 91234 22700
rect 91234 22660 91255 22700
rect 91337 22660 91358 22700
rect 91358 22660 91398 22700
rect 91398 22660 91423 22700
rect 91169 22637 91255 22660
rect 91337 22637 91423 22660
rect 95169 22700 95255 22723
rect 95337 22700 95423 22723
rect 95169 22660 95194 22700
rect 95194 22660 95234 22700
rect 95234 22660 95255 22700
rect 95337 22660 95358 22700
rect 95358 22660 95398 22700
rect 95398 22660 95423 22700
rect 95169 22637 95255 22660
rect 95337 22637 95423 22660
rect 99169 22700 99255 22723
rect 99337 22700 99423 22723
rect 99169 22660 99194 22700
rect 99194 22660 99234 22700
rect 99234 22660 99255 22700
rect 99337 22660 99358 22700
rect 99358 22660 99398 22700
rect 99398 22660 99423 22700
rect 99169 22637 99255 22660
rect 99337 22637 99423 22660
rect 4409 21944 4495 21967
rect 4577 21944 4663 21967
rect 4409 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4495 21944
rect 4577 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4663 21944
rect 4409 21881 4495 21904
rect 4577 21881 4663 21904
rect 8409 21944 8495 21967
rect 8577 21944 8663 21967
rect 8409 21904 8434 21944
rect 8434 21904 8474 21944
rect 8474 21904 8495 21944
rect 8577 21904 8598 21944
rect 8598 21904 8638 21944
rect 8638 21904 8663 21944
rect 8409 21881 8495 21904
rect 8577 21881 8663 21904
rect 12409 21944 12495 21967
rect 12577 21944 12663 21967
rect 12409 21904 12434 21944
rect 12434 21904 12474 21944
rect 12474 21904 12495 21944
rect 12577 21904 12598 21944
rect 12598 21904 12638 21944
rect 12638 21904 12663 21944
rect 12409 21881 12495 21904
rect 12577 21881 12663 21904
rect 16409 21944 16495 21967
rect 16577 21944 16663 21967
rect 16409 21904 16434 21944
rect 16434 21904 16474 21944
rect 16474 21904 16495 21944
rect 16577 21904 16598 21944
rect 16598 21904 16638 21944
rect 16638 21904 16663 21944
rect 16409 21881 16495 21904
rect 16577 21881 16663 21904
rect 20409 21944 20495 21967
rect 20577 21944 20663 21967
rect 20409 21904 20434 21944
rect 20434 21904 20474 21944
rect 20474 21904 20495 21944
rect 20577 21904 20598 21944
rect 20598 21904 20638 21944
rect 20638 21904 20663 21944
rect 20409 21881 20495 21904
rect 20577 21881 20663 21904
rect 24409 21944 24495 21967
rect 24577 21944 24663 21967
rect 24409 21904 24434 21944
rect 24434 21904 24474 21944
rect 24474 21904 24495 21944
rect 24577 21904 24598 21944
rect 24598 21904 24638 21944
rect 24638 21904 24663 21944
rect 24409 21881 24495 21904
rect 24577 21881 24663 21904
rect 28409 21944 28495 21967
rect 28577 21944 28663 21967
rect 28409 21904 28434 21944
rect 28434 21904 28474 21944
rect 28474 21904 28495 21944
rect 28577 21904 28598 21944
rect 28598 21904 28638 21944
rect 28638 21904 28663 21944
rect 28409 21881 28495 21904
rect 28577 21881 28663 21904
rect 32409 21944 32495 21967
rect 32577 21944 32663 21967
rect 32409 21904 32434 21944
rect 32434 21904 32474 21944
rect 32474 21904 32495 21944
rect 32577 21904 32598 21944
rect 32598 21904 32638 21944
rect 32638 21904 32663 21944
rect 32409 21881 32495 21904
rect 32577 21881 32663 21904
rect 36409 21944 36495 21967
rect 36577 21944 36663 21967
rect 36409 21904 36434 21944
rect 36434 21904 36474 21944
rect 36474 21904 36495 21944
rect 36577 21904 36598 21944
rect 36598 21904 36638 21944
rect 36638 21904 36663 21944
rect 36409 21881 36495 21904
rect 36577 21881 36663 21904
rect 40409 21944 40495 21967
rect 40577 21944 40663 21967
rect 40409 21904 40434 21944
rect 40434 21904 40474 21944
rect 40474 21904 40495 21944
rect 40577 21904 40598 21944
rect 40598 21904 40638 21944
rect 40638 21904 40663 21944
rect 40409 21881 40495 21904
rect 40577 21881 40663 21904
rect 44409 21944 44495 21967
rect 44577 21944 44663 21967
rect 44409 21904 44434 21944
rect 44434 21904 44474 21944
rect 44474 21904 44495 21944
rect 44577 21904 44598 21944
rect 44598 21904 44638 21944
rect 44638 21904 44663 21944
rect 44409 21881 44495 21904
rect 44577 21881 44663 21904
rect 48409 21944 48495 21967
rect 48577 21944 48663 21967
rect 48409 21904 48434 21944
rect 48434 21904 48474 21944
rect 48474 21904 48495 21944
rect 48577 21904 48598 21944
rect 48598 21904 48638 21944
rect 48638 21904 48663 21944
rect 48409 21881 48495 21904
rect 48577 21881 48663 21904
rect 52409 21944 52495 21967
rect 52577 21944 52663 21967
rect 52409 21904 52434 21944
rect 52434 21904 52474 21944
rect 52474 21904 52495 21944
rect 52577 21904 52598 21944
rect 52598 21904 52638 21944
rect 52638 21904 52663 21944
rect 52409 21881 52495 21904
rect 52577 21881 52663 21904
rect 56409 21944 56495 21967
rect 56577 21944 56663 21967
rect 56409 21904 56434 21944
rect 56434 21904 56474 21944
rect 56474 21904 56495 21944
rect 56577 21904 56598 21944
rect 56598 21904 56638 21944
rect 56638 21904 56663 21944
rect 56409 21881 56495 21904
rect 56577 21881 56663 21904
rect 60409 21944 60495 21967
rect 60577 21944 60663 21967
rect 60409 21904 60434 21944
rect 60434 21904 60474 21944
rect 60474 21904 60495 21944
rect 60577 21904 60598 21944
rect 60598 21904 60638 21944
rect 60638 21904 60663 21944
rect 60409 21881 60495 21904
rect 60577 21881 60663 21904
rect 64409 21944 64495 21967
rect 64577 21944 64663 21967
rect 64409 21904 64434 21944
rect 64434 21904 64474 21944
rect 64474 21904 64495 21944
rect 64577 21904 64598 21944
rect 64598 21904 64638 21944
rect 64638 21904 64663 21944
rect 64409 21881 64495 21904
rect 64577 21881 64663 21904
rect 68409 21944 68495 21967
rect 68577 21944 68663 21967
rect 68409 21904 68434 21944
rect 68434 21904 68474 21944
rect 68474 21904 68495 21944
rect 68577 21904 68598 21944
rect 68598 21904 68638 21944
rect 68638 21904 68663 21944
rect 68409 21881 68495 21904
rect 68577 21881 68663 21904
rect 72409 21944 72495 21967
rect 72577 21944 72663 21967
rect 72409 21904 72434 21944
rect 72434 21904 72474 21944
rect 72474 21904 72495 21944
rect 72577 21904 72598 21944
rect 72598 21904 72638 21944
rect 72638 21904 72663 21944
rect 72409 21881 72495 21904
rect 72577 21881 72663 21904
rect 76409 21944 76495 21967
rect 76577 21944 76663 21967
rect 76409 21904 76434 21944
rect 76434 21904 76474 21944
rect 76474 21904 76495 21944
rect 76577 21904 76598 21944
rect 76598 21904 76638 21944
rect 76638 21904 76663 21944
rect 76409 21881 76495 21904
rect 76577 21881 76663 21904
rect 80409 21944 80495 21967
rect 80577 21944 80663 21967
rect 80409 21904 80434 21944
rect 80434 21904 80474 21944
rect 80474 21904 80495 21944
rect 80577 21904 80598 21944
rect 80598 21904 80638 21944
rect 80638 21904 80663 21944
rect 80409 21881 80495 21904
rect 80577 21881 80663 21904
rect 84409 21944 84495 21967
rect 84577 21944 84663 21967
rect 84409 21904 84434 21944
rect 84434 21904 84474 21944
rect 84474 21904 84495 21944
rect 84577 21904 84598 21944
rect 84598 21904 84638 21944
rect 84638 21904 84663 21944
rect 84409 21881 84495 21904
rect 84577 21881 84663 21904
rect 88409 21944 88495 21967
rect 88577 21944 88663 21967
rect 88409 21904 88434 21944
rect 88434 21904 88474 21944
rect 88474 21904 88495 21944
rect 88577 21904 88598 21944
rect 88598 21904 88638 21944
rect 88638 21904 88663 21944
rect 88409 21881 88495 21904
rect 88577 21881 88663 21904
rect 92409 21944 92495 21967
rect 92577 21944 92663 21967
rect 92409 21904 92434 21944
rect 92434 21904 92474 21944
rect 92474 21904 92495 21944
rect 92577 21904 92598 21944
rect 92598 21904 92638 21944
rect 92638 21904 92663 21944
rect 92409 21881 92495 21904
rect 92577 21881 92663 21904
rect 96409 21944 96495 21967
rect 96577 21944 96663 21967
rect 96409 21904 96434 21944
rect 96434 21904 96474 21944
rect 96474 21904 96495 21944
rect 96577 21904 96598 21944
rect 96598 21904 96638 21944
rect 96638 21904 96663 21944
rect 96409 21881 96495 21904
rect 96577 21881 96663 21904
rect 3169 21188 3255 21211
rect 3337 21188 3423 21211
rect 3169 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3255 21188
rect 3337 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3423 21188
rect 3169 21125 3255 21148
rect 3337 21125 3423 21148
rect 7169 21188 7255 21211
rect 7337 21188 7423 21211
rect 7169 21148 7194 21188
rect 7194 21148 7234 21188
rect 7234 21148 7255 21188
rect 7337 21148 7358 21188
rect 7358 21148 7398 21188
rect 7398 21148 7423 21188
rect 7169 21125 7255 21148
rect 7337 21125 7423 21148
rect 11169 21188 11255 21211
rect 11337 21188 11423 21211
rect 11169 21148 11194 21188
rect 11194 21148 11234 21188
rect 11234 21148 11255 21188
rect 11337 21148 11358 21188
rect 11358 21148 11398 21188
rect 11398 21148 11423 21188
rect 11169 21125 11255 21148
rect 11337 21125 11423 21148
rect 15169 21188 15255 21211
rect 15337 21188 15423 21211
rect 15169 21148 15194 21188
rect 15194 21148 15234 21188
rect 15234 21148 15255 21188
rect 15337 21148 15358 21188
rect 15358 21148 15398 21188
rect 15398 21148 15423 21188
rect 15169 21125 15255 21148
rect 15337 21125 15423 21148
rect 19169 21188 19255 21211
rect 19337 21188 19423 21211
rect 19169 21148 19194 21188
rect 19194 21148 19234 21188
rect 19234 21148 19255 21188
rect 19337 21148 19358 21188
rect 19358 21148 19398 21188
rect 19398 21148 19423 21188
rect 19169 21125 19255 21148
rect 19337 21125 19423 21148
rect 23169 21188 23255 21211
rect 23337 21188 23423 21211
rect 23169 21148 23194 21188
rect 23194 21148 23234 21188
rect 23234 21148 23255 21188
rect 23337 21148 23358 21188
rect 23358 21148 23398 21188
rect 23398 21148 23423 21188
rect 23169 21125 23255 21148
rect 23337 21125 23423 21148
rect 27169 21188 27255 21211
rect 27337 21188 27423 21211
rect 27169 21148 27194 21188
rect 27194 21148 27234 21188
rect 27234 21148 27255 21188
rect 27337 21148 27358 21188
rect 27358 21148 27398 21188
rect 27398 21148 27423 21188
rect 27169 21125 27255 21148
rect 27337 21125 27423 21148
rect 31169 21188 31255 21211
rect 31337 21188 31423 21211
rect 31169 21148 31194 21188
rect 31194 21148 31234 21188
rect 31234 21148 31255 21188
rect 31337 21148 31358 21188
rect 31358 21148 31398 21188
rect 31398 21148 31423 21188
rect 31169 21125 31255 21148
rect 31337 21125 31423 21148
rect 35169 21188 35255 21211
rect 35337 21188 35423 21211
rect 35169 21148 35194 21188
rect 35194 21148 35234 21188
rect 35234 21148 35255 21188
rect 35337 21148 35358 21188
rect 35358 21148 35398 21188
rect 35398 21148 35423 21188
rect 35169 21125 35255 21148
rect 35337 21125 35423 21148
rect 39169 21188 39255 21211
rect 39337 21188 39423 21211
rect 39169 21148 39194 21188
rect 39194 21148 39234 21188
rect 39234 21148 39255 21188
rect 39337 21148 39358 21188
rect 39358 21148 39398 21188
rect 39398 21148 39423 21188
rect 39169 21125 39255 21148
rect 39337 21125 39423 21148
rect 43169 21188 43255 21211
rect 43337 21188 43423 21211
rect 43169 21148 43194 21188
rect 43194 21148 43234 21188
rect 43234 21148 43255 21188
rect 43337 21148 43358 21188
rect 43358 21148 43398 21188
rect 43398 21148 43423 21188
rect 43169 21125 43255 21148
rect 43337 21125 43423 21148
rect 47169 21188 47255 21211
rect 47337 21188 47423 21211
rect 47169 21148 47194 21188
rect 47194 21148 47234 21188
rect 47234 21148 47255 21188
rect 47337 21148 47358 21188
rect 47358 21148 47398 21188
rect 47398 21148 47423 21188
rect 47169 21125 47255 21148
rect 47337 21125 47423 21148
rect 51169 21188 51255 21211
rect 51337 21188 51423 21211
rect 51169 21148 51194 21188
rect 51194 21148 51234 21188
rect 51234 21148 51255 21188
rect 51337 21148 51358 21188
rect 51358 21148 51398 21188
rect 51398 21148 51423 21188
rect 51169 21125 51255 21148
rect 51337 21125 51423 21148
rect 55169 21188 55255 21211
rect 55337 21188 55423 21211
rect 55169 21148 55194 21188
rect 55194 21148 55234 21188
rect 55234 21148 55255 21188
rect 55337 21148 55358 21188
rect 55358 21148 55398 21188
rect 55398 21148 55423 21188
rect 55169 21125 55255 21148
rect 55337 21125 55423 21148
rect 59169 21188 59255 21211
rect 59337 21188 59423 21211
rect 59169 21148 59194 21188
rect 59194 21148 59234 21188
rect 59234 21148 59255 21188
rect 59337 21148 59358 21188
rect 59358 21148 59398 21188
rect 59398 21148 59423 21188
rect 59169 21125 59255 21148
rect 59337 21125 59423 21148
rect 63169 21188 63255 21211
rect 63337 21188 63423 21211
rect 63169 21148 63194 21188
rect 63194 21148 63234 21188
rect 63234 21148 63255 21188
rect 63337 21148 63358 21188
rect 63358 21148 63398 21188
rect 63398 21148 63423 21188
rect 63169 21125 63255 21148
rect 63337 21125 63423 21148
rect 67169 21188 67255 21211
rect 67337 21188 67423 21211
rect 67169 21148 67194 21188
rect 67194 21148 67234 21188
rect 67234 21148 67255 21188
rect 67337 21148 67358 21188
rect 67358 21148 67398 21188
rect 67398 21148 67423 21188
rect 67169 21125 67255 21148
rect 67337 21125 67423 21148
rect 71169 21188 71255 21211
rect 71337 21188 71423 21211
rect 71169 21148 71194 21188
rect 71194 21148 71234 21188
rect 71234 21148 71255 21188
rect 71337 21148 71358 21188
rect 71358 21148 71398 21188
rect 71398 21148 71423 21188
rect 71169 21125 71255 21148
rect 71337 21125 71423 21148
rect 75169 21188 75255 21211
rect 75337 21188 75423 21211
rect 75169 21148 75194 21188
rect 75194 21148 75234 21188
rect 75234 21148 75255 21188
rect 75337 21148 75358 21188
rect 75358 21148 75398 21188
rect 75398 21148 75423 21188
rect 75169 21125 75255 21148
rect 75337 21125 75423 21148
rect 79169 21188 79255 21211
rect 79337 21188 79423 21211
rect 79169 21148 79194 21188
rect 79194 21148 79234 21188
rect 79234 21148 79255 21188
rect 79337 21148 79358 21188
rect 79358 21148 79398 21188
rect 79398 21148 79423 21188
rect 79169 21125 79255 21148
rect 79337 21125 79423 21148
rect 83169 21188 83255 21211
rect 83337 21188 83423 21211
rect 83169 21148 83194 21188
rect 83194 21148 83234 21188
rect 83234 21148 83255 21188
rect 83337 21148 83358 21188
rect 83358 21148 83398 21188
rect 83398 21148 83423 21188
rect 83169 21125 83255 21148
rect 83337 21125 83423 21148
rect 87169 21188 87255 21211
rect 87337 21188 87423 21211
rect 87169 21148 87194 21188
rect 87194 21148 87234 21188
rect 87234 21148 87255 21188
rect 87337 21148 87358 21188
rect 87358 21148 87398 21188
rect 87398 21148 87423 21188
rect 87169 21125 87255 21148
rect 87337 21125 87423 21148
rect 91169 21188 91255 21211
rect 91337 21188 91423 21211
rect 91169 21148 91194 21188
rect 91194 21148 91234 21188
rect 91234 21148 91255 21188
rect 91337 21148 91358 21188
rect 91358 21148 91398 21188
rect 91398 21148 91423 21188
rect 91169 21125 91255 21148
rect 91337 21125 91423 21148
rect 95169 21188 95255 21211
rect 95337 21188 95423 21211
rect 95169 21148 95194 21188
rect 95194 21148 95234 21188
rect 95234 21148 95255 21188
rect 95337 21148 95358 21188
rect 95358 21148 95398 21188
rect 95398 21148 95423 21188
rect 95169 21125 95255 21148
rect 95337 21125 95423 21148
rect 99169 21188 99255 21211
rect 99337 21188 99423 21211
rect 99169 21148 99194 21188
rect 99194 21148 99234 21188
rect 99234 21148 99255 21188
rect 99337 21148 99358 21188
rect 99358 21148 99398 21188
rect 99398 21148 99423 21188
rect 99169 21125 99255 21148
rect 99337 21125 99423 21148
rect 4409 20432 4495 20455
rect 4577 20432 4663 20455
rect 4409 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4495 20432
rect 4577 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4663 20432
rect 4409 20369 4495 20392
rect 4577 20369 4663 20392
rect 8409 20432 8495 20455
rect 8577 20432 8663 20455
rect 8409 20392 8434 20432
rect 8434 20392 8474 20432
rect 8474 20392 8495 20432
rect 8577 20392 8598 20432
rect 8598 20392 8638 20432
rect 8638 20392 8663 20432
rect 8409 20369 8495 20392
rect 8577 20369 8663 20392
rect 12409 20432 12495 20455
rect 12577 20432 12663 20455
rect 12409 20392 12434 20432
rect 12434 20392 12474 20432
rect 12474 20392 12495 20432
rect 12577 20392 12598 20432
rect 12598 20392 12638 20432
rect 12638 20392 12663 20432
rect 12409 20369 12495 20392
rect 12577 20369 12663 20392
rect 16409 20432 16495 20455
rect 16577 20432 16663 20455
rect 16409 20392 16434 20432
rect 16434 20392 16474 20432
rect 16474 20392 16495 20432
rect 16577 20392 16598 20432
rect 16598 20392 16638 20432
rect 16638 20392 16663 20432
rect 16409 20369 16495 20392
rect 16577 20369 16663 20392
rect 20409 20432 20495 20455
rect 20577 20432 20663 20455
rect 20409 20392 20434 20432
rect 20434 20392 20474 20432
rect 20474 20392 20495 20432
rect 20577 20392 20598 20432
rect 20598 20392 20638 20432
rect 20638 20392 20663 20432
rect 20409 20369 20495 20392
rect 20577 20369 20663 20392
rect 24409 20432 24495 20455
rect 24577 20432 24663 20455
rect 24409 20392 24434 20432
rect 24434 20392 24474 20432
rect 24474 20392 24495 20432
rect 24577 20392 24598 20432
rect 24598 20392 24638 20432
rect 24638 20392 24663 20432
rect 24409 20369 24495 20392
rect 24577 20369 24663 20392
rect 28409 20432 28495 20455
rect 28577 20432 28663 20455
rect 28409 20392 28434 20432
rect 28434 20392 28474 20432
rect 28474 20392 28495 20432
rect 28577 20392 28598 20432
rect 28598 20392 28638 20432
rect 28638 20392 28663 20432
rect 28409 20369 28495 20392
rect 28577 20369 28663 20392
rect 32409 20432 32495 20455
rect 32577 20432 32663 20455
rect 32409 20392 32434 20432
rect 32434 20392 32474 20432
rect 32474 20392 32495 20432
rect 32577 20392 32598 20432
rect 32598 20392 32638 20432
rect 32638 20392 32663 20432
rect 32409 20369 32495 20392
rect 32577 20369 32663 20392
rect 36409 20432 36495 20455
rect 36577 20432 36663 20455
rect 36409 20392 36434 20432
rect 36434 20392 36474 20432
rect 36474 20392 36495 20432
rect 36577 20392 36598 20432
rect 36598 20392 36638 20432
rect 36638 20392 36663 20432
rect 36409 20369 36495 20392
rect 36577 20369 36663 20392
rect 40409 20432 40495 20455
rect 40577 20432 40663 20455
rect 40409 20392 40434 20432
rect 40434 20392 40474 20432
rect 40474 20392 40495 20432
rect 40577 20392 40598 20432
rect 40598 20392 40638 20432
rect 40638 20392 40663 20432
rect 40409 20369 40495 20392
rect 40577 20369 40663 20392
rect 44409 20432 44495 20455
rect 44577 20432 44663 20455
rect 44409 20392 44434 20432
rect 44434 20392 44474 20432
rect 44474 20392 44495 20432
rect 44577 20392 44598 20432
rect 44598 20392 44638 20432
rect 44638 20392 44663 20432
rect 44409 20369 44495 20392
rect 44577 20369 44663 20392
rect 48409 20432 48495 20455
rect 48577 20432 48663 20455
rect 48409 20392 48434 20432
rect 48434 20392 48474 20432
rect 48474 20392 48495 20432
rect 48577 20392 48598 20432
rect 48598 20392 48638 20432
rect 48638 20392 48663 20432
rect 48409 20369 48495 20392
rect 48577 20369 48663 20392
rect 52409 20432 52495 20455
rect 52577 20432 52663 20455
rect 52409 20392 52434 20432
rect 52434 20392 52474 20432
rect 52474 20392 52495 20432
rect 52577 20392 52598 20432
rect 52598 20392 52638 20432
rect 52638 20392 52663 20432
rect 52409 20369 52495 20392
rect 52577 20369 52663 20392
rect 56409 20432 56495 20455
rect 56577 20432 56663 20455
rect 56409 20392 56434 20432
rect 56434 20392 56474 20432
rect 56474 20392 56495 20432
rect 56577 20392 56598 20432
rect 56598 20392 56638 20432
rect 56638 20392 56663 20432
rect 56409 20369 56495 20392
rect 56577 20369 56663 20392
rect 60409 20432 60495 20455
rect 60577 20432 60663 20455
rect 60409 20392 60434 20432
rect 60434 20392 60474 20432
rect 60474 20392 60495 20432
rect 60577 20392 60598 20432
rect 60598 20392 60638 20432
rect 60638 20392 60663 20432
rect 60409 20369 60495 20392
rect 60577 20369 60663 20392
rect 64409 20432 64495 20455
rect 64577 20432 64663 20455
rect 64409 20392 64434 20432
rect 64434 20392 64474 20432
rect 64474 20392 64495 20432
rect 64577 20392 64598 20432
rect 64598 20392 64638 20432
rect 64638 20392 64663 20432
rect 64409 20369 64495 20392
rect 64577 20369 64663 20392
rect 68409 20432 68495 20455
rect 68577 20432 68663 20455
rect 68409 20392 68434 20432
rect 68434 20392 68474 20432
rect 68474 20392 68495 20432
rect 68577 20392 68598 20432
rect 68598 20392 68638 20432
rect 68638 20392 68663 20432
rect 68409 20369 68495 20392
rect 68577 20369 68663 20392
rect 72409 20432 72495 20455
rect 72577 20432 72663 20455
rect 72409 20392 72434 20432
rect 72434 20392 72474 20432
rect 72474 20392 72495 20432
rect 72577 20392 72598 20432
rect 72598 20392 72638 20432
rect 72638 20392 72663 20432
rect 72409 20369 72495 20392
rect 72577 20369 72663 20392
rect 76409 20432 76495 20455
rect 76577 20432 76663 20455
rect 76409 20392 76434 20432
rect 76434 20392 76474 20432
rect 76474 20392 76495 20432
rect 76577 20392 76598 20432
rect 76598 20392 76638 20432
rect 76638 20392 76663 20432
rect 76409 20369 76495 20392
rect 76577 20369 76663 20392
rect 80409 20432 80495 20455
rect 80577 20432 80663 20455
rect 80409 20392 80434 20432
rect 80434 20392 80474 20432
rect 80474 20392 80495 20432
rect 80577 20392 80598 20432
rect 80598 20392 80638 20432
rect 80638 20392 80663 20432
rect 80409 20369 80495 20392
rect 80577 20369 80663 20392
rect 84409 20432 84495 20455
rect 84577 20432 84663 20455
rect 84409 20392 84434 20432
rect 84434 20392 84474 20432
rect 84474 20392 84495 20432
rect 84577 20392 84598 20432
rect 84598 20392 84638 20432
rect 84638 20392 84663 20432
rect 84409 20369 84495 20392
rect 84577 20369 84663 20392
rect 88409 20432 88495 20455
rect 88577 20432 88663 20455
rect 88409 20392 88434 20432
rect 88434 20392 88474 20432
rect 88474 20392 88495 20432
rect 88577 20392 88598 20432
rect 88598 20392 88638 20432
rect 88638 20392 88663 20432
rect 88409 20369 88495 20392
rect 88577 20369 88663 20392
rect 92409 20432 92495 20455
rect 92577 20432 92663 20455
rect 92409 20392 92434 20432
rect 92434 20392 92474 20432
rect 92474 20392 92495 20432
rect 92577 20392 92598 20432
rect 92598 20392 92638 20432
rect 92638 20392 92663 20432
rect 92409 20369 92495 20392
rect 92577 20369 92663 20392
rect 96409 20432 96495 20455
rect 96577 20432 96663 20455
rect 96409 20392 96434 20432
rect 96434 20392 96474 20432
rect 96474 20392 96495 20432
rect 96577 20392 96598 20432
rect 96598 20392 96638 20432
rect 96638 20392 96663 20432
rect 96409 20369 96495 20392
rect 96577 20369 96663 20392
rect 3169 19676 3255 19699
rect 3337 19676 3423 19699
rect 3169 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3255 19676
rect 3337 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3423 19676
rect 3169 19613 3255 19636
rect 3337 19613 3423 19636
rect 7169 19676 7255 19699
rect 7337 19676 7423 19699
rect 7169 19636 7194 19676
rect 7194 19636 7234 19676
rect 7234 19636 7255 19676
rect 7337 19636 7358 19676
rect 7358 19636 7398 19676
rect 7398 19636 7423 19676
rect 7169 19613 7255 19636
rect 7337 19613 7423 19636
rect 11169 19676 11255 19699
rect 11337 19676 11423 19699
rect 11169 19636 11194 19676
rect 11194 19636 11234 19676
rect 11234 19636 11255 19676
rect 11337 19636 11358 19676
rect 11358 19636 11398 19676
rect 11398 19636 11423 19676
rect 11169 19613 11255 19636
rect 11337 19613 11423 19636
rect 15169 19676 15255 19699
rect 15337 19676 15423 19699
rect 15169 19636 15194 19676
rect 15194 19636 15234 19676
rect 15234 19636 15255 19676
rect 15337 19636 15358 19676
rect 15358 19636 15398 19676
rect 15398 19636 15423 19676
rect 15169 19613 15255 19636
rect 15337 19613 15423 19636
rect 19169 19676 19255 19699
rect 19337 19676 19423 19699
rect 19169 19636 19194 19676
rect 19194 19636 19234 19676
rect 19234 19636 19255 19676
rect 19337 19636 19358 19676
rect 19358 19636 19398 19676
rect 19398 19636 19423 19676
rect 19169 19613 19255 19636
rect 19337 19613 19423 19636
rect 23169 19676 23255 19699
rect 23337 19676 23423 19699
rect 23169 19636 23194 19676
rect 23194 19636 23234 19676
rect 23234 19636 23255 19676
rect 23337 19636 23358 19676
rect 23358 19636 23398 19676
rect 23398 19636 23423 19676
rect 23169 19613 23255 19636
rect 23337 19613 23423 19636
rect 27169 19676 27255 19699
rect 27337 19676 27423 19699
rect 27169 19636 27194 19676
rect 27194 19636 27234 19676
rect 27234 19636 27255 19676
rect 27337 19636 27358 19676
rect 27358 19636 27398 19676
rect 27398 19636 27423 19676
rect 27169 19613 27255 19636
rect 27337 19613 27423 19636
rect 31169 19676 31255 19699
rect 31337 19676 31423 19699
rect 31169 19636 31194 19676
rect 31194 19636 31234 19676
rect 31234 19636 31255 19676
rect 31337 19636 31358 19676
rect 31358 19636 31398 19676
rect 31398 19636 31423 19676
rect 31169 19613 31255 19636
rect 31337 19613 31423 19636
rect 35169 19676 35255 19699
rect 35337 19676 35423 19699
rect 35169 19636 35194 19676
rect 35194 19636 35234 19676
rect 35234 19636 35255 19676
rect 35337 19636 35358 19676
rect 35358 19636 35398 19676
rect 35398 19636 35423 19676
rect 35169 19613 35255 19636
rect 35337 19613 35423 19636
rect 39169 19676 39255 19699
rect 39337 19676 39423 19699
rect 39169 19636 39194 19676
rect 39194 19636 39234 19676
rect 39234 19636 39255 19676
rect 39337 19636 39358 19676
rect 39358 19636 39398 19676
rect 39398 19636 39423 19676
rect 39169 19613 39255 19636
rect 39337 19613 39423 19636
rect 43169 19676 43255 19699
rect 43337 19676 43423 19699
rect 43169 19636 43194 19676
rect 43194 19636 43234 19676
rect 43234 19636 43255 19676
rect 43337 19636 43358 19676
rect 43358 19636 43398 19676
rect 43398 19636 43423 19676
rect 43169 19613 43255 19636
rect 43337 19613 43423 19636
rect 47169 19676 47255 19699
rect 47337 19676 47423 19699
rect 47169 19636 47194 19676
rect 47194 19636 47234 19676
rect 47234 19636 47255 19676
rect 47337 19636 47358 19676
rect 47358 19636 47398 19676
rect 47398 19636 47423 19676
rect 47169 19613 47255 19636
rect 47337 19613 47423 19636
rect 51169 19676 51255 19699
rect 51337 19676 51423 19699
rect 51169 19636 51194 19676
rect 51194 19636 51234 19676
rect 51234 19636 51255 19676
rect 51337 19636 51358 19676
rect 51358 19636 51398 19676
rect 51398 19636 51423 19676
rect 51169 19613 51255 19636
rect 51337 19613 51423 19636
rect 55169 19676 55255 19699
rect 55337 19676 55423 19699
rect 55169 19636 55194 19676
rect 55194 19636 55234 19676
rect 55234 19636 55255 19676
rect 55337 19636 55358 19676
rect 55358 19636 55398 19676
rect 55398 19636 55423 19676
rect 55169 19613 55255 19636
rect 55337 19613 55423 19636
rect 59169 19676 59255 19699
rect 59337 19676 59423 19699
rect 59169 19636 59194 19676
rect 59194 19636 59234 19676
rect 59234 19636 59255 19676
rect 59337 19636 59358 19676
rect 59358 19636 59398 19676
rect 59398 19636 59423 19676
rect 59169 19613 59255 19636
rect 59337 19613 59423 19636
rect 63169 19676 63255 19699
rect 63337 19676 63423 19699
rect 63169 19636 63194 19676
rect 63194 19636 63234 19676
rect 63234 19636 63255 19676
rect 63337 19636 63358 19676
rect 63358 19636 63398 19676
rect 63398 19636 63423 19676
rect 63169 19613 63255 19636
rect 63337 19613 63423 19636
rect 67169 19676 67255 19699
rect 67337 19676 67423 19699
rect 67169 19636 67194 19676
rect 67194 19636 67234 19676
rect 67234 19636 67255 19676
rect 67337 19636 67358 19676
rect 67358 19636 67398 19676
rect 67398 19636 67423 19676
rect 67169 19613 67255 19636
rect 67337 19613 67423 19636
rect 71169 19676 71255 19699
rect 71337 19676 71423 19699
rect 71169 19636 71194 19676
rect 71194 19636 71234 19676
rect 71234 19636 71255 19676
rect 71337 19636 71358 19676
rect 71358 19636 71398 19676
rect 71398 19636 71423 19676
rect 71169 19613 71255 19636
rect 71337 19613 71423 19636
rect 75169 19676 75255 19699
rect 75337 19676 75423 19699
rect 75169 19636 75194 19676
rect 75194 19636 75234 19676
rect 75234 19636 75255 19676
rect 75337 19636 75358 19676
rect 75358 19636 75398 19676
rect 75398 19636 75423 19676
rect 75169 19613 75255 19636
rect 75337 19613 75423 19636
rect 79169 19676 79255 19699
rect 79337 19676 79423 19699
rect 79169 19636 79194 19676
rect 79194 19636 79234 19676
rect 79234 19636 79255 19676
rect 79337 19636 79358 19676
rect 79358 19636 79398 19676
rect 79398 19636 79423 19676
rect 79169 19613 79255 19636
rect 79337 19613 79423 19636
rect 83169 19676 83255 19699
rect 83337 19676 83423 19699
rect 83169 19636 83194 19676
rect 83194 19636 83234 19676
rect 83234 19636 83255 19676
rect 83337 19636 83358 19676
rect 83358 19636 83398 19676
rect 83398 19636 83423 19676
rect 83169 19613 83255 19636
rect 83337 19613 83423 19636
rect 87169 19676 87255 19699
rect 87337 19676 87423 19699
rect 87169 19636 87194 19676
rect 87194 19636 87234 19676
rect 87234 19636 87255 19676
rect 87337 19636 87358 19676
rect 87358 19636 87398 19676
rect 87398 19636 87423 19676
rect 87169 19613 87255 19636
rect 87337 19613 87423 19636
rect 91169 19676 91255 19699
rect 91337 19676 91423 19699
rect 91169 19636 91194 19676
rect 91194 19636 91234 19676
rect 91234 19636 91255 19676
rect 91337 19636 91358 19676
rect 91358 19636 91398 19676
rect 91398 19636 91423 19676
rect 91169 19613 91255 19636
rect 91337 19613 91423 19636
rect 95169 19676 95255 19699
rect 95337 19676 95423 19699
rect 95169 19636 95194 19676
rect 95194 19636 95234 19676
rect 95234 19636 95255 19676
rect 95337 19636 95358 19676
rect 95358 19636 95398 19676
rect 95398 19636 95423 19676
rect 95169 19613 95255 19636
rect 95337 19613 95423 19636
rect 99169 19676 99255 19699
rect 99337 19676 99423 19699
rect 99169 19636 99194 19676
rect 99194 19636 99234 19676
rect 99234 19636 99255 19676
rect 99337 19636 99358 19676
rect 99358 19636 99398 19676
rect 99398 19636 99423 19676
rect 99169 19613 99255 19636
rect 99337 19613 99423 19636
rect 86469 19277 86555 19363
rect 4409 18920 4495 18943
rect 4577 18920 4663 18943
rect 4409 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4495 18920
rect 4577 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4663 18920
rect 4409 18857 4495 18880
rect 4577 18857 4663 18880
rect 8409 18920 8495 18943
rect 8577 18920 8663 18943
rect 8409 18880 8434 18920
rect 8434 18880 8474 18920
rect 8474 18880 8495 18920
rect 8577 18880 8598 18920
rect 8598 18880 8638 18920
rect 8638 18880 8663 18920
rect 8409 18857 8495 18880
rect 8577 18857 8663 18880
rect 12409 18920 12495 18943
rect 12577 18920 12663 18943
rect 12409 18880 12434 18920
rect 12434 18880 12474 18920
rect 12474 18880 12495 18920
rect 12577 18880 12598 18920
rect 12598 18880 12638 18920
rect 12638 18880 12663 18920
rect 12409 18857 12495 18880
rect 12577 18857 12663 18880
rect 16409 18920 16495 18943
rect 16577 18920 16663 18943
rect 16409 18880 16434 18920
rect 16434 18880 16474 18920
rect 16474 18880 16495 18920
rect 16577 18880 16598 18920
rect 16598 18880 16638 18920
rect 16638 18880 16663 18920
rect 16409 18857 16495 18880
rect 16577 18857 16663 18880
rect 20409 18920 20495 18943
rect 20577 18920 20663 18943
rect 20409 18880 20434 18920
rect 20434 18880 20474 18920
rect 20474 18880 20495 18920
rect 20577 18880 20598 18920
rect 20598 18880 20638 18920
rect 20638 18880 20663 18920
rect 20409 18857 20495 18880
rect 20577 18857 20663 18880
rect 24409 18920 24495 18943
rect 24577 18920 24663 18943
rect 24409 18880 24434 18920
rect 24434 18880 24474 18920
rect 24474 18880 24495 18920
rect 24577 18880 24598 18920
rect 24598 18880 24638 18920
rect 24638 18880 24663 18920
rect 24409 18857 24495 18880
rect 24577 18857 24663 18880
rect 28409 18920 28495 18943
rect 28577 18920 28663 18943
rect 28409 18880 28434 18920
rect 28434 18880 28474 18920
rect 28474 18880 28495 18920
rect 28577 18880 28598 18920
rect 28598 18880 28638 18920
rect 28638 18880 28663 18920
rect 28409 18857 28495 18880
rect 28577 18857 28663 18880
rect 32409 18920 32495 18943
rect 32577 18920 32663 18943
rect 32409 18880 32434 18920
rect 32434 18880 32474 18920
rect 32474 18880 32495 18920
rect 32577 18880 32598 18920
rect 32598 18880 32638 18920
rect 32638 18880 32663 18920
rect 32409 18857 32495 18880
rect 32577 18857 32663 18880
rect 36409 18920 36495 18943
rect 36577 18920 36663 18943
rect 36409 18880 36434 18920
rect 36434 18880 36474 18920
rect 36474 18880 36495 18920
rect 36577 18880 36598 18920
rect 36598 18880 36638 18920
rect 36638 18880 36663 18920
rect 36409 18857 36495 18880
rect 36577 18857 36663 18880
rect 40409 18920 40495 18943
rect 40577 18920 40663 18943
rect 40409 18880 40434 18920
rect 40434 18880 40474 18920
rect 40474 18880 40495 18920
rect 40577 18880 40598 18920
rect 40598 18880 40638 18920
rect 40638 18880 40663 18920
rect 40409 18857 40495 18880
rect 40577 18857 40663 18880
rect 44409 18920 44495 18943
rect 44577 18920 44663 18943
rect 44409 18880 44434 18920
rect 44434 18880 44474 18920
rect 44474 18880 44495 18920
rect 44577 18880 44598 18920
rect 44598 18880 44638 18920
rect 44638 18880 44663 18920
rect 44409 18857 44495 18880
rect 44577 18857 44663 18880
rect 48409 18920 48495 18943
rect 48577 18920 48663 18943
rect 48409 18880 48434 18920
rect 48434 18880 48474 18920
rect 48474 18880 48495 18920
rect 48577 18880 48598 18920
rect 48598 18880 48638 18920
rect 48638 18880 48663 18920
rect 48409 18857 48495 18880
rect 48577 18857 48663 18880
rect 52409 18920 52495 18943
rect 52577 18920 52663 18943
rect 52409 18880 52434 18920
rect 52434 18880 52474 18920
rect 52474 18880 52495 18920
rect 52577 18880 52598 18920
rect 52598 18880 52638 18920
rect 52638 18880 52663 18920
rect 52409 18857 52495 18880
rect 52577 18857 52663 18880
rect 56409 18920 56495 18943
rect 56577 18920 56663 18943
rect 56409 18880 56434 18920
rect 56434 18880 56474 18920
rect 56474 18880 56495 18920
rect 56577 18880 56598 18920
rect 56598 18880 56638 18920
rect 56638 18880 56663 18920
rect 56409 18857 56495 18880
rect 56577 18857 56663 18880
rect 60409 18920 60495 18943
rect 60577 18920 60663 18943
rect 60409 18880 60434 18920
rect 60434 18880 60474 18920
rect 60474 18880 60495 18920
rect 60577 18880 60598 18920
rect 60598 18880 60638 18920
rect 60638 18880 60663 18920
rect 60409 18857 60495 18880
rect 60577 18857 60663 18880
rect 64409 18920 64495 18943
rect 64577 18920 64663 18943
rect 64409 18880 64434 18920
rect 64434 18880 64474 18920
rect 64474 18880 64495 18920
rect 64577 18880 64598 18920
rect 64598 18880 64638 18920
rect 64638 18880 64663 18920
rect 64409 18857 64495 18880
rect 64577 18857 64663 18880
rect 68409 18920 68495 18943
rect 68577 18920 68663 18943
rect 68409 18880 68434 18920
rect 68434 18880 68474 18920
rect 68474 18880 68495 18920
rect 68577 18880 68598 18920
rect 68598 18880 68638 18920
rect 68638 18880 68663 18920
rect 68409 18857 68495 18880
rect 68577 18857 68663 18880
rect 72409 18920 72495 18943
rect 72577 18920 72663 18943
rect 72409 18880 72434 18920
rect 72434 18880 72474 18920
rect 72474 18880 72495 18920
rect 72577 18880 72598 18920
rect 72598 18880 72638 18920
rect 72638 18880 72663 18920
rect 72409 18857 72495 18880
rect 72577 18857 72663 18880
rect 76409 18920 76495 18943
rect 76577 18920 76663 18943
rect 76409 18880 76434 18920
rect 76434 18880 76474 18920
rect 76474 18880 76495 18920
rect 76577 18880 76598 18920
rect 76598 18880 76638 18920
rect 76638 18880 76663 18920
rect 76409 18857 76495 18880
rect 76577 18857 76663 18880
rect 80409 18920 80495 18943
rect 80577 18920 80663 18943
rect 80409 18880 80434 18920
rect 80434 18880 80474 18920
rect 80474 18880 80495 18920
rect 80577 18880 80598 18920
rect 80598 18880 80638 18920
rect 80638 18880 80663 18920
rect 80409 18857 80495 18880
rect 80577 18857 80663 18880
rect 84409 18920 84495 18943
rect 84577 18920 84663 18943
rect 84409 18880 84434 18920
rect 84434 18880 84474 18920
rect 84474 18880 84495 18920
rect 84577 18880 84598 18920
rect 84598 18880 84638 18920
rect 84638 18880 84663 18920
rect 84409 18857 84495 18880
rect 84577 18857 84663 18880
rect 88409 18920 88495 18943
rect 88577 18920 88663 18943
rect 88409 18880 88434 18920
rect 88434 18880 88474 18920
rect 88474 18880 88495 18920
rect 88577 18880 88598 18920
rect 88598 18880 88638 18920
rect 88638 18880 88663 18920
rect 88409 18857 88495 18880
rect 88577 18857 88663 18880
rect 92409 18920 92495 18943
rect 92577 18920 92663 18943
rect 92409 18880 92434 18920
rect 92434 18880 92474 18920
rect 92474 18880 92495 18920
rect 92577 18880 92598 18920
rect 92598 18880 92638 18920
rect 92638 18880 92663 18920
rect 92409 18857 92495 18880
rect 92577 18857 92663 18880
rect 96409 18920 96495 18943
rect 96577 18920 96663 18943
rect 96409 18880 96434 18920
rect 96434 18880 96474 18920
rect 96474 18880 96495 18920
rect 96577 18880 96598 18920
rect 96598 18880 96638 18920
rect 96638 18880 96663 18920
rect 96409 18857 96495 18880
rect 96577 18857 96663 18880
rect 3169 18164 3255 18187
rect 3337 18164 3423 18187
rect 3169 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3255 18164
rect 3337 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3423 18164
rect 3169 18101 3255 18124
rect 3337 18101 3423 18124
rect 7169 18164 7255 18187
rect 7337 18164 7423 18187
rect 7169 18124 7194 18164
rect 7194 18124 7234 18164
rect 7234 18124 7255 18164
rect 7337 18124 7358 18164
rect 7358 18124 7398 18164
rect 7398 18124 7423 18164
rect 7169 18101 7255 18124
rect 7337 18101 7423 18124
rect 11169 18164 11255 18187
rect 11337 18164 11423 18187
rect 11169 18124 11194 18164
rect 11194 18124 11234 18164
rect 11234 18124 11255 18164
rect 11337 18124 11358 18164
rect 11358 18124 11398 18164
rect 11398 18124 11423 18164
rect 11169 18101 11255 18124
rect 11337 18101 11423 18124
rect 15169 18164 15255 18187
rect 15337 18164 15423 18187
rect 15169 18124 15194 18164
rect 15194 18124 15234 18164
rect 15234 18124 15255 18164
rect 15337 18124 15358 18164
rect 15358 18124 15398 18164
rect 15398 18124 15423 18164
rect 15169 18101 15255 18124
rect 15337 18101 15423 18124
rect 19169 18164 19255 18187
rect 19337 18164 19423 18187
rect 19169 18124 19194 18164
rect 19194 18124 19234 18164
rect 19234 18124 19255 18164
rect 19337 18124 19358 18164
rect 19358 18124 19398 18164
rect 19398 18124 19423 18164
rect 19169 18101 19255 18124
rect 19337 18101 19423 18124
rect 23169 18164 23255 18187
rect 23337 18164 23423 18187
rect 23169 18124 23194 18164
rect 23194 18124 23234 18164
rect 23234 18124 23255 18164
rect 23337 18124 23358 18164
rect 23358 18124 23398 18164
rect 23398 18124 23423 18164
rect 23169 18101 23255 18124
rect 23337 18101 23423 18124
rect 27169 18164 27255 18187
rect 27337 18164 27423 18187
rect 27169 18124 27194 18164
rect 27194 18124 27234 18164
rect 27234 18124 27255 18164
rect 27337 18124 27358 18164
rect 27358 18124 27398 18164
rect 27398 18124 27423 18164
rect 27169 18101 27255 18124
rect 27337 18101 27423 18124
rect 31169 18164 31255 18187
rect 31337 18164 31423 18187
rect 31169 18124 31194 18164
rect 31194 18124 31234 18164
rect 31234 18124 31255 18164
rect 31337 18124 31358 18164
rect 31358 18124 31398 18164
rect 31398 18124 31423 18164
rect 31169 18101 31255 18124
rect 31337 18101 31423 18124
rect 35169 18164 35255 18187
rect 35337 18164 35423 18187
rect 35169 18124 35194 18164
rect 35194 18124 35234 18164
rect 35234 18124 35255 18164
rect 35337 18124 35358 18164
rect 35358 18124 35398 18164
rect 35398 18124 35423 18164
rect 35169 18101 35255 18124
rect 35337 18101 35423 18124
rect 39169 18164 39255 18187
rect 39337 18164 39423 18187
rect 39169 18124 39194 18164
rect 39194 18124 39234 18164
rect 39234 18124 39255 18164
rect 39337 18124 39358 18164
rect 39358 18124 39398 18164
rect 39398 18124 39423 18164
rect 39169 18101 39255 18124
rect 39337 18101 39423 18124
rect 43169 18164 43255 18187
rect 43337 18164 43423 18187
rect 43169 18124 43194 18164
rect 43194 18124 43234 18164
rect 43234 18124 43255 18164
rect 43337 18124 43358 18164
rect 43358 18124 43398 18164
rect 43398 18124 43423 18164
rect 43169 18101 43255 18124
rect 43337 18101 43423 18124
rect 47169 18164 47255 18187
rect 47337 18164 47423 18187
rect 47169 18124 47194 18164
rect 47194 18124 47234 18164
rect 47234 18124 47255 18164
rect 47337 18124 47358 18164
rect 47358 18124 47398 18164
rect 47398 18124 47423 18164
rect 47169 18101 47255 18124
rect 47337 18101 47423 18124
rect 51169 18164 51255 18187
rect 51337 18164 51423 18187
rect 51169 18124 51194 18164
rect 51194 18124 51234 18164
rect 51234 18124 51255 18164
rect 51337 18124 51358 18164
rect 51358 18124 51398 18164
rect 51398 18124 51423 18164
rect 51169 18101 51255 18124
rect 51337 18101 51423 18124
rect 55169 18164 55255 18187
rect 55337 18164 55423 18187
rect 55169 18124 55194 18164
rect 55194 18124 55234 18164
rect 55234 18124 55255 18164
rect 55337 18124 55358 18164
rect 55358 18124 55398 18164
rect 55398 18124 55423 18164
rect 55169 18101 55255 18124
rect 55337 18101 55423 18124
rect 59169 18164 59255 18187
rect 59337 18164 59423 18187
rect 59169 18124 59194 18164
rect 59194 18124 59234 18164
rect 59234 18124 59255 18164
rect 59337 18124 59358 18164
rect 59358 18124 59398 18164
rect 59398 18124 59423 18164
rect 59169 18101 59255 18124
rect 59337 18101 59423 18124
rect 63169 18164 63255 18187
rect 63337 18164 63423 18187
rect 63169 18124 63194 18164
rect 63194 18124 63234 18164
rect 63234 18124 63255 18164
rect 63337 18124 63358 18164
rect 63358 18124 63398 18164
rect 63398 18124 63423 18164
rect 63169 18101 63255 18124
rect 63337 18101 63423 18124
rect 67169 18164 67255 18187
rect 67337 18164 67423 18187
rect 67169 18124 67194 18164
rect 67194 18124 67234 18164
rect 67234 18124 67255 18164
rect 67337 18124 67358 18164
rect 67358 18124 67398 18164
rect 67398 18124 67423 18164
rect 67169 18101 67255 18124
rect 67337 18101 67423 18124
rect 71169 18164 71255 18187
rect 71337 18164 71423 18187
rect 71169 18124 71194 18164
rect 71194 18124 71234 18164
rect 71234 18124 71255 18164
rect 71337 18124 71358 18164
rect 71358 18124 71398 18164
rect 71398 18124 71423 18164
rect 71169 18101 71255 18124
rect 71337 18101 71423 18124
rect 75169 18164 75255 18187
rect 75337 18164 75423 18187
rect 75169 18124 75194 18164
rect 75194 18124 75234 18164
rect 75234 18124 75255 18164
rect 75337 18124 75358 18164
rect 75358 18124 75398 18164
rect 75398 18124 75423 18164
rect 75169 18101 75255 18124
rect 75337 18101 75423 18124
rect 79169 18164 79255 18187
rect 79337 18164 79423 18187
rect 79169 18124 79194 18164
rect 79194 18124 79234 18164
rect 79234 18124 79255 18164
rect 79337 18124 79358 18164
rect 79358 18124 79398 18164
rect 79398 18124 79423 18164
rect 79169 18101 79255 18124
rect 79337 18101 79423 18124
rect 83169 18164 83255 18187
rect 83337 18164 83423 18187
rect 83169 18124 83194 18164
rect 83194 18124 83234 18164
rect 83234 18124 83255 18164
rect 83337 18124 83358 18164
rect 83358 18124 83398 18164
rect 83398 18124 83423 18164
rect 83169 18101 83255 18124
rect 83337 18101 83423 18124
rect 87169 18164 87255 18187
rect 87337 18164 87423 18187
rect 87169 18124 87194 18164
rect 87194 18124 87234 18164
rect 87234 18124 87255 18164
rect 87337 18124 87358 18164
rect 87358 18124 87398 18164
rect 87398 18124 87423 18164
rect 87169 18101 87255 18124
rect 87337 18101 87423 18124
rect 91169 18164 91255 18187
rect 91337 18164 91423 18187
rect 91169 18124 91194 18164
rect 91194 18124 91234 18164
rect 91234 18124 91255 18164
rect 91337 18124 91358 18164
rect 91358 18124 91398 18164
rect 91398 18124 91423 18164
rect 91169 18101 91255 18124
rect 91337 18101 91423 18124
rect 95169 18164 95255 18187
rect 95337 18164 95423 18187
rect 95169 18124 95194 18164
rect 95194 18124 95234 18164
rect 95234 18124 95255 18164
rect 95337 18124 95358 18164
rect 95358 18124 95398 18164
rect 95398 18124 95423 18164
rect 95169 18101 95255 18124
rect 95337 18101 95423 18124
rect 99169 18164 99255 18187
rect 99337 18164 99423 18187
rect 99169 18124 99194 18164
rect 99194 18124 99234 18164
rect 99234 18124 99255 18164
rect 99337 18124 99358 18164
rect 99358 18124 99398 18164
rect 99398 18124 99423 18164
rect 99169 18101 99255 18124
rect 99337 18101 99423 18124
rect 4409 17408 4495 17431
rect 4577 17408 4663 17431
rect 4409 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4495 17408
rect 4577 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4663 17408
rect 4409 17345 4495 17368
rect 4577 17345 4663 17368
rect 8409 17408 8495 17431
rect 8577 17408 8663 17431
rect 8409 17368 8434 17408
rect 8434 17368 8474 17408
rect 8474 17368 8495 17408
rect 8577 17368 8598 17408
rect 8598 17368 8638 17408
rect 8638 17368 8663 17408
rect 8409 17345 8495 17368
rect 8577 17345 8663 17368
rect 12409 17408 12495 17431
rect 12577 17408 12663 17431
rect 12409 17368 12434 17408
rect 12434 17368 12474 17408
rect 12474 17368 12495 17408
rect 12577 17368 12598 17408
rect 12598 17368 12638 17408
rect 12638 17368 12663 17408
rect 12409 17345 12495 17368
rect 12577 17345 12663 17368
rect 16409 17408 16495 17431
rect 16577 17408 16663 17431
rect 16409 17368 16434 17408
rect 16434 17368 16474 17408
rect 16474 17368 16495 17408
rect 16577 17368 16598 17408
rect 16598 17368 16638 17408
rect 16638 17368 16663 17408
rect 16409 17345 16495 17368
rect 16577 17345 16663 17368
rect 20409 17408 20495 17431
rect 20577 17408 20663 17431
rect 20409 17368 20434 17408
rect 20434 17368 20474 17408
rect 20474 17368 20495 17408
rect 20577 17368 20598 17408
rect 20598 17368 20638 17408
rect 20638 17368 20663 17408
rect 20409 17345 20495 17368
rect 20577 17345 20663 17368
rect 24409 17408 24495 17431
rect 24577 17408 24663 17431
rect 24409 17368 24434 17408
rect 24434 17368 24474 17408
rect 24474 17368 24495 17408
rect 24577 17368 24598 17408
rect 24598 17368 24638 17408
rect 24638 17368 24663 17408
rect 24409 17345 24495 17368
rect 24577 17345 24663 17368
rect 28409 17408 28495 17431
rect 28577 17408 28663 17431
rect 28409 17368 28434 17408
rect 28434 17368 28474 17408
rect 28474 17368 28495 17408
rect 28577 17368 28598 17408
rect 28598 17368 28638 17408
rect 28638 17368 28663 17408
rect 28409 17345 28495 17368
rect 28577 17345 28663 17368
rect 32409 17408 32495 17431
rect 32577 17408 32663 17431
rect 32409 17368 32434 17408
rect 32434 17368 32474 17408
rect 32474 17368 32495 17408
rect 32577 17368 32598 17408
rect 32598 17368 32638 17408
rect 32638 17368 32663 17408
rect 32409 17345 32495 17368
rect 32577 17345 32663 17368
rect 36409 17408 36495 17431
rect 36577 17408 36663 17431
rect 36409 17368 36434 17408
rect 36434 17368 36474 17408
rect 36474 17368 36495 17408
rect 36577 17368 36598 17408
rect 36598 17368 36638 17408
rect 36638 17368 36663 17408
rect 36409 17345 36495 17368
rect 36577 17345 36663 17368
rect 40409 17408 40495 17431
rect 40577 17408 40663 17431
rect 40409 17368 40434 17408
rect 40434 17368 40474 17408
rect 40474 17368 40495 17408
rect 40577 17368 40598 17408
rect 40598 17368 40638 17408
rect 40638 17368 40663 17408
rect 40409 17345 40495 17368
rect 40577 17345 40663 17368
rect 44409 17408 44495 17431
rect 44577 17408 44663 17431
rect 44409 17368 44434 17408
rect 44434 17368 44474 17408
rect 44474 17368 44495 17408
rect 44577 17368 44598 17408
rect 44598 17368 44638 17408
rect 44638 17368 44663 17408
rect 44409 17345 44495 17368
rect 44577 17345 44663 17368
rect 48409 17408 48495 17431
rect 48577 17408 48663 17431
rect 48409 17368 48434 17408
rect 48434 17368 48474 17408
rect 48474 17368 48495 17408
rect 48577 17368 48598 17408
rect 48598 17368 48638 17408
rect 48638 17368 48663 17408
rect 48409 17345 48495 17368
rect 48577 17345 48663 17368
rect 52409 17408 52495 17431
rect 52577 17408 52663 17431
rect 52409 17368 52434 17408
rect 52434 17368 52474 17408
rect 52474 17368 52495 17408
rect 52577 17368 52598 17408
rect 52598 17368 52638 17408
rect 52638 17368 52663 17408
rect 52409 17345 52495 17368
rect 52577 17345 52663 17368
rect 56409 17408 56495 17431
rect 56577 17408 56663 17431
rect 56409 17368 56434 17408
rect 56434 17368 56474 17408
rect 56474 17368 56495 17408
rect 56577 17368 56598 17408
rect 56598 17368 56638 17408
rect 56638 17368 56663 17408
rect 56409 17345 56495 17368
rect 56577 17345 56663 17368
rect 60409 17408 60495 17431
rect 60577 17408 60663 17431
rect 60409 17368 60434 17408
rect 60434 17368 60474 17408
rect 60474 17368 60495 17408
rect 60577 17368 60598 17408
rect 60598 17368 60638 17408
rect 60638 17368 60663 17408
rect 60409 17345 60495 17368
rect 60577 17345 60663 17368
rect 64409 17408 64495 17431
rect 64577 17408 64663 17431
rect 64409 17368 64434 17408
rect 64434 17368 64474 17408
rect 64474 17368 64495 17408
rect 64577 17368 64598 17408
rect 64598 17368 64638 17408
rect 64638 17368 64663 17408
rect 64409 17345 64495 17368
rect 64577 17345 64663 17368
rect 68409 17408 68495 17431
rect 68577 17408 68663 17431
rect 68409 17368 68434 17408
rect 68434 17368 68474 17408
rect 68474 17368 68495 17408
rect 68577 17368 68598 17408
rect 68598 17368 68638 17408
rect 68638 17368 68663 17408
rect 68409 17345 68495 17368
rect 68577 17345 68663 17368
rect 72409 17408 72495 17431
rect 72577 17408 72663 17431
rect 72409 17368 72434 17408
rect 72434 17368 72474 17408
rect 72474 17368 72495 17408
rect 72577 17368 72598 17408
rect 72598 17368 72638 17408
rect 72638 17368 72663 17408
rect 72409 17345 72495 17368
rect 72577 17345 72663 17368
rect 76409 17408 76495 17431
rect 76577 17408 76663 17431
rect 76409 17368 76434 17408
rect 76434 17368 76474 17408
rect 76474 17368 76495 17408
rect 76577 17368 76598 17408
rect 76598 17368 76638 17408
rect 76638 17368 76663 17408
rect 76409 17345 76495 17368
rect 76577 17345 76663 17368
rect 80409 17408 80495 17431
rect 80577 17408 80663 17431
rect 80409 17368 80434 17408
rect 80434 17368 80474 17408
rect 80474 17368 80495 17408
rect 80577 17368 80598 17408
rect 80598 17368 80638 17408
rect 80638 17368 80663 17408
rect 80409 17345 80495 17368
rect 80577 17345 80663 17368
rect 84409 17408 84495 17431
rect 84577 17408 84663 17431
rect 84409 17368 84434 17408
rect 84434 17368 84474 17408
rect 84474 17368 84495 17408
rect 84577 17368 84598 17408
rect 84598 17368 84638 17408
rect 84638 17368 84663 17408
rect 84409 17345 84495 17368
rect 84577 17345 84663 17368
rect 88409 17408 88495 17431
rect 88577 17408 88663 17431
rect 88409 17368 88434 17408
rect 88434 17368 88474 17408
rect 88474 17368 88495 17408
rect 88577 17368 88598 17408
rect 88598 17368 88638 17408
rect 88638 17368 88663 17408
rect 88409 17345 88495 17368
rect 88577 17345 88663 17368
rect 92409 17408 92495 17431
rect 92577 17408 92663 17431
rect 92409 17368 92434 17408
rect 92434 17368 92474 17408
rect 92474 17368 92495 17408
rect 92577 17368 92598 17408
rect 92598 17368 92638 17408
rect 92638 17368 92663 17408
rect 92409 17345 92495 17368
rect 92577 17345 92663 17368
rect 96409 17408 96495 17431
rect 96577 17408 96663 17431
rect 96409 17368 96434 17408
rect 96434 17368 96474 17408
rect 96474 17368 96495 17408
rect 96577 17368 96598 17408
rect 96598 17368 96638 17408
rect 96638 17368 96663 17408
rect 96409 17345 96495 17368
rect 96577 17345 96663 17368
rect 3169 16652 3255 16675
rect 3337 16652 3423 16675
rect 3169 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3255 16652
rect 3337 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3423 16652
rect 3169 16589 3255 16612
rect 3337 16589 3423 16612
rect 7169 16652 7255 16675
rect 7337 16652 7423 16675
rect 7169 16612 7194 16652
rect 7194 16612 7234 16652
rect 7234 16612 7255 16652
rect 7337 16612 7358 16652
rect 7358 16612 7398 16652
rect 7398 16612 7423 16652
rect 7169 16589 7255 16612
rect 7337 16589 7423 16612
rect 11169 16652 11255 16675
rect 11337 16652 11423 16675
rect 11169 16612 11194 16652
rect 11194 16612 11234 16652
rect 11234 16612 11255 16652
rect 11337 16612 11358 16652
rect 11358 16612 11398 16652
rect 11398 16612 11423 16652
rect 11169 16589 11255 16612
rect 11337 16589 11423 16612
rect 15169 16652 15255 16675
rect 15337 16652 15423 16675
rect 15169 16612 15194 16652
rect 15194 16612 15234 16652
rect 15234 16612 15255 16652
rect 15337 16612 15358 16652
rect 15358 16612 15398 16652
rect 15398 16612 15423 16652
rect 15169 16589 15255 16612
rect 15337 16589 15423 16612
rect 19169 16652 19255 16675
rect 19337 16652 19423 16675
rect 19169 16612 19194 16652
rect 19194 16612 19234 16652
rect 19234 16612 19255 16652
rect 19337 16612 19358 16652
rect 19358 16612 19398 16652
rect 19398 16612 19423 16652
rect 19169 16589 19255 16612
rect 19337 16589 19423 16612
rect 23169 16652 23255 16675
rect 23337 16652 23423 16675
rect 23169 16612 23194 16652
rect 23194 16612 23234 16652
rect 23234 16612 23255 16652
rect 23337 16612 23358 16652
rect 23358 16612 23398 16652
rect 23398 16612 23423 16652
rect 23169 16589 23255 16612
rect 23337 16589 23423 16612
rect 27169 16652 27255 16675
rect 27337 16652 27423 16675
rect 27169 16612 27194 16652
rect 27194 16612 27234 16652
rect 27234 16612 27255 16652
rect 27337 16612 27358 16652
rect 27358 16612 27398 16652
rect 27398 16612 27423 16652
rect 27169 16589 27255 16612
rect 27337 16589 27423 16612
rect 31169 16652 31255 16675
rect 31337 16652 31423 16675
rect 31169 16612 31194 16652
rect 31194 16612 31234 16652
rect 31234 16612 31255 16652
rect 31337 16612 31358 16652
rect 31358 16612 31398 16652
rect 31398 16612 31423 16652
rect 31169 16589 31255 16612
rect 31337 16589 31423 16612
rect 35169 16652 35255 16675
rect 35337 16652 35423 16675
rect 35169 16612 35194 16652
rect 35194 16612 35234 16652
rect 35234 16612 35255 16652
rect 35337 16612 35358 16652
rect 35358 16612 35398 16652
rect 35398 16612 35423 16652
rect 35169 16589 35255 16612
rect 35337 16589 35423 16612
rect 39169 16652 39255 16675
rect 39337 16652 39423 16675
rect 39169 16612 39194 16652
rect 39194 16612 39234 16652
rect 39234 16612 39255 16652
rect 39337 16612 39358 16652
rect 39358 16612 39398 16652
rect 39398 16612 39423 16652
rect 39169 16589 39255 16612
rect 39337 16589 39423 16612
rect 43169 16652 43255 16675
rect 43337 16652 43423 16675
rect 43169 16612 43194 16652
rect 43194 16612 43234 16652
rect 43234 16612 43255 16652
rect 43337 16612 43358 16652
rect 43358 16612 43398 16652
rect 43398 16612 43423 16652
rect 43169 16589 43255 16612
rect 43337 16589 43423 16612
rect 47169 16652 47255 16675
rect 47337 16652 47423 16675
rect 47169 16612 47194 16652
rect 47194 16612 47234 16652
rect 47234 16612 47255 16652
rect 47337 16612 47358 16652
rect 47358 16612 47398 16652
rect 47398 16612 47423 16652
rect 47169 16589 47255 16612
rect 47337 16589 47423 16612
rect 51169 16652 51255 16675
rect 51337 16652 51423 16675
rect 51169 16612 51194 16652
rect 51194 16612 51234 16652
rect 51234 16612 51255 16652
rect 51337 16612 51358 16652
rect 51358 16612 51398 16652
rect 51398 16612 51423 16652
rect 51169 16589 51255 16612
rect 51337 16589 51423 16612
rect 55169 16652 55255 16675
rect 55337 16652 55423 16675
rect 55169 16612 55194 16652
rect 55194 16612 55234 16652
rect 55234 16612 55255 16652
rect 55337 16612 55358 16652
rect 55358 16612 55398 16652
rect 55398 16612 55423 16652
rect 55169 16589 55255 16612
rect 55337 16589 55423 16612
rect 59169 16652 59255 16675
rect 59337 16652 59423 16675
rect 59169 16612 59194 16652
rect 59194 16612 59234 16652
rect 59234 16612 59255 16652
rect 59337 16612 59358 16652
rect 59358 16612 59398 16652
rect 59398 16612 59423 16652
rect 59169 16589 59255 16612
rect 59337 16589 59423 16612
rect 63169 16652 63255 16675
rect 63337 16652 63423 16675
rect 63169 16612 63194 16652
rect 63194 16612 63234 16652
rect 63234 16612 63255 16652
rect 63337 16612 63358 16652
rect 63358 16612 63398 16652
rect 63398 16612 63423 16652
rect 63169 16589 63255 16612
rect 63337 16589 63423 16612
rect 67169 16652 67255 16675
rect 67337 16652 67423 16675
rect 67169 16612 67194 16652
rect 67194 16612 67234 16652
rect 67234 16612 67255 16652
rect 67337 16612 67358 16652
rect 67358 16612 67398 16652
rect 67398 16612 67423 16652
rect 67169 16589 67255 16612
rect 67337 16589 67423 16612
rect 4409 15896 4495 15919
rect 4577 15896 4663 15919
rect 4409 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4495 15896
rect 4577 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4663 15896
rect 4409 15833 4495 15856
rect 4577 15833 4663 15856
rect 8409 15896 8495 15919
rect 8577 15896 8663 15919
rect 8409 15856 8434 15896
rect 8434 15856 8474 15896
rect 8474 15856 8495 15896
rect 8577 15856 8598 15896
rect 8598 15856 8638 15896
rect 8638 15856 8663 15896
rect 8409 15833 8495 15856
rect 8577 15833 8663 15856
rect 12409 15896 12495 15919
rect 12577 15896 12663 15919
rect 12409 15856 12434 15896
rect 12434 15856 12474 15896
rect 12474 15856 12495 15896
rect 12577 15856 12598 15896
rect 12598 15856 12638 15896
rect 12638 15856 12663 15896
rect 12409 15833 12495 15856
rect 12577 15833 12663 15856
rect 16409 15896 16495 15919
rect 16577 15896 16663 15919
rect 16409 15856 16434 15896
rect 16434 15856 16474 15896
rect 16474 15856 16495 15896
rect 16577 15856 16598 15896
rect 16598 15856 16638 15896
rect 16638 15856 16663 15896
rect 16409 15833 16495 15856
rect 16577 15833 16663 15856
rect 20409 15896 20495 15919
rect 20577 15896 20663 15919
rect 20409 15856 20434 15896
rect 20434 15856 20474 15896
rect 20474 15856 20495 15896
rect 20577 15856 20598 15896
rect 20598 15856 20638 15896
rect 20638 15856 20663 15896
rect 20409 15833 20495 15856
rect 20577 15833 20663 15856
rect 24409 15896 24495 15919
rect 24577 15896 24663 15919
rect 24409 15856 24434 15896
rect 24434 15856 24474 15896
rect 24474 15856 24495 15896
rect 24577 15856 24598 15896
rect 24598 15856 24638 15896
rect 24638 15856 24663 15896
rect 24409 15833 24495 15856
rect 24577 15833 24663 15856
rect 28409 15896 28495 15919
rect 28577 15896 28663 15919
rect 28409 15856 28434 15896
rect 28434 15856 28474 15896
rect 28474 15856 28495 15896
rect 28577 15856 28598 15896
rect 28598 15856 28638 15896
rect 28638 15856 28663 15896
rect 28409 15833 28495 15856
rect 28577 15833 28663 15856
rect 32409 15896 32495 15919
rect 32577 15896 32663 15919
rect 32409 15856 32434 15896
rect 32434 15856 32474 15896
rect 32474 15856 32495 15896
rect 32577 15856 32598 15896
rect 32598 15856 32638 15896
rect 32638 15856 32663 15896
rect 32409 15833 32495 15856
rect 32577 15833 32663 15856
rect 36409 15896 36495 15919
rect 36577 15896 36663 15919
rect 36409 15856 36434 15896
rect 36434 15856 36474 15896
rect 36474 15856 36495 15896
rect 36577 15856 36598 15896
rect 36598 15856 36638 15896
rect 36638 15856 36663 15896
rect 36409 15833 36495 15856
rect 36577 15833 36663 15856
rect 40409 15896 40495 15919
rect 40577 15896 40663 15919
rect 40409 15856 40434 15896
rect 40434 15856 40474 15896
rect 40474 15856 40495 15896
rect 40577 15856 40598 15896
rect 40598 15856 40638 15896
rect 40638 15856 40663 15896
rect 40409 15833 40495 15856
rect 40577 15833 40663 15856
rect 44409 15896 44495 15919
rect 44577 15896 44663 15919
rect 44409 15856 44434 15896
rect 44434 15856 44474 15896
rect 44474 15856 44495 15896
rect 44577 15856 44598 15896
rect 44598 15856 44638 15896
rect 44638 15856 44663 15896
rect 44409 15833 44495 15856
rect 44577 15833 44663 15856
rect 48409 15896 48495 15919
rect 48577 15896 48663 15919
rect 48409 15856 48434 15896
rect 48434 15856 48474 15896
rect 48474 15856 48495 15896
rect 48577 15856 48598 15896
rect 48598 15856 48638 15896
rect 48638 15856 48663 15896
rect 48409 15833 48495 15856
rect 48577 15833 48663 15856
rect 52409 15896 52495 15919
rect 52577 15896 52663 15919
rect 52409 15856 52434 15896
rect 52434 15856 52474 15896
rect 52474 15856 52495 15896
rect 52577 15856 52598 15896
rect 52598 15856 52638 15896
rect 52638 15856 52663 15896
rect 52409 15833 52495 15856
rect 52577 15833 52663 15856
rect 56409 15896 56495 15919
rect 56577 15896 56663 15919
rect 56409 15856 56434 15896
rect 56434 15856 56474 15896
rect 56474 15856 56495 15896
rect 56577 15856 56598 15896
rect 56598 15856 56638 15896
rect 56638 15856 56663 15896
rect 56409 15833 56495 15856
rect 56577 15833 56663 15856
rect 60409 15896 60495 15919
rect 60577 15896 60663 15919
rect 60409 15856 60434 15896
rect 60434 15856 60474 15896
rect 60474 15856 60495 15896
rect 60577 15856 60598 15896
rect 60598 15856 60638 15896
rect 60638 15856 60663 15896
rect 60409 15833 60495 15856
rect 60577 15833 60663 15856
rect 64409 15896 64495 15919
rect 64577 15896 64663 15919
rect 64409 15856 64434 15896
rect 64434 15856 64474 15896
rect 64474 15856 64495 15896
rect 64577 15856 64598 15896
rect 64598 15856 64638 15896
rect 64638 15856 64663 15896
rect 64409 15833 64495 15856
rect 64577 15833 64663 15856
rect 68409 15896 68495 15919
rect 68577 15896 68663 15919
rect 68409 15856 68434 15896
rect 68434 15856 68474 15896
rect 68474 15856 68495 15896
rect 68577 15856 68598 15896
rect 68598 15856 68638 15896
rect 68638 15856 68663 15896
rect 68409 15833 68495 15856
rect 68577 15833 68663 15856
rect 3169 15140 3255 15163
rect 3337 15140 3423 15163
rect 3169 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3255 15140
rect 3337 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3423 15140
rect 3169 15077 3255 15100
rect 3337 15077 3423 15100
rect 7169 15140 7255 15163
rect 7337 15140 7423 15163
rect 7169 15100 7194 15140
rect 7194 15100 7234 15140
rect 7234 15100 7255 15140
rect 7337 15100 7358 15140
rect 7358 15100 7398 15140
rect 7398 15100 7423 15140
rect 7169 15077 7255 15100
rect 7337 15077 7423 15100
rect 11169 15140 11255 15163
rect 11337 15140 11423 15163
rect 11169 15100 11194 15140
rect 11194 15100 11234 15140
rect 11234 15100 11255 15140
rect 11337 15100 11358 15140
rect 11358 15100 11398 15140
rect 11398 15100 11423 15140
rect 11169 15077 11255 15100
rect 11337 15077 11423 15100
rect 15169 15140 15255 15163
rect 15337 15140 15423 15163
rect 15169 15100 15194 15140
rect 15194 15100 15234 15140
rect 15234 15100 15255 15140
rect 15337 15100 15358 15140
rect 15358 15100 15398 15140
rect 15398 15100 15423 15140
rect 15169 15077 15255 15100
rect 15337 15077 15423 15100
rect 19169 15140 19255 15163
rect 19337 15140 19423 15163
rect 19169 15100 19194 15140
rect 19194 15100 19234 15140
rect 19234 15100 19255 15140
rect 19337 15100 19358 15140
rect 19358 15100 19398 15140
rect 19398 15100 19423 15140
rect 19169 15077 19255 15100
rect 19337 15077 19423 15100
rect 23169 15140 23255 15163
rect 23337 15140 23423 15163
rect 23169 15100 23194 15140
rect 23194 15100 23234 15140
rect 23234 15100 23255 15140
rect 23337 15100 23358 15140
rect 23358 15100 23398 15140
rect 23398 15100 23423 15140
rect 23169 15077 23255 15100
rect 23337 15077 23423 15100
rect 27169 15140 27255 15163
rect 27337 15140 27423 15163
rect 27169 15100 27194 15140
rect 27194 15100 27234 15140
rect 27234 15100 27255 15140
rect 27337 15100 27358 15140
rect 27358 15100 27398 15140
rect 27398 15100 27423 15140
rect 27169 15077 27255 15100
rect 27337 15077 27423 15100
rect 31169 15140 31255 15163
rect 31337 15140 31423 15163
rect 31169 15100 31194 15140
rect 31194 15100 31234 15140
rect 31234 15100 31255 15140
rect 31337 15100 31358 15140
rect 31358 15100 31398 15140
rect 31398 15100 31423 15140
rect 31169 15077 31255 15100
rect 31337 15077 31423 15100
rect 35169 15140 35255 15163
rect 35337 15140 35423 15163
rect 35169 15100 35194 15140
rect 35194 15100 35234 15140
rect 35234 15100 35255 15140
rect 35337 15100 35358 15140
rect 35358 15100 35398 15140
rect 35398 15100 35423 15140
rect 35169 15077 35255 15100
rect 35337 15077 35423 15100
rect 39169 15140 39255 15163
rect 39337 15140 39423 15163
rect 39169 15100 39194 15140
rect 39194 15100 39234 15140
rect 39234 15100 39255 15140
rect 39337 15100 39358 15140
rect 39358 15100 39398 15140
rect 39398 15100 39423 15140
rect 39169 15077 39255 15100
rect 39337 15077 39423 15100
rect 43169 15140 43255 15163
rect 43337 15140 43423 15163
rect 43169 15100 43194 15140
rect 43194 15100 43234 15140
rect 43234 15100 43255 15140
rect 43337 15100 43358 15140
rect 43358 15100 43398 15140
rect 43398 15100 43423 15140
rect 43169 15077 43255 15100
rect 43337 15077 43423 15100
rect 47169 15140 47255 15163
rect 47337 15140 47423 15163
rect 47169 15100 47194 15140
rect 47194 15100 47234 15140
rect 47234 15100 47255 15140
rect 47337 15100 47358 15140
rect 47358 15100 47398 15140
rect 47398 15100 47423 15140
rect 47169 15077 47255 15100
rect 47337 15077 47423 15100
rect 51169 15140 51255 15163
rect 51337 15140 51423 15163
rect 51169 15100 51194 15140
rect 51194 15100 51234 15140
rect 51234 15100 51255 15140
rect 51337 15100 51358 15140
rect 51358 15100 51398 15140
rect 51398 15100 51423 15140
rect 51169 15077 51255 15100
rect 51337 15077 51423 15100
rect 55169 15140 55255 15163
rect 55337 15140 55423 15163
rect 55169 15100 55194 15140
rect 55194 15100 55234 15140
rect 55234 15100 55255 15140
rect 55337 15100 55358 15140
rect 55358 15100 55398 15140
rect 55398 15100 55423 15140
rect 55169 15077 55255 15100
rect 55337 15077 55423 15100
rect 59169 15140 59255 15163
rect 59337 15140 59423 15163
rect 59169 15100 59194 15140
rect 59194 15100 59234 15140
rect 59234 15100 59255 15140
rect 59337 15100 59358 15140
rect 59358 15100 59398 15140
rect 59398 15100 59423 15140
rect 59169 15077 59255 15100
rect 59337 15077 59423 15100
rect 63169 15140 63255 15163
rect 63337 15140 63423 15163
rect 63169 15100 63194 15140
rect 63194 15100 63234 15140
rect 63234 15100 63255 15140
rect 63337 15100 63358 15140
rect 63358 15100 63398 15140
rect 63398 15100 63423 15140
rect 63169 15077 63255 15100
rect 63337 15077 63423 15100
rect 67169 15140 67255 15163
rect 67337 15140 67423 15163
rect 67169 15100 67194 15140
rect 67194 15100 67234 15140
rect 67234 15100 67255 15140
rect 67337 15100 67358 15140
rect 67358 15100 67398 15140
rect 67398 15100 67423 15140
rect 67169 15077 67255 15100
rect 67337 15077 67423 15100
rect 72409 15036 72495 15122
rect 72577 15036 72663 15122
rect 72409 14868 72495 14954
rect 72577 14868 72663 14954
rect 72409 14700 72495 14786
rect 72577 14700 72663 14786
rect 72409 14532 72495 14618
rect 72577 14532 72663 14618
rect 4409 14384 4495 14407
rect 4577 14384 4663 14407
rect 4409 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4495 14384
rect 4577 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4663 14384
rect 4409 14321 4495 14344
rect 4577 14321 4663 14344
rect 8409 14384 8495 14407
rect 8577 14384 8663 14407
rect 8409 14344 8434 14384
rect 8434 14344 8474 14384
rect 8474 14344 8495 14384
rect 8577 14344 8598 14384
rect 8598 14344 8638 14384
rect 8638 14344 8663 14384
rect 8409 14321 8495 14344
rect 8577 14321 8663 14344
rect 12409 14384 12495 14407
rect 12577 14384 12663 14407
rect 12409 14344 12434 14384
rect 12434 14344 12474 14384
rect 12474 14344 12495 14384
rect 12577 14344 12598 14384
rect 12598 14344 12638 14384
rect 12638 14344 12663 14384
rect 12409 14321 12495 14344
rect 12577 14321 12663 14344
rect 16409 14384 16495 14407
rect 16577 14384 16663 14407
rect 16409 14344 16434 14384
rect 16434 14344 16474 14384
rect 16474 14344 16495 14384
rect 16577 14344 16598 14384
rect 16598 14344 16638 14384
rect 16638 14344 16663 14384
rect 16409 14321 16495 14344
rect 16577 14321 16663 14344
rect 20409 14384 20495 14407
rect 20577 14384 20663 14407
rect 20409 14344 20434 14384
rect 20434 14344 20474 14384
rect 20474 14344 20495 14384
rect 20577 14344 20598 14384
rect 20598 14344 20638 14384
rect 20638 14344 20663 14384
rect 20409 14321 20495 14344
rect 20577 14321 20663 14344
rect 24409 14384 24495 14407
rect 24577 14384 24663 14407
rect 24409 14344 24434 14384
rect 24434 14344 24474 14384
rect 24474 14344 24495 14384
rect 24577 14344 24598 14384
rect 24598 14344 24638 14384
rect 24638 14344 24663 14384
rect 24409 14321 24495 14344
rect 24577 14321 24663 14344
rect 28409 14384 28495 14407
rect 28577 14384 28663 14407
rect 28409 14344 28434 14384
rect 28434 14344 28474 14384
rect 28474 14344 28495 14384
rect 28577 14344 28598 14384
rect 28598 14344 28638 14384
rect 28638 14344 28663 14384
rect 28409 14321 28495 14344
rect 28577 14321 28663 14344
rect 32409 14384 32495 14407
rect 32577 14384 32663 14407
rect 32409 14344 32434 14384
rect 32434 14344 32474 14384
rect 32474 14344 32495 14384
rect 32577 14344 32598 14384
rect 32598 14344 32638 14384
rect 32638 14344 32663 14384
rect 32409 14321 32495 14344
rect 32577 14321 32663 14344
rect 36409 14384 36495 14407
rect 36577 14384 36663 14407
rect 36409 14344 36434 14384
rect 36434 14344 36474 14384
rect 36474 14344 36495 14384
rect 36577 14344 36598 14384
rect 36598 14344 36638 14384
rect 36638 14344 36663 14384
rect 36409 14321 36495 14344
rect 36577 14321 36663 14344
rect 40409 14384 40495 14407
rect 40577 14384 40663 14407
rect 40409 14344 40434 14384
rect 40434 14344 40474 14384
rect 40474 14344 40495 14384
rect 40577 14344 40598 14384
rect 40598 14344 40638 14384
rect 40638 14344 40663 14384
rect 40409 14321 40495 14344
rect 40577 14321 40663 14344
rect 44409 14384 44495 14407
rect 44577 14384 44663 14407
rect 44409 14344 44434 14384
rect 44434 14344 44474 14384
rect 44474 14344 44495 14384
rect 44577 14344 44598 14384
rect 44598 14344 44638 14384
rect 44638 14344 44663 14384
rect 44409 14321 44495 14344
rect 44577 14321 44663 14344
rect 48409 14384 48495 14407
rect 48577 14384 48663 14407
rect 48409 14344 48434 14384
rect 48434 14344 48474 14384
rect 48474 14344 48495 14384
rect 48577 14344 48598 14384
rect 48598 14344 48638 14384
rect 48638 14344 48663 14384
rect 48409 14321 48495 14344
rect 48577 14321 48663 14344
rect 52409 14384 52495 14407
rect 52577 14384 52663 14407
rect 52409 14344 52434 14384
rect 52434 14344 52474 14384
rect 52474 14344 52495 14384
rect 52577 14344 52598 14384
rect 52598 14344 52638 14384
rect 52638 14344 52663 14384
rect 52409 14321 52495 14344
rect 52577 14321 52663 14344
rect 56409 14384 56495 14407
rect 56577 14384 56663 14407
rect 56409 14344 56434 14384
rect 56434 14344 56474 14384
rect 56474 14344 56495 14384
rect 56577 14344 56598 14384
rect 56598 14344 56638 14384
rect 56638 14344 56663 14384
rect 56409 14321 56495 14344
rect 56577 14321 56663 14344
rect 60409 14384 60495 14407
rect 60577 14384 60663 14407
rect 60409 14344 60434 14384
rect 60434 14344 60474 14384
rect 60474 14344 60495 14384
rect 60577 14344 60598 14384
rect 60598 14344 60638 14384
rect 60638 14344 60663 14384
rect 60409 14321 60495 14344
rect 60577 14321 60663 14344
rect 64409 14384 64495 14407
rect 64577 14384 64663 14407
rect 64409 14344 64434 14384
rect 64434 14344 64474 14384
rect 64474 14344 64495 14384
rect 64577 14344 64598 14384
rect 64598 14344 64638 14384
rect 64638 14344 64663 14384
rect 64409 14321 64495 14344
rect 64577 14321 64663 14344
rect 68409 14384 68495 14407
rect 68577 14384 68663 14407
rect 68409 14344 68434 14384
rect 68434 14344 68474 14384
rect 68474 14344 68495 14384
rect 68577 14344 68598 14384
rect 68598 14344 68638 14384
rect 68638 14344 68663 14384
rect 68409 14321 68495 14344
rect 68577 14321 68663 14344
rect 72409 14364 72495 14450
rect 72577 14364 72663 14450
rect 72409 14196 72495 14282
rect 72577 14196 72663 14282
rect 72409 14028 72495 14114
rect 72577 14028 72663 14114
rect 72409 13860 72495 13946
rect 72577 13860 72663 13946
rect 72409 13692 72495 13778
rect 72577 13692 72663 13778
rect 3169 13628 3255 13651
rect 3337 13628 3423 13651
rect 3169 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3255 13628
rect 3337 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3423 13628
rect 3169 13565 3255 13588
rect 3337 13565 3423 13588
rect 7169 13628 7255 13651
rect 7337 13628 7423 13651
rect 7169 13588 7194 13628
rect 7194 13588 7234 13628
rect 7234 13588 7255 13628
rect 7337 13588 7358 13628
rect 7358 13588 7398 13628
rect 7398 13588 7423 13628
rect 7169 13565 7255 13588
rect 7337 13565 7423 13588
rect 11169 13628 11255 13651
rect 11337 13628 11423 13651
rect 11169 13588 11194 13628
rect 11194 13588 11234 13628
rect 11234 13588 11255 13628
rect 11337 13588 11358 13628
rect 11358 13588 11398 13628
rect 11398 13588 11423 13628
rect 11169 13565 11255 13588
rect 11337 13565 11423 13588
rect 15169 13628 15255 13651
rect 15337 13628 15423 13651
rect 15169 13588 15194 13628
rect 15194 13588 15234 13628
rect 15234 13588 15255 13628
rect 15337 13588 15358 13628
rect 15358 13588 15398 13628
rect 15398 13588 15423 13628
rect 15169 13565 15255 13588
rect 15337 13565 15423 13588
rect 19169 13628 19255 13651
rect 19337 13628 19423 13651
rect 19169 13588 19194 13628
rect 19194 13588 19234 13628
rect 19234 13588 19255 13628
rect 19337 13588 19358 13628
rect 19358 13588 19398 13628
rect 19398 13588 19423 13628
rect 19169 13565 19255 13588
rect 19337 13565 19423 13588
rect 23169 13628 23255 13651
rect 23337 13628 23423 13651
rect 23169 13588 23194 13628
rect 23194 13588 23234 13628
rect 23234 13588 23255 13628
rect 23337 13588 23358 13628
rect 23358 13588 23398 13628
rect 23398 13588 23423 13628
rect 23169 13565 23255 13588
rect 23337 13565 23423 13588
rect 27169 13628 27255 13651
rect 27337 13628 27423 13651
rect 27169 13588 27194 13628
rect 27194 13588 27234 13628
rect 27234 13588 27255 13628
rect 27337 13588 27358 13628
rect 27358 13588 27398 13628
rect 27398 13588 27423 13628
rect 27169 13565 27255 13588
rect 27337 13565 27423 13588
rect 31169 13628 31255 13651
rect 31337 13628 31423 13651
rect 31169 13588 31194 13628
rect 31194 13588 31234 13628
rect 31234 13588 31255 13628
rect 31337 13588 31358 13628
rect 31358 13588 31398 13628
rect 31398 13588 31423 13628
rect 31169 13565 31255 13588
rect 31337 13565 31423 13588
rect 35169 13628 35255 13651
rect 35337 13628 35423 13651
rect 35169 13588 35194 13628
rect 35194 13588 35234 13628
rect 35234 13588 35255 13628
rect 35337 13588 35358 13628
rect 35358 13588 35398 13628
rect 35398 13588 35423 13628
rect 35169 13565 35255 13588
rect 35337 13565 35423 13588
rect 39169 13628 39255 13651
rect 39337 13628 39423 13651
rect 39169 13588 39194 13628
rect 39194 13588 39234 13628
rect 39234 13588 39255 13628
rect 39337 13588 39358 13628
rect 39358 13588 39398 13628
rect 39398 13588 39423 13628
rect 39169 13565 39255 13588
rect 39337 13565 39423 13588
rect 43169 13628 43255 13651
rect 43337 13628 43423 13651
rect 43169 13588 43194 13628
rect 43194 13588 43234 13628
rect 43234 13588 43255 13628
rect 43337 13588 43358 13628
rect 43358 13588 43398 13628
rect 43398 13588 43423 13628
rect 43169 13565 43255 13588
rect 43337 13565 43423 13588
rect 47169 13628 47255 13651
rect 47337 13628 47423 13651
rect 47169 13588 47194 13628
rect 47194 13588 47234 13628
rect 47234 13588 47255 13628
rect 47337 13588 47358 13628
rect 47358 13588 47398 13628
rect 47398 13588 47423 13628
rect 47169 13565 47255 13588
rect 47337 13565 47423 13588
rect 51169 13628 51255 13651
rect 51337 13628 51423 13651
rect 51169 13588 51194 13628
rect 51194 13588 51234 13628
rect 51234 13588 51255 13628
rect 51337 13588 51358 13628
rect 51358 13588 51398 13628
rect 51398 13588 51423 13628
rect 51169 13565 51255 13588
rect 51337 13565 51423 13588
rect 55169 13628 55255 13651
rect 55337 13628 55423 13651
rect 55169 13588 55194 13628
rect 55194 13588 55234 13628
rect 55234 13588 55255 13628
rect 55337 13588 55358 13628
rect 55358 13588 55398 13628
rect 55398 13588 55423 13628
rect 55169 13565 55255 13588
rect 55337 13565 55423 13588
rect 59169 13628 59255 13651
rect 59337 13628 59423 13651
rect 59169 13588 59194 13628
rect 59194 13588 59234 13628
rect 59234 13588 59255 13628
rect 59337 13588 59358 13628
rect 59358 13588 59398 13628
rect 59398 13588 59423 13628
rect 59169 13565 59255 13588
rect 59337 13565 59423 13588
rect 63169 13628 63255 13651
rect 63337 13628 63423 13651
rect 63169 13588 63194 13628
rect 63194 13588 63234 13628
rect 63234 13588 63255 13628
rect 63337 13588 63358 13628
rect 63358 13588 63398 13628
rect 63398 13588 63423 13628
rect 63169 13565 63255 13588
rect 63337 13565 63423 13588
rect 67169 13628 67255 13651
rect 67337 13628 67423 13651
rect 67169 13588 67194 13628
rect 67194 13588 67234 13628
rect 67234 13588 67255 13628
rect 67337 13588 67358 13628
rect 67358 13588 67398 13628
rect 67398 13588 67423 13628
rect 67169 13565 67255 13588
rect 67337 13565 67423 13588
rect 72409 13524 72495 13610
rect 72577 13524 72663 13610
rect 72409 13356 72495 13442
rect 72577 13356 72663 13442
rect 72409 13188 72495 13274
rect 72577 13188 72663 13274
rect 72409 13020 72495 13106
rect 72577 13020 72663 13106
rect 4409 12872 4495 12895
rect 4577 12872 4663 12895
rect 4409 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4495 12872
rect 4577 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4663 12872
rect 4409 12809 4495 12832
rect 4577 12809 4663 12832
rect 8409 12872 8495 12895
rect 8577 12872 8663 12895
rect 8409 12832 8434 12872
rect 8434 12832 8474 12872
rect 8474 12832 8495 12872
rect 8577 12832 8598 12872
rect 8598 12832 8638 12872
rect 8638 12832 8663 12872
rect 8409 12809 8495 12832
rect 8577 12809 8663 12832
rect 12409 12872 12495 12895
rect 12577 12872 12663 12895
rect 12409 12832 12434 12872
rect 12434 12832 12474 12872
rect 12474 12832 12495 12872
rect 12577 12832 12598 12872
rect 12598 12832 12638 12872
rect 12638 12832 12663 12872
rect 12409 12809 12495 12832
rect 12577 12809 12663 12832
rect 16409 12872 16495 12895
rect 16577 12872 16663 12895
rect 16409 12832 16434 12872
rect 16434 12832 16474 12872
rect 16474 12832 16495 12872
rect 16577 12832 16598 12872
rect 16598 12832 16638 12872
rect 16638 12832 16663 12872
rect 16409 12809 16495 12832
rect 16577 12809 16663 12832
rect 20409 12872 20495 12895
rect 20577 12872 20663 12895
rect 20409 12832 20434 12872
rect 20434 12832 20474 12872
rect 20474 12832 20495 12872
rect 20577 12832 20598 12872
rect 20598 12832 20638 12872
rect 20638 12832 20663 12872
rect 20409 12809 20495 12832
rect 20577 12809 20663 12832
rect 24409 12872 24495 12895
rect 24577 12872 24663 12895
rect 24409 12832 24434 12872
rect 24434 12832 24474 12872
rect 24474 12832 24495 12872
rect 24577 12832 24598 12872
rect 24598 12832 24638 12872
rect 24638 12832 24663 12872
rect 24409 12809 24495 12832
rect 24577 12809 24663 12832
rect 28409 12872 28495 12895
rect 28577 12872 28663 12895
rect 28409 12832 28434 12872
rect 28434 12832 28474 12872
rect 28474 12832 28495 12872
rect 28577 12832 28598 12872
rect 28598 12832 28638 12872
rect 28638 12832 28663 12872
rect 28409 12809 28495 12832
rect 28577 12809 28663 12832
rect 32409 12872 32495 12895
rect 32577 12872 32663 12895
rect 32409 12832 32434 12872
rect 32434 12832 32474 12872
rect 32474 12832 32495 12872
rect 32577 12832 32598 12872
rect 32598 12832 32638 12872
rect 32638 12832 32663 12872
rect 32409 12809 32495 12832
rect 32577 12809 32663 12832
rect 36409 12872 36495 12895
rect 36577 12872 36663 12895
rect 36409 12832 36434 12872
rect 36434 12832 36474 12872
rect 36474 12832 36495 12872
rect 36577 12832 36598 12872
rect 36598 12832 36638 12872
rect 36638 12832 36663 12872
rect 36409 12809 36495 12832
rect 36577 12809 36663 12832
rect 40409 12872 40495 12895
rect 40577 12872 40663 12895
rect 40409 12832 40434 12872
rect 40434 12832 40474 12872
rect 40474 12832 40495 12872
rect 40577 12832 40598 12872
rect 40598 12832 40638 12872
rect 40638 12832 40663 12872
rect 40409 12809 40495 12832
rect 40577 12809 40663 12832
rect 44409 12872 44495 12895
rect 44577 12872 44663 12895
rect 44409 12832 44434 12872
rect 44434 12832 44474 12872
rect 44474 12832 44495 12872
rect 44577 12832 44598 12872
rect 44598 12832 44638 12872
rect 44638 12832 44663 12872
rect 44409 12809 44495 12832
rect 44577 12809 44663 12832
rect 48409 12872 48495 12895
rect 48577 12872 48663 12895
rect 48409 12832 48434 12872
rect 48434 12832 48474 12872
rect 48474 12832 48495 12872
rect 48577 12832 48598 12872
rect 48598 12832 48638 12872
rect 48638 12832 48663 12872
rect 48409 12809 48495 12832
rect 48577 12809 48663 12832
rect 52409 12872 52495 12895
rect 52577 12872 52663 12895
rect 52409 12832 52434 12872
rect 52434 12832 52474 12872
rect 52474 12832 52495 12872
rect 52577 12832 52598 12872
rect 52598 12832 52638 12872
rect 52638 12832 52663 12872
rect 52409 12809 52495 12832
rect 52577 12809 52663 12832
rect 56409 12872 56495 12895
rect 56577 12872 56663 12895
rect 56409 12832 56434 12872
rect 56434 12832 56474 12872
rect 56474 12832 56495 12872
rect 56577 12832 56598 12872
rect 56598 12832 56638 12872
rect 56638 12832 56663 12872
rect 56409 12809 56495 12832
rect 56577 12809 56663 12832
rect 60409 12872 60495 12895
rect 60577 12872 60663 12895
rect 60409 12832 60434 12872
rect 60434 12832 60474 12872
rect 60474 12832 60495 12872
rect 60577 12832 60598 12872
rect 60598 12832 60638 12872
rect 60638 12832 60663 12872
rect 60409 12809 60495 12832
rect 60577 12809 60663 12832
rect 64409 12872 64495 12895
rect 64577 12872 64663 12895
rect 64409 12832 64434 12872
rect 64434 12832 64474 12872
rect 64474 12832 64495 12872
rect 64577 12832 64598 12872
rect 64598 12832 64638 12872
rect 64638 12832 64663 12872
rect 64409 12809 64495 12832
rect 64577 12809 64663 12832
rect 68409 12872 68495 12895
rect 68577 12872 68663 12895
rect 76409 15036 76495 15122
rect 76577 15036 76663 15122
rect 76409 14868 76495 14954
rect 76577 14868 76663 14954
rect 76409 14700 76495 14786
rect 76577 14700 76663 14786
rect 76409 14532 76495 14618
rect 76577 14532 76663 14618
rect 76409 14364 76495 14450
rect 76577 14364 76663 14450
rect 76409 14196 76495 14282
rect 76577 14196 76663 14282
rect 76409 14028 76495 14114
rect 76577 14028 76663 14114
rect 76409 13860 76495 13946
rect 76577 13860 76663 13946
rect 76409 13692 76495 13778
rect 76577 13692 76663 13778
rect 76409 13524 76495 13610
rect 76577 13524 76663 13610
rect 76409 13356 76495 13442
rect 76577 13356 76663 13442
rect 76409 13188 76495 13274
rect 76577 13188 76663 13274
rect 76409 13020 76495 13106
rect 76577 13020 76663 13106
rect 80409 15036 80495 15122
rect 80577 15036 80663 15122
rect 80409 14868 80495 14954
rect 80577 14868 80663 14954
rect 80409 14700 80495 14786
rect 80577 14700 80663 14786
rect 80409 14532 80495 14618
rect 80577 14532 80663 14618
rect 80409 14364 80495 14450
rect 80577 14364 80663 14450
rect 80409 14196 80495 14282
rect 80577 14196 80663 14282
rect 80409 14028 80495 14114
rect 80577 14028 80663 14114
rect 80409 13860 80495 13946
rect 80577 13860 80663 13946
rect 80409 13692 80495 13778
rect 80577 13692 80663 13778
rect 80409 13524 80495 13610
rect 80577 13524 80663 13610
rect 80409 13356 80495 13442
rect 80577 13356 80663 13442
rect 80409 13188 80495 13274
rect 80577 13188 80663 13274
rect 80409 13020 80495 13106
rect 80577 13020 80663 13106
rect 84409 15036 84495 15122
rect 84577 15036 84663 15122
rect 84409 14868 84495 14954
rect 84577 14868 84663 14954
rect 84409 14700 84495 14786
rect 84577 14700 84663 14786
rect 84409 14532 84495 14618
rect 84577 14532 84663 14618
rect 84409 14364 84495 14450
rect 84577 14364 84663 14450
rect 84409 14196 84495 14282
rect 84577 14196 84663 14282
rect 84409 14028 84495 14114
rect 84577 14028 84663 14114
rect 84409 13860 84495 13946
rect 84577 13860 84663 13946
rect 84409 13692 84495 13778
rect 84577 13692 84663 13778
rect 84409 13524 84495 13610
rect 84577 13524 84663 13610
rect 84409 13356 84495 13442
rect 84577 13356 84663 13442
rect 84409 13188 84495 13274
rect 84577 13188 84663 13274
rect 84409 13020 84495 13106
rect 84577 13020 84663 13106
rect 88409 15036 88495 15122
rect 88577 15036 88663 15122
rect 88409 14868 88495 14954
rect 88577 14868 88663 14954
rect 88409 14700 88495 14786
rect 88577 14700 88663 14786
rect 88409 14532 88495 14618
rect 88577 14532 88663 14618
rect 88409 14364 88495 14450
rect 88577 14364 88663 14450
rect 88409 14196 88495 14282
rect 88577 14196 88663 14282
rect 88409 14028 88495 14114
rect 88577 14028 88663 14114
rect 88409 13860 88495 13946
rect 88577 13860 88663 13946
rect 88409 13692 88495 13778
rect 88577 13692 88663 13778
rect 88409 13524 88495 13610
rect 88577 13524 88663 13610
rect 88409 13356 88495 13442
rect 88577 13356 88663 13442
rect 88409 13188 88495 13274
rect 88577 13188 88663 13274
rect 88409 13020 88495 13106
rect 88577 13020 88663 13106
rect 92409 15036 92495 15122
rect 92577 15036 92663 15122
rect 92409 14868 92495 14954
rect 92577 14868 92663 14954
rect 92409 14700 92495 14786
rect 92577 14700 92663 14786
rect 92409 14532 92495 14618
rect 92577 14532 92663 14618
rect 92409 14364 92495 14450
rect 92577 14364 92663 14450
rect 92409 14196 92495 14282
rect 92577 14196 92663 14282
rect 92409 14028 92495 14114
rect 92577 14028 92663 14114
rect 92409 13860 92495 13946
rect 92577 13860 92663 13946
rect 92409 13692 92495 13778
rect 92577 13692 92663 13778
rect 92409 13524 92495 13610
rect 92577 13524 92663 13610
rect 92409 13356 92495 13442
rect 92577 13356 92663 13442
rect 92409 13188 92495 13274
rect 92577 13188 92663 13274
rect 92409 13020 92495 13106
rect 92577 13020 92663 13106
rect 96409 15036 96495 15122
rect 96577 15036 96663 15122
rect 96409 14868 96495 14954
rect 96577 14868 96663 14954
rect 96409 14700 96495 14786
rect 96577 14700 96663 14786
rect 96409 14532 96495 14618
rect 96577 14532 96663 14618
rect 96409 14364 96495 14450
rect 96577 14364 96663 14450
rect 96409 14196 96495 14282
rect 96577 14196 96663 14282
rect 96409 14028 96495 14114
rect 96577 14028 96663 14114
rect 96409 13860 96495 13946
rect 96577 13860 96663 13946
rect 96409 13692 96495 13778
rect 96577 13692 96663 13778
rect 96409 13524 96495 13610
rect 96577 13524 96663 13610
rect 96409 13356 96495 13442
rect 96577 13356 96663 13442
rect 96409 13188 96495 13274
rect 96577 13188 96663 13274
rect 96409 13020 96495 13106
rect 96577 13020 96663 13106
rect 68409 12832 68434 12872
rect 68434 12832 68474 12872
rect 68474 12832 68495 12872
rect 68577 12832 68598 12872
rect 68598 12832 68638 12872
rect 68638 12832 68663 12872
rect 68409 12809 68495 12832
rect 68577 12809 68663 12832
rect 75169 12160 75255 12246
rect 75337 12160 75423 12246
rect 3169 12116 3255 12139
rect 3337 12116 3423 12139
rect 3169 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3255 12116
rect 3337 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3423 12116
rect 3169 12053 3255 12076
rect 3337 12053 3423 12076
rect 7169 12116 7255 12139
rect 7337 12116 7423 12139
rect 7169 12076 7194 12116
rect 7194 12076 7234 12116
rect 7234 12076 7255 12116
rect 7337 12076 7358 12116
rect 7358 12076 7398 12116
rect 7398 12076 7423 12116
rect 7169 12053 7255 12076
rect 7337 12053 7423 12076
rect 11169 12116 11255 12139
rect 11337 12116 11423 12139
rect 11169 12076 11194 12116
rect 11194 12076 11234 12116
rect 11234 12076 11255 12116
rect 11337 12076 11358 12116
rect 11358 12076 11398 12116
rect 11398 12076 11423 12116
rect 11169 12053 11255 12076
rect 11337 12053 11423 12076
rect 15169 12116 15255 12139
rect 15337 12116 15423 12139
rect 15169 12076 15194 12116
rect 15194 12076 15234 12116
rect 15234 12076 15255 12116
rect 15337 12076 15358 12116
rect 15358 12076 15398 12116
rect 15398 12076 15423 12116
rect 15169 12053 15255 12076
rect 15337 12053 15423 12076
rect 19169 12116 19255 12139
rect 19337 12116 19423 12139
rect 19169 12076 19194 12116
rect 19194 12076 19234 12116
rect 19234 12076 19255 12116
rect 19337 12076 19358 12116
rect 19358 12076 19398 12116
rect 19398 12076 19423 12116
rect 19169 12053 19255 12076
rect 19337 12053 19423 12076
rect 23169 12116 23255 12139
rect 23337 12116 23423 12139
rect 23169 12076 23194 12116
rect 23194 12076 23234 12116
rect 23234 12076 23255 12116
rect 23337 12076 23358 12116
rect 23358 12076 23398 12116
rect 23398 12076 23423 12116
rect 23169 12053 23255 12076
rect 23337 12053 23423 12076
rect 27169 12116 27255 12139
rect 27337 12116 27423 12139
rect 27169 12076 27194 12116
rect 27194 12076 27234 12116
rect 27234 12076 27255 12116
rect 27337 12076 27358 12116
rect 27358 12076 27398 12116
rect 27398 12076 27423 12116
rect 27169 12053 27255 12076
rect 27337 12053 27423 12076
rect 31169 12116 31255 12139
rect 31337 12116 31423 12139
rect 31169 12076 31194 12116
rect 31194 12076 31234 12116
rect 31234 12076 31255 12116
rect 31337 12076 31358 12116
rect 31358 12076 31398 12116
rect 31398 12076 31423 12116
rect 31169 12053 31255 12076
rect 31337 12053 31423 12076
rect 35169 12116 35255 12139
rect 35337 12116 35423 12139
rect 35169 12076 35194 12116
rect 35194 12076 35234 12116
rect 35234 12076 35255 12116
rect 35337 12076 35358 12116
rect 35358 12076 35398 12116
rect 35398 12076 35423 12116
rect 35169 12053 35255 12076
rect 35337 12053 35423 12076
rect 39169 12116 39255 12139
rect 39337 12116 39423 12139
rect 39169 12076 39194 12116
rect 39194 12076 39234 12116
rect 39234 12076 39255 12116
rect 39337 12076 39358 12116
rect 39358 12076 39398 12116
rect 39398 12076 39423 12116
rect 39169 12053 39255 12076
rect 39337 12053 39423 12076
rect 43169 12116 43255 12139
rect 43337 12116 43423 12139
rect 43169 12076 43194 12116
rect 43194 12076 43234 12116
rect 43234 12076 43255 12116
rect 43337 12076 43358 12116
rect 43358 12076 43398 12116
rect 43398 12076 43423 12116
rect 43169 12053 43255 12076
rect 43337 12053 43423 12076
rect 47169 12116 47255 12139
rect 47337 12116 47423 12139
rect 47169 12076 47194 12116
rect 47194 12076 47234 12116
rect 47234 12076 47255 12116
rect 47337 12076 47358 12116
rect 47358 12076 47398 12116
rect 47398 12076 47423 12116
rect 47169 12053 47255 12076
rect 47337 12053 47423 12076
rect 51169 12116 51255 12139
rect 51337 12116 51423 12139
rect 51169 12076 51194 12116
rect 51194 12076 51234 12116
rect 51234 12076 51255 12116
rect 51337 12076 51358 12116
rect 51358 12076 51398 12116
rect 51398 12076 51423 12116
rect 51169 12053 51255 12076
rect 51337 12053 51423 12076
rect 55169 12116 55255 12139
rect 55337 12116 55423 12139
rect 55169 12076 55194 12116
rect 55194 12076 55234 12116
rect 55234 12076 55255 12116
rect 55337 12076 55358 12116
rect 55358 12076 55398 12116
rect 55398 12076 55423 12116
rect 55169 12053 55255 12076
rect 55337 12053 55423 12076
rect 59169 12116 59255 12139
rect 59337 12116 59423 12139
rect 59169 12076 59194 12116
rect 59194 12076 59234 12116
rect 59234 12076 59255 12116
rect 59337 12076 59358 12116
rect 59358 12076 59398 12116
rect 59398 12076 59423 12116
rect 59169 12053 59255 12076
rect 59337 12053 59423 12076
rect 63169 12116 63255 12139
rect 63337 12116 63423 12139
rect 63169 12076 63194 12116
rect 63194 12076 63234 12116
rect 63234 12076 63255 12116
rect 63337 12076 63358 12116
rect 63358 12076 63398 12116
rect 63398 12076 63423 12116
rect 63169 12053 63255 12076
rect 63337 12053 63423 12076
rect 67169 12116 67255 12139
rect 67337 12116 67423 12139
rect 67169 12076 67194 12116
rect 67194 12076 67234 12116
rect 67234 12076 67255 12116
rect 67337 12076 67358 12116
rect 67358 12076 67398 12116
rect 67398 12076 67423 12116
rect 67169 12053 67255 12076
rect 67337 12053 67423 12076
rect 75169 11992 75255 12078
rect 75337 11992 75423 12078
rect 75169 11824 75255 11910
rect 75337 11824 75423 11910
rect 75169 11656 75255 11742
rect 75337 11656 75423 11742
rect 75169 11488 75255 11574
rect 75337 11488 75423 11574
rect 4409 11360 4495 11383
rect 4577 11360 4663 11383
rect 4409 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4495 11360
rect 4577 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4663 11360
rect 4409 11297 4495 11320
rect 4577 11297 4663 11320
rect 8409 11360 8495 11383
rect 8577 11360 8663 11383
rect 8409 11320 8434 11360
rect 8434 11320 8474 11360
rect 8474 11320 8495 11360
rect 8577 11320 8598 11360
rect 8598 11320 8638 11360
rect 8638 11320 8663 11360
rect 8409 11297 8495 11320
rect 8577 11297 8663 11320
rect 12409 11360 12495 11383
rect 12577 11360 12663 11383
rect 12409 11320 12434 11360
rect 12434 11320 12474 11360
rect 12474 11320 12495 11360
rect 12577 11320 12598 11360
rect 12598 11320 12638 11360
rect 12638 11320 12663 11360
rect 12409 11297 12495 11320
rect 12577 11297 12663 11320
rect 16409 11360 16495 11383
rect 16577 11360 16663 11383
rect 16409 11320 16434 11360
rect 16434 11320 16474 11360
rect 16474 11320 16495 11360
rect 16577 11320 16598 11360
rect 16598 11320 16638 11360
rect 16638 11320 16663 11360
rect 16409 11297 16495 11320
rect 16577 11297 16663 11320
rect 20409 11360 20495 11383
rect 20577 11360 20663 11383
rect 20409 11320 20434 11360
rect 20434 11320 20474 11360
rect 20474 11320 20495 11360
rect 20577 11320 20598 11360
rect 20598 11320 20638 11360
rect 20638 11320 20663 11360
rect 20409 11297 20495 11320
rect 20577 11297 20663 11320
rect 24409 11360 24495 11383
rect 24577 11360 24663 11383
rect 24409 11320 24434 11360
rect 24434 11320 24474 11360
rect 24474 11320 24495 11360
rect 24577 11320 24598 11360
rect 24598 11320 24638 11360
rect 24638 11320 24663 11360
rect 24409 11297 24495 11320
rect 24577 11297 24663 11320
rect 28409 11360 28495 11383
rect 28577 11360 28663 11383
rect 28409 11320 28434 11360
rect 28434 11320 28474 11360
rect 28474 11320 28495 11360
rect 28577 11320 28598 11360
rect 28598 11320 28638 11360
rect 28638 11320 28663 11360
rect 28409 11297 28495 11320
rect 28577 11297 28663 11320
rect 32409 11360 32495 11383
rect 32577 11360 32663 11383
rect 32409 11320 32434 11360
rect 32434 11320 32474 11360
rect 32474 11320 32495 11360
rect 32577 11320 32598 11360
rect 32598 11320 32638 11360
rect 32638 11320 32663 11360
rect 32409 11297 32495 11320
rect 32577 11297 32663 11320
rect 36409 11360 36495 11383
rect 36577 11360 36663 11383
rect 36409 11320 36434 11360
rect 36434 11320 36474 11360
rect 36474 11320 36495 11360
rect 36577 11320 36598 11360
rect 36598 11320 36638 11360
rect 36638 11320 36663 11360
rect 36409 11297 36495 11320
rect 36577 11297 36663 11320
rect 40409 11360 40495 11383
rect 40577 11360 40663 11383
rect 40409 11320 40434 11360
rect 40434 11320 40474 11360
rect 40474 11320 40495 11360
rect 40577 11320 40598 11360
rect 40598 11320 40638 11360
rect 40638 11320 40663 11360
rect 40409 11297 40495 11320
rect 40577 11297 40663 11320
rect 44409 11360 44495 11383
rect 44577 11360 44663 11383
rect 44409 11320 44434 11360
rect 44434 11320 44474 11360
rect 44474 11320 44495 11360
rect 44577 11320 44598 11360
rect 44598 11320 44638 11360
rect 44638 11320 44663 11360
rect 44409 11297 44495 11320
rect 44577 11297 44663 11320
rect 48409 11360 48495 11383
rect 48577 11360 48663 11383
rect 48409 11320 48434 11360
rect 48434 11320 48474 11360
rect 48474 11320 48495 11360
rect 48577 11320 48598 11360
rect 48598 11320 48638 11360
rect 48638 11320 48663 11360
rect 48409 11297 48495 11320
rect 48577 11297 48663 11320
rect 52409 11360 52495 11383
rect 52577 11360 52663 11383
rect 52409 11320 52434 11360
rect 52434 11320 52474 11360
rect 52474 11320 52495 11360
rect 52577 11320 52598 11360
rect 52598 11320 52638 11360
rect 52638 11320 52663 11360
rect 52409 11297 52495 11320
rect 52577 11297 52663 11320
rect 56409 11360 56495 11383
rect 56577 11360 56663 11383
rect 56409 11320 56434 11360
rect 56434 11320 56474 11360
rect 56474 11320 56495 11360
rect 56577 11320 56598 11360
rect 56598 11320 56638 11360
rect 56638 11320 56663 11360
rect 56409 11297 56495 11320
rect 56577 11297 56663 11320
rect 60409 11360 60495 11383
rect 60577 11360 60663 11383
rect 60409 11320 60434 11360
rect 60434 11320 60474 11360
rect 60474 11320 60495 11360
rect 60577 11320 60598 11360
rect 60598 11320 60638 11360
rect 60638 11320 60663 11360
rect 60409 11297 60495 11320
rect 60577 11297 60663 11320
rect 64409 11360 64495 11383
rect 64577 11360 64663 11383
rect 64409 11320 64434 11360
rect 64434 11320 64474 11360
rect 64474 11320 64495 11360
rect 64577 11320 64598 11360
rect 64598 11320 64638 11360
rect 64638 11320 64663 11360
rect 64409 11297 64495 11320
rect 64577 11297 64663 11320
rect 68409 11360 68495 11383
rect 68577 11360 68663 11383
rect 68409 11320 68434 11360
rect 68434 11320 68474 11360
rect 68474 11320 68495 11360
rect 68577 11320 68598 11360
rect 68598 11320 68638 11360
rect 68638 11320 68663 11360
rect 68409 11297 68495 11320
rect 68577 11297 68663 11320
rect 75169 11320 75255 11406
rect 75337 11320 75423 11406
rect 75169 11152 75255 11238
rect 75337 11152 75423 11238
rect 75169 10984 75255 11070
rect 75337 10984 75423 11070
rect 75169 10816 75255 10902
rect 75337 10816 75423 10902
rect 75169 10648 75255 10734
rect 75337 10648 75423 10734
rect 3169 10604 3255 10627
rect 3337 10604 3423 10627
rect 3169 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3255 10604
rect 3337 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3423 10604
rect 3169 10541 3255 10564
rect 3337 10541 3423 10564
rect 7169 10604 7255 10627
rect 7337 10604 7423 10627
rect 7169 10564 7194 10604
rect 7194 10564 7234 10604
rect 7234 10564 7255 10604
rect 7337 10564 7358 10604
rect 7358 10564 7398 10604
rect 7398 10564 7423 10604
rect 7169 10541 7255 10564
rect 7337 10541 7423 10564
rect 11169 10604 11255 10627
rect 11337 10604 11423 10627
rect 11169 10564 11194 10604
rect 11194 10564 11234 10604
rect 11234 10564 11255 10604
rect 11337 10564 11358 10604
rect 11358 10564 11398 10604
rect 11398 10564 11423 10604
rect 11169 10541 11255 10564
rect 11337 10541 11423 10564
rect 15169 10604 15255 10627
rect 15337 10604 15423 10627
rect 15169 10564 15194 10604
rect 15194 10564 15234 10604
rect 15234 10564 15255 10604
rect 15337 10564 15358 10604
rect 15358 10564 15398 10604
rect 15398 10564 15423 10604
rect 15169 10541 15255 10564
rect 15337 10541 15423 10564
rect 19169 10604 19255 10627
rect 19337 10604 19423 10627
rect 19169 10564 19194 10604
rect 19194 10564 19234 10604
rect 19234 10564 19255 10604
rect 19337 10564 19358 10604
rect 19358 10564 19398 10604
rect 19398 10564 19423 10604
rect 19169 10541 19255 10564
rect 19337 10541 19423 10564
rect 23169 10604 23255 10627
rect 23337 10604 23423 10627
rect 23169 10564 23194 10604
rect 23194 10564 23234 10604
rect 23234 10564 23255 10604
rect 23337 10564 23358 10604
rect 23358 10564 23398 10604
rect 23398 10564 23423 10604
rect 23169 10541 23255 10564
rect 23337 10541 23423 10564
rect 27169 10604 27255 10627
rect 27337 10604 27423 10627
rect 27169 10564 27194 10604
rect 27194 10564 27234 10604
rect 27234 10564 27255 10604
rect 27337 10564 27358 10604
rect 27358 10564 27398 10604
rect 27398 10564 27423 10604
rect 27169 10541 27255 10564
rect 27337 10541 27423 10564
rect 31169 10604 31255 10627
rect 31337 10604 31423 10627
rect 31169 10564 31194 10604
rect 31194 10564 31234 10604
rect 31234 10564 31255 10604
rect 31337 10564 31358 10604
rect 31358 10564 31398 10604
rect 31398 10564 31423 10604
rect 31169 10541 31255 10564
rect 31337 10541 31423 10564
rect 35169 10604 35255 10627
rect 35337 10604 35423 10627
rect 35169 10564 35194 10604
rect 35194 10564 35234 10604
rect 35234 10564 35255 10604
rect 35337 10564 35358 10604
rect 35358 10564 35398 10604
rect 35398 10564 35423 10604
rect 35169 10541 35255 10564
rect 35337 10541 35423 10564
rect 39169 10604 39255 10627
rect 39337 10604 39423 10627
rect 39169 10564 39194 10604
rect 39194 10564 39234 10604
rect 39234 10564 39255 10604
rect 39337 10564 39358 10604
rect 39358 10564 39398 10604
rect 39398 10564 39423 10604
rect 39169 10541 39255 10564
rect 39337 10541 39423 10564
rect 43169 10604 43255 10627
rect 43337 10604 43423 10627
rect 43169 10564 43194 10604
rect 43194 10564 43234 10604
rect 43234 10564 43255 10604
rect 43337 10564 43358 10604
rect 43358 10564 43398 10604
rect 43398 10564 43423 10604
rect 43169 10541 43255 10564
rect 43337 10541 43423 10564
rect 47169 10604 47255 10627
rect 47337 10604 47423 10627
rect 47169 10564 47194 10604
rect 47194 10564 47234 10604
rect 47234 10564 47255 10604
rect 47337 10564 47358 10604
rect 47358 10564 47398 10604
rect 47398 10564 47423 10604
rect 47169 10541 47255 10564
rect 47337 10541 47423 10564
rect 51169 10604 51255 10627
rect 51337 10604 51423 10627
rect 51169 10564 51194 10604
rect 51194 10564 51234 10604
rect 51234 10564 51255 10604
rect 51337 10564 51358 10604
rect 51358 10564 51398 10604
rect 51398 10564 51423 10604
rect 51169 10541 51255 10564
rect 51337 10541 51423 10564
rect 55169 10604 55255 10627
rect 55337 10604 55423 10627
rect 55169 10564 55194 10604
rect 55194 10564 55234 10604
rect 55234 10564 55255 10604
rect 55337 10564 55358 10604
rect 55358 10564 55398 10604
rect 55398 10564 55423 10604
rect 55169 10541 55255 10564
rect 55337 10541 55423 10564
rect 59169 10604 59255 10627
rect 59337 10604 59423 10627
rect 59169 10564 59194 10604
rect 59194 10564 59234 10604
rect 59234 10564 59255 10604
rect 59337 10564 59358 10604
rect 59358 10564 59398 10604
rect 59398 10564 59423 10604
rect 59169 10541 59255 10564
rect 59337 10541 59423 10564
rect 63169 10604 63255 10627
rect 63337 10604 63423 10627
rect 63169 10564 63194 10604
rect 63194 10564 63234 10604
rect 63234 10564 63255 10604
rect 63337 10564 63358 10604
rect 63358 10564 63398 10604
rect 63398 10564 63423 10604
rect 63169 10541 63255 10564
rect 63337 10541 63423 10564
rect 67169 10604 67255 10627
rect 67337 10604 67423 10627
rect 67169 10564 67194 10604
rect 67194 10564 67234 10604
rect 67234 10564 67255 10604
rect 67337 10564 67358 10604
rect 67358 10564 67398 10604
rect 67398 10564 67423 10604
rect 67169 10541 67255 10564
rect 67337 10541 67423 10564
rect 75169 10480 75255 10566
rect 75337 10480 75423 10566
rect 75169 10312 75255 10398
rect 75337 10312 75423 10398
rect 75169 10144 75255 10230
rect 75337 10144 75423 10230
rect 79169 12160 79255 12246
rect 79337 12160 79423 12246
rect 79169 11992 79255 12078
rect 79337 11992 79423 12078
rect 79169 11824 79255 11910
rect 79337 11824 79423 11910
rect 79169 11656 79255 11742
rect 79337 11656 79423 11742
rect 79169 11488 79255 11574
rect 79337 11488 79423 11574
rect 79169 11320 79255 11406
rect 79337 11320 79423 11406
rect 79169 11152 79255 11238
rect 79337 11152 79423 11238
rect 79169 10984 79255 11070
rect 79337 10984 79423 11070
rect 79169 10816 79255 10902
rect 79337 10816 79423 10902
rect 79169 10648 79255 10734
rect 79337 10648 79423 10734
rect 79169 10480 79255 10566
rect 79337 10480 79423 10566
rect 79169 10312 79255 10398
rect 79337 10312 79423 10398
rect 79169 10144 79255 10230
rect 79337 10144 79423 10230
rect 83169 12160 83255 12246
rect 83337 12160 83423 12246
rect 83169 11992 83255 12078
rect 83337 11992 83423 12078
rect 83169 11824 83255 11910
rect 83337 11824 83423 11910
rect 83169 11656 83255 11742
rect 83337 11656 83423 11742
rect 83169 11488 83255 11574
rect 83337 11488 83423 11574
rect 83169 11320 83255 11406
rect 83337 11320 83423 11406
rect 83169 11152 83255 11238
rect 83337 11152 83423 11238
rect 83169 10984 83255 11070
rect 83337 10984 83423 11070
rect 83169 10816 83255 10902
rect 83337 10816 83423 10902
rect 83169 10648 83255 10734
rect 83337 10648 83423 10734
rect 83169 10480 83255 10566
rect 83337 10480 83423 10566
rect 83169 10312 83255 10398
rect 83337 10312 83423 10398
rect 83169 10144 83255 10230
rect 83337 10144 83423 10230
rect 87169 12160 87255 12246
rect 87337 12160 87423 12246
rect 87169 11992 87255 12078
rect 87337 11992 87423 12078
rect 87169 11824 87255 11910
rect 87337 11824 87423 11910
rect 87169 11656 87255 11742
rect 87337 11656 87423 11742
rect 87169 11488 87255 11574
rect 87337 11488 87423 11574
rect 87169 11320 87255 11406
rect 87337 11320 87423 11406
rect 87169 11152 87255 11238
rect 87337 11152 87423 11238
rect 87169 10984 87255 11070
rect 87337 10984 87423 11070
rect 87169 10816 87255 10902
rect 87337 10816 87423 10902
rect 87169 10648 87255 10734
rect 87337 10648 87423 10734
rect 87169 10480 87255 10566
rect 87337 10480 87423 10566
rect 87169 10312 87255 10398
rect 87337 10312 87423 10398
rect 87169 10144 87255 10230
rect 87337 10144 87423 10230
rect 91169 12160 91255 12246
rect 91337 12160 91423 12246
rect 91169 11992 91255 12078
rect 91337 11992 91423 12078
rect 91169 11824 91255 11910
rect 91337 11824 91423 11910
rect 91169 11656 91255 11742
rect 91337 11656 91423 11742
rect 91169 11488 91255 11574
rect 91337 11488 91423 11574
rect 91169 11320 91255 11406
rect 91337 11320 91423 11406
rect 91169 11152 91255 11238
rect 91337 11152 91423 11238
rect 91169 10984 91255 11070
rect 91337 10984 91423 11070
rect 91169 10816 91255 10902
rect 91337 10816 91423 10902
rect 91169 10648 91255 10734
rect 91337 10648 91423 10734
rect 91169 10480 91255 10566
rect 91337 10480 91423 10566
rect 91169 10312 91255 10398
rect 91337 10312 91423 10398
rect 91169 10144 91255 10230
rect 91337 10144 91423 10230
rect 95169 12160 95255 12246
rect 95337 12160 95423 12246
rect 95169 11992 95255 12078
rect 95337 11992 95423 12078
rect 95169 11824 95255 11910
rect 95337 11824 95423 11910
rect 95169 11656 95255 11742
rect 95337 11656 95423 11742
rect 95169 11488 95255 11574
rect 95337 11488 95423 11574
rect 95169 11320 95255 11406
rect 95337 11320 95423 11406
rect 95169 11152 95255 11238
rect 95337 11152 95423 11238
rect 95169 10984 95255 11070
rect 95337 10984 95423 11070
rect 95169 10816 95255 10902
rect 95337 10816 95423 10902
rect 95169 10648 95255 10734
rect 95337 10648 95423 10734
rect 95169 10480 95255 10566
rect 95337 10480 95423 10566
rect 95169 10312 95255 10398
rect 95337 10312 95423 10398
rect 95169 10144 95255 10230
rect 95337 10144 95423 10230
rect 4409 9848 4495 9871
rect 4577 9848 4663 9871
rect 4409 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4495 9848
rect 4577 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4663 9848
rect 4409 9785 4495 9808
rect 4577 9785 4663 9808
rect 8409 9848 8495 9871
rect 8577 9848 8663 9871
rect 8409 9808 8434 9848
rect 8434 9808 8474 9848
rect 8474 9808 8495 9848
rect 8577 9808 8598 9848
rect 8598 9808 8638 9848
rect 8638 9808 8663 9848
rect 8409 9785 8495 9808
rect 8577 9785 8663 9808
rect 12409 9848 12495 9871
rect 12577 9848 12663 9871
rect 12409 9808 12434 9848
rect 12434 9808 12474 9848
rect 12474 9808 12495 9848
rect 12577 9808 12598 9848
rect 12598 9808 12638 9848
rect 12638 9808 12663 9848
rect 12409 9785 12495 9808
rect 12577 9785 12663 9808
rect 16409 9848 16495 9871
rect 16577 9848 16663 9871
rect 16409 9808 16434 9848
rect 16434 9808 16474 9848
rect 16474 9808 16495 9848
rect 16577 9808 16598 9848
rect 16598 9808 16638 9848
rect 16638 9808 16663 9848
rect 16409 9785 16495 9808
rect 16577 9785 16663 9808
rect 20409 9848 20495 9871
rect 20577 9848 20663 9871
rect 20409 9808 20434 9848
rect 20434 9808 20474 9848
rect 20474 9808 20495 9848
rect 20577 9808 20598 9848
rect 20598 9808 20638 9848
rect 20638 9808 20663 9848
rect 20409 9785 20495 9808
rect 20577 9785 20663 9808
rect 24409 9848 24495 9871
rect 24577 9848 24663 9871
rect 24409 9808 24434 9848
rect 24434 9808 24474 9848
rect 24474 9808 24495 9848
rect 24577 9808 24598 9848
rect 24598 9808 24638 9848
rect 24638 9808 24663 9848
rect 24409 9785 24495 9808
rect 24577 9785 24663 9808
rect 28409 9848 28495 9871
rect 28577 9848 28663 9871
rect 28409 9808 28434 9848
rect 28434 9808 28474 9848
rect 28474 9808 28495 9848
rect 28577 9808 28598 9848
rect 28598 9808 28638 9848
rect 28638 9808 28663 9848
rect 28409 9785 28495 9808
rect 28577 9785 28663 9808
rect 32409 9848 32495 9871
rect 32577 9848 32663 9871
rect 32409 9808 32434 9848
rect 32434 9808 32474 9848
rect 32474 9808 32495 9848
rect 32577 9808 32598 9848
rect 32598 9808 32638 9848
rect 32638 9808 32663 9848
rect 32409 9785 32495 9808
rect 32577 9785 32663 9808
rect 36409 9848 36495 9871
rect 36577 9848 36663 9871
rect 36409 9808 36434 9848
rect 36434 9808 36474 9848
rect 36474 9808 36495 9848
rect 36577 9808 36598 9848
rect 36598 9808 36638 9848
rect 36638 9808 36663 9848
rect 36409 9785 36495 9808
rect 36577 9785 36663 9808
rect 40409 9848 40495 9871
rect 40577 9848 40663 9871
rect 40409 9808 40434 9848
rect 40434 9808 40474 9848
rect 40474 9808 40495 9848
rect 40577 9808 40598 9848
rect 40598 9808 40638 9848
rect 40638 9808 40663 9848
rect 40409 9785 40495 9808
rect 40577 9785 40663 9808
rect 44409 9848 44495 9871
rect 44577 9848 44663 9871
rect 44409 9808 44434 9848
rect 44434 9808 44474 9848
rect 44474 9808 44495 9848
rect 44577 9808 44598 9848
rect 44598 9808 44638 9848
rect 44638 9808 44663 9848
rect 44409 9785 44495 9808
rect 44577 9785 44663 9808
rect 48409 9848 48495 9871
rect 48577 9848 48663 9871
rect 48409 9808 48434 9848
rect 48434 9808 48474 9848
rect 48474 9808 48495 9848
rect 48577 9808 48598 9848
rect 48598 9808 48638 9848
rect 48638 9808 48663 9848
rect 48409 9785 48495 9808
rect 48577 9785 48663 9808
rect 52409 9848 52495 9871
rect 52577 9848 52663 9871
rect 52409 9808 52434 9848
rect 52434 9808 52474 9848
rect 52474 9808 52495 9848
rect 52577 9808 52598 9848
rect 52598 9808 52638 9848
rect 52638 9808 52663 9848
rect 52409 9785 52495 9808
rect 52577 9785 52663 9808
rect 56409 9848 56495 9871
rect 56577 9848 56663 9871
rect 56409 9808 56434 9848
rect 56434 9808 56474 9848
rect 56474 9808 56495 9848
rect 56577 9808 56598 9848
rect 56598 9808 56638 9848
rect 56638 9808 56663 9848
rect 56409 9785 56495 9808
rect 56577 9785 56663 9808
rect 60409 9848 60495 9871
rect 60577 9848 60663 9871
rect 60409 9808 60434 9848
rect 60434 9808 60474 9848
rect 60474 9808 60495 9848
rect 60577 9808 60598 9848
rect 60598 9808 60638 9848
rect 60638 9808 60663 9848
rect 60409 9785 60495 9808
rect 60577 9785 60663 9808
rect 64409 9848 64495 9871
rect 64577 9848 64663 9871
rect 64409 9808 64434 9848
rect 64434 9808 64474 9848
rect 64474 9808 64495 9848
rect 64577 9808 64598 9848
rect 64598 9808 64638 9848
rect 64638 9808 64663 9848
rect 64409 9785 64495 9808
rect 64577 9785 64663 9808
rect 68409 9848 68495 9871
rect 68577 9848 68663 9871
rect 68409 9808 68434 9848
rect 68434 9808 68474 9848
rect 68474 9808 68495 9848
rect 68577 9808 68598 9848
rect 68598 9808 68638 9848
rect 68638 9808 68663 9848
rect 68409 9785 68495 9808
rect 68577 9785 68663 9808
rect 3169 9092 3255 9115
rect 3337 9092 3423 9115
rect 3169 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3255 9092
rect 3337 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3423 9092
rect 3169 9029 3255 9052
rect 3337 9029 3423 9052
rect 7169 9092 7255 9115
rect 7337 9092 7423 9115
rect 7169 9052 7194 9092
rect 7194 9052 7234 9092
rect 7234 9052 7255 9092
rect 7337 9052 7358 9092
rect 7358 9052 7398 9092
rect 7398 9052 7423 9092
rect 7169 9029 7255 9052
rect 7337 9029 7423 9052
rect 11169 9092 11255 9115
rect 11337 9092 11423 9115
rect 11169 9052 11194 9092
rect 11194 9052 11234 9092
rect 11234 9052 11255 9092
rect 11337 9052 11358 9092
rect 11358 9052 11398 9092
rect 11398 9052 11423 9092
rect 11169 9029 11255 9052
rect 11337 9029 11423 9052
rect 15169 9092 15255 9115
rect 15337 9092 15423 9115
rect 15169 9052 15194 9092
rect 15194 9052 15234 9092
rect 15234 9052 15255 9092
rect 15337 9052 15358 9092
rect 15358 9052 15398 9092
rect 15398 9052 15423 9092
rect 15169 9029 15255 9052
rect 15337 9029 15423 9052
rect 19169 9092 19255 9115
rect 19337 9092 19423 9115
rect 19169 9052 19194 9092
rect 19194 9052 19234 9092
rect 19234 9052 19255 9092
rect 19337 9052 19358 9092
rect 19358 9052 19398 9092
rect 19398 9052 19423 9092
rect 19169 9029 19255 9052
rect 19337 9029 19423 9052
rect 23169 9092 23255 9115
rect 23337 9092 23423 9115
rect 23169 9052 23194 9092
rect 23194 9052 23234 9092
rect 23234 9052 23255 9092
rect 23337 9052 23358 9092
rect 23358 9052 23398 9092
rect 23398 9052 23423 9092
rect 23169 9029 23255 9052
rect 23337 9029 23423 9052
rect 27169 9092 27255 9115
rect 27337 9092 27423 9115
rect 27169 9052 27194 9092
rect 27194 9052 27234 9092
rect 27234 9052 27255 9092
rect 27337 9052 27358 9092
rect 27358 9052 27398 9092
rect 27398 9052 27423 9092
rect 27169 9029 27255 9052
rect 27337 9029 27423 9052
rect 31169 9092 31255 9115
rect 31337 9092 31423 9115
rect 31169 9052 31194 9092
rect 31194 9052 31234 9092
rect 31234 9052 31255 9092
rect 31337 9052 31358 9092
rect 31358 9052 31398 9092
rect 31398 9052 31423 9092
rect 31169 9029 31255 9052
rect 31337 9029 31423 9052
rect 35169 9092 35255 9115
rect 35337 9092 35423 9115
rect 35169 9052 35194 9092
rect 35194 9052 35234 9092
rect 35234 9052 35255 9092
rect 35337 9052 35358 9092
rect 35358 9052 35398 9092
rect 35398 9052 35423 9092
rect 35169 9029 35255 9052
rect 35337 9029 35423 9052
rect 39169 9092 39255 9115
rect 39337 9092 39423 9115
rect 39169 9052 39194 9092
rect 39194 9052 39234 9092
rect 39234 9052 39255 9092
rect 39337 9052 39358 9092
rect 39358 9052 39398 9092
rect 39398 9052 39423 9092
rect 39169 9029 39255 9052
rect 39337 9029 39423 9052
rect 43169 9092 43255 9115
rect 43337 9092 43423 9115
rect 43169 9052 43194 9092
rect 43194 9052 43234 9092
rect 43234 9052 43255 9092
rect 43337 9052 43358 9092
rect 43358 9052 43398 9092
rect 43398 9052 43423 9092
rect 43169 9029 43255 9052
rect 43337 9029 43423 9052
rect 47169 9092 47255 9115
rect 47337 9092 47423 9115
rect 47169 9052 47194 9092
rect 47194 9052 47234 9092
rect 47234 9052 47255 9092
rect 47337 9052 47358 9092
rect 47358 9052 47398 9092
rect 47398 9052 47423 9092
rect 47169 9029 47255 9052
rect 47337 9029 47423 9052
rect 51169 9092 51255 9115
rect 51337 9092 51423 9115
rect 51169 9052 51194 9092
rect 51194 9052 51234 9092
rect 51234 9052 51255 9092
rect 51337 9052 51358 9092
rect 51358 9052 51398 9092
rect 51398 9052 51423 9092
rect 51169 9029 51255 9052
rect 51337 9029 51423 9052
rect 55169 9092 55255 9115
rect 55337 9092 55423 9115
rect 55169 9052 55194 9092
rect 55194 9052 55234 9092
rect 55234 9052 55255 9092
rect 55337 9052 55358 9092
rect 55358 9052 55398 9092
rect 55398 9052 55423 9092
rect 55169 9029 55255 9052
rect 55337 9029 55423 9052
rect 59169 9092 59255 9115
rect 59337 9092 59423 9115
rect 59169 9052 59194 9092
rect 59194 9052 59234 9092
rect 59234 9052 59255 9092
rect 59337 9052 59358 9092
rect 59358 9052 59398 9092
rect 59398 9052 59423 9092
rect 59169 9029 59255 9052
rect 59337 9029 59423 9052
rect 63169 9092 63255 9115
rect 63337 9092 63423 9115
rect 63169 9052 63194 9092
rect 63194 9052 63234 9092
rect 63234 9052 63255 9092
rect 63337 9052 63358 9092
rect 63358 9052 63398 9092
rect 63398 9052 63423 9092
rect 63169 9029 63255 9052
rect 63337 9029 63423 9052
rect 67169 9092 67255 9115
rect 67337 9092 67423 9115
rect 67169 9052 67194 9092
rect 67194 9052 67234 9092
rect 67234 9052 67255 9092
rect 67337 9052 67358 9092
rect 67358 9052 67398 9092
rect 67398 9052 67423 9092
rect 67169 9029 67255 9052
rect 67337 9029 67423 9052
rect 4409 8336 4495 8359
rect 4577 8336 4663 8359
rect 4409 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4495 8336
rect 4577 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4663 8336
rect 4409 8273 4495 8296
rect 4577 8273 4663 8296
rect 8409 8336 8495 8359
rect 8577 8336 8663 8359
rect 8409 8296 8434 8336
rect 8434 8296 8474 8336
rect 8474 8296 8495 8336
rect 8577 8296 8598 8336
rect 8598 8296 8638 8336
rect 8638 8296 8663 8336
rect 8409 8273 8495 8296
rect 8577 8273 8663 8296
rect 12409 8336 12495 8359
rect 12577 8336 12663 8359
rect 12409 8296 12434 8336
rect 12434 8296 12474 8336
rect 12474 8296 12495 8336
rect 12577 8296 12598 8336
rect 12598 8296 12638 8336
rect 12638 8296 12663 8336
rect 12409 8273 12495 8296
rect 12577 8273 12663 8296
rect 16409 8336 16495 8359
rect 16577 8336 16663 8359
rect 16409 8296 16434 8336
rect 16434 8296 16474 8336
rect 16474 8296 16495 8336
rect 16577 8296 16598 8336
rect 16598 8296 16638 8336
rect 16638 8296 16663 8336
rect 16409 8273 16495 8296
rect 16577 8273 16663 8296
rect 20409 8336 20495 8359
rect 20577 8336 20663 8359
rect 20409 8296 20434 8336
rect 20434 8296 20474 8336
rect 20474 8296 20495 8336
rect 20577 8296 20598 8336
rect 20598 8296 20638 8336
rect 20638 8296 20663 8336
rect 20409 8273 20495 8296
rect 20577 8273 20663 8296
rect 24409 8336 24495 8359
rect 24577 8336 24663 8359
rect 24409 8296 24434 8336
rect 24434 8296 24474 8336
rect 24474 8296 24495 8336
rect 24577 8296 24598 8336
rect 24598 8296 24638 8336
rect 24638 8296 24663 8336
rect 24409 8273 24495 8296
rect 24577 8273 24663 8296
rect 28409 8336 28495 8359
rect 28577 8336 28663 8359
rect 28409 8296 28434 8336
rect 28434 8296 28474 8336
rect 28474 8296 28495 8336
rect 28577 8296 28598 8336
rect 28598 8296 28638 8336
rect 28638 8296 28663 8336
rect 28409 8273 28495 8296
rect 28577 8273 28663 8296
rect 32409 8336 32495 8359
rect 32577 8336 32663 8359
rect 32409 8296 32434 8336
rect 32434 8296 32474 8336
rect 32474 8296 32495 8336
rect 32577 8296 32598 8336
rect 32598 8296 32638 8336
rect 32638 8296 32663 8336
rect 32409 8273 32495 8296
rect 32577 8273 32663 8296
rect 36409 8336 36495 8359
rect 36577 8336 36663 8359
rect 36409 8296 36434 8336
rect 36434 8296 36474 8336
rect 36474 8296 36495 8336
rect 36577 8296 36598 8336
rect 36598 8296 36638 8336
rect 36638 8296 36663 8336
rect 36409 8273 36495 8296
rect 36577 8273 36663 8296
rect 40409 8336 40495 8359
rect 40577 8336 40663 8359
rect 40409 8296 40434 8336
rect 40434 8296 40474 8336
rect 40474 8296 40495 8336
rect 40577 8296 40598 8336
rect 40598 8296 40638 8336
rect 40638 8296 40663 8336
rect 40409 8273 40495 8296
rect 40577 8273 40663 8296
rect 44409 8336 44495 8359
rect 44577 8336 44663 8359
rect 44409 8296 44434 8336
rect 44434 8296 44474 8336
rect 44474 8296 44495 8336
rect 44577 8296 44598 8336
rect 44598 8296 44638 8336
rect 44638 8296 44663 8336
rect 44409 8273 44495 8296
rect 44577 8273 44663 8296
rect 48409 8336 48495 8359
rect 48577 8336 48663 8359
rect 48409 8296 48434 8336
rect 48434 8296 48474 8336
rect 48474 8296 48495 8336
rect 48577 8296 48598 8336
rect 48598 8296 48638 8336
rect 48638 8296 48663 8336
rect 48409 8273 48495 8296
rect 48577 8273 48663 8296
rect 52409 8336 52495 8359
rect 52577 8336 52663 8359
rect 52409 8296 52434 8336
rect 52434 8296 52474 8336
rect 52474 8296 52495 8336
rect 52577 8296 52598 8336
rect 52598 8296 52638 8336
rect 52638 8296 52663 8336
rect 52409 8273 52495 8296
rect 52577 8273 52663 8296
rect 56409 8336 56495 8359
rect 56577 8336 56663 8359
rect 56409 8296 56434 8336
rect 56434 8296 56474 8336
rect 56474 8296 56495 8336
rect 56577 8296 56598 8336
rect 56598 8296 56638 8336
rect 56638 8296 56663 8336
rect 56409 8273 56495 8296
rect 56577 8273 56663 8296
rect 60409 8336 60495 8359
rect 60577 8336 60663 8359
rect 60409 8296 60434 8336
rect 60434 8296 60474 8336
rect 60474 8296 60495 8336
rect 60577 8296 60598 8336
rect 60598 8296 60638 8336
rect 60638 8296 60663 8336
rect 60409 8273 60495 8296
rect 60577 8273 60663 8296
rect 64409 8336 64495 8359
rect 64577 8336 64663 8359
rect 64409 8296 64434 8336
rect 64434 8296 64474 8336
rect 64474 8296 64495 8336
rect 64577 8296 64598 8336
rect 64598 8296 64638 8336
rect 64638 8296 64663 8336
rect 64409 8273 64495 8296
rect 64577 8273 64663 8296
rect 68409 8336 68495 8359
rect 68577 8336 68663 8359
rect 68409 8296 68434 8336
rect 68434 8296 68474 8336
rect 68474 8296 68495 8336
rect 68577 8296 68598 8336
rect 68598 8296 68638 8336
rect 68638 8296 68663 8336
rect 68409 8273 68495 8296
rect 68577 8273 68663 8296
rect 3169 7580 3255 7603
rect 3337 7580 3423 7603
rect 3169 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3255 7580
rect 3337 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3423 7580
rect 3169 7517 3255 7540
rect 3337 7517 3423 7540
rect 7169 7580 7255 7603
rect 7337 7580 7423 7603
rect 7169 7540 7194 7580
rect 7194 7540 7234 7580
rect 7234 7540 7255 7580
rect 7337 7540 7358 7580
rect 7358 7540 7398 7580
rect 7398 7540 7423 7580
rect 7169 7517 7255 7540
rect 7337 7517 7423 7540
rect 11169 7580 11255 7603
rect 11337 7580 11423 7603
rect 11169 7540 11194 7580
rect 11194 7540 11234 7580
rect 11234 7540 11255 7580
rect 11337 7540 11358 7580
rect 11358 7540 11398 7580
rect 11398 7540 11423 7580
rect 11169 7517 11255 7540
rect 11337 7517 11423 7540
rect 15169 7580 15255 7603
rect 15337 7580 15423 7603
rect 15169 7540 15194 7580
rect 15194 7540 15234 7580
rect 15234 7540 15255 7580
rect 15337 7540 15358 7580
rect 15358 7540 15398 7580
rect 15398 7540 15423 7580
rect 15169 7517 15255 7540
rect 15337 7517 15423 7540
rect 19169 7580 19255 7603
rect 19337 7580 19423 7603
rect 19169 7540 19194 7580
rect 19194 7540 19234 7580
rect 19234 7540 19255 7580
rect 19337 7540 19358 7580
rect 19358 7540 19398 7580
rect 19398 7540 19423 7580
rect 19169 7517 19255 7540
rect 19337 7517 19423 7540
rect 23169 7580 23255 7603
rect 23337 7580 23423 7603
rect 23169 7540 23194 7580
rect 23194 7540 23234 7580
rect 23234 7540 23255 7580
rect 23337 7540 23358 7580
rect 23358 7540 23398 7580
rect 23398 7540 23423 7580
rect 23169 7517 23255 7540
rect 23337 7517 23423 7540
rect 27169 7580 27255 7603
rect 27337 7580 27423 7603
rect 27169 7540 27194 7580
rect 27194 7540 27234 7580
rect 27234 7540 27255 7580
rect 27337 7540 27358 7580
rect 27358 7540 27398 7580
rect 27398 7540 27423 7580
rect 27169 7517 27255 7540
rect 27337 7517 27423 7540
rect 31169 7580 31255 7603
rect 31337 7580 31423 7603
rect 31169 7540 31194 7580
rect 31194 7540 31234 7580
rect 31234 7540 31255 7580
rect 31337 7540 31358 7580
rect 31358 7540 31398 7580
rect 31398 7540 31423 7580
rect 31169 7517 31255 7540
rect 31337 7517 31423 7540
rect 35169 7580 35255 7603
rect 35337 7580 35423 7603
rect 35169 7540 35194 7580
rect 35194 7540 35234 7580
rect 35234 7540 35255 7580
rect 35337 7540 35358 7580
rect 35358 7540 35398 7580
rect 35398 7540 35423 7580
rect 35169 7517 35255 7540
rect 35337 7517 35423 7540
rect 39169 7580 39255 7603
rect 39337 7580 39423 7603
rect 39169 7540 39194 7580
rect 39194 7540 39234 7580
rect 39234 7540 39255 7580
rect 39337 7540 39358 7580
rect 39358 7540 39398 7580
rect 39398 7540 39423 7580
rect 39169 7517 39255 7540
rect 39337 7517 39423 7540
rect 43169 7580 43255 7603
rect 43337 7580 43423 7603
rect 43169 7540 43194 7580
rect 43194 7540 43234 7580
rect 43234 7540 43255 7580
rect 43337 7540 43358 7580
rect 43358 7540 43398 7580
rect 43398 7540 43423 7580
rect 43169 7517 43255 7540
rect 43337 7517 43423 7540
rect 47169 7580 47255 7603
rect 47337 7580 47423 7603
rect 47169 7540 47194 7580
rect 47194 7540 47234 7580
rect 47234 7540 47255 7580
rect 47337 7540 47358 7580
rect 47358 7540 47398 7580
rect 47398 7540 47423 7580
rect 47169 7517 47255 7540
rect 47337 7517 47423 7540
rect 51169 7580 51255 7603
rect 51337 7580 51423 7603
rect 51169 7540 51194 7580
rect 51194 7540 51234 7580
rect 51234 7540 51255 7580
rect 51337 7540 51358 7580
rect 51358 7540 51398 7580
rect 51398 7540 51423 7580
rect 51169 7517 51255 7540
rect 51337 7517 51423 7540
rect 55169 7580 55255 7603
rect 55337 7580 55423 7603
rect 55169 7540 55194 7580
rect 55194 7540 55234 7580
rect 55234 7540 55255 7580
rect 55337 7540 55358 7580
rect 55358 7540 55398 7580
rect 55398 7540 55423 7580
rect 55169 7517 55255 7540
rect 55337 7517 55423 7540
rect 59169 7580 59255 7603
rect 59337 7580 59423 7603
rect 59169 7540 59194 7580
rect 59194 7540 59234 7580
rect 59234 7540 59255 7580
rect 59337 7540 59358 7580
rect 59358 7540 59398 7580
rect 59398 7540 59423 7580
rect 59169 7517 59255 7540
rect 59337 7517 59423 7540
rect 63169 7580 63255 7603
rect 63337 7580 63423 7603
rect 63169 7540 63194 7580
rect 63194 7540 63234 7580
rect 63234 7540 63255 7580
rect 63337 7540 63358 7580
rect 63358 7540 63398 7580
rect 63398 7540 63423 7580
rect 63169 7517 63255 7540
rect 63337 7517 63423 7540
rect 67169 7580 67255 7603
rect 67337 7580 67423 7603
rect 67169 7540 67194 7580
rect 67194 7540 67234 7580
rect 67234 7540 67255 7580
rect 67337 7540 67358 7580
rect 67358 7540 67398 7580
rect 67398 7540 67423 7580
rect 67169 7517 67255 7540
rect 67337 7517 67423 7540
rect 71169 7580 71255 7603
rect 71337 7580 71423 7603
rect 71169 7540 71194 7580
rect 71194 7540 71234 7580
rect 71234 7540 71255 7580
rect 71337 7540 71358 7580
rect 71358 7540 71398 7580
rect 71398 7540 71423 7580
rect 71169 7517 71255 7540
rect 71337 7517 71423 7540
rect 75169 7580 75255 7603
rect 75337 7580 75423 7603
rect 75169 7540 75194 7580
rect 75194 7540 75234 7580
rect 75234 7540 75255 7580
rect 75337 7540 75358 7580
rect 75358 7540 75398 7580
rect 75398 7540 75423 7580
rect 75169 7517 75255 7540
rect 75337 7517 75423 7540
rect 79169 7580 79255 7603
rect 79337 7580 79423 7603
rect 79169 7540 79194 7580
rect 79194 7540 79234 7580
rect 79234 7540 79255 7580
rect 79337 7540 79358 7580
rect 79358 7540 79398 7580
rect 79398 7540 79423 7580
rect 79169 7517 79255 7540
rect 79337 7517 79423 7540
rect 83169 7580 83255 7603
rect 83337 7580 83423 7603
rect 83169 7540 83194 7580
rect 83194 7540 83234 7580
rect 83234 7540 83255 7580
rect 83337 7540 83358 7580
rect 83358 7540 83398 7580
rect 83398 7540 83423 7580
rect 83169 7517 83255 7540
rect 83337 7517 83423 7540
rect 87169 7580 87255 7603
rect 87337 7580 87423 7603
rect 87169 7540 87194 7580
rect 87194 7540 87234 7580
rect 87234 7540 87255 7580
rect 87337 7540 87358 7580
rect 87358 7540 87398 7580
rect 87398 7540 87423 7580
rect 87169 7517 87255 7540
rect 87337 7517 87423 7540
rect 91169 7580 91255 7603
rect 91337 7580 91423 7603
rect 91169 7540 91194 7580
rect 91194 7540 91234 7580
rect 91234 7540 91255 7580
rect 91337 7540 91358 7580
rect 91358 7540 91398 7580
rect 91398 7540 91423 7580
rect 91169 7517 91255 7540
rect 91337 7517 91423 7540
rect 95169 7580 95255 7603
rect 95337 7580 95423 7603
rect 95169 7540 95194 7580
rect 95194 7540 95234 7580
rect 95234 7540 95255 7580
rect 95337 7540 95358 7580
rect 95358 7540 95398 7580
rect 95398 7540 95423 7580
rect 95169 7517 95255 7540
rect 95337 7517 95423 7540
rect 99169 7580 99255 7603
rect 99337 7580 99423 7603
rect 99169 7540 99194 7580
rect 99194 7540 99234 7580
rect 99234 7540 99255 7580
rect 99337 7540 99358 7580
rect 99358 7540 99398 7580
rect 99398 7540 99423 7580
rect 99169 7517 99255 7540
rect 99337 7517 99423 7540
rect 86469 7349 86555 7435
rect 4409 6824 4495 6847
rect 4577 6824 4663 6847
rect 4409 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4495 6824
rect 4577 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4663 6824
rect 4409 6761 4495 6784
rect 4577 6761 4663 6784
rect 8409 6824 8495 6847
rect 8577 6824 8663 6847
rect 8409 6784 8434 6824
rect 8434 6784 8474 6824
rect 8474 6784 8495 6824
rect 8577 6784 8598 6824
rect 8598 6784 8638 6824
rect 8638 6784 8663 6824
rect 8409 6761 8495 6784
rect 8577 6761 8663 6784
rect 12409 6824 12495 6847
rect 12577 6824 12663 6847
rect 12409 6784 12434 6824
rect 12434 6784 12474 6824
rect 12474 6784 12495 6824
rect 12577 6784 12598 6824
rect 12598 6784 12638 6824
rect 12638 6784 12663 6824
rect 12409 6761 12495 6784
rect 12577 6761 12663 6784
rect 16409 6824 16495 6847
rect 16577 6824 16663 6847
rect 16409 6784 16434 6824
rect 16434 6784 16474 6824
rect 16474 6784 16495 6824
rect 16577 6784 16598 6824
rect 16598 6784 16638 6824
rect 16638 6784 16663 6824
rect 16409 6761 16495 6784
rect 16577 6761 16663 6784
rect 20409 6824 20495 6847
rect 20577 6824 20663 6847
rect 20409 6784 20434 6824
rect 20434 6784 20474 6824
rect 20474 6784 20495 6824
rect 20577 6784 20598 6824
rect 20598 6784 20638 6824
rect 20638 6784 20663 6824
rect 20409 6761 20495 6784
rect 20577 6761 20663 6784
rect 24409 6824 24495 6847
rect 24577 6824 24663 6847
rect 24409 6784 24434 6824
rect 24434 6784 24474 6824
rect 24474 6784 24495 6824
rect 24577 6784 24598 6824
rect 24598 6784 24638 6824
rect 24638 6784 24663 6824
rect 24409 6761 24495 6784
rect 24577 6761 24663 6784
rect 28409 6824 28495 6847
rect 28577 6824 28663 6847
rect 28409 6784 28434 6824
rect 28434 6784 28474 6824
rect 28474 6784 28495 6824
rect 28577 6784 28598 6824
rect 28598 6784 28638 6824
rect 28638 6784 28663 6824
rect 28409 6761 28495 6784
rect 28577 6761 28663 6784
rect 32409 6824 32495 6847
rect 32577 6824 32663 6847
rect 32409 6784 32434 6824
rect 32434 6784 32474 6824
rect 32474 6784 32495 6824
rect 32577 6784 32598 6824
rect 32598 6784 32638 6824
rect 32638 6784 32663 6824
rect 32409 6761 32495 6784
rect 32577 6761 32663 6784
rect 36409 6824 36495 6847
rect 36577 6824 36663 6847
rect 36409 6784 36434 6824
rect 36434 6784 36474 6824
rect 36474 6784 36495 6824
rect 36577 6784 36598 6824
rect 36598 6784 36638 6824
rect 36638 6784 36663 6824
rect 36409 6761 36495 6784
rect 36577 6761 36663 6784
rect 40409 6824 40495 6847
rect 40577 6824 40663 6847
rect 40409 6784 40434 6824
rect 40434 6784 40474 6824
rect 40474 6784 40495 6824
rect 40577 6784 40598 6824
rect 40598 6784 40638 6824
rect 40638 6784 40663 6824
rect 40409 6761 40495 6784
rect 40577 6761 40663 6784
rect 44409 6824 44495 6847
rect 44577 6824 44663 6847
rect 44409 6784 44434 6824
rect 44434 6784 44474 6824
rect 44474 6784 44495 6824
rect 44577 6784 44598 6824
rect 44598 6784 44638 6824
rect 44638 6784 44663 6824
rect 44409 6761 44495 6784
rect 44577 6761 44663 6784
rect 48409 6824 48495 6847
rect 48577 6824 48663 6847
rect 48409 6784 48434 6824
rect 48434 6784 48474 6824
rect 48474 6784 48495 6824
rect 48577 6784 48598 6824
rect 48598 6784 48638 6824
rect 48638 6784 48663 6824
rect 48409 6761 48495 6784
rect 48577 6761 48663 6784
rect 52409 6824 52495 6847
rect 52577 6824 52663 6847
rect 52409 6784 52434 6824
rect 52434 6784 52474 6824
rect 52474 6784 52495 6824
rect 52577 6784 52598 6824
rect 52598 6784 52638 6824
rect 52638 6784 52663 6824
rect 52409 6761 52495 6784
rect 52577 6761 52663 6784
rect 56409 6824 56495 6847
rect 56577 6824 56663 6847
rect 56409 6784 56434 6824
rect 56434 6784 56474 6824
rect 56474 6784 56495 6824
rect 56577 6784 56598 6824
rect 56598 6784 56638 6824
rect 56638 6784 56663 6824
rect 56409 6761 56495 6784
rect 56577 6761 56663 6784
rect 60409 6824 60495 6847
rect 60577 6824 60663 6847
rect 60409 6784 60434 6824
rect 60434 6784 60474 6824
rect 60474 6784 60495 6824
rect 60577 6784 60598 6824
rect 60598 6784 60638 6824
rect 60638 6784 60663 6824
rect 60409 6761 60495 6784
rect 60577 6761 60663 6784
rect 64409 6824 64495 6847
rect 64577 6824 64663 6847
rect 64409 6784 64434 6824
rect 64434 6784 64474 6824
rect 64474 6784 64495 6824
rect 64577 6784 64598 6824
rect 64598 6784 64638 6824
rect 64638 6784 64663 6824
rect 64409 6761 64495 6784
rect 64577 6761 64663 6784
rect 68409 6824 68495 6847
rect 68577 6824 68663 6847
rect 68409 6784 68434 6824
rect 68434 6784 68474 6824
rect 68474 6784 68495 6824
rect 68577 6784 68598 6824
rect 68598 6784 68638 6824
rect 68638 6784 68663 6824
rect 68409 6761 68495 6784
rect 68577 6761 68663 6784
rect 72409 6824 72495 6847
rect 72577 6824 72663 6847
rect 72409 6784 72434 6824
rect 72434 6784 72474 6824
rect 72474 6784 72495 6824
rect 72577 6784 72598 6824
rect 72598 6784 72638 6824
rect 72638 6784 72663 6824
rect 72409 6761 72495 6784
rect 72577 6761 72663 6784
rect 76409 6824 76495 6847
rect 76577 6824 76663 6847
rect 76409 6784 76434 6824
rect 76434 6784 76474 6824
rect 76474 6784 76495 6824
rect 76577 6784 76598 6824
rect 76598 6784 76638 6824
rect 76638 6784 76663 6824
rect 76409 6761 76495 6784
rect 76577 6761 76663 6784
rect 80409 6824 80495 6847
rect 80577 6824 80663 6847
rect 80409 6784 80434 6824
rect 80434 6784 80474 6824
rect 80474 6784 80495 6824
rect 80577 6784 80598 6824
rect 80598 6784 80638 6824
rect 80638 6784 80663 6824
rect 80409 6761 80495 6784
rect 80577 6761 80663 6784
rect 84409 6824 84495 6847
rect 84577 6824 84663 6847
rect 84409 6784 84434 6824
rect 84434 6784 84474 6824
rect 84474 6784 84495 6824
rect 84577 6784 84598 6824
rect 84598 6784 84638 6824
rect 84638 6784 84663 6824
rect 84409 6761 84495 6784
rect 84577 6761 84663 6784
rect 88409 6824 88495 6847
rect 88577 6824 88663 6847
rect 88409 6784 88434 6824
rect 88434 6784 88474 6824
rect 88474 6784 88495 6824
rect 88577 6784 88598 6824
rect 88598 6784 88638 6824
rect 88638 6784 88663 6824
rect 88409 6761 88495 6784
rect 88577 6761 88663 6784
rect 92409 6824 92495 6847
rect 92577 6824 92663 6847
rect 92409 6784 92434 6824
rect 92434 6784 92474 6824
rect 92474 6784 92495 6824
rect 92577 6784 92598 6824
rect 92598 6784 92638 6824
rect 92638 6784 92663 6824
rect 92409 6761 92495 6784
rect 92577 6761 92663 6784
rect 96409 6824 96495 6847
rect 96577 6824 96663 6847
rect 96409 6784 96434 6824
rect 96434 6784 96474 6824
rect 96474 6784 96495 6824
rect 96577 6784 96598 6824
rect 96598 6784 96638 6824
rect 96638 6784 96663 6824
rect 96409 6761 96495 6784
rect 96577 6761 96663 6784
rect 3169 6068 3255 6091
rect 3337 6068 3423 6091
rect 3169 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3255 6068
rect 3337 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3423 6068
rect 3169 6005 3255 6028
rect 3337 6005 3423 6028
rect 7169 6068 7255 6091
rect 7337 6068 7423 6091
rect 7169 6028 7194 6068
rect 7194 6028 7234 6068
rect 7234 6028 7255 6068
rect 7337 6028 7358 6068
rect 7358 6028 7398 6068
rect 7398 6028 7423 6068
rect 7169 6005 7255 6028
rect 7337 6005 7423 6028
rect 11169 6068 11255 6091
rect 11337 6068 11423 6091
rect 11169 6028 11194 6068
rect 11194 6028 11234 6068
rect 11234 6028 11255 6068
rect 11337 6028 11358 6068
rect 11358 6028 11398 6068
rect 11398 6028 11423 6068
rect 11169 6005 11255 6028
rect 11337 6005 11423 6028
rect 15169 6068 15255 6091
rect 15337 6068 15423 6091
rect 15169 6028 15194 6068
rect 15194 6028 15234 6068
rect 15234 6028 15255 6068
rect 15337 6028 15358 6068
rect 15358 6028 15398 6068
rect 15398 6028 15423 6068
rect 15169 6005 15255 6028
rect 15337 6005 15423 6028
rect 19169 6068 19255 6091
rect 19337 6068 19423 6091
rect 19169 6028 19194 6068
rect 19194 6028 19234 6068
rect 19234 6028 19255 6068
rect 19337 6028 19358 6068
rect 19358 6028 19398 6068
rect 19398 6028 19423 6068
rect 19169 6005 19255 6028
rect 19337 6005 19423 6028
rect 23169 6068 23255 6091
rect 23337 6068 23423 6091
rect 23169 6028 23194 6068
rect 23194 6028 23234 6068
rect 23234 6028 23255 6068
rect 23337 6028 23358 6068
rect 23358 6028 23398 6068
rect 23398 6028 23423 6068
rect 23169 6005 23255 6028
rect 23337 6005 23423 6028
rect 27169 6068 27255 6091
rect 27337 6068 27423 6091
rect 27169 6028 27194 6068
rect 27194 6028 27234 6068
rect 27234 6028 27255 6068
rect 27337 6028 27358 6068
rect 27358 6028 27398 6068
rect 27398 6028 27423 6068
rect 27169 6005 27255 6028
rect 27337 6005 27423 6028
rect 31169 6068 31255 6091
rect 31337 6068 31423 6091
rect 31169 6028 31194 6068
rect 31194 6028 31234 6068
rect 31234 6028 31255 6068
rect 31337 6028 31358 6068
rect 31358 6028 31398 6068
rect 31398 6028 31423 6068
rect 31169 6005 31255 6028
rect 31337 6005 31423 6028
rect 35169 6068 35255 6091
rect 35337 6068 35423 6091
rect 35169 6028 35194 6068
rect 35194 6028 35234 6068
rect 35234 6028 35255 6068
rect 35337 6028 35358 6068
rect 35358 6028 35398 6068
rect 35398 6028 35423 6068
rect 35169 6005 35255 6028
rect 35337 6005 35423 6028
rect 39169 6068 39255 6091
rect 39337 6068 39423 6091
rect 39169 6028 39194 6068
rect 39194 6028 39234 6068
rect 39234 6028 39255 6068
rect 39337 6028 39358 6068
rect 39358 6028 39398 6068
rect 39398 6028 39423 6068
rect 39169 6005 39255 6028
rect 39337 6005 39423 6028
rect 43169 6068 43255 6091
rect 43337 6068 43423 6091
rect 43169 6028 43194 6068
rect 43194 6028 43234 6068
rect 43234 6028 43255 6068
rect 43337 6028 43358 6068
rect 43358 6028 43398 6068
rect 43398 6028 43423 6068
rect 43169 6005 43255 6028
rect 43337 6005 43423 6028
rect 47169 6068 47255 6091
rect 47337 6068 47423 6091
rect 47169 6028 47194 6068
rect 47194 6028 47234 6068
rect 47234 6028 47255 6068
rect 47337 6028 47358 6068
rect 47358 6028 47398 6068
rect 47398 6028 47423 6068
rect 47169 6005 47255 6028
rect 47337 6005 47423 6028
rect 51169 6068 51255 6091
rect 51337 6068 51423 6091
rect 51169 6028 51194 6068
rect 51194 6028 51234 6068
rect 51234 6028 51255 6068
rect 51337 6028 51358 6068
rect 51358 6028 51398 6068
rect 51398 6028 51423 6068
rect 51169 6005 51255 6028
rect 51337 6005 51423 6028
rect 55169 6068 55255 6091
rect 55337 6068 55423 6091
rect 55169 6028 55194 6068
rect 55194 6028 55234 6068
rect 55234 6028 55255 6068
rect 55337 6028 55358 6068
rect 55358 6028 55398 6068
rect 55398 6028 55423 6068
rect 55169 6005 55255 6028
rect 55337 6005 55423 6028
rect 59169 6068 59255 6091
rect 59337 6068 59423 6091
rect 59169 6028 59194 6068
rect 59194 6028 59234 6068
rect 59234 6028 59255 6068
rect 59337 6028 59358 6068
rect 59358 6028 59398 6068
rect 59398 6028 59423 6068
rect 59169 6005 59255 6028
rect 59337 6005 59423 6028
rect 63169 6068 63255 6091
rect 63337 6068 63423 6091
rect 63169 6028 63194 6068
rect 63194 6028 63234 6068
rect 63234 6028 63255 6068
rect 63337 6028 63358 6068
rect 63358 6028 63398 6068
rect 63398 6028 63423 6068
rect 63169 6005 63255 6028
rect 63337 6005 63423 6028
rect 67169 6068 67255 6091
rect 67337 6068 67423 6091
rect 67169 6028 67194 6068
rect 67194 6028 67234 6068
rect 67234 6028 67255 6068
rect 67337 6028 67358 6068
rect 67358 6028 67398 6068
rect 67398 6028 67423 6068
rect 67169 6005 67255 6028
rect 67337 6005 67423 6028
rect 71169 6068 71255 6091
rect 71337 6068 71423 6091
rect 71169 6028 71194 6068
rect 71194 6028 71234 6068
rect 71234 6028 71255 6068
rect 71337 6028 71358 6068
rect 71358 6028 71398 6068
rect 71398 6028 71423 6068
rect 71169 6005 71255 6028
rect 71337 6005 71423 6028
rect 75169 6068 75255 6091
rect 75337 6068 75423 6091
rect 75169 6028 75194 6068
rect 75194 6028 75234 6068
rect 75234 6028 75255 6068
rect 75337 6028 75358 6068
rect 75358 6028 75398 6068
rect 75398 6028 75423 6068
rect 75169 6005 75255 6028
rect 75337 6005 75423 6028
rect 79169 6068 79255 6091
rect 79337 6068 79423 6091
rect 79169 6028 79194 6068
rect 79194 6028 79234 6068
rect 79234 6028 79255 6068
rect 79337 6028 79358 6068
rect 79358 6028 79398 6068
rect 79398 6028 79423 6068
rect 79169 6005 79255 6028
rect 79337 6005 79423 6028
rect 83169 6068 83255 6091
rect 83337 6068 83423 6091
rect 83169 6028 83194 6068
rect 83194 6028 83234 6068
rect 83234 6028 83255 6068
rect 83337 6028 83358 6068
rect 83358 6028 83398 6068
rect 83398 6028 83423 6068
rect 83169 6005 83255 6028
rect 83337 6005 83423 6028
rect 87169 6068 87255 6091
rect 87337 6068 87423 6091
rect 87169 6028 87194 6068
rect 87194 6028 87234 6068
rect 87234 6028 87255 6068
rect 87337 6028 87358 6068
rect 87358 6028 87398 6068
rect 87398 6028 87423 6068
rect 87169 6005 87255 6028
rect 87337 6005 87423 6028
rect 91169 6068 91255 6091
rect 91337 6068 91423 6091
rect 91169 6028 91194 6068
rect 91194 6028 91234 6068
rect 91234 6028 91255 6068
rect 91337 6028 91358 6068
rect 91358 6028 91398 6068
rect 91398 6028 91423 6068
rect 91169 6005 91255 6028
rect 91337 6005 91423 6028
rect 95169 6068 95255 6091
rect 95337 6068 95423 6091
rect 95169 6028 95194 6068
rect 95194 6028 95234 6068
rect 95234 6028 95255 6068
rect 95337 6028 95358 6068
rect 95358 6028 95398 6068
rect 95398 6028 95423 6068
rect 95169 6005 95255 6028
rect 95337 6005 95423 6028
rect 99169 6068 99255 6091
rect 99337 6068 99423 6091
rect 99169 6028 99194 6068
rect 99194 6028 99234 6068
rect 99234 6028 99255 6068
rect 99337 6028 99358 6068
rect 99358 6028 99398 6068
rect 99398 6028 99423 6068
rect 99169 6005 99255 6028
rect 99337 6005 99423 6028
rect 4409 5312 4495 5335
rect 4577 5312 4663 5335
rect 4409 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4495 5312
rect 4577 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4663 5312
rect 4409 5249 4495 5272
rect 4577 5249 4663 5272
rect 8409 5312 8495 5335
rect 8577 5312 8663 5335
rect 8409 5272 8434 5312
rect 8434 5272 8474 5312
rect 8474 5272 8495 5312
rect 8577 5272 8598 5312
rect 8598 5272 8638 5312
rect 8638 5272 8663 5312
rect 8409 5249 8495 5272
rect 8577 5249 8663 5272
rect 12409 5312 12495 5335
rect 12577 5312 12663 5335
rect 12409 5272 12434 5312
rect 12434 5272 12474 5312
rect 12474 5272 12495 5312
rect 12577 5272 12598 5312
rect 12598 5272 12638 5312
rect 12638 5272 12663 5312
rect 12409 5249 12495 5272
rect 12577 5249 12663 5272
rect 16409 5312 16495 5335
rect 16577 5312 16663 5335
rect 16409 5272 16434 5312
rect 16434 5272 16474 5312
rect 16474 5272 16495 5312
rect 16577 5272 16598 5312
rect 16598 5272 16638 5312
rect 16638 5272 16663 5312
rect 16409 5249 16495 5272
rect 16577 5249 16663 5272
rect 20409 5312 20495 5335
rect 20577 5312 20663 5335
rect 20409 5272 20434 5312
rect 20434 5272 20474 5312
rect 20474 5272 20495 5312
rect 20577 5272 20598 5312
rect 20598 5272 20638 5312
rect 20638 5272 20663 5312
rect 20409 5249 20495 5272
rect 20577 5249 20663 5272
rect 24409 5312 24495 5335
rect 24577 5312 24663 5335
rect 24409 5272 24434 5312
rect 24434 5272 24474 5312
rect 24474 5272 24495 5312
rect 24577 5272 24598 5312
rect 24598 5272 24638 5312
rect 24638 5272 24663 5312
rect 24409 5249 24495 5272
rect 24577 5249 24663 5272
rect 28409 5312 28495 5335
rect 28577 5312 28663 5335
rect 28409 5272 28434 5312
rect 28434 5272 28474 5312
rect 28474 5272 28495 5312
rect 28577 5272 28598 5312
rect 28598 5272 28638 5312
rect 28638 5272 28663 5312
rect 28409 5249 28495 5272
rect 28577 5249 28663 5272
rect 32409 5312 32495 5335
rect 32577 5312 32663 5335
rect 32409 5272 32434 5312
rect 32434 5272 32474 5312
rect 32474 5272 32495 5312
rect 32577 5272 32598 5312
rect 32598 5272 32638 5312
rect 32638 5272 32663 5312
rect 32409 5249 32495 5272
rect 32577 5249 32663 5272
rect 36409 5312 36495 5335
rect 36577 5312 36663 5335
rect 36409 5272 36434 5312
rect 36434 5272 36474 5312
rect 36474 5272 36495 5312
rect 36577 5272 36598 5312
rect 36598 5272 36638 5312
rect 36638 5272 36663 5312
rect 36409 5249 36495 5272
rect 36577 5249 36663 5272
rect 40409 5312 40495 5335
rect 40577 5312 40663 5335
rect 40409 5272 40434 5312
rect 40434 5272 40474 5312
rect 40474 5272 40495 5312
rect 40577 5272 40598 5312
rect 40598 5272 40638 5312
rect 40638 5272 40663 5312
rect 40409 5249 40495 5272
rect 40577 5249 40663 5272
rect 44409 5312 44495 5335
rect 44577 5312 44663 5335
rect 44409 5272 44434 5312
rect 44434 5272 44474 5312
rect 44474 5272 44495 5312
rect 44577 5272 44598 5312
rect 44598 5272 44638 5312
rect 44638 5272 44663 5312
rect 44409 5249 44495 5272
rect 44577 5249 44663 5272
rect 48409 5312 48495 5335
rect 48577 5312 48663 5335
rect 48409 5272 48434 5312
rect 48434 5272 48474 5312
rect 48474 5272 48495 5312
rect 48577 5272 48598 5312
rect 48598 5272 48638 5312
rect 48638 5272 48663 5312
rect 48409 5249 48495 5272
rect 48577 5249 48663 5272
rect 52409 5312 52495 5335
rect 52577 5312 52663 5335
rect 52409 5272 52434 5312
rect 52434 5272 52474 5312
rect 52474 5272 52495 5312
rect 52577 5272 52598 5312
rect 52598 5272 52638 5312
rect 52638 5272 52663 5312
rect 52409 5249 52495 5272
rect 52577 5249 52663 5272
rect 56409 5312 56495 5335
rect 56577 5312 56663 5335
rect 56409 5272 56434 5312
rect 56434 5272 56474 5312
rect 56474 5272 56495 5312
rect 56577 5272 56598 5312
rect 56598 5272 56638 5312
rect 56638 5272 56663 5312
rect 56409 5249 56495 5272
rect 56577 5249 56663 5272
rect 60409 5312 60495 5335
rect 60577 5312 60663 5335
rect 60409 5272 60434 5312
rect 60434 5272 60474 5312
rect 60474 5272 60495 5312
rect 60577 5272 60598 5312
rect 60598 5272 60638 5312
rect 60638 5272 60663 5312
rect 60409 5249 60495 5272
rect 60577 5249 60663 5272
rect 64409 5312 64495 5335
rect 64577 5312 64663 5335
rect 64409 5272 64434 5312
rect 64434 5272 64474 5312
rect 64474 5272 64495 5312
rect 64577 5272 64598 5312
rect 64598 5272 64638 5312
rect 64638 5272 64663 5312
rect 64409 5249 64495 5272
rect 64577 5249 64663 5272
rect 68409 5312 68495 5335
rect 68577 5312 68663 5335
rect 68409 5272 68434 5312
rect 68434 5272 68474 5312
rect 68474 5272 68495 5312
rect 68577 5272 68598 5312
rect 68598 5272 68638 5312
rect 68638 5272 68663 5312
rect 68409 5249 68495 5272
rect 68577 5249 68663 5272
rect 72409 5312 72495 5335
rect 72577 5312 72663 5335
rect 72409 5272 72434 5312
rect 72434 5272 72474 5312
rect 72474 5272 72495 5312
rect 72577 5272 72598 5312
rect 72598 5272 72638 5312
rect 72638 5272 72663 5312
rect 72409 5249 72495 5272
rect 72577 5249 72663 5272
rect 76409 5312 76495 5335
rect 76577 5312 76663 5335
rect 76409 5272 76434 5312
rect 76434 5272 76474 5312
rect 76474 5272 76495 5312
rect 76577 5272 76598 5312
rect 76598 5272 76638 5312
rect 76638 5272 76663 5312
rect 76409 5249 76495 5272
rect 76577 5249 76663 5272
rect 80409 5312 80495 5335
rect 80577 5312 80663 5335
rect 80409 5272 80434 5312
rect 80434 5272 80474 5312
rect 80474 5272 80495 5312
rect 80577 5272 80598 5312
rect 80598 5272 80638 5312
rect 80638 5272 80663 5312
rect 80409 5249 80495 5272
rect 80577 5249 80663 5272
rect 84409 5312 84495 5335
rect 84577 5312 84663 5335
rect 84409 5272 84434 5312
rect 84434 5272 84474 5312
rect 84474 5272 84495 5312
rect 84577 5272 84598 5312
rect 84598 5272 84638 5312
rect 84638 5272 84663 5312
rect 84409 5249 84495 5272
rect 84577 5249 84663 5272
rect 88409 5312 88495 5335
rect 88577 5312 88663 5335
rect 88409 5272 88434 5312
rect 88434 5272 88474 5312
rect 88474 5272 88495 5312
rect 88577 5272 88598 5312
rect 88598 5272 88638 5312
rect 88638 5272 88663 5312
rect 88409 5249 88495 5272
rect 88577 5249 88663 5272
rect 92409 5312 92495 5335
rect 92577 5312 92663 5335
rect 92409 5272 92434 5312
rect 92434 5272 92474 5312
rect 92474 5272 92495 5312
rect 92577 5272 92598 5312
rect 92598 5272 92638 5312
rect 92638 5272 92663 5312
rect 92409 5249 92495 5272
rect 92577 5249 92663 5272
rect 96409 5312 96495 5335
rect 96577 5312 96663 5335
rect 96409 5272 96434 5312
rect 96434 5272 96474 5312
rect 96474 5272 96495 5312
rect 96577 5272 96598 5312
rect 96598 5272 96638 5312
rect 96638 5272 96663 5312
rect 96409 5249 96495 5272
rect 96577 5249 96663 5272
rect 3169 4556 3255 4579
rect 3337 4556 3423 4579
rect 3169 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3255 4556
rect 3337 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3423 4556
rect 3169 4493 3255 4516
rect 3337 4493 3423 4516
rect 7169 4556 7255 4579
rect 7337 4556 7423 4579
rect 7169 4516 7194 4556
rect 7194 4516 7234 4556
rect 7234 4516 7255 4556
rect 7337 4516 7358 4556
rect 7358 4516 7398 4556
rect 7398 4516 7423 4556
rect 7169 4493 7255 4516
rect 7337 4493 7423 4516
rect 11169 4556 11255 4579
rect 11337 4556 11423 4579
rect 11169 4516 11194 4556
rect 11194 4516 11234 4556
rect 11234 4516 11255 4556
rect 11337 4516 11358 4556
rect 11358 4516 11398 4556
rect 11398 4516 11423 4556
rect 11169 4493 11255 4516
rect 11337 4493 11423 4516
rect 15169 4556 15255 4579
rect 15337 4556 15423 4579
rect 15169 4516 15194 4556
rect 15194 4516 15234 4556
rect 15234 4516 15255 4556
rect 15337 4516 15358 4556
rect 15358 4516 15398 4556
rect 15398 4516 15423 4556
rect 15169 4493 15255 4516
rect 15337 4493 15423 4516
rect 19169 4556 19255 4579
rect 19337 4556 19423 4579
rect 19169 4516 19194 4556
rect 19194 4516 19234 4556
rect 19234 4516 19255 4556
rect 19337 4516 19358 4556
rect 19358 4516 19398 4556
rect 19398 4516 19423 4556
rect 19169 4493 19255 4516
rect 19337 4493 19423 4516
rect 23169 4556 23255 4579
rect 23337 4556 23423 4579
rect 23169 4516 23194 4556
rect 23194 4516 23234 4556
rect 23234 4516 23255 4556
rect 23337 4516 23358 4556
rect 23358 4516 23398 4556
rect 23398 4516 23423 4556
rect 23169 4493 23255 4516
rect 23337 4493 23423 4516
rect 27169 4556 27255 4579
rect 27337 4556 27423 4579
rect 27169 4516 27194 4556
rect 27194 4516 27234 4556
rect 27234 4516 27255 4556
rect 27337 4516 27358 4556
rect 27358 4516 27398 4556
rect 27398 4516 27423 4556
rect 27169 4493 27255 4516
rect 27337 4493 27423 4516
rect 31169 4556 31255 4579
rect 31337 4556 31423 4579
rect 31169 4516 31194 4556
rect 31194 4516 31234 4556
rect 31234 4516 31255 4556
rect 31337 4516 31358 4556
rect 31358 4516 31398 4556
rect 31398 4516 31423 4556
rect 31169 4493 31255 4516
rect 31337 4493 31423 4516
rect 35169 4556 35255 4579
rect 35337 4556 35423 4579
rect 35169 4516 35194 4556
rect 35194 4516 35234 4556
rect 35234 4516 35255 4556
rect 35337 4516 35358 4556
rect 35358 4516 35398 4556
rect 35398 4516 35423 4556
rect 35169 4493 35255 4516
rect 35337 4493 35423 4516
rect 39169 4556 39255 4579
rect 39337 4556 39423 4579
rect 39169 4516 39194 4556
rect 39194 4516 39234 4556
rect 39234 4516 39255 4556
rect 39337 4516 39358 4556
rect 39358 4516 39398 4556
rect 39398 4516 39423 4556
rect 39169 4493 39255 4516
rect 39337 4493 39423 4516
rect 43169 4556 43255 4579
rect 43337 4556 43423 4579
rect 43169 4516 43194 4556
rect 43194 4516 43234 4556
rect 43234 4516 43255 4556
rect 43337 4516 43358 4556
rect 43358 4516 43398 4556
rect 43398 4516 43423 4556
rect 43169 4493 43255 4516
rect 43337 4493 43423 4516
rect 47169 4556 47255 4579
rect 47337 4556 47423 4579
rect 47169 4516 47194 4556
rect 47194 4516 47234 4556
rect 47234 4516 47255 4556
rect 47337 4516 47358 4556
rect 47358 4516 47398 4556
rect 47398 4516 47423 4556
rect 47169 4493 47255 4516
rect 47337 4493 47423 4516
rect 51169 4556 51255 4579
rect 51337 4556 51423 4579
rect 51169 4516 51194 4556
rect 51194 4516 51234 4556
rect 51234 4516 51255 4556
rect 51337 4516 51358 4556
rect 51358 4516 51398 4556
rect 51398 4516 51423 4556
rect 51169 4493 51255 4516
rect 51337 4493 51423 4516
rect 55169 4556 55255 4579
rect 55337 4556 55423 4579
rect 55169 4516 55194 4556
rect 55194 4516 55234 4556
rect 55234 4516 55255 4556
rect 55337 4516 55358 4556
rect 55358 4516 55398 4556
rect 55398 4516 55423 4556
rect 55169 4493 55255 4516
rect 55337 4493 55423 4516
rect 59169 4556 59255 4579
rect 59337 4556 59423 4579
rect 59169 4516 59194 4556
rect 59194 4516 59234 4556
rect 59234 4516 59255 4556
rect 59337 4516 59358 4556
rect 59358 4516 59398 4556
rect 59398 4516 59423 4556
rect 59169 4493 59255 4516
rect 59337 4493 59423 4516
rect 63169 4556 63255 4579
rect 63337 4556 63423 4579
rect 63169 4516 63194 4556
rect 63194 4516 63234 4556
rect 63234 4516 63255 4556
rect 63337 4516 63358 4556
rect 63358 4516 63398 4556
rect 63398 4516 63423 4556
rect 63169 4493 63255 4516
rect 63337 4493 63423 4516
rect 67169 4556 67255 4579
rect 67337 4556 67423 4579
rect 67169 4516 67194 4556
rect 67194 4516 67234 4556
rect 67234 4516 67255 4556
rect 67337 4516 67358 4556
rect 67358 4516 67398 4556
rect 67398 4516 67423 4556
rect 67169 4493 67255 4516
rect 67337 4493 67423 4516
rect 71169 4556 71255 4579
rect 71337 4556 71423 4579
rect 71169 4516 71194 4556
rect 71194 4516 71234 4556
rect 71234 4516 71255 4556
rect 71337 4516 71358 4556
rect 71358 4516 71398 4556
rect 71398 4516 71423 4556
rect 71169 4493 71255 4516
rect 71337 4493 71423 4516
rect 75169 4556 75255 4579
rect 75337 4556 75423 4579
rect 75169 4516 75194 4556
rect 75194 4516 75234 4556
rect 75234 4516 75255 4556
rect 75337 4516 75358 4556
rect 75358 4516 75398 4556
rect 75398 4516 75423 4556
rect 75169 4493 75255 4516
rect 75337 4493 75423 4516
rect 79169 4556 79255 4579
rect 79337 4556 79423 4579
rect 79169 4516 79194 4556
rect 79194 4516 79234 4556
rect 79234 4516 79255 4556
rect 79337 4516 79358 4556
rect 79358 4516 79398 4556
rect 79398 4516 79423 4556
rect 79169 4493 79255 4516
rect 79337 4493 79423 4516
rect 83169 4556 83255 4579
rect 83337 4556 83423 4579
rect 83169 4516 83194 4556
rect 83194 4516 83234 4556
rect 83234 4516 83255 4556
rect 83337 4516 83358 4556
rect 83358 4516 83398 4556
rect 83398 4516 83423 4556
rect 83169 4493 83255 4516
rect 83337 4493 83423 4516
rect 87169 4556 87255 4579
rect 87337 4556 87423 4579
rect 87169 4516 87194 4556
rect 87194 4516 87234 4556
rect 87234 4516 87255 4556
rect 87337 4516 87358 4556
rect 87358 4516 87398 4556
rect 87398 4516 87423 4556
rect 87169 4493 87255 4516
rect 87337 4493 87423 4516
rect 91169 4556 91255 4579
rect 91337 4556 91423 4579
rect 91169 4516 91194 4556
rect 91194 4516 91234 4556
rect 91234 4516 91255 4556
rect 91337 4516 91358 4556
rect 91358 4516 91398 4556
rect 91398 4516 91423 4556
rect 91169 4493 91255 4516
rect 91337 4493 91423 4516
rect 95169 4556 95255 4579
rect 95337 4556 95423 4579
rect 95169 4516 95194 4556
rect 95194 4516 95234 4556
rect 95234 4516 95255 4556
rect 95337 4516 95358 4556
rect 95358 4516 95398 4556
rect 95398 4516 95423 4556
rect 95169 4493 95255 4516
rect 95337 4493 95423 4516
rect 99169 4556 99255 4579
rect 99337 4556 99423 4579
rect 99169 4516 99194 4556
rect 99194 4516 99234 4556
rect 99234 4516 99255 4556
rect 99337 4516 99358 4556
rect 99358 4516 99398 4556
rect 99398 4516 99423 4556
rect 99169 4493 99255 4516
rect 99337 4493 99423 4516
rect 4409 3800 4495 3823
rect 4577 3800 4663 3823
rect 4409 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4495 3800
rect 4577 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4663 3800
rect 4409 3737 4495 3760
rect 4577 3737 4663 3760
rect 8409 3800 8495 3823
rect 8577 3800 8663 3823
rect 8409 3760 8434 3800
rect 8434 3760 8474 3800
rect 8474 3760 8495 3800
rect 8577 3760 8598 3800
rect 8598 3760 8638 3800
rect 8638 3760 8663 3800
rect 8409 3737 8495 3760
rect 8577 3737 8663 3760
rect 12409 3800 12495 3823
rect 12577 3800 12663 3823
rect 12409 3760 12434 3800
rect 12434 3760 12474 3800
rect 12474 3760 12495 3800
rect 12577 3760 12598 3800
rect 12598 3760 12638 3800
rect 12638 3760 12663 3800
rect 12409 3737 12495 3760
rect 12577 3737 12663 3760
rect 16409 3800 16495 3823
rect 16577 3800 16663 3823
rect 16409 3760 16434 3800
rect 16434 3760 16474 3800
rect 16474 3760 16495 3800
rect 16577 3760 16598 3800
rect 16598 3760 16638 3800
rect 16638 3760 16663 3800
rect 16409 3737 16495 3760
rect 16577 3737 16663 3760
rect 20409 3800 20495 3823
rect 20577 3800 20663 3823
rect 20409 3760 20434 3800
rect 20434 3760 20474 3800
rect 20474 3760 20495 3800
rect 20577 3760 20598 3800
rect 20598 3760 20638 3800
rect 20638 3760 20663 3800
rect 20409 3737 20495 3760
rect 20577 3737 20663 3760
rect 24409 3800 24495 3823
rect 24577 3800 24663 3823
rect 24409 3760 24434 3800
rect 24434 3760 24474 3800
rect 24474 3760 24495 3800
rect 24577 3760 24598 3800
rect 24598 3760 24638 3800
rect 24638 3760 24663 3800
rect 24409 3737 24495 3760
rect 24577 3737 24663 3760
rect 28409 3800 28495 3823
rect 28577 3800 28663 3823
rect 28409 3760 28434 3800
rect 28434 3760 28474 3800
rect 28474 3760 28495 3800
rect 28577 3760 28598 3800
rect 28598 3760 28638 3800
rect 28638 3760 28663 3800
rect 28409 3737 28495 3760
rect 28577 3737 28663 3760
rect 32409 3800 32495 3823
rect 32577 3800 32663 3823
rect 32409 3760 32434 3800
rect 32434 3760 32474 3800
rect 32474 3760 32495 3800
rect 32577 3760 32598 3800
rect 32598 3760 32638 3800
rect 32638 3760 32663 3800
rect 32409 3737 32495 3760
rect 32577 3737 32663 3760
rect 36409 3800 36495 3823
rect 36577 3800 36663 3823
rect 36409 3760 36434 3800
rect 36434 3760 36474 3800
rect 36474 3760 36495 3800
rect 36577 3760 36598 3800
rect 36598 3760 36638 3800
rect 36638 3760 36663 3800
rect 36409 3737 36495 3760
rect 36577 3737 36663 3760
rect 40409 3800 40495 3823
rect 40577 3800 40663 3823
rect 40409 3760 40434 3800
rect 40434 3760 40474 3800
rect 40474 3760 40495 3800
rect 40577 3760 40598 3800
rect 40598 3760 40638 3800
rect 40638 3760 40663 3800
rect 40409 3737 40495 3760
rect 40577 3737 40663 3760
rect 44409 3800 44495 3823
rect 44577 3800 44663 3823
rect 44409 3760 44434 3800
rect 44434 3760 44474 3800
rect 44474 3760 44495 3800
rect 44577 3760 44598 3800
rect 44598 3760 44638 3800
rect 44638 3760 44663 3800
rect 44409 3737 44495 3760
rect 44577 3737 44663 3760
rect 48409 3800 48495 3823
rect 48577 3800 48663 3823
rect 48409 3760 48434 3800
rect 48434 3760 48474 3800
rect 48474 3760 48495 3800
rect 48577 3760 48598 3800
rect 48598 3760 48638 3800
rect 48638 3760 48663 3800
rect 48409 3737 48495 3760
rect 48577 3737 48663 3760
rect 52409 3800 52495 3823
rect 52577 3800 52663 3823
rect 52409 3760 52434 3800
rect 52434 3760 52474 3800
rect 52474 3760 52495 3800
rect 52577 3760 52598 3800
rect 52598 3760 52638 3800
rect 52638 3760 52663 3800
rect 52409 3737 52495 3760
rect 52577 3737 52663 3760
rect 56409 3800 56495 3823
rect 56577 3800 56663 3823
rect 56409 3760 56434 3800
rect 56434 3760 56474 3800
rect 56474 3760 56495 3800
rect 56577 3760 56598 3800
rect 56598 3760 56638 3800
rect 56638 3760 56663 3800
rect 56409 3737 56495 3760
rect 56577 3737 56663 3760
rect 60409 3800 60495 3823
rect 60577 3800 60663 3823
rect 60409 3760 60434 3800
rect 60434 3760 60474 3800
rect 60474 3760 60495 3800
rect 60577 3760 60598 3800
rect 60598 3760 60638 3800
rect 60638 3760 60663 3800
rect 60409 3737 60495 3760
rect 60577 3737 60663 3760
rect 64409 3800 64495 3823
rect 64577 3800 64663 3823
rect 64409 3760 64434 3800
rect 64434 3760 64474 3800
rect 64474 3760 64495 3800
rect 64577 3760 64598 3800
rect 64598 3760 64638 3800
rect 64638 3760 64663 3800
rect 64409 3737 64495 3760
rect 64577 3737 64663 3760
rect 68409 3800 68495 3823
rect 68577 3800 68663 3823
rect 68409 3760 68434 3800
rect 68434 3760 68474 3800
rect 68474 3760 68495 3800
rect 68577 3760 68598 3800
rect 68598 3760 68638 3800
rect 68638 3760 68663 3800
rect 68409 3737 68495 3760
rect 68577 3737 68663 3760
rect 72409 3800 72495 3823
rect 72577 3800 72663 3823
rect 72409 3760 72434 3800
rect 72434 3760 72474 3800
rect 72474 3760 72495 3800
rect 72577 3760 72598 3800
rect 72598 3760 72638 3800
rect 72638 3760 72663 3800
rect 72409 3737 72495 3760
rect 72577 3737 72663 3760
rect 76409 3800 76495 3823
rect 76577 3800 76663 3823
rect 76409 3760 76434 3800
rect 76434 3760 76474 3800
rect 76474 3760 76495 3800
rect 76577 3760 76598 3800
rect 76598 3760 76638 3800
rect 76638 3760 76663 3800
rect 76409 3737 76495 3760
rect 76577 3737 76663 3760
rect 80409 3800 80495 3823
rect 80577 3800 80663 3823
rect 80409 3760 80434 3800
rect 80434 3760 80474 3800
rect 80474 3760 80495 3800
rect 80577 3760 80598 3800
rect 80598 3760 80638 3800
rect 80638 3760 80663 3800
rect 80409 3737 80495 3760
rect 80577 3737 80663 3760
rect 84409 3800 84495 3823
rect 84577 3800 84663 3823
rect 84409 3760 84434 3800
rect 84434 3760 84474 3800
rect 84474 3760 84495 3800
rect 84577 3760 84598 3800
rect 84598 3760 84638 3800
rect 84638 3760 84663 3800
rect 84409 3737 84495 3760
rect 84577 3737 84663 3760
rect 88409 3800 88495 3823
rect 88577 3800 88663 3823
rect 88409 3760 88434 3800
rect 88434 3760 88474 3800
rect 88474 3760 88495 3800
rect 88577 3760 88598 3800
rect 88598 3760 88638 3800
rect 88638 3760 88663 3800
rect 88409 3737 88495 3760
rect 88577 3737 88663 3760
rect 92409 3800 92495 3823
rect 92577 3800 92663 3823
rect 92409 3760 92434 3800
rect 92434 3760 92474 3800
rect 92474 3760 92495 3800
rect 92577 3760 92598 3800
rect 92598 3760 92638 3800
rect 92638 3760 92663 3800
rect 92409 3737 92495 3760
rect 92577 3737 92663 3760
rect 96409 3800 96495 3823
rect 96577 3800 96663 3823
rect 96409 3760 96434 3800
rect 96434 3760 96474 3800
rect 96474 3760 96495 3800
rect 96577 3760 96598 3800
rect 96598 3760 96638 3800
rect 96638 3760 96663 3800
rect 96409 3737 96495 3760
rect 96577 3737 96663 3760
rect 3169 3044 3255 3067
rect 3337 3044 3423 3067
rect 3169 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3255 3044
rect 3337 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3423 3044
rect 3169 2981 3255 3004
rect 3337 2981 3423 3004
rect 7169 3044 7255 3067
rect 7337 3044 7423 3067
rect 7169 3004 7194 3044
rect 7194 3004 7234 3044
rect 7234 3004 7255 3044
rect 7337 3004 7358 3044
rect 7358 3004 7398 3044
rect 7398 3004 7423 3044
rect 7169 2981 7255 3004
rect 7337 2981 7423 3004
rect 11169 3044 11255 3067
rect 11337 3044 11423 3067
rect 11169 3004 11194 3044
rect 11194 3004 11234 3044
rect 11234 3004 11255 3044
rect 11337 3004 11358 3044
rect 11358 3004 11398 3044
rect 11398 3004 11423 3044
rect 11169 2981 11255 3004
rect 11337 2981 11423 3004
rect 15169 3044 15255 3067
rect 15337 3044 15423 3067
rect 15169 3004 15194 3044
rect 15194 3004 15234 3044
rect 15234 3004 15255 3044
rect 15337 3004 15358 3044
rect 15358 3004 15398 3044
rect 15398 3004 15423 3044
rect 15169 2981 15255 3004
rect 15337 2981 15423 3004
rect 19169 3044 19255 3067
rect 19337 3044 19423 3067
rect 19169 3004 19194 3044
rect 19194 3004 19234 3044
rect 19234 3004 19255 3044
rect 19337 3004 19358 3044
rect 19358 3004 19398 3044
rect 19398 3004 19423 3044
rect 19169 2981 19255 3004
rect 19337 2981 19423 3004
rect 23169 3044 23255 3067
rect 23337 3044 23423 3067
rect 23169 3004 23194 3044
rect 23194 3004 23234 3044
rect 23234 3004 23255 3044
rect 23337 3004 23358 3044
rect 23358 3004 23398 3044
rect 23398 3004 23423 3044
rect 23169 2981 23255 3004
rect 23337 2981 23423 3004
rect 27169 3044 27255 3067
rect 27337 3044 27423 3067
rect 27169 3004 27194 3044
rect 27194 3004 27234 3044
rect 27234 3004 27255 3044
rect 27337 3004 27358 3044
rect 27358 3004 27398 3044
rect 27398 3004 27423 3044
rect 27169 2981 27255 3004
rect 27337 2981 27423 3004
rect 31169 3044 31255 3067
rect 31337 3044 31423 3067
rect 31169 3004 31194 3044
rect 31194 3004 31234 3044
rect 31234 3004 31255 3044
rect 31337 3004 31358 3044
rect 31358 3004 31398 3044
rect 31398 3004 31423 3044
rect 31169 2981 31255 3004
rect 31337 2981 31423 3004
rect 35169 3044 35255 3067
rect 35337 3044 35423 3067
rect 35169 3004 35194 3044
rect 35194 3004 35234 3044
rect 35234 3004 35255 3044
rect 35337 3004 35358 3044
rect 35358 3004 35398 3044
rect 35398 3004 35423 3044
rect 35169 2981 35255 3004
rect 35337 2981 35423 3004
rect 39169 3044 39255 3067
rect 39337 3044 39423 3067
rect 39169 3004 39194 3044
rect 39194 3004 39234 3044
rect 39234 3004 39255 3044
rect 39337 3004 39358 3044
rect 39358 3004 39398 3044
rect 39398 3004 39423 3044
rect 39169 2981 39255 3004
rect 39337 2981 39423 3004
rect 43169 3044 43255 3067
rect 43337 3044 43423 3067
rect 43169 3004 43194 3044
rect 43194 3004 43234 3044
rect 43234 3004 43255 3044
rect 43337 3004 43358 3044
rect 43358 3004 43398 3044
rect 43398 3004 43423 3044
rect 43169 2981 43255 3004
rect 43337 2981 43423 3004
rect 47169 3044 47255 3067
rect 47337 3044 47423 3067
rect 47169 3004 47194 3044
rect 47194 3004 47234 3044
rect 47234 3004 47255 3044
rect 47337 3004 47358 3044
rect 47358 3004 47398 3044
rect 47398 3004 47423 3044
rect 47169 2981 47255 3004
rect 47337 2981 47423 3004
rect 51169 3044 51255 3067
rect 51337 3044 51423 3067
rect 51169 3004 51194 3044
rect 51194 3004 51234 3044
rect 51234 3004 51255 3044
rect 51337 3004 51358 3044
rect 51358 3004 51398 3044
rect 51398 3004 51423 3044
rect 51169 2981 51255 3004
rect 51337 2981 51423 3004
rect 55169 3044 55255 3067
rect 55337 3044 55423 3067
rect 55169 3004 55194 3044
rect 55194 3004 55234 3044
rect 55234 3004 55255 3044
rect 55337 3004 55358 3044
rect 55358 3004 55398 3044
rect 55398 3004 55423 3044
rect 55169 2981 55255 3004
rect 55337 2981 55423 3004
rect 59169 3044 59255 3067
rect 59337 3044 59423 3067
rect 59169 3004 59194 3044
rect 59194 3004 59234 3044
rect 59234 3004 59255 3044
rect 59337 3004 59358 3044
rect 59358 3004 59398 3044
rect 59398 3004 59423 3044
rect 59169 2981 59255 3004
rect 59337 2981 59423 3004
rect 63169 3044 63255 3067
rect 63337 3044 63423 3067
rect 63169 3004 63194 3044
rect 63194 3004 63234 3044
rect 63234 3004 63255 3044
rect 63337 3004 63358 3044
rect 63358 3004 63398 3044
rect 63398 3004 63423 3044
rect 63169 2981 63255 3004
rect 63337 2981 63423 3004
rect 67169 3044 67255 3067
rect 67337 3044 67423 3067
rect 67169 3004 67194 3044
rect 67194 3004 67234 3044
rect 67234 3004 67255 3044
rect 67337 3004 67358 3044
rect 67358 3004 67398 3044
rect 67398 3004 67423 3044
rect 67169 2981 67255 3004
rect 67337 2981 67423 3004
rect 71169 3044 71255 3067
rect 71337 3044 71423 3067
rect 71169 3004 71194 3044
rect 71194 3004 71234 3044
rect 71234 3004 71255 3044
rect 71337 3004 71358 3044
rect 71358 3004 71398 3044
rect 71398 3004 71423 3044
rect 71169 2981 71255 3004
rect 71337 2981 71423 3004
rect 75169 3044 75255 3067
rect 75337 3044 75423 3067
rect 75169 3004 75194 3044
rect 75194 3004 75234 3044
rect 75234 3004 75255 3044
rect 75337 3004 75358 3044
rect 75358 3004 75398 3044
rect 75398 3004 75423 3044
rect 75169 2981 75255 3004
rect 75337 2981 75423 3004
rect 79169 3044 79255 3067
rect 79337 3044 79423 3067
rect 79169 3004 79194 3044
rect 79194 3004 79234 3044
rect 79234 3004 79255 3044
rect 79337 3004 79358 3044
rect 79358 3004 79398 3044
rect 79398 3004 79423 3044
rect 79169 2981 79255 3004
rect 79337 2981 79423 3004
rect 83169 3044 83255 3067
rect 83337 3044 83423 3067
rect 83169 3004 83194 3044
rect 83194 3004 83234 3044
rect 83234 3004 83255 3044
rect 83337 3004 83358 3044
rect 83358 3004 83398 3044
rect 83398 3004 83423 3044
rect 83169 2981 83255 3004
rect 83337 2981 83423 3004
rect 87169 3044 87255 3067
rect 87337 3044 87423 3067
rect 87169 3004 87194 3044
rect 87194 3004 87234 3044
rect 87234 3004 87255 3044
rect 87337 3004 87358 3044
rect 87358 3004 87398 3044
rect 87398 3004 87423 3044
rect 87169 2981 87255 3004
rect 87337 2981 87423 3004
rect 91169 3044 91255 3067
rect 91337 3044 91423 3067
rect 91169 3004 91194 3044
rect 91194 3004 91234 3044
rect 91234 3004 91255 3044
rect 91337 3004 91358 3044
rect 91358 3004 91398 3044
rect 91398 3004 91423 3044
rect 91169 2981 91255 3004
rect 91337 2981 91423 3004
rect 95169 3044 95255 3067
rect 95337 3044 95423 3067
rect 95169 3004 95194 3044
rect 95194 3004 95234 3044
rect 95234 3004 95255 3044
rect 95337 3004 95358 3044
rect 95358 3004 95398 3044
rect 95398 3004 95423 3044
rect 95169 2981 95255 3004
rect 95337 2981 95423 3004
rect 99169 3044 99255 3067
rect 99337 3044 99423 3067
rect 99169 3004 99194 3044
rect 99194 3004 99234 3044
rect 99234 3004 99255 3044
rect 99337 3004 99358 3044
rect 99358 3004 99398 3044
rect 99398 3004 99423 3044
rect 99169 2981 99255 3004
rect 99337 2981 99423 3004
rect 4409 2288 4495 2311
rect 4577 2288 4663 2311
rect 4409 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4495 2288
rect 4577 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4663 2288
rect 4409 2225 4495 2248
rect 4577 2225 4663 2248
rect 8409 2288 8495 2311
rect 8577 2288 8663 2311
rect 8409 2248 8434 2288
rect 8434 2248 8474 2288
rect 8474 2248 8495 2288
rect 8577 2248 8598 2288
rect 8598 2248 8638 2288
rect 8638 2248 8663 2288
rect 8409 2225 8495 2248
rect 8577 2225 8663 2248
rect 12409 2288 12495 2311
rect 12577 2288 12663 2311
rect 12409 2248 12434 2288
rect 12434 2248 12474 2288
rect 12474 2248 12495 2288
rect 12577 2248 12598 2288
rect 12598 2248 12638 2288
rect 12638 2248 12663 2288
rect 12409 2225 12495 2248
rect 12577 2225 12663 2248
rect 16409 2288 16495 2311
rect 16577 2288 16663 2311
rect 16409 2248 16434 2288
rect 16434 2248 16474 2288
rect 16474 2248 16495 2288
rect 16577 2248 16598 2288
rect 16598 2248 16638 2288
rect 16638 2248 16663 2288
rect 16409 2225 16495 2248
rect 16577 2225 16663 2248
rect 20409 2288 20495 2311
rect 20577 2288 20663 2311
rect 20409 2248 20434 2288
rect 20434 2248 20474 2288
rect 20474 2248 20495 2288
rect 20577 2248 20598 2288
rect 20598 2248 20638 2288
rect 20638 2248 20663 2288
rect 20409 2225 20495 2248
rect 20577 2225 20663 2248
rect 24409 2288 24495 2311
rect 24577 2288 24663 2311
rect 24409 2248 24434 2288
rect 24434 2248 24474 2288
rect 24474 2248 24495 2288
rect 24577 2248 24598 2288
rect 24598 2248 24638 2288
rect 24638 2248 24663 2288
rect 24409 2225 24495 2248
rect 24577 2225 24663 2248
rect 28409 2288 28495 2311
rect 28577 2288 28663 2311
rect 28409 2248 28434 2288
rect 28434 2248 28474 2288
rect 28474 2248 28495 2288
rect 28577 2248 28598 2288
rect 28598 2248 28638 2288
rect 28638 2248 28663 2288
rect 28409 2225 28495 2248
rect 28577 2225 28663 2248
rect 32409 2288 32495 2311
rect 32577 2288 32663 2311
rect 32409 2248 32434 2288
rect 32434 2248 32474 2288
rect 32474 2248 32495 2288
rect 32577 2248 32598 2288
rect 32598 2248 32638 2288
rect 32638 2248 32663 2288
rect 32409 2225 32495 2248
rect 32577 2225 32663 2248
rect 36409 2288 36495 2311
rect 36577 2288 36663 2311
rect 36409 2248 36434 2288
rect 36434 2248 36474 2288
rect 36474 2248 36495 2288
rect 36577 2248 36598 2288
rect 36598 2248 36638 2288
rect 36638 2248 36663 2288
rect 36409 2225 36495 2248
rect 36577 2225 36663 2248
rect 40409 2288 40495 2311
rect 40577 2288 40663 2311
rect 40409 2248 40434 2288
rect 40434 2248 40474 2288
rect 40474 2248 40495 2288
rect 40577 2248 40598 2288
rect 40598 2248 40638 2288
rect 40638 2248 40663 2288
rect 40409 2225 40495 2248
rect 40577 2225 40663 2248
rect 44409 2288 44495 2311
rect 44577 2288 44663 2311
rect 44409 2248 44434 2288
rect 44434 2248 44474 2288
rect 44474 2248 44495 2288
rect 44577 2248 44598 2288
rect 44598 2248 44638 2288
rect 44638 2248 44663 2288
rect 44409 2225 44495 2248
rect 44577 2225 44663 2248
rect 48409 2288 48495 2311
rect 48577 2288 48663 2311
rect 48409 2248 48434 2288
rect 48434 2248 48474 2288
rect 48474 2248 48495 2288
rect 48577 2248 48598 2288
rect 48598 2248 48638 2288
rect 48638 2248 48663 2288
rect 48409 2225 48495 2248
rect 48577 2225 48663 2248
rect 52409 2288 52495 2311
rect 52577 2288 52663 2311
rect 52409 2248 52434 2288
rect 52434 2248 52474 2288
rect 52474 2248 52495 2288
rect 52577 2248 52598 2288
rect 52598 2248 52638 2288
rect 52638 2248 52663 2288
rect 52409 2225 52495 2248
rect 52577 2225 52663 2248
rect 56409 2288 56495 2311
rect 56577 2288 56663 2311
rect 56409 2248 56434 2288
rect 56434 2248 56474 2288
rect 56474 2248 56495 2288
rect 56577 2248 56598 2288
rect 56598 2248 56638 2288
rect 56638 2248 56663 2288
rect 56409 2225 56495 2248
rect 56577 2225 56663 2248
rect 60409 2288 60495 2311
rect 60577 2288 60663 2311
rect 60409 2248 60434 2288
rect 60434 2248 60474 2288
rect 60474 2248 60495 2288
rect 60577 2248 60598 2288
rect 60598 2248 60638 2288
rect 60638 2248 60663 2288
rect 60409 2225 60495 2248
rect 60577 2225 60663 2248
rect 64409 2288 64495 2311
rect 64577 2288 64663 2311
rect 64409 2248 64434 2288
rect 64434 2248 64474 2288
rect 64474 2248 64495 2288
rect 64577 2248 64598 2288
rect 64598 2248 64638 2288
rect 64638 2248 64663 2288
rect 64409 2225 64495 2248
rect 64577 2225 64663 2248
rect 68409 2288 68495 2311
rect 68577 2288 68663 2311
rect 68409 2248 68434 2288
rect 68434 2248 68474 2288
rect 68474 2248 68495 2288
rect 68577 2248 68598 2288
rect 68598 2248 68638 2288
rect 68638 2248 68663 2288
rect 68409 2225 68495 2248
rect 68577 2225 68663 2248
rect 72409 2288 72495 2311
rect 72577 2288 72663 2311
rect 72409 2248 72434 2288
rect 72434 2248 72474 2288
rect 72474 2248 72495 2288
rect 72577 2248 72598 2288
rect 72598 2248 72638 2288
rect 72638 2248 72663 2288
rect 72409 2225 72495 2248
rect 72577 2225 72663 2248
rect 76409 2288 76495 2311
rect 76577 2288 76663 2311
rect 76409 2248 76434 2288
rect 76434 2248 76474 2288
rect 76474 2248 76495 2288
rect 76577 2248 76598 2288
rect 76598 2248 76638 2288
rect 76638 2248 76663 2288
rect 76409 2225 76495 2248
rect 76577 2225 76663 2248
rect 80409 2288 80495 2311
rect 80577 2288 80663 2311
rect 80409 2248 80434 2288
rect 80434 2248 80474 2288
rect 80474 2248 80495 2288
rect 80577 2248 80598 2288
rect 80598 2248 80638 2288
rect 80638 2248 80663 2288
rect 80409 2225 80495 2248
rect 80577 2225 80663 2248
rect 84409 2288 84495 2311
rect 84577 2288 84663 2311
rect 84409 2248 84434 2288
rect 84434 2248 84474 2288
rect 84474 2248 84495 2288
rect 84577 2248 84598 2288
rect 84598 2248 84638 2288
rect 84638 2248 84663 2288
rect 84409 2225 84495 2248
rect 84577 2225 84663 2248
rect 88409 2288 88495 2311
rect 88577 2288 88663 2311
rect 88409 2248 88434 2288
rect 88434 2248 88474 2288
rect 88474 2248 88495 2288
rect 88577 2248 88598 2288
rect 88598 2248 88638 2288
rect 88638 2248 88663 2288
rect 88409 2225 88495 2248
rect 88577 2225 88663 2248
rect 92409 2288 92495 2311
rect 92577 2288 92663 2311
rect 92409 2248 92434 2288
rect 92434 2248 92474 2288
rect 92474 2248 92495 2288
rect 92577 2248 92598 2288
rect 92598 2248 92638 2288
rect 92638 2248 92663 2288
rect 92409 2225 92495 2248
rect 92577 2225 92663 2248
rect 96409 2288 96495 2311
rect 96577 2288 96663 2311
rect 96409 2248 96434 2288
rect 96434 2248 96474 2288
rect 96474 2248 96495 2288
rect 96577 2248 96598 2288
rect 96598 2248 96638 2288
rect 96638 2248 96663 2288
rect 96409 2225 96495 2248
rect 96577 2225 96663 2248
rect 3169 1532 3255 1555
rect 3337 1532 3423 1555
rect 3169 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3255 1532
rect 3337 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3423 1532
rect 3169 1469 3255 1492
rect 3337 1469 3423 1492
rect 7169 1532 7255 1555
rect 7337 1532 7423 1555
rect 7169 1492 7194 1532
rect 7194 1492 7234 1532
rect 7234 1492 7255 1532
rect 7337 1492 7358 1532
rect 7358 1492 7398 1532
rect 7398 1492 7423 1532
rect 7169 1469 7255 1492
rect 7337 1469 7423 1492
rect 11169 1532 11255 1555
rect 11337 1532 11423 1555
rect 11169 1492 11194 1532
rect 11194 1492 11234 1532
rect 11234 1492 11255 1532
rect 11337 1492 11358 1532
rect 11358 1492 11398 1532
rect 11398 1492 11423 1532
rect 11169 1469 11255 1492
rect 11337 1469 11423 1492
rect 15169 1532 15255 1555
rect 15337 1532 15423 1555
rect 15169 1492 15194 1532
rect 15194 1492 15234 1532
rect 15234 1492 15255 1532
rect 15337 1492 15358 1532
rect 15358 1492 15398 1532
rect 15398 1492 15423 1532
rect 15169 1469 15255 1492
rect 15337 1469 15423 1492
rect 19169 1532 19255 1555
rect 19337 1532 19423 1555
rect 19169 1492 19194 1532
rect 19194 1492 19234 1532
rect 19234 1492 19255 1532
rect 19337 1492 19358 1532
rect 19358 1492 19398 1532
rect 19398 1492 19423 1532
rect 19169 1469 19255 1492
rect 19337 1469 19423 1492
rect 23169 1532 23255 1555
rect 23337 1532 23423 1555
rect 23169 1492 23194 1532
rect 23194 1492 23234 1532
rect 23234 1492 23255 1532
rect 23337 1492 23358 1532
rect 23358 1492 23398 1532
rect 23398 1492 23423 1532
rect 23169 1469 23255 1492
rect 23337 1469 23423 1492
rect 27169 1532 27255 1555
rect 27337 1532 27423 1555
rect 27169 1492 27194 1532
rect 27194 1492 27234 1532
rect 27234 1492 27255 1532
rect 27337 1492 27358 1532
rect 27358 1492 27398 1532
rect 27398 1492 27423 1532
rect 27169 1469 27255 1492
rect 27337 1469 27423 1492
rect 31169 1532 31255 1555
rect 31337 1532 31423 1555
rect 31169 1492 31194 1532
rect 31194 1492 31234 1532
rect 31234 1492 31255 1532
rect 31337 1492 31358 1532
rect 31358 1492 31398 1532
rect 31398 1492 31423 1532
rect 31169 1469 31255 1492
rect 31337 1469 31423 1492
rect 35169 1532 35255 1555
rect 35337 1532 35423 1555
rect 35169 1492 35194 1532
rect 35194 1492 35234 1532
rect 35234 1492 35255 1532
rect 35337 1492 35358 1532
rect 35358 1492 35398 1532
rect 35398 1492 35423 1532
rect 35169 1469 35255 1492
rect 35337 1469 35423 1492
rect 39169 1532 39255 1555
rect 39337 1532 39423 1555
rect 39169 1492 39194 1532
rect 39194 1492 39234 1532
rect 39234 1492 39255 1532
rect 39337 1492 39358 1532
rect 39358 1492 39398 1532
rect 39398 1492 39423 1532
rect 39169 1469 39255 1492
rect 39337 1469 39423 1492
rect 43169 1532 43255 1555
rect 43337 1532 43423 1555
rect 43169 1492 43194 1532
rect 43194 1492 43234 1532
rect 43234 1492 43255 1532
rect 43337 1492 43358 1532
rect 43358 1492 43398 1532
rect 43398 1492 43423 1532
rect 43169 1469 43255 1492
rect 43337 1469 43423 1492
rect 47169 1532 47255 1555
rect 47337 1532 47423 1555
rect 47169 1492 47194 1532
rect 47194 1492 47234 1532
rect 47234 1492 47255 1532
rect 47337 1492 47358 1532
rect 47358 1492 47398 1532
rect 47398 1492 47423 1532
rect 47169 1469 47255 1492
rect 47337 1469 47423 1492
rect 51169 1532 51255 1555
rect 51337 1532 51423 1555
rect 51169 1492 51194 1532
rect 51194 1492 51234 1532
rect 51234 1492 51255 1532
rect 51337 1492 51358 1532
rect 51358 1492 51398 1532
rect 51398 1492 51423 1532
rect 51169 1469 51255 1492
rect 51337 1469 51423 1492
rect 55169 1532 55255 1555
rect 55337 1532 55423 1555
rect 55169 1492 55194 1532
rect 55194 1492 55234 1532
rect 55234 1492 55255 1532
rect 55337 1492 55358 1532
rect 55358 1492 55398 1532
rect 55398 1492 55423 1532
rect 55169 1469 55255 1492
rect 55337 1469 55423 1492
rect 59169 1532 59255 1555
rect 59337 1532 59423 1555
rect 59169 1492 59194 1532
rect 59194 1492 59234 1532
rect 59234 1492 59255 1532
rect 59337 1492 59358 1532
rect 59358 1492 59398 1532
rect 59398 1492 59423 1532
rect 59169 1469 59255 1492
rect 59337 1469 59423 1492
rect 63169 1532 63255 1555
rect 63337 1532 63423 1555
rect 63169 1492 63194 1532
rect 63194 1492 63234 1532
rect 63234 1492 63255 1532
rect 63337 1492 63358 1532
rect 63358 1492 63398 1532
rect 63398 1492 63423 1532
rect 63169 1469 63255 1492
rect 63337 1469 63423 1492
rect 67169 1532 67255 1555
rect 67337 1532 67423 1555
rect 67169 1492 67194 1532
rect 67194 1492 67234 1532
rect 67234 1492 67255 1532
rect 67337 1492 67358 1532
rect 67358 1492 67398 1532
rect 67398 1492 67423 1532
rect 67169 1469 67255 1492
rect 67337 1469 67423 1492
rect 71169 1532 71255 1555
rect 71337 1532 71423 1555
rect 71169 1492 71194 1532
rect 71194 1492 71234 1532
rect 71234 1492 71255 1532
rect 71337 1492 71358 1532
rect 71358 1492 71398 1532
rect 71398 1492 71423 1532
rect 71169 1469 71255 1492
rect 71337 1469 71423 1492
rect 75169 1532 75255 1555
rect 75337 1532 75423 1555
rect 75169 1492 75194 1532
rect 75194 1492 75234 1532
rect 75234 1492 75255 1532
rect 75337 1492 75358 1532
rect 75358 1492 75398 1532
rect 75398 1492 75423 1532
rect 75169 1469 75255 1492
rect 75337 1469 75423 1492
rect 79169 1532 79255 1555
rect 79337 1532 79423 1555
rect 79169 1492 79194 1532
rect 79194 1492 79234 1532
rect 79234 1492 79255 1532
rect 79337 1492 79358 1532
rect 79358 1492 79398 1532
rect 79398 1492 79423 1532
rect 79169 1469 79255 1492
rect 79337 1469 79423 1492
rect 83169 1532 83255 1555
rect 83337 1532 83423 1555
rect 83169 1492 83194 1532
rect 83194 1492 83234 1532
rect 83234 1492 83255 1532
rect 83337 1492 83358 1532
rect 83358 1492 83398 1532
rect 83398 1492 83423 1532
rect 83169 1469 83255 1492
rect 83337 1469 83423 1492
rect 87169 1532 87255 1555
rect 87337 1532 87423 1555
rect 87169 1492 87194 1532
rect 87194 1492 87234 1532
rect 87234 1492 87255 1532
rect 87337 1492 87358 1532
rect 87358 1492 87398 1532
rect 87398 1492 87423 1532
rect 87169 1469 87255 1492
rect 87337 1469 87423 1492
rect 91169 1532 91255 1555
rect 91337 1532 91423 1555
rect 91169 1492 91194 1532
rect 91194 1492 91234 1532
rect 91234 1492 91255 1532
rect 91337 1492 91358 1532
rect 91358 1492 91398 1532
rect 91398 1492 91423 1532
rect 91169 1469 91255 1492
rect 91337 1469 91423 1492
rect 95169 1532 95255 1555
rect 95337 1532 95423 1555
rect 95169 1492 95194 1532
rect 95194 1492 95234 1532
rect 95234 1492 95255 1532
rect 95337 1492 95358 1532
rect 95358 1492 95398 1532
rect 95398 1492 95423 1532
rect 95169 1469 95255 1492
rect 95337 1469 95423 1492
rect 99169 1532 99255 1555
rect 99337 1532 99423 1555
rect 99169 1492 99194 1532
rect 99194 1492 99234 1532
rect 99234 1492 99255 1532
rect 99337 1492 99358 1532
rect 99358 1492 99398 1532
rect 99398 1492 99423 1532
rect 99169 1469 99255 1492
rect 99337 1469 99423 1492
rect 4409 776 4495 799
rect 4577 776 4663 799
rect 4409 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4495 776
rect 4577 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4663 776
rect 4409 713 4495 736
rect 4577 713 4663 736
rect 8409 776 8495 799
rect 8577 776 8663 799
rect 8409 736 8434 776
rect 8434 736 8474 776
rect 8474 736 8495 776
rect 8577 736 8598 776
rect 8598 736 8638 776
rect 8638 736 8663 776
rect 8409 713 8495 736
rect 8577 713 8663 736
rect 12409 776 12495 799
rect 12577 776 12663 799
rect 12409 736 12434 776
rect 12434 736 12474 776
rect 12474 736 12495 776
rect 12577 736 12598 776
rect 12598 736 12638 776
rect 12638 736 12663 776
rect 12409 713 12495 736
rect 12577 713 12663 736
rect 16409 776 16495 799
rect 16577 776 16663 799
rect 16409 736 16434 776
rect 16434 736 16474 776
rect 16474 736 16495 776
rect 16577 736 16598 776
rect 16598 736 16638 776
rect 16638 736 16663 776
rect 16409 713 16495 736
rect 16577 713 16663 736
rect 20409 776 20495 799
rect 20577 776 20663 799
rect 20409 736 20434 776
rect 20434 736 20474 776
rect 20474 736 20495 776
rect 20577 736 20598 776
rect 20598 736 20638 776
rect 20638 736 20663 776
rect 20409 713 20495 736
rect 20577 713 20663 736
rect 24409 776 24495 799
rect 24577 776 24663 799
rect 24409 736 24434 776
rect 24434 736 24474 776
rect 24474 736 24495 776
rect 24577 736 24598 776
rect 24598 736 24638 776
rect 24638 736 24663 776
rect 24409 713 24495 736
rect 24577 713 24663 736
rect 28409 776 28495 799
rect 28577 776 28663 799
rect 28409 736 28434 776
rect 28434 736 28474 776
rect 28474 736 28495 776
rect 28577 736 28598 776
rect 28598 736 28638 776
rect 28638 736 28663 776
rect 28409 713 28495 736
rect 28577 713 28663 736
rect 32409 776 32495 799
rect 32577 776 32663 799
rect 32409 736 32434 776
rect 32434 736 32474 776
rect 32474 736 32495 776
rect 32577 736 32598 776
rect 32598 736 32638 776
rect 32638 736 32663 776
rect 32409 713 32495 736
rect 32577 713 32663 736
rect 36409 776 36495 799
rect 36577 776 36663 799
rect 36409 736 36434 776
rect 36434 736 36474 776
rect 36474 736 36495 776
rect 36577 736 36598 776
rect 36598 736 36638 776
rect 36638 736 36663 776
rect 36409 713 36495 736
rect 36577 713 36663 736
rect 40409 776 40495 799
rect 40577 776 40663 799
rect 40409 736 40434 776
rect 40434 736 40474 776
rect 40474 736 40495 776
rect 40577 736 40598 776
rect 40598 736 40638 776
rect 40638 736 40663 776
rect 40409 713 40495 736
rect 40577 713 40663 736
rect 44409 776 44495 799
rect 44577 776 44663 799
rect 44409 736 44434 776
rect 44434 736 44474 776
rect 44474 736 44495 776
rect 44577 736 44598 776
rect 44598 736 44638 776
rect 44638 736 44663 776
rect 44409 713 44495 736
rect 44577 713 44663 736
rect 48409 776 48495 799
rect 48577 776 48663 799
rect 48409 736 48434 776
rect 48434 736 48474 776
rect 48474 736 48495 776
rect 48577 736 48598 776
rect 48598 736 48638 776
rect 48638 736 48663 776
rect 48409 713 48495 736
rect 48577 713 48663 736
rect 52409 776 52495 799
rect 52577 776 52663 799
rect 52409 736 52434 776
rect 52434 736 52474 776
rect 52474 736 52495 776
rect 52577 736 52598 776
rect 52598 736 52638 776
rect 52638 736 52663 776
rect 52409 713 52495 736
rect 52577 713 52663 736
rect 56409 776 56495 799
rect 56577 776 56663 799
rect 56409 736 56434 776
rect 56434 736 56474 776
rect 56474 736 56495 776
rect 56577 736 56598 776
rect 56598 736 56638 776
rect 56638 736 56663 776
rect 56409 713 56495 736
rect 56577 713 56663 736
rect 60409 776 60495 799
rect 60577 776 60663 799
rect 60409 736 60434 776
rect 60434 736 60474 776
rect 60474 736 60495 776
rect 60577 736 60598 776
rect 60598 736 60638 776
rect 60638 736 60663 776
rect 60409 713 60495 736
rect 60577 713 60663 736
rect 64409 776 64495 799
rect 64577 776 64663 799
rect 64409 736 64434 776
rect 64434 736 64474 776
rect 64474 736 64495 776
rect 64577 736 64598 776
rect 64598 736 64638 776
rect 64638 736 64663 776
rect 64409 713 64495 736
rect 64577 713 64663 736
rect 68409 776 68495 799
rect 68577 776 68663 799
rect 68409 736 68434 776
rect 68434 736 68474 776
rect 68474 736 68495 776
rect 68577 736 68598 776
rect 68598 736 68638 776
rect 68638 736 68663 776
rect 68409 713 68495 736
rect 68577 713 68663 736
rect 72409 776 72495 799
rect 72577 776 72663 799
rect 72409 736 72434 776
rect 72434 736 72474 776
rect 72474 736 72495 776
rect 72577 736 72598 776
rect 72598 736 72638 776
rect 72638 736 72663 776
rect 72409 713 72495 736
rect 72577 713 72663 736
rect 76409 776 76495 799
rect 76577 776 76663 799
rect 76409 736 76434 776
rect 76434 736 76474 776
rect 76474 736 76495 776
rect 76577 736 76598 776
rect 76598 736 76638 776
rect 76638 736 76663 776
rect 76409 713 76495 736
rect 76577 713 76663 736
rect 80409 776 80495 799
rect 80577 776 80663 799
rect 80409 736 80434 776
rect 80434 736 80474 776
rect 80474 736 80495 776
rect 80577 736 80598 776
rect 80598 736 80638 776
rect 80638 736 80663 776
rect 80409 713 80495 736
rect 80577 713 80663 736
rect 84409 776 84495 799
rect 84577 776 84663 799
rect 84409 736 84434 776
rect 84434 736 84474 776
rect 84474 736 84495 776
rect 84577 736 84598 776
rect 84598 736 84638 776
rect 84638 736 84663 776
rect 84409 713 84495 736
rect 84577 713 84663 736
rect 88409 776 88495 799
rect 88577 776 88663 799
rect 88409 736 88434 776
rect 88434 736 88474 776
rect 88474 736 88495 776
rect 88577 736 88598 776
rect 88598 736 88638 776
rect 88638 736 88663 776
rect 88409 713 88495 736
rect 88577 713 88663 736
rect 92409 776 92495 799
rect 92577 776 92663 799
rect 92409 736 92434 776
rect 92434 736 92474 776
rect 92474 736 92495 776
rect 92577 736 92598 776
rect 92598 736 92638 776
rect 92638 736 92663 776
rect 92409 713 92495 736
rect 92577 713 92663 736
rect 96409 776 96495 799
rect 96577 776 96663 799
rect 96409 736 96434 776
rect 96434 736 96474 776
rect 96474 736 96495 776
rect 96577 736 96598 776
rect 96598 736 96638 776
rect 96638 736 96663 776
rect 96409 713 96495 736
rect 96577 713 96663 736
<< metal6 >>
rect 3076 37843 3516 38600
rect 3076 37757 3169 37843
rect 3255 37757 3337 37843
rect 3423 37757 3516 37843
rect 3076 36331 3516 37757
rect 3076 36245 3169 36331
rect 3255 36245 3337 36331
rect 3423 36245 3516 36331
rect 3076 35666 3516 36245
rect 3076 35286 3106 35666
rect 3486 35286 3516 35666
rect 3076 34819 3516 35286
rect 3076 34733 3169 34819
rect 3255 34733 3337 34819
rect 3423 34733 3516 34819
rect 3076 33307 3516 34733
rect 3076 33221 3169 33307
rect 3255 33221 3337 33307
rect 3423 33221 3516 33307
rect 3076 31795 3516 33221
rect 3076 31709 3169 31795
rect 3255 31709 3337 31795
rect 3423 31709 3516 31795
rect 3076 31666 3516 31709
rect 3076 31286 3106 31666
rect 3486 31286 3516 31666
rect 3076 30283 3516 31286
rect 3076 30197 3169 30283
rect 3255 30197 3337 30283
rect 3423 30197 3516 30283
rect 3076 28771 3516 30197
rect 3076 28685 3169 28771
rect 3255 28685 3337 28771
rect 3423 28685 3516 28771
rect 3076 27666 3516 28685
rect 3076 27286 3106 27666
rect 3486 27286 3516 27666
rect 3076 27259 3516 27286
rect 3076 27173 3169 27259
rect 3255 27173 3337 27259
rect 3423 27173 3516 27259
rect 3076 25747 3516 27173
rect 3076 25661 3169 25747
rect 3255 25661 3337 25747
rect 3423 25661 3516 25747
rect 3076 24235 3516 25661
rect 3076 24149 3169 24235
rect 3255 24149 3337 24235
rect 3423 24149 3516 24235
rect 3076 23666 3516 24149
rect 3076 23286 3106 23666
rect 3486 23286 3516 23666
rect 3076 22723 3516 23286
rect 3076 22637 3169 22723
rect 3255 22637 3337 22723
rect 3423 22637 3516 22723
rect 3076 21211 3516 22637
rect 3076 21125 3169 21211
rect 3255 21125 3337 21211
rect 3423 21125 3516 21211
rect 3076 19699 3516 21125
rect 3076 19666 3169 19699
rect 3255 19666 3337 19699
rect 3423 19666 3516 19699
rect 3076 19286 3106 19666
rect 3486 19286 3516 19666
rect 3076 18187 3516 19286
rect 3076 18101 3169 18187
rect 3255 18101 3337 18187
rect 3423 18101 3516 18187
rect 3076 16675 3516 18101
rect 3076 16589 3169 16675
rect 3255 16589 3337 16675
rect 3423 16589 3516 16675
rect 3076 15666 3516 16589
rect 3076 15286 3106 15666
rect 3486 15286 3516 15666
rect 3076 15163 3516 15286
rect 3076 15077 3169 15163
rect 3255 15077 3337 15163
rect 3423 15077 3516 15163
rect 3076 13651 3516 15077
rect 3076 13565 3169 13651
rect 3255 13565 3337 13651
rect 3423 13565 3516 13651
rect 3076 12139 3516 13565
rect 3076 12053 3169 12139
rect 3255 12053 3337 12139
rect 3423 12053 3516 12139
rect 3076 11666 3516 12053
rect 3076 11286 3106 11666
rect 3486 11286 3516 11666
rect 3076 10627 3516 11286
rect 3076 10541 3169 10627
rect 3255 10541 3337 10627
rect 3423 10541 3516 10627
rect 3076 9115 3516 10541
rect 3076 9029 3169 9115
rect 3255 9029 3337 9115
rect 3423 9029 3516 9115
rect 3076 7666 3516 9029
rect 3076 7286 3106 7666
rect 3486 7286 3516 7666
rect 3076 6091 3516 7286
rect 3076 6005 3169 6091
rect 3255 6005 3337 6091
rect 3423 6005 3516 6091
rect 3076 4579 3516 6005
rect 3076 4493 3169 4579
rect 3255 4493 3337 4579
rect 3423 4493 3516 4579
rect 3076 3666 3516 4493
rect 3076 3286 3106 3666
rect 3486 3286 3516 3666
rect 3076 3067 3516 3286
rect 3076 2981 3169 3067
rect 3255 2981 3337 3067
rect 3423 2981 3516 3067
rect 3076 1555 3516 2981
rect 3076 1469 3169 1555
rect 3255 1469 3337 1555
rect 3423 1469 3516 1555
rect 3076 712 3516 1469
rect 4316 38599 4756 38682
rect 4316 38513 4409 38599
rect 4495 38513 4577 38599
rect 4663 38513 4756 38599
rect 4316 37087 4756 38513
rect 4316 37001 4409 37087
rect 4495 37001 4577 37087
rect 4663 37001 4756 37087
rect 4316 36906 4756 37001
rect 4316 36526 4346 36906
rect 4726 36526 4756 36906
rect 4316 35575 4756 36526
rect 4316 35489 4409 35575
rect 4495 35489 4577 35575
rect 4663 35489 4756 35575
rect 4316 34063 4756 35489
rect 4316 33977 4409 34063
rect 4495 33977 4577 34063
rect 4663 33977 4756 34063
rect 4316 32906 4756 33977
rect 4316 32526 4346 32906
rect 4726 32526 4756 32906
rect 4316 32465 4409 32526
rect 4495 32465 4577 32526
rect 4663 32465 4756 32526
rect 4316 31039 4756 32465
rect 4316 30953 4409 31039
rect 4495 30953 4577 31039
rect 4663 30953 4756 31039
rect 4316 29527 4756 30953
rect 4316 29441 4409 29527
rect 4495 29441 4577 29527
rect 4663 29441 4756 29527
rect 4316 28906 4756 29441
rect 4316 28526 4346 28906
rect 4726 28526 4756 28906
rect 4316 28015 4756 28526
rect 4316 27929 4409 28015
rect 4495 27929 4577 28015
rect 4663 27929 4756 28015
rect 4316 26503 4756 27929
rect 4316 26417 4409 26503
rect 4495 26417 4577 26503
rect 4663 26417 4756 26503
rect 4316 24991 4756 26417
rect 4316 24906 4409 24991
rect 4495 24906 4577 24991
rect 4663 24906 4756 24991
rect 4316 24526 4346 24906
rect 4726 24526 4756 24906
rect 4316 23479 4756 24526
rect 4316 23393 4409 23479
rect 4495 23393 4577 23479
rect 4663 23393 4756 23479
rect 4316 21967 4756 23393
rect 4316 21881 4409 21967
rect 4495 21881 4577 21967
rect 4663 21881 4756 21967
rect 4316 20906 4756 21881
rect 4316 20526 4346 20906
rect 4726 20526 4756 20906
rect 4316 20455 4756 20526
rect 4316 20369 4409 20455
rect 4495 20369 4577 20455
rect 4663 20369 4756 20455
rect 4316 18943 4756 20369
rect 4316 18857 4409 18943
rect 4495 18857 4577 18943
rect 4663 18857 4756 18943
rect 4316 17431 4756 18857
rect 4316 17345 4409 17431
rect 4495 17345 4577 17431
rect 4663 17345 4756 17431
rect 4316 16906 4756 17345
rect 4316 16526 4346 16906
rect 4726 16526 4756 16906
rect 4316 15919 4756 16526
rect 4316 15833 4409 15919
rect 4495 15833 4577 15919
rect 4663 15833 4756 15919
rect 4316 14407 4756 15833
rect 4316 14321 4409 14407
rect 4495 14321 4577 14407
rect 4663 14321 4756 14407
rect 4316 12906 4756 14321
rect 4316 12526 4346 12906
rect 4726 12526 4756 12906
rect 4316 11383 4756 12526
rect 4316 11297 4409 11383
rect 4495 11297 4577 11383
rect 4663 11297 4756 11383
rect 4316 9871 4756 11297
rect 4316 9785 4409 9871
rect 4495 9785 4577 9871
rect 4663 9785 4756 9871
rect 4316 8906 4756 9785
rect 4316 8526 4346 8906
rect 4726 8526 4756 8906
rect 4316 8359 4756 8526
rect 4316 8273 4409 8359
rect 4495 8273 4577 8359
rect 4663 8273 4756 8359
rect 4316 6847 4756 8273
rect 4316 6761 4409 6847
rect 4495 6761 4577 6847
rect 4663 6761 4756 6847
rect 4316 5335 4756 6761
rect 4316 5249 4409 5335
rect 4495 5249 4577 5335
rect 4663 5249 4756 5335
rect 4316 4906 4756 5249
rect 4316 4526 4346 4906
rect 4726 4526 4756 4906
rect 4316 3823 4756 4526
rect 4316 3737 4409 3823
rect 4495 3737 4577 3823
rect 4663 3737 4756 3823
rect 4316 2311 4756 3737
rect 4316 2225 4409 2311
rect 4495 2225 4577 2311
rect 4663 2225 4756 2311
rect 4316 799 4756 2225
rect 4316 713 4409 799
rect 4495 713 4577 799
rect 4663 713 4756 799
rect 4316 630 4756 713
rect 7076 37843 7516 38600
rect 7076 37757 7169 37843
rect 7255 37757 7337 37843
rect 7423 37757 7516 37843
rect 7076 36331 7516 37757
rect 7076 36245 7169 36331
rect 7255 36245 7337 36331
rect 7423 36245 7516 36331
rect 7076 35666 7516 36245
rect 7076 35286 7106 35666
rect 7486 35286 7516 35666
rect 7076 34819 7516 35286
rect 7076 34733 7169 34819
rect 7255 34733 7337 34819
rect 7423 34733 7516 34819
rect 7076 33307 7516 34733
rect 7076 33221 7169 33307
rect 7255 33221 7337 33307
rect 7423 33221 7516 33307
rect 7076 31795 7516 33221
rect 7076 31709 7169 31795
rect 7255 31709 7337 31795
rect 7423 31709 7516 31795
rect 7076 31666 7516 31709
rect 7076 31286 7106 31666
rect 7486 31286 7516 31666
rect 7076 30283 7516 31286
rect 7076 30197 7169 30283
rect 7255 30197 7337 30283
rect 7423 30197 7516 30283
rect 7076 28771 7516 30197
rect 7076 28685 7169 28771
rect 7255 28685 7337 28771
rect 7423 28685 7516 28771
rect 7076 27666 7516 28685
rect 7076 27286 7106 27666
rect 7486 27286 7516 27666
rect 7076 27259 7516 27286
rect 7076 27173 7169 27259
rect 7255 27173 7337 27259
rect 7423 27173 7516 27259
rect 7076 25747 7516 27173
rect 7076 25661 7169 25747
rect 7255 25661 7337 25747
rect 7423 25661 7516 25747
rect 7076 24235 7516 25661
rect 7076 24149 7169 24235
rect 7255 24149 7337 24235
rect 7423 24149 7516 24235
rect 7076 23666 7516 24149
rect 7076 23286 7106 23666
rect 7486 23286 7516 23666
rect 7076 22723 7516 23286
rect 7076 22637 7169 22723
rect 7255 22637 7337 22723
rect 7423 22637 7516 22723
rect 7076 21211 7516 22637
rect 7076 21125 7169 21211
rect 7255 21125 7337 21211
rect 7423 21125 7516 21211
rect 7076 19699 7516 21125
rect 7076 19666 7169 19699
rect 7255 19666 7337 19699
rect 7423 19666 7516 19699
rect 7076 19286 7106 19666
rect 7486 19286 7516 19666
rect 7076 18187 7516 19286
rect 7076 18101 7169 18187
rect 7255 18101 7337 18187
rect 7423 18101 7516 18187
rect 7076 16675 7516 18101
rect 7076 16589 7169 16675
rect 7255 16589 7337 16675
rect 7423 16589 7516 16675
rect 7076 15666 7516 16589
rect 7076 15286 7106 15666
rect 7486 15286 7516 15666
rect 7076 15163 7516 15286
rect 7076 15077 7169 15163
rect 7255 15077 7337 15163
rect 7423 15077 7516 15163
rect 7076 13651 7516 15077
rect 7076 13565 7169 13651
rect 7255 13565 7337 13651
rect 7423 13565 7516 13651
rect 7076 12139 7516 13565
rect 7076 12053 7169 12139
rect 7255 12053 7337 12139
rect 7423 12053 7516 12139
rect 7076 11666 7516 12053
rect 7076 11286 7106 11666
rect 7486 11286 7516 11666
rect 7076 10627 7516 11286
rect 7076 10541 7169 10627
rect 7255 10541 7337 10627
rect 7423 10541 7516 10627
rect 7076 9115 7516 10541
rect 7076 9029 7169 9115
rect 7255 9029 7337 9115
rect 7423 9029 7516 9115
rect 7076 7666 7516 9029
rect 7076 7286 7106 7666
rect 7486 7286 7516 7666
rect 7076 6091 7516 7286
rect 7076 6005 7169 6091
rect 7255 6005 7337 6091
rect 7423 6005 7516 6091
rect 7076 4579 7516 6005
rect 7076 4493 7169 4579
rect 7255 4493 7337 4579
rect 7423 4493 7516 4579
rect 7076 3666 7516 4493
rect 7076 3286 7106 3666
rect 7486 3286 7516 3666
rect 7076 3067 7516 3286
rect 7076 2981 7169 3067
rect 7255 2981 7337 3067
rect 7423 2981 7516 3067
rect 7076 1555 7516 2981
rect 7076 1469 7169 1555
rect 7255 1469 7337 1555
rect 7423 1469 7516 1555
rect 7076 712 7516 1469
rect 8316 38599 8756 38682
rect 8316 38513 8409 38599
rect 8495 38513 8577 38599
rect 8663 38513 8756 38599
rect 8316 37087 8756 38513
rect 8316 37001 8409 37087
rect 8495 37001 8577 37087
rect 8663 37001 8756 37087
rect 8316 36906 8756 37001
rect 8316 36526 8346 36906
rect 8726 36526 8756 36906
rect 8316 35575 8756 36526
rect 8316 35489 8409 35575
rect 8495 35489 8577 35575
rect 8663 35489 8756 35575
rect 8316 34063 8756 35489
rect 8316 33977 8409 34063
rect 8495 33977 8577 34063
rect 8663 33977 8756 34063
rect 8316 32906 8756 33977
rect 8316 32526 8346 32906
rect 8726 32526 8756 32906
rect 8316 32465 8409 32526
rect 8495 32465 8577 32526
rect 8663 32465 8756 32526
rect 8316 31039 8756 32465
rect 8316 30953 8409 31039
rect 8495 30953 8577 31039
rect 8663 30953 8756 31039
rect 8316 29527 8756 30953
rect 8316 29441 8409 29527
rect 8495 29441 8577 29527
rect 8663 29441 8756 29527
rect 8316 28906 8756 29441
rect 8316 28526 8346 28906
rect 8726 28526 8756 28906
rect 8316 28015 8756 28526
rect 8316 27929 8409 28015
rect 8495 27929 8577 28015
rect 8663 27929 8756 28015
rect 8316 26503 8756 27929
rect 8316 26417 8409 26503
rect 8495 26417 8577 26503
rect 8663 26417 8756 26503
rect 8316 24991 8756 26417
rect 8316 24906 8409 24991
rect 8495 24906 8577 24991
rect 8663 24906 8756 24991
rect 8316 24526 8346 24906
rect 8726 24526 8756 24906
rect 8316 23479 8756 24526
rect 8316 23393 8409 23479
rect 8495 23393 8577 23479
rect 8663 23393 8756 23479
rect 8316 21967 8756 23393
rect 8316 21881 8409 21967
rect 8495 21881 8577 21967
rect 8663 21881 8756 21967
rect 8316 20906 8756 21881
rect 8316 20526 8346 20906
rect 8726 20526 8756 20906
rect 8316 20455 8756 20526
rect 8316 20369 8409 20455
rect 8495 20369 8577 20455
rect 8663 20369 8756 20455
rect 8316 18943 8756 20369
rect 8316 18857 8409 18943
rect 8495 18857 8577 18943
rect 8663 18857 8756 18943
rect 8316 17431 8756 18857
rect 8316 17345 8409 17431
rect 8495 17345 8577 17431
rect 8663 17345 8756 17431
rect 8316 16906 8756 17345
rect 8316 16526 8346 16906
rect 8726 16526 8756 16906
rect 8316 15919 8756 16526
rect 8316 15833 8409 15919
rect 8495 15833 8577 15919
rect 8663 15833 8756 15919
rect 8316 14407 8756 15833
rect 8316 14321 8409 14407
rect 8495 14321 8577 14407
rect 8663 14321 8756 14407
rect 8316 12906 8756 14321
rect 8316 12526 8346 12906
rect 8726 12526 8756 12906
rect 8316 11383 8756 12526
rect 8316 11297 8409 11383
rect 8495 11297 8577 11383
rect 8663 11297 8756 11383
rect 8316 9871 8756 11297
rect 8316 9785 8409 9871
rect 8495 9785 8577 9871
rect 8663 9785 8756 9871
rect 8316 8906 8756 9785
rect 8316 8526 8346 8906
rect 8726 8526 8756 8906
rect 8316 8359 8756 8526
rect 8316 8273 8409 8359
rect 8495 8273 8577 8359
rect 8663 8273 8756 8359
rect 8316 6847 8756 8273
rect 8316 6761 8409 6847
rect 8495 6761 8577 6847
rect 8663 6761 8756 6847
rect 8316 5335 8756 6761
rect 8316 5249 8409 5335
rect 8495 5249 8577 5335
rect 8663 5249 8756 5335
rect 8316 4906 8756 5249
rect 8316 4526 8346 4906
rect 8726 4526 8756 4906
rect 8316 3823 8756 4526
rect 8316 3737 8409 3823
rect 8495 3737 8577 3823
rect 8663 3737 8756 3823
rect 8316 2311 8756 3737
rect 8316 2225 8409 2311
rect 8495 2225 8577 2311
rect 8663 2225 8756 2311
rect 8316 799 8756 2225
rect 8316 713 8409 799
rect 8495 713 8577 799
rect 8663 713 8756 799
rect 8316 630 8756 713
rect 11076 37843 11516 38600
rect 11076 37757 11169 37843
rect 11255 37757 11337 37843
rect 11423 37757 11516 37843
rect 11076 36331 11516 37757
rect 11076 36245 11169 36331
rect 11255 36245 11337 36331
rect 11423 36245 11516 36331
rect 11076 35666 11516 36245
rect 11076 35286 11106 35666
rect 11486 35286 11516 35666
rect 11076 34819 11516 35286
rect 11076 34733 11169 34819
rect 11255 34733 11337 34819
rect 11423 34733 11516 34819
rect 11076 33307 11516 34733
rect 11076 33221 11169 33307
rect 11255 33221 11337 33307
rect 11423 33221 11516 33307
rect 11076 31795 11516 33221
rect 11076 31709 11169 31795
rect 11255 31709 11337 31795
rect 11423 31709 11516 31795
rect 11076 31666 11516 31709
rect 11076 31286 11106 31666
rect 11486 31286 11516 31666
rect 11076 30283 11516 31286
rect 11076 30197 11169 30283
rect 11255 30197 11337 30283
rect 11423 30197 11516 30283
rect 11076 28771 11516 30197
rect 11076 28685 11169 28771
rect 11255 28685 11337 28771
rect 11423 28685 11516 28771
rect 11076 27666 11516 28685
rect 11076 27286 11106 27666
rect 11486 27286 11516 27666
rect 11076 27259 11516 27286
rect 11076 27173 11169 27259
rect 11255 27173 11337 27259
rect 11423 27173 11516 27259
rect 11076 25747 11516 27173
rect 11076 25661 11169 25747
rect 11255 25661 11337 25747
rect 11423 25661 11516 25747
rect 11076 24235 11516 25661
rect 11076 24149 11169 24235
rect 11255 24149 11337 24235
rect 11423 24149 11516 24235
rect 11076 23666 11516 24149
rect 11076 23286 11106 23666
rect 11486 23286 11516 23666
rect 11076 22723 11516 23286
rect 11076 22637 11169 22723
rect 11255 22637 11337 22723
rect 11423 22637 11516 22723
rect 11076 21211 11516 22637
rect 11076 21125 11169 21211
rect 11255 21125 11337 21211
rect 11423 21125 11516 21211
rect 11076 19699 11516 21125
rect 11076 19666 11169 19699
rect 11255 19666 11337 19699
rect 11423 19666 11516 19699
rect 11076 19286 11106 19666
rect 11486 19286 11516 19666
rect 11076 18187 11516 19286
rect 11076 18101 11169 18187
rect 11255 18101 11337 18187
rect 11423 18101 11516 18187
rect 11076 16675 11516 18101
rect 11076 16589 11169 16675
rect 11255 16589 11337 16675
rect 11423 16589 11516 16675
rect 11076 15666 11516 16589
rect 11076 15286 11106 15666
rect 11486 15286 11516 15666
rect 11076 15163 11516 15286
rect 11076 15077 11169 15163
rect 11255 15077 11337 15163
rect 11423 15077 11516 15163
rect 11076 13651 11516 15077
rect 11076 13565 11169 13651
rect 11255 13565 11337 13651
rect 11423 13565 11516 13651
rect 11076 12139 11516 13565
rect 11076 12053 11169 12139
rect 11255 12053 11337 12139
rect 11423 12053 11516 12139
rect 11076 11666 11516 12053
rect 11076 11286 11106 11666
rect 11486 11286 11516 11666
rect 11076 10627 11516 11286
rect 11076 10541 11169 10627
rect 11255 10541 11337 10627
rect 11423 10541 11516 10627
rect 11076 9115 11516 10541
rect 11076 9029 11169 9115
rect 11255 9029 11337 9115
rect 11423 9029 11516 9115
rect 11076 7666 11516 9029
rect 11076 7286 11106 7666
rect 11486 7286 11516 7666
rect 11076 6091 11516 7286
rect 11076 6005 11169 6091
rect 11255 6005 11337 6091
rect 11423 6005 11516 6091
rect 11076 4579 11516 6005
rect 11076 4493 11169 4579
rect 11255 4493 11337 4579
rect 11423 4493 11516 4579
rect 11076 3666 11516 4493
rect 11076 3286 11106 3666
rect 11486 3286 11516 3666
rect 11076 3067 11516 3286
rect 11076 2981 11169 3067
rect 11255 2981 11337 3067
rect 11423 2981 11516 3067
rect 11076 1555 11516 2981
rect 11076 1469 11169 1555
rect 11255 1469 11337 1555
rect 11423 1469 11516 1555
rect 11076 712 11516 1469
rect 12316 38599 12756 38682
rect 12316 38513 12409 38599
rect 12495 38513 12577 38599
rect 12663 38513 12756 38599
rect 12316 37087 12756 38513
rect 12316 37001 12409 37087
rect 12495 37001 12577 37087
rect 12663 37001 12756 37087
rect 12316 36906 12756 37001
rect 12316 36526 12346 36906
rect 12726 36526 12756 36906
rect 12316 35575 12756 36526
rect 12316 35489 12409 35575
rect 12495 35489 12577 35575
rect 12663 35489 12756 35575
rect 12316 34063 12756 35489
rect 12316 33977 12409 34063
rect 12495 33977 12577 34063
rect 12663 33977 12756 34063
rect 12316 32906 12756 33977
rect 12316 32526 12346 32906
rect 12726 32526 12756 32906
rect 12316 32465 12409 32526
rect 12495 32465 12577 32526
rect 12663 32465 12756 32526
rect 12316 31039 12756 32465
rect 12316 30953 12409 31039
rect 12495 30953 12577 31039
rect 12663 30953 12756 31039
rect 12316 29527 12756 30953
rect 12316 29441 12409 29527
rect 12495 29441 12577 29527
rect 12663 29441 12756 29527
rect 12316 28906 12756 29441
rect 12316 28526 12346 28906
rect 12726 28526 12756 28906
rect 12316 28015 12756 28526
rect 12316 27929 12409 28015
rect 12495 27929 12577 28015
rect 12663 27929 12756 28015
rect 12316 26503 12756 27929
rect 12316 26417 12409 26503
rect 12495 26417 12577 26503
rect 12663 26417 12756 26503
rect 12316 24991 12756 26417
rect 12316 24906 12409 24991
rect 12495 24906 12577 24991
rect 12663 24906 12756 24991
rect 12316 24526 12346 24906
rect 12726 24526 12756 24906
rect 12316 23479 12756 24526
rect 12316 23393 12409 23479
rect 12495 23393 12577 23479
rect 12663 23393 12756 23479
rect 12316 21967 12756 23393
rect 12316 21881 12409 21967
rect 12495 21881 12577 21967
rect 12663 21881 12756 21967
rect 12316 20906 12756 21881
rect 12316 20526 12346 20906
rect 12726 20526 12756 20906
rect 12316 20455 12756 20526
rect 12316 20369 12409 20455
rect 12495 20369 12577 20455
rect 12663 20369 12756 20455
rect 12316 18943 12756 20369
rect 12316 18857 12409 18943
rect 12495 18857 12577 18943
rect 12663 18857 12756 18943
rect 12316 17431 12756 18857
rect 12316 17345 12409 17431
rect 12495 17345 12577 17431
rect 12663 17345 12756 17431
rect 12316 16906 12756 17345
rect 12316 16526 12346 16906
rect 12726 16526 12756 16906
rect 12316 15919 12756 16526
rect 12316 15833 12409 15919
rect 12495 15833 12577 15919
rect 12663 15833 12756 15919
rect 12316 14407 12756 15833
rect 12316 14321 12409 14407
rect 12495 14321 12577 14407
rect 12663 14321 12756 14407
rect 12316 12906 12756 14321
rect 12316 12526 12346 12906
rect 12726 12526 12756 12906
rect 12316 11383 12756 12526
rect 12316 11297 12409 11383
rect 12495 11297 12577 11383
rect 12663 11297 12756 11383
rect 12316 9871 12756 11297
rect 12316 9785 12409 9871
rect 12495 9785 12577 9871
rect 12663 9785 12756 9871
rect 12316 8906 12756 9785
rect 12316 8526 12346 8906
rect 12726 8526 12756 8906
rect 12316 8359 12756 8526
rect 12316 8273 12409 8359
rect 12495 8273 12577 8359
rect 12663 8273 12756 8359
rect 12316 6847 12756 8273
rect 12316 6761 12409 6847
rect 12495 6761 12577 6847
rect 12663 6761 12756 6847
rect 12316 5335 12756 6761
rect 12316 5249 12409 5335
rect 12495 5249 12577 5335
rect 12663 5249 12756 5335
rect 12316 4906 12756 5249
rect 12316 4526 12346 4906
rect 12726 4526 12756 4906
rect 12316 3823 12756 4526
rect 12316 3737 12409 3823
rect 12495 3737 12577 3823
rect 12663 3737 12756 3823
rect 12316 2311 12756 3737
rect 12316 2225 12409 2311
rect 12495 2225 12577 2311
rect 12663 2225 12756 2311
rect 12316 799 12756 2225
rect 12316 713 12409 799
rect 12495 713 12577 799
rect 12663 713 12756 799
rect 12316 630 12756 713
rect 15076 37843 15516 38600
rect 15076 37757 15169 37843
rect 15255 37757 15337 37843
rect 15423 37757 15516 37843
rect 15076 36331 15516 37757
rect 15076 36245 15169 36331
rect 15255 36245 15337 36331
rect 15423 36245 15516 36331
rect 15076 35666 15516 36245
rect 15076 35286 15106 35666
rect 15486 35286 15516 35666
rect 15076 34819 15516 35286
rect 15076 34733 15169 34819
rect 15255 34733 15337 34819
rect 15423 34733 15516 34819
rect 15076 33307 15516 34733
rect 15076 33221 15169 33307
rect 15255 33221 15337 33307
rect 15423 33221 15516 33307
rect 15076 31795 15516 33221
rect 15076 31709 15169 31795
rect 15255 31709 15337 31795
rect 15423 31709 15516 31795
rect 15076 31666 15516 31709
rect 15076 31286 15106 31666
rect 15486 31286 15516 31666
rect 15076 30283 15516 31286
rect 15076 30197 15169 30283
rect 15255 30197 15337 30283
rect 15423 30197 15516 30283
rect 15076 28771 15516 30197
rect 15076 28685 15169 28771
rect 15255 28685 15337 28771
rect 15423 28685 15516 28771
rect 15076 27666 15516 28685
rect 15076 27286 15106 27666
rect 15486 27286 15516 27666
rect 15076 27259 15516 27286
rect 15076 27173 15169 27259
rect 15255 27173 15337 27259
rect 15423 27173 15516 27259
rect 15076 25747 15516 27173
rect 15076 25661 15169 25747
rect 15255 25661 15337 25747
rect 15423 25661 15516 25747
rect 15076 24235 15516 25661
rect 15076 24149 15169 24235
rect 15255 24149 15337 24235
rect 15423 24149 15516 24235
rect 15076 23666 15516 24149
rect 15076 23286 15106 23666
rect 15486 23286 15516 23666
rect 15076 22723 15516 23286
rect 15076 22637 15169 22723
rect 15255 22637 15337 22723
rect 15423 22637 15516 22723
rect 15076 21211 15516 22637
rect 15076 21125 15169 21211
rect 15255 21125 15337 21211
rect 15423 21125 15516 21211
rect 15076 19699 15516 21125
rect 15076 19666 15169 19699
rect 15255 19666 15337 19699
rect 15423 19666 15516 19699
rect 15076 19286 15106 19666
rect 15486 19286 15516 19666
rect 15076 18187 15516 19286
rect 15076 18101 15169 18187
rect 15255 18101 15337 18187
rect 15423 18101 15516 18187
rect 15076 16675 15516 18101
rect 15076 16589 15169 16675
rect 15255 16589 15337 16675
rect 15423 16589 15516 16675
rect 15076 15666 15516 16589
rect 15076 15286 15106 15666
rect 15486 15286 15516 15666
rect 15076 15163 15516 15286
rect 15076 15077 15169 15163
rect 15255 15077 15337 15163
rect 15423 15077 15516 15163
rect 15076 13651 15516 15077
rect 15076 13565 15169 13651
rect 15255 13565 15337 13651
rect 15423 13565 15516 13651
rect 15076 12139 15516 13565
rect 15076 12053 15169 12139
rect 15255 12053 15337 12139
rect 15423 12053 15516 12139
rect 15076 11666 15516 12053
rect 15076 11286 15106 11666
rect 15486 11286 15516 11666
rect 15076 10627 15516 11286
rect 15076 10541 15169 10627
rect 15255 10541 15337 10627
rect 15423 10541 15516 10627
rect 15076 9115 15516 10541
rect 15076 9029 15169 9115
rect 15255 9029 15337 9115
rect 15423 9029 15516 9115
rect 15076 7666 15516 9029
rect 15076 7286 15106 7666
rect 15486 7286 15516 7666
rect 15076 6091 15516 7286
rect 15076 6005 15169 6091
rect 15255 6005 15337 6091
rect 15423 6005 15516 6091
rect 15076 4579 15516 6005
rect 15076 4493 15169 4579
rect 15255 4493 15337 4579
rect 15423 4493 15516 4579
rect 15076 3666 15516 4493
rect 15076 3286 15106 3666
rect 15486 3286 15516 3666
rect 15076 3067 15516 3286
rect 15076 2981 15169 3067
rect 15255 2981 15337 3067
rect 15423 2981 15516 3067
rect 15076 1555 15516 2981
rect 15076 1469 15169 1555
rect 15255 1469 15337 1555
rect 15423 1469 15516 1555
rect 15076 712 15516 1469
rect 16316 38599 16756 38682
rect 16316 38513 16409 38599
rect 16495 38513 16577 38599
rect 16663 38513 16756 38599
rect 16316 37087 16756 38513
rect 16316 37001 16409 37087
rect 16495 37001 16577 37087
rect 16663 37001 16756 37087
rect 16316 36906 16756 37001
rect 16316 36526 16346 36906
rect 16726 36526 16756 36906
rect 16316 35575 16756 36526
rect 16316 35489 16409 35575
rect 16495 35489 16577 35575
rect 16663 35489 16756 35575
rect 16316 34063 16756 35489
rect 16316 33977 16409 34063
rect 16495 33977 16577 34063
rect 16663 33977 16756 34063
rect 16316 32906 16756 33977
rect 16316 32526 16346 32906
rect 16726 32526 16756 32906
rect 16316 32465 16409 32526
rect 16495 32465 16577 32526
rect 16663 32465 16756 32526
rect 16316 31039 16756 32465
rect 16316 30953 16409 31039
rect 16495 30953 16577 31039
rect 16663 30953 16756 31039
rect 16316 29527 16756 30953
rect 16316 29441 16409 29527
rect 16495 29441 16577 29527
rect 16663 29441 16756 29527
rect 16316 28906 16756 29441
rect 16316 28526 16346 28906
rect 16726 28526 16756 28906
rect 16316 28015 16756 28526
rect 16316 27929 16409 28015
rect 16495 27929 16577 28015
rect 16663 27929 16756 28015
rect 16316 26503 16756 27929
rect 16316 26417 16409 26503
rect 16495 26417 16577 26503
rect 16663 26417 16756 26503
rect 16316 24991 16756 26417
rect 16316 24906 16409 24991
rect 16495 24906 16577 24991
rect 16663 24906 16756 24991
rect 16316 24526 16346 24906
rect 16726 24526 16756 24906
rect 16316 23479 16756 24526
rect 16316 23393 16409 23479
rect 16495 23393 16577 23479
rect 16663 23393 16756 23479
rect 16316 21967 16756 23393
rect 16316 21881 16409 21967
rect 16495 21881 16577 21967
rect 16663 21881 16756 21967
rect 16316 20906 16756 21881
rect 16316 20526 16346 20906
rect 16726 20526 16756 20906
rect 16316 20455 16756 20526
rect 16316 20369 16409 20455
rect 16495 20369 16577 20455
rect 16663 20369 16756 20455
rect 16316 18943 16756 20369
rect 16316 18857 16409 18943
rect 16495 18857 16577 18943
rect 16663 18857 16756 18943
rect 16316 17431 16756 18857
rect 16316 17345 16409 17431
rect 16495 17345 16577 17431
rect 16663 17345 16756 17431
rect 16316 16906 16756 17345
rect 16316 16526 16346 16906
rect 16726 16526 16756 16906
rect 16316 15919 16756 16526
rect 16316 15833 16409 15919
rect 16495 15833 16577 15919
rect 16663 15833 16756 15919
rect 16316 14407 16756 15833
rect 16316 14321 16409 14407
rect 16495 14321 16577 14407
rect 16663 14321 16756 14407
rect 16316 12906 16756 14321
rect 16316 12526 16346 12906
rect 16726 12526 16756 12906
rect 16316 11383 16756 12526
rect 16316 11297 16409 11383
rect 16495 11297 16577 11383
rect 16663 11297 16756 11383
rect 16316 9871 16756 11297
rect 16316 9785 16409 9871
rect 16495 9785 16577 9871
rect 16663 9785 16756 9871
rect 16316 8906 16756 9785
rect 16316 8526 16346 8906
rect 16726 8526 16756 8906
rect 16316 8359 16756 8526
rect 16316 8273 16409 8359
rect 16495 8273 16577 8359
rect 16663 8273 16756 8359
rect 16316 6847 16756 8273
rect 16316 6761 16409 6847
rect 16495 6761 16577 6847
rect 16663 6761 16756 6847
rect 16316 5335 16756 6761
rect 16316 5249 16409 5335
rect 16495 5249 16577 5335
rect 16663 5249 16756 5335
rect 16316 4906 16756 5249
rect 16316 4526 16346 4906
rect 16726 4526 16756 4906
rect 16316 3823 16756 4526
rect 16316 3737 16409 3823
rect 16495 3737 16577 3823
rect 16663 3737 16756 3823
rect 16316 2311 16756 3737
rect 16316 2225 16409 2311
rect 16495 2225 16577 2311
rect 16663 2225 16756 2311
rect 16316 799 16756 2225
rect 16316 713 16409 799
rect 16495 713 16577 799
rect 16663 713 16756 799
rect 16316 630 16756 713
rect 19076 37843 19516 38600
rect 19076 37757 19169 37843
rect 19255 37757 19337 37843
rect 19423 37757 19516 37843
rect 19076 36331 19516 37757
rect 19076 36245 19169 36331
rect 19255 36245 19337 36331
rect 19423 36245 19516 36331
rect 19076 35666 19516 36245
rect 19076 35286 19106 35666
rect 19486 35286 19516 35666
rect 19076 34819 19516 35286
rect 19076 34733 19169 34819
rect 19255 34733 19337 34819
rect 19423 34733 19516 34819
rect 19076 33307 19516 34733
rect 19076 33221 19169 33307
rect 19255 33221 19337 33307
rect 19423 33221 19516 33307
rect 19076 31795 19516 33221
rect 19076 31709 19169 31795
rect 19255 31709 19337 31795
rect 19423 31709 19516 31795
rect 19076 31666 19516 31709
rect 19076 31286 19106 31666
rect 19486 31286 19516 31666
rect 19076 30283 19516 31286
rect 19076 30197 19169 30283
rect 19255 30197 19337 30283
rect 19423 30197 19516 30283
rect 19076 28771 19516 30197
rect 19076 28685 19169 28771
rect 19255 28685 19337 28771
rect 19423 28685 19516 28771
rect 19076 27666 19516 28685
rect 19076 27286 19106 27666
rect 19486 27286 19516 27666
rect 19076 27259 19516 27286
rect 19076 27173 19169 27259
rect 19255 27173 19337 27259
rect 19423 27173 19516 27259
rect 19076 25747 19516 27173
rect 19076 25661 19169 25747
rect 19255 25661 19337 25747
rect 19423 25661 19516 25747
rect 19076 24235 19516 25661
rect 19076 24149 19169 24235
rect 19255 24149 19337 24235
rect 19423 24149 19516 24235
rect 19076 23666 19516 24149
rect 19076 23286 19106 23666
rect 19486 23286 19516 23666
rect 19076 22723 19516 23286
rect 19076 22637 19169 22723
rect 19255 22637 19337 22723
rect 19423 22637 19516 22723
rect 19076 21211 19516 22637
rect 19076 21125 19169 21211
rect 19255 21125 19337 21211
rect 19423 21125 19516 21211
rect 19076 19699 19516 21125
rect 19076 19666 19169 19699
rect 19255 19666 19337 19699
rect 19423 19666 19516 19699
rect 19076 19286 19106 19666
rect 19486 19286 19516 19666
rect 19076 18187 19516 19286
rect 19076 18101 19169 18187
rect 19255 18101 19337 18187
rect 19423 18101 19516 18187
rect 19076 16675 19516 18101
rect 19076 16589 19169 16675
rect 19255 16589 19337 16675
rect 19423 16589 19516 16675
rect 19076 15666 19516 16589
rect 19076 15286 19106 15666
rect 19486 15286 19516 15666
rect 19076 15163 19516 15286
rect 19076 15077 19169 15163
rect 19255 15077 19337 15163
rect 19423 15077 19516 15163
rect 19076 13651 19516 15077
rect 19076 13565 19169 13651
rect 19255 13565 19337 13651
rect 19423 13565 19516 13651
rect 19076 12139 19516 13565
rect 19076 12053 19169 12139
rect 19255 12053 19337 12139
rect 19423 12053 19516 12139
rect 19076 11666 19516 12053
rect 19076 11286 19106 11666
rect 19486 11286 19516 11666
rect 19076 10627 19516 11286
rect 19076 10541 19169 10627
rect 19255 10541 19337 10627
rect 19423 10541 19516 10627
rect 19076 9115 19516 10541
rect 19076 9029 19169 9115
rect 19255 9029 19337 9115
rect 19423 9029 19516 9115
rect 19076 7666 19516 9029
rect 19076 7286 19106 7666
rect 19486 7286 19516 7666
rect 19076 6091 19516 7286
rect 19076 6005 19169 6091
rect 19255 6005 19337 6091
rect 19423 6005 19516 6091
rect 19076 4579 19516 6005
rect 19076 4493 19169 4579
rect 19255 4493 19337 4579
rect 19423 4493 19516 4579
rect 19076 3666 19516 4493
rect 19076 3286 19106 3666
rect 19486 3286 19516 3666
rect 19076 3067 19516 3286
rect 19076 2981 19169 3067
rect 19255 2981 19337 3067
rect 19423 2981 19516 3067
rect 19076 1555 19516 2981
rect 19076 1469 19169 1555
rect 19255 1469 19337 1555
rect 19423 1469 19516 1555
rect 19076 712 19516 1469
rect 20316 38599 20756 38682
rect 20316 38513 20409 38599
rect 20495 38513 20577 38599
rect 20663 38513 20756 38599
rect 20316 37087 20756 38513
rect 20316 37001 20409 37087
rect 20495 37001 20577 37087
rect 20663 37001 20756 37087
rect 20316 36906 20756 37001
rect 20316 36526 20346 36906
rect 20726 36526 20756 36906
rect 20316 35575 20756 36526
rect 20316 35489 20409 35575
rect 20495 35489 20577 35575
rect 20663 35489 20756 35575
rect 20316 34063 20756 35489
rect 20316 33977 20409 34063
rect 20495 33977 20577 34063
rect 20663 33977 20756 34063
rect 20316 32906 20756 33977
rect 20316 32526 20346 32906
rect 20726 32526 20756 32906
rect 20316 32465 20409 32526
rect 20495 32465 20577 32526
rect 20663 32465 20756 32526
rect 20316 31039 20756 32465
rect 20316 30953 20409 31039
rect 20495 30953 20577 31039
rect 20663 30953 20756 31039
rect 20316 29527 20756 30953
rect 20316 29441 20409 29527
rect 20495 29441 20577 29527
rect 20663 29441 20756 29527
rect 20316 28906 20756 29441
rect 20316 28526 20346 28906
rect 20726 28526 20756 28906
rect 20316 28015 20756 28526
rect 20316 27929 20409 28015
rect 20495 27929 20577 28015
rect 20663 27929 20756 28015
rect 20316 26503 20756 27929
rect 20316 26417 20409 26503
rect 20495 26417 20577 26503
rect 20663 26417 20756 26503
rect 20316 24991 20756 26417
rect 20316 24906 20409 24991
rect 20495 24906 20577 24991
rect 20663 24906 20756 24991
rect 20316 24526 20346 24906
rect 20726 24526 20756 24906
rect 20316 23479 20756 24526
rect 20316 23393 20409 23479
rect 20495 23393 20577 23479
rect 20663 23393 20756 23479
rect 20316 21967 20756 23393
rect 20316 21881 20409 21967
rect 20495 21881 20577 21967
rect 20663 21881 20756 21967
rect 20316 20906 20756 21881
rect 20316 20526 20346 20906
rect 20726 20526 20756 20906
rect 20316 20455 20756 20526
rect 20316 20369 20409 20455
rect 20495 20369 20577 20455
rect 20663 20369 20756 20455
rect 20316 18943 20756 20369
rect 20316 18857 20409 18943
rect 20495 18857 20577 18943
rect 20663 18857 20756 18943
rect 20316 17431 20756 18857
rect 20316 17345 20409 17431
rect 20495 17345 20577 17431
rect 20663 17345 20756 17431
rect 20316 16906 20756 17345
rect 20316 16526 20346 16906
rect 20726 16526 20756 16906
rect 20316 15919 20756 16526
rect 20316 15833 20409 15919
rect 20495 15833 20577 15919
rect 20663 15833 20756 15919
rect 20316 14407 20756 15833
rect 20316 14321 20409 14407
rect 20495 14321 20577 14407
rect 20663 14321 20756 14407
rect 20316 12906 20756 14321
rect 20316 12526 20346 12906
rect 20726 12526 20756 12906
rect 20316 11383 20756 12526
rect 20316 11297 20409 11383
rect 20495 11297 20577 11383
rect 20663 11297 20756 11383
rect 20316 9871 20756 11297
rect 20316 9785 20409 9871
rect 20495 9785 20577 9871
rect 20663 9785 20756 9871
rect 20316 8906 20756 9785
rect 20316 8526 20346 8906
rect 20726 8526 20756 8906
rect 20316 8359 20756 8526
rect 20316 8273 20409 8359
rect 20495 8273 20577 8359
rect 20663 8273 20756 8359
rect 20316 6847 20756 8273
rect 20316 6761 20409 6847
rect 20495 6761 20577 6847
rect 20663 6761 20756 6847
rect 20316 5335 20756 6761
rect 20316 5249 20409 5335
rect 20495 5249 20577 5335
rect 20663 5249 20756 5335
rect 20316 4906 20756 5249
rect 20316 4526 20346 4906
rect 20726 4526 20756 4906
rect 20316 3823 20756 4526
rect 20316 3737 20409 3823
rect 20495 3737 20577 3823
rect 20663 3737 20756 3823
rect 20316 2311 20756 3737
rect 20316 2225 20409 2311
rect 20495 2225 20577 2311
rect 20663 2225 20756 2311
rect 20316 799 20756 2225
rect 20316 713 20409 799
rect 20495 713 20577 799
rect 20663 713 20756 799
rect 20316 630 20756 713
rect 23076 37843 23516 38600
rect 23076 37757 23169 37843
rect 23255 37757 23337 37843
rect 23423 37757 23516 37843
rect 23076 36331 23516 37757
rect 23076 36245 23169 36331
rect 23255 36245 23337 36331
rect 23423 36245 23516 36331
rect 23076 35666 23516 36245
rect 23076 35286 23106 35666
rect 23486 35286 23516 35666
rect 23076 34819 23516 35286
rect 23076 34733 23169 34819
rect 23255 34733 23337 34819
rect 23423 34733 23516 34819
rect 23076 33307 23516 34733
rect 23076 33221 23169 33307
rect 23255 33221 23337 33307
rect 23423 33221 23516 33307
rect 23076 31795 23516 33221
rect 23076 31709 23169 31795
rect 23255 31709 23337 31795
rect 23423 31709 23516 31795
rect 23076 31666 23516 31709
rect 23076 31286 23106 31666
rect 23486 31286 23516 31666
rect 23076 30283 23516 31286
rect 23076 30197 23169 30283
rect 23255 30197 23337 30283
rect 23423 30197 23516 30283
rect 23076 28771 23516 30197
rect 23076 28685 23169 28771
rect 23255 28685 23337 28771
rect 23423 28685 23516 28771
rect 23076 27666 23516 28685
rect 23076 27286 23106 27666
rect 23486 27286 23516 27666
rect 23076 27259 23516 27286
rect 23076 27173 23169 27259
rect 23255 27173 23337 27259
rect 23423 27173 23516 27259
rect 23076 25747 23516 27173
rect 23076 25661 23169 25747
rect 23255 25661 23337 25747
rect 23423 25661 23516 25747
rect 23076 24235 23516 25661
rect 23076 24149 23169 24235
rect 23255 24149 23337 24235
rect 23423 24149 23516 24235
rect 23076 23666 23516 24149
rect 23076 23286 23106 23666
rect 23486 23286 23516 23666
rect 23076 22723 23516 23286
rect 23076 22637 23169 22723
rect 23255 22637 23337 22723
rect 23423 22637 23516 22723
rect 23076 21211 23516 22637
rect 23076 21125 23169 21211
rect 23255 21125 23337 21211
rect 23423 21125 23516 21211
rect 23076 19699 23516 21125
rect 23076 19666 23169 19699
rect 23255 19666 23337 19699
rect 23423 19666 23516 19699
rect 23076 19286 23106 19666
rect 23486 19286 23516 19666
rect 23076 18187 23516 19286
rect 23076 18101 23169 18187
rect 23255 18101 23337 18187
rect 23423 18101 23516 18187
rect 23076 16675 23516 18101
rect 23076 16589 23169 16675
rect 23255 16589 23337 16675
rect 23423 16589 23516 16675
rect 23076 15666 23516 16589
rect 23076 15286 23106 15666
rect 23486 15286 23516 15666
rect 23076 15163 23516 15286
rect 23076 15077 23169 15163
rect 23255 15077 23337 15163
rect 23423 15077 23516 15163
rect 23076 13651 23516 15077
rect 23076 13565 23169 13651
rect 23255 13565 23337 13651
rect 23423 13565 23516 13651
rect 23076 12139 23516 13565
rect 23076 12053 23169 12139
rect 23255 12053 23337 12139
rect 23423 12053 23516 12139
rect 23076 11666 23516 12053
rect 23076 11286 23106 11666
rect 23486 11286 23516 11666
rect 23076 10627 23516 11286
rect 23076 10541 23169 10627
rect 23255 10541 23337 10627
rect 23423 10541 23516 10627
rect 23076 9115 23516 10541
rect 23076 9029 23169 9115
rect 23255 9029 23337 9115
rect 23423 9029 23516 9115
rect 23076 7666 23516 9029
rect 23076 7286 23106 7666
rect 23486 7286 23516 7666
rect 23076 6091 23516 7286
rect 23076 6005 23169 6091
rect 23255 6005 23337 6091
rect 23423 6005 23516 6091
rect 23076 4579 23516 6005
rect 23076 4493 23169 4579
rect 23255 4493 23337 4579
rect 23423 4493 23516 4579
rect 23076 3666 23516 4493
rect 23076 3286 23106 3666
rect 23486 3286 23516 3666
rect 23076 3067 23516 3286
rect 23076 2981 23169 3067
rect 23255 2981 23337 3067
rect 23423 2981 23516 3067
rect 23076 1555 23516 2981
rect 23076 1469 23169 1555
rect 23255 1469 23337 1555
rect 23423 1469 23516 1555
rect 23076 712 23516 1469
rect 24316 38599 24756 38682
rect 24316 38513 24409 38599
rect 24495 38513 24577 38599
rect 24663 38513 24756 38599
rect 24316 37087 24756 38513
rect 24316 37001 24409 37087
rect 24495 37001 24577 37087
rect 24663 37001 24756 37087
rect 24316 36906 24756 37001
rect 24316 36526 24346 36906
rect 24726 36526 24756 36906
rect 24316 35575 24756 36526
rect 24316 35489 24409 35575
rect 24495 35489 24577 35575
rect 24663 35489 24756 35575
rect 24316 34063 24756 35489
rect 24316 33977 24409 34063
rect 24495 33977 24577 34063
rect 24663 33977 24756 34063
rect 24316 32906 24756 33977
rect 24316 32526 24346 32906
rect 24726 32526 24756 32906
rect 24316 32465 24409 32526
rect 24495 32465 24577 32526
rect 24663 32465 24756 32526
rect 24316 31039 24756 32465
rect 24316 30953 24409 31039
rect 24495 30953 24577 31039
rect 24663 30953 24756 31039
rect 24316 29527 24756 30953
rect 24316 29441 24409 29527
rect 24495 29441 24577 29527
rect 24663 29441 24756 29527
rect 24316 28906 24756 29441
rect 24316 28526 24346 28906
rect 24726 28526 24756 28906
rect 24316 28015 24756 28526
rect 24316 27929 24409 28015
rect 24495 27929 24577 28015
rect 24663 27929 24756 28015
rect 24316 26503 24756 27929
rect 24316 26417 24409 26503
rect 24495 26417 24577 26503
rect 24663 26417 24756 26503
rect 24316 24991 24756 26417
rect 24316 24906 24409 24991
rect 24495 24906 24577 24991
rect 24663 24906 24756 24991
rect 24316 24526 24346 24906
rect 24726 24526 24756 24906
rect 24316 23479 24756 24526
rect 24316 23393 24409 23479
rect 24495 23393 24577 23479
rect 24663 23393 24756 23479
rect 24316 21967 24756 23393
rect 24316 21881 24409 21967
rect 24495 21881 24577 21967
rect 24663 21881 24756 21967
rect 24316 20906 24756 21881
rect 24316 20526 24346 20906
rect 24726 20526 24756 20906
rect 24316 20455 24756 20526
rect 24316 20369 24409 20455
rect 24495 20369 24577 20455
rect 24663 20369 24756 20455
rect 24316 18943 24756 20369
rect 24316 18857 24409 18943
rect 24495 18857 24577 18943
rect 24663 18857 24756 18943
rect 24316 17431 24756 18857
rect 24316 17345 24409 17431
rect 24495 17345 24577 17431
rect 24663 17345 24756 17431
rect 24316 16906 24756 17345
rect 24316 16526 24346 16906
rect 24726 16526 24756 16906
rect 24316 15919 24756 16526
rect 24316 15833 24409 15919
rect 24495 15833 24577 15919
rect 24663 15833 24756 15919
rect 24316 14407 24756 15833
rect 24316 14321 24409 14407
rect 24495 14321 24577 14407
rect 24663 14321 24756 14407
rect 24316 12906 24756 14321
rect 24316 12526 24346 12906
rect 24726 12526 24756 12906
rect 24316 11383 24756 12526
rect 24316 11297 24409 11383
rect 24495 11297 24577 11383
rect 24663 11297 24756 11383
rect 24316 9871 24756 11297
rect 24316 9785 24409 9871
rect 24495 9785 24577 9871
rect 24663 9785 24756 9871
rect 24316 8906 24756 9785
rect 24316 8526 24346 8906
rect 24726 8526 24756 8906
rect 24316 8359 24756 8526
rect 24316 8273 24409 8359
rect 24495 8273 24577 8359
rect 24663 8273 24756 8359
rect 24316 6847 24756 8273
rect 24316 6761 24409 6847
rect 24495 6761 24577 6847
rect 24663 6761 24756 6847
rect 24316 5335 24756 6761
rect 24316 5249 24409 5335
rect 24495 5249 24577 5335
rect 24663 5249 24756 5335
rect 24316 4906 24756 5249
rect 24316 4526 24346 4906
rect 24726 4526 24756 4906
rect 24316 3823 24756 4526
rect 24316 3737 24409 3823
rect 24495 3737 24577 3823
rect 24663 3737 24756 3823
rect 24316 2311 24756 3737
rect 24316 2225 24409 2311
rect 24495 2225 24577 2311
rect 24663 2225 24756 2311
rect 24316 799 24756 2225
rect 24316 713 24409 799
rect 24495 713 24577 799
rect 24663 713 24756 799
rect 24316 630 24756 713
rect 27076 37843 27516 38600
rect 27076 37757 27169 37843
rect 27255 37757 27337 37843
rect 27423 37757 27516 37843
rect 27076 36331 27516 37757
rect 27076 36245 27169 36331
rect 27255 36245 27337 36331
rect 27423 36245 27516 36331
rect 27076 35666 27516 36245
rect 27076 35286 27106 35666
rect 27486 35286 27516 35666
rect 27076 34819 27516 35286
rect 27076 34733 27169 34819
rect 27255 34733 27337 34819
rect 27423 34733 27516 34819
rect 27076 33307 27516 34733
rect 27076 33221 27169 33307
rect 27255 33221 27337 33307
rect 27423 33221 27516 33307
rect 27076 31795 27516 33221
rect 27076 31709 27169 31795
rect 27255 31709 27337 31795
rect 27423 31709 27516 31795
rect 27076 31666 27516 31709
rect 27076 31286 27106 31666
rect 27486 31286 27516 31666
rect 27076 30283 27516 31286
rect 27076 30197 27169 30283
rect 27255 30197 27337 30283
rect 27423 30197 27516 30283
rect 27076 28771 27516 30197
rect 27076 28685 27169 28771
rect 27255 28685 27337 28771
rect 27423 28685 27516 28771
rect 27076 27666 27516 28685
rect 27076 27286 27106 27666
rect 27486 27286 27516 27666
rect 27076 27259 27516 27286
rect 27076 27173 27169 27259
rect 27255 27173 27337 27259
rect 27423 27173 27516 27259
rect 27076 25747 27516 27173
rect 27076 25661 27169 25747
rect 27255 25661 27337 25747
rect 27423 25661 27516 25747
rect 27076 24235 27516 25661
rect 27076 24149 27169 24235
rect 27255 24149 27337 24235
rect 27423 24149 27516 24235
rect 27076 23666 27516 24149
rect 27076 23286 27106 23666
rect 27486 23286 27516 23666
rect 27076 22723 27516 23286
rect 27076 22637 27169 22723
rect 27255 22637 27337 22723
rect 27423 22637 27516 22723
rect 27076 21211 27516 22637
rect 27076 21125 27169 21211
rect 27255 21125 27337 21211
rect 27423 21125 27516 21211
rect 27076 19699 27516 21125
rect 27076 19666 27169 19699
rect 27255 19666 27337 19699
rect 27423 19666 27516 19699
rect 27076 19286 27106 19666
rect 27486 19286 27516 19666
rect 27076 18187 27516 19286
rect 27076 18101 27169 18187
rect 27255 18101 27337 18187
rect 27423 18101 27516 18187
rect 27076 16675 27516 18101
rect 27076 16589 27169 16675
rect 27255 16589 27337 16675
rect 27423 16589 27516 16675
rect 27076 15666 27516 16589
rect 27076 15286 27106 15666
rect 27486 15286 27516 15666
rect 27076 15163 27516 15286
rect 27076 15077 27169 15163
rect 27255 15077 27337 15163
rect 27423 15077 27516 15163
rect 27076 13651 27516 15077
rect 27076 13565 27169 13651
rect 27255 13565 27337 13651
rect 27423 13565 27516 13651
rect 27076 12139 27516 13565
rect 27076 12053 27169 12139
rect 27255 12053 27337 12139
rect 27423 12053 27516 12139
rect 27076 11666 27516 12053
rect 27076 11286 27106 11666
rect 27486 11286 27516 11666
rect 27076 10627 27516 11286
rect 27076 10541 27169 10627
rect 27255 10541 27337 10627
rect 27423 10541 27516 10627
rect 27076 9115 27516 10541
rect 27076 9029 27169 9115
rect 27255 9029 27337 9115
rect 27423 9029 27516 9115
rect 27076 7666 27516 9029
rect 27076 7286 27106 7666
rect 27486 7286 27516 7666
rect 27076 6091 27516 7286
rect 27076 6005 27169 6091
rect 27255 6005 27337 6091
rect 27423 6005 27516 6091
rect 27076 4579 27516 6005
rect 27076 4493 27169 4579
rect 27255 4493 27337 4579
rect 27423 4493 27516 4579
rect 27076 3666 27516 4493
rect 27076 3286 27106 3666
rect 27486 3286 27516 3666
rect 27076 3067 27516 3286
rect 27076 2981 27169 3067
rect 27255 2981 27337 3067
rect 27423 2981 27516 3067
rect 27076 1555 27516 2981
rect 27076 1469 27169 1555
rect 27255 1469 27337 1555
rect 27423 1469 27516 1555
rect 27076 712 27516 1469
rect 28316 38599 28756 38682
rect 28316 38513 28409 38599
rect 28495 38513 28577 38599
rect 28663 38513 28756 38599
rect 28316 37087 28756 38513
rect 28316 37001 28409 37087
rect 28495 37001 28577 37087
rect 28663 37001 28756 37087
rect 28316 36906 28756 37001
rect 28316 36526 28346 36906
rect 28726 36526 28756 36906
rect 28316 35575 28756 36526
rect 28316 35489 28409 35575
rect 28495 35489 28577 35575
rect 28663 35489 28756 35575
rect 28316 34063 28756 35489
rect 28316 33977 28409 34063
rect 28495 33977 28577 34063
rect 28663 33977 28756 34063
rect 28316 32906 28756 33977
rect 28316 32526 28346 32906
rect 28726 32526 28756 32906
rect 28316 32465 28409 32526
rect 28495 32465 28577 32526
rect 28663 32465 28756 32526
rect 28316 31039 28756 32465
rect 28316 30953 28409 31039
rect 28495 30953 28577 31039
rect 28663 30953 28756 31039
rect 28316 29527 28756 30953
rect 28316 29441 28409 29527
rect 28495 29441 28577 29527
rect 28663 29441 28756 29527
rect 28316 28906 28756 29441
rect 28316 28526 28346 28906
rect 28726 28526 28756 28906
rect 28316 28015 28756 28526
rect 28316 27929 28409 28015
rect 28495 27929 28577 28015
rect 28663 27929 28756 28015
rect 28316 26503 28756 27929
rect 28316 26417 28409 26503
rect 28495 26417 28577 26503
rect 28663 26417 28756 26503
rect 28316 24991 28756 26417
rect 28316 24906 28409 24991
rect 28495 24906 28577 24991
rect 28663 24906 28756 24991
rect 28316 24526 28346 24906
rect 28726 24526 28756 24906
rect 28316 23479 28756 24526
rect 28316 23393 28409 23479
rect 28495 23393 28577 23479
rect 28663 23393 28756 23479
rect 28316 21967 28756 23393
rect 28316 21881 28409 21967
rect 28495 21881 28577 21967
rect 28663 21881 28756 21967
rect 28316 20906 28756 21881
rect 28316 20526 28346 20906
rect 28726 20526 28756 20906
rect 28316 20455 28756 20526
rect 28316 20369 28409 20455
rect 28495 20369 28577 20455
rect 28663 20369 28756 20455
rect 28316 18943 28756 20369
rect 28316 18857 28409 18943
rect 28495 18857 28577 18943
rect 28663 18857 28756 18943
rect 28316 17431 28756 18857
rect 28316 17345 28409 17431
rect 28495 17345 28577 17431
rect 28663 17345 28756 17431
rect 28316 16906 28756 17345
rect 28316 16526 28346 16906
rect 28726 16526 28756 16906
rect 28316 15919 28756 16526
rect 28316 15833 28409 15919
rect 28495 15833 28577 15919
rect 28663 15833 28756 15919
rect 28316 14407 28756 15833
rect 28316 14321 28409 14407
rect 28495 14321 28577 14407
rect 28663 14321 28756 14407
rect 28316 12906 28756 14321
rect 28316 12526 28346 12906
rect 28726 12526 28756 12906
rect 28316 11383 28756 12526
rect 28316 11297 28409 11383
rect 28495 11297 28577 11383
rect 28663 11297 28756 11383
rect 28316 9871 28756 11297
rect 28316 9785 28409 9871
rect 28495 9785 28577 9871
rect 28663 9785 28756 9871
rect 28316 8906 28756 9785
rect 28316 8526 28346 8906
rect 28726 8526 28756 8906
rect 28316 8359 28756 8526
rect 28316 8273 28409 8359
rect 28495 8273 28577 8359
rect 28663 8273 28756 8359
rect 28316 6847 28756 8273
rect 28316 6761 28409 6847
rect 28495 6761 28577 6847
rect 28663 6761 28756 6847
rect 28316 5335 28756 6761
rect 28316 5249 28409 5335
rect 28495 5249 28577 5335
rect 28663 5249 28756 5335
rect 28316 4906 28756 5249
rect 28316 4526 28346 4906
rect 28726 4526 28756 4906
rect 28316 3823 28756 4526
rect 28316 3737 28409 3823
rect 28495 3737 28577 3823
rect 28663 3737 28756 3823
rect 28316 2311 28756 3737
rect 28316 2225 28409 2311
rect 28495 2225 28577 2311
rect 28663 2225 28756 2311
rect 28316 799 28756 2225
rect 28316 713 28409 799
rect 28495 713 28577 799
rect 28663 713 28756 799
rect 28316 630 28756 713
rect 31076 37843 31516 38600
rect 31076 37757 31169 37843
rect 31255 37757 31337 37843
rect 31423 37757 31516 37843
rect 31076 36331 31516 37757
rect 31076 36245 31169 36331
rect 31255 36245 31337 36331
rect 31423 36245 31516 36331
rect 31076 35666 31516 36245
rect 31076 35286 31106 35666
rect 31486 35286 31516 35666
rect 31076 34819 31516 35286
rect 31076 34733 31169 34819
rect 31255 34733 31337 34819
rect 31423 34733 31516 34819
rect 31076 33307 31516 34733
rect 31076 33221 31169 33307
rect 31255 33221 31337 33307
rect 31423 33221 31516 33307
rect 31076 31795 31516 33221
rect 31076 31709 31169 31795
rect 31255 31709 31337 31795
rect 31423 31709 31516 31795
rect 31076 31666 31516 31709
rect 31076 31286 31106 31666
rect 31486 31286 31516 31666
rect 31076 30283 31516 31286
rect 31076 30197 31169 30283
rect 31255 30197 31337 30283
rect 31423 30197 31516 30283
rect 31076 28771 31516 30197
rect 31076 28685 31169 28771
rect 31255 28685 31337 28771
rect 31423 28685 31516 28771
rect 31076 27666 31516 28685
rect 31076 27286 31106 27666
rect 31486 27286 31516 27666
rect 31076 27259 31516 27286
rect 31076 27173 31169 27259
rect 31255 27173 31337 27259
rect 31423 27173 31516 27259
rect 31076 25747 31516 27173
rect 31076 25661 31169 25747
rect 31255 25661 31337 25747
rect 31423 25661 31516 25747
rect 31076 24235 31516 25661
rect 31076 24149 31169 24235
rect 31255 24149 31337 24235
rect 31423 24149 31516 24235
rect 31076 23666 31516 24149
rect 31076 23286 31106 23666
rect 31486 23286 31516 23666
rect 31076 22723 31516 23286
rect 31076 22637 31169 22723
rect 31255 22637 31337 22723
rect 31423 22637 31516 22723
rect 31076 21211 31516 22637
rect 31076 21125 31169 21211
rect 31255 21125 31337 21211
rect 31423 21125 31516 21211
rect 31076 19699 31516 21125
rect 31076 19666 31169 19699
rect 31255 19666 31337 19699
rect 31423 19666 31516 19699
rect 31076 19286 31106 19666
rect 31486 19286 31516 19666
rect 31076 18187 31516 19286
rect 31076 18101 31169 18187
rect 31255 18101 31337 18187
rect 31423 18101 31516 18187
rect 31076 16675 31516 18101
rect 31076 16589 31169 16675
rect 31255 16589 31337 16675
rect 31423 16589 31516 16675
rect 31076 15666 31516 16589
rect 31076 15286 31106 15666
rect 31486 15286 31516 15666
rect 31076 15163 31516 15286
rect 31076 15077 31169 15163
rect 31255 15077 31337 15163
rect 31423 15077 31516 15163
rect 31076 13651 31516 15077
rect 31076 13565 31169 13651
rect 31255 13565 31337 13651
rect 31423 13565 31516 13651
rect 31076 12139 31516 13565
rect 31076 12053 31169 12139
rect 31255 12053 31337 12139
rect 31423 12053 31516 12139
rect 31076 11666 31516 12053
rect 31076 11286 31106 11666
rect 31486 11286 31516 11666
rect 31076 10627 31516 11286
rect 31076 10541 31169 10627
rect 31255 10541 31337 10627
rect 31423 10541 31516 10627
rect 31076 9115 31516 10541
rect 31076 9029 31169 9115
rect 31255 9029 31337 9115
rect 31423 9029 31516 9115
rect 31076 7666 31516 9029
rect 31076 7286 31106 7666
rect 31486 7286 31516 7666
rect 31076 6091 31516 7286
rect 31076 6005 31169 6091
rect 31255 6005 31337 6091
rect 31423 6005 31516 6091
rect 31076 4579 31516 6005
rect 31076 4493 31169 4579
rect 31255 4493 31337 4579
rect 31423 4493 31516 4579
rect 31076 3666 31516 4493
rect 31076 3286 31106 3666
rect 31486 3286 31516 3666
rect 31076 3067 31516 3286
rect 31076 2981 31169 3067
rect 31255 2981 31337 3067
rect 31423 2981 31516 3067
rect 31076 1555 31516 2981
rect 31076 1469 31169 1555
rect 31255 1469 31337 1555
rect 31423 1469 31516 1555
rect 31076 712 31516 1469
rect 32316 38599 32756 38682
rect 32316 38513 32409 38599
rect 32495 38513 32577 38599
rect 32663 38513 32756 38599
rect 32316 37087 32756 38513
rect 32316 37001 32409 37087
rect 32495 37001 32577 37087
rect 32663 37001 32756 37087
rect 32316 36906 32756 37001
rect 32316 36526 32346 36906
rect 32726 36526 32756 36906
rect 32316 35575 32756 36526
rect 32316 35489 32409 35575
rect 32495 35489 32577 35575
rect 32663 35489 32756 35575
rect 32316 34063 32756 35489
rect 32316 33977 32409 34063
rect 32495 33977 32577 34063
rect 32663 33977 32756 34063
rect 32316 32906 32756 33977
rect 32316 32526 32346 32906
rect 32726 32526 32756 32906
rect 32316 32465 32409 32526
rect 32495 32465 32577 32526
rect 32663 32465 32756 32526
rect 32316 31039 32756 32465
rect 32316 30953 32409 31039
rect 32495 30953 32577 31039
rect 32663 30953 32756 31039
rect 32316 29527 32756 30953
rect 32316 29441 32409 29527
rect 32495 29441 32577 29527
rect 32663 29441 32756 29527
rect 32316 28906 32756 29441
rect 32316 28526 32346 28906
rect 32726 28526 32756 28906
rect 32316 28015 32756 28526
rect 32316 27929 32409 28015
rect 32495 27929 32577 28015
rect 32663 27929 32756 28015
rect 32316 26503 32756 27929
rect 32316 26417 32409 26503
rect 32495 26417 32577 26503
rect 32663 26417 32756 26503
rect 32316 24991 32756 26417
rect 32316 24906 32409 24991
rect 32495 24906 32577 24991
rect 32663 24906 32756 24991
rect 32316 24526 32346 24906
rect 32726 24526 32756 24906
rect 32316 23479 32756 24526
rect 32316 23393 32409 23479
rect 32495 23393 32577 23479
rect 32663 23393 32756 23479
rect 32316 21967 32756 23393
rect 32316 21881 32409 21967
rect 32495 21881 32577 21967
rect 32663 21881 32756 21967
rect 32316 20906 32756 21881
rect 32316 20526 32346 20906
rect 32726 20526 32756 20906
rect 32316 20455 32756 20526
rect 32316 20369 32409 20455
rect 32495 20369 32577 20455
rect 32663 20369 32756 20455
rect 32316 18943 32756 20369
rect 32316 18857 32409 18943
rect 32495 18857 32577 18943
rect 32663 18857 32756 18943
rect 32316 17431 32756 18857
rect 32316 17345 32409 17431
rect 32495 17345 32577 17431
rect 32663 17345 32756 17431
rect 32316 16906 32756 17345
rect 32316 16526 32346 16906
rect 32726 16526 32756 16906
rect 32316 15919 32756 16526
rect 32316 15833 32409 15919
rect 32495 15833 32577 15919
rect 32663 15833 32756 15919
rect 32316 14407 32756 15833
rect 32316 14321 32409 14407
rect 32495 14321 32577 14407
rect 32663 14321 32756 14407
rect 32316 12906 32756 14321
rect 32316 12526 32346 12906
rect 32726 12526 32756 12906
rect 32316 11383 32756 12526
rect 32316 11297 32409 11383
rect 32495 11297 32577 11383
rect 32663 11297 32756 11383
rect 32316 9871 32756 11297
rect 32316 9785 32409 9871
rect 32495 9785 32577 9871
rect 32663 9785 32756 9871
rect 32316 8906 32756 9785
rect 32316 8526 32346 8906
rect 32726 8526 32756 8906
rect 32316 8359 32756 8526
rect 32316 8273 32409 8359
rect 32495 8273 32577 8359
rect 32663 8273 32756 8359
rect 32316 6847 32756 8273
rect 32316 6761 32409 6847
rect 32495 6761 32577 6847
rect 32663 6761 32756 6847
rect 32316 5335 32756 6761
rect 32316 5249 32409 5335
rect 32495 5249 32577 5335
rect 32663 5249 32756 5335
rect 32316 4906 32756 5249
rect 32316 4526 32346 4906
rect 32726 4526 32756 4906
rect 32316 3823 32756 4526
rect 32316 3737 32409 3823
rect 32495 3737 32577 3823
rect 32663 3737 32756 3823
rect 32316 2311 32756 3737
rect 32316 2225 32409 2311
rect 32495 2225 32577 2311
rect 32663 2225 32756 2311
rect 32316 799 32756 2225
rect 32316 713 32409 799
rect 32495 713 32577 799
rect 32663 713 32756 799
rect 32316 630 32756 713
rect 35076 37843 35516 38600
rect 35076 37757 35169 37843
rect 35255 37757 35337 37843
rect 35423 37757 35516 37843
rect 35076 36331 35516 37757
rect 35076 36245 35169 36331
rect 35255 36245 35337 36331
rect 35423 36245 35516 36331
rect 35076 35666 35516 36245
rect 35076 35286 35106 35666
rect 35486 35286 35516 35666
rect 35076 34819 35516 35286
rect 35076 34733 35169 34819
rect 35255 34733 35337 34819
rect 35423 34733 35516 34819
rect 35076 33307 35516 34733
rect 35076 33221 35169 33307
rect 35255 33221 35337 33307
rect 35423 33221 35516 33307
rect 35076 31795 35516 33221
rect 35076 31709 35169 31795
rect 35255 31709 35337 31795
rect 35423 31709 35516 31795
rect 35076 31666 35516 31709
rect 35076 31286 35106 31666
rect 35486 31286 35516 31666
rect 35076 30283 35516 31286
rect 35076 30197 35169 30283
rect 35255 30197 35337 30283
rect 35423 30197 35516 30283
rect 35076 28771 35516 30197
rect 35076 28685 35169 28771
rect 35255 28685 35337 28771
rect 35423 28685 35516 28771
rect 35076 27666 35516 28685
rect 35076 27286 35106 27666
rect 35486 27286 35516 27666
rect 35076 27259 35516 27286
rect 35076 27173 35169 27259
rect 35255 27173 35337 27259
rect 35423 27173 35516 27259
rect 35076 25747 35516 27173
rect 35076 25661 35169 25747
rect 35255 25661 35337 25747
rect 35423 25661 35516 25747
rect 35076 24235 35516 25661
rect 35076 24149 35169 24235
rect 35255 24149 35337 24235
rect 35423 24149 35516 24235
rect 35076 23666 35516 24149
rect 35076 23286 35106 23666
rect 35486 23286 35516 23666
rect 35076 22723 35516 23286
rect 35076 22637 35169 22723
rect 35255 22637 35337 22723
rect 35423 22637 35516 22723
rect 35076 21211 35516 22637
rect 35076 21125 35169 21211
rect 35255 21125 35337 21211
rect 35423 21125 35516 21211
rect 35076 19699 35516 21125
rect 35076 19666 35169 19699
rect 35255 19666 35337 19699
rect 35423 19666 35516 19699
rect 35076 19286 35106 19666
rect 35486 19286 35516 19666
rect 35076 18187 35516 19286
rect 35076 18101 35169 18187
rect 35255 18101 35337 18187
rect 35423 18101 35516 18187
rect 35076 16675 35516 18101
rect 35076 16589 35169 16675
rect 35255 16589 35337 16675
rect 35423 16589 35516 16675
rect 35076 15666 35516 16589
rect 35076 15286 35106 15666
rect 35486 15286 35516 15666
rect 35076 15163 35516 15286
rect 35076 15077 35169 15163
rect 35255 15077 35337 15163
rect 35423 15077 35516 15163
rect 35076 13651 35516 15077
rect 35076 13565 35169 13651
rect 35255 13565 35337 13651
rect 35423 13565 35516 13651
rect 35076 12139 35516 13565
rect 35076 12053 35169 12139
rect 35255 12053 35337 12139
rect 35423 12053 35516 12139
rect 35076 11666 35516 12053
rect 35076 11286 35106 11666
rect 35486 11286 35516 11666
rect 35076 10627 35516 11286
rect 35076 10541 35169 10627
rect 35255 10541 35337 10627
rect 35423 10541 35516 10627
rect 35076 9115 35516 10541
rect 35076 9029 35169 9115
rect 35255 9029 35337 9115
rect 35423 9029 35516 9115
rect 35076 7666 35516 9029
rect 35076 7286 35106 7666
rect 35486 7286 35516 7666
rect 35076 6091 35516 7286
rect 35076 6005 35169 6091
rect 35255 6005 35337 6091
rect 35423 6005 35516 6091
rect 35076 4579 35516 6005
rect 35076 4493 35169 4579
rect 35255 4493 35337 4579
rect 35423 4493 35516 4579
rect 35076 3666 35516 4493
rect 35076 3286 35106 3666
rect 35486 3286 35516 3666
rect 35076 3067 35516 3286
rect 35076 2981 35169 3067
rect 35255 2981 35337 3067
rect 35423 2981 35516 3067
rect 35076 1555 35516 2981
rect 35076 1469 35169 1555
rect 35255 1469 35337 1555
rect 35423 1469 35516 1555
rect 35076 712 35516 1469
rect 36316 38599 36756 38682
rect 36316 38513 36409 38599
rect 36495 38513 36577 38599
rect 36663 38513 36756 38599
rect 36316 37087 36756 38513
rect 36316 37001 36409 37087
rect 36495 37001 36577 37087
rect 36663 37001 36756 37087
rect 36316 36906 36756 37001
rect 36316 36526 36346 36906
rect 36726 36526 36756 36906
rect 36316 35575 36756 36526
rect 36316 35489 36409 35575
rect 36495 35489 36577 35575
rect 36663 35489 36756 35575
rect 36316 34063 36756 35489
rect 36316 33977 36409 34063
rect 36495 33977 36577 34063
rect 36663 33977 36756 34063
rect 36316 32906 36756 33977
rect 36316 32526 36346 32906
rect 36726 32526 36756 32906
rect 36316 32465 36409 32526
rect 36495 32465 36577 32526
rect 36663 32465 36756 32526
rect 36316 31039 36756 32465
rect 36316 30953 36409 31039
rect 36495 30953 36577 31039
rect 36663 30953 36756 31039
rect 36316 29527 36756 30953
rect 36316 29441 36409 29527
rect 36495 29441 36577 29527
rect 36663 29441 36756 29527
rect 36316 28906 36756 29441
rect 36316 28526 36346 28906
rect 36726 28526 36756 28906
rect 36316 28015 36756 28526
rect 36316 27929 36409 28015
rect 36495 27929 36577 28015
rect 36663 27929 36756 28015
rect 36316 26503 36756 27929
rect 36316 26417 36409 26503
rect 36495 26417 36577 26503
rect 36663 26417 36756 26503
rect 36316 24991 36756 26417
rect 36316 24906 36409 24991
rect 36495 24906 36577 24991
rect 36663 24906 36756 24991
rect 36316 24526 36346 24906
rect 36726 24526 36756 24906
rect 36316 23479 36756 24526
rect 36316 23393 36409 23479
rect 36495 23393 36577 23479
rect 36663 23393 36756 23479
rect 36316 21967 36756 23393
rect 36316 21881 36409 21967
rect 36495 21881 36577 21967
rect 36663 21881 36756 21967
rect 36316 20906 36756 21881
rect 36316 20526 36346 20906
rect 36726 20526 36756 20906
rect 36316 20455 36756 20526
rect 36316 20369 36409 20455
rect 36495 20369 36577 20455
rect 36663 20369 36756 20455
rect 36316 18943 36756 20369
rect 36316 18857 36409 18943
rect 36495 18857 36577 18943
rect 36663 18857 36756 18943
rect 36316 17431 36756 18857
rect 36316 17345 36409 17431
rect 36495 17345 36577 17431
rect 36663 17345 36756 17431
rect 36316 16906 36756 17345
rect 36316 16526 36346 16906
rect 36726 16526 36756 16906
rect 36316 15919 36756 16526
rect 36316 15833 36409 15919
rect 36495 15833 36577 15919
rect 36663 15833 36756 15919
rect 36316 14407 36756 15833
rect 36316 14321 36409 14407
rect 36495 14321 36577 14407
rect 36663 14321 36756 14407
rect 36316 12906 36756 14321
rect 36316 12526 36346 12906
rect 36726 12526 36756 12906
rect 36316 11383 36756 12526
rect 36316 11297 36409 11383
rect 36495 11297 36577 11383
rect 36663 11297 36756 11383
rect 36316 9871 36756 11297
rect 36316 9785 36409 9871
rect 36495 9785 36577 9871
rect 36663 9785 36756 9871
rect 36316 8906 36756 9785
rect 36316 8526 36346 8906
rect 36726 8526 36756 8906
rect 36316 8359 36756 8526
rect 36316 8273 36409 8359
rect 36495 8273 36577 8359
rect 36663 8273 36756 8359
rect 36316 6847 36756 8273
rect 36316 6761 36409 6847
rect 36495 6761 36577 6847
rect 36663 6761 36756 6847
rect 36316 5335 36756 6761
rect 36316 5249 36409 5335
rect 36495 5249 36577 5335
rect 36663 5249 36756 5335
rect 36316 4906 36756 5249
rect 36316 4526 36346 4906
rect 36726 4526 36756 4906
rect 36316 3823 36756 4526
rect 36316 3737 36409 3823
rect 36495 3737 36577 3823
rect 36663 3737 36756 3823
rect 36316 2311 36756 3737
rect 36316 2225 36409 2311
rect 36495 2225 36577 2311
rect 36663 2225 36756 2311
rect 36316 799 36756 2225
rect 36316 713 36409 799
rect 36495 713 36577 799
rect 36663 713 36756 799
rect 36316 630 36756 713
rect 39076 37843 39516 38600
rect 39076 37757 39169 37843
rect 39255 37757 39337 37843
rect 39423 37757 39516 37843
rect 39076 36331 39516 37757
rect 39076 36245 39169 36331
rect 39255 36245 39337 36331
rect 39423 36245 39516 36331
rect 39076 35666 39516 36245
rect 39076 35286 39106 35666
rect 39486 35286 39516 35666
rect 39076 34819 39516 35286
rect 39076 34733 39169 34819
rect 39255 34733 39337 34819
rect 39423 34733 39516 34819
rect 39076 33307 39516 34733
rect 39076 33221 39169 33307
rect 39255 33221 39337 33307
rect 39423 33221 39516 33307
rect 39076 31795 39516 33221
rect 39076 31709 39169 31795
rect 39255 31709 39337 31795
rect 39423 31709 39516 31795
rect 39076 31666 39516 31709
rect 39076 31286 39106 31666
rect 39486 31286 39516 31666
rect 39076 30283 39516 31286
rect 39076 30197 39169 30283
rect 39255 30197 39337 30283
rect 39423 30197 39516 30283
rect 39076 28771 39516 30197
rect 39076 28685 39169 28771
rect 39255 28685 39337 28771
rect 39423 28685 39516 28771
rect 39076 27666 39516 28685
rect 39076 27286 39106 27666
rect 39486 27286 39516 27666
rect 39076 27259 39516 27286
rect 39076 27173 39169 27259
rect 39255 27173 39337 27259
rect 39423 27173 39516 27259
rect 39076 25747 39516 27173
rect 39076 25661 39169 25747
rect 39255 25661 39337 25747
rect 39423 25661 39516 25747
rect 39076 24235 39516 25661
rect 39076 24149 39169 24235
rect 39255 24149 39337 24235
rect 39423 24149 39516 24235
rect 39076 23666 39516 24149
rect 39076 23286 39106 23666
rect 39486 23286 39516 23666
rect 39076 22723 39516 23286
rect 39076 22637 39169 22723
rect 39255 22637 39337 22723
rect 39423 22637 39516 22723
rect 39076 21211 39516 22637
rect 39076 21125 39169 21211
rect 39255 21125 39337 21211
rect 39423 21125 39516 21211
rect 39076 19699 39516 21125
rect 39076 19666 39169 19699
rect 39255 19666 39337 19699
rect 39423 19666 39516 19699
rect 39076 19286 39106 19666
rect 39486 19286 39516 19666
rect 39076 18187 39516 19286
rect 39076 18101 39169 18187
rect 39255 18101 39337 18187
rect 39423 18101 39516 18187
rect 39076 16675 39516 18101
rect 39076 16589 39169 16675
rect 39255 16589 39337 16675
rect 39423 16589 39516 16675
rect 39076 15666 39516 16589
rect 39076 15286 39106 15666
rect 39486 15286 39516 15666
rect 39076 15163 39516 15286
rect 39076 15077 39169 15163
rect 39255 15077 39337 15163
rect 39423 15077 39516 15163
rect 39076 13651 39516 15077
rect 39076 13565 39169 13651
rect 39255 13565 39337 13651
rect 39423 13565 39516 13651
rect 39076 12139 39516 13565
rect 39076 12053 39169 12139
rect 39255 12053 39337 12139
rect 39423 12053 39516 12139
rect 39076 11666 39516 12053
rect 39076 11286 39106 11666
rect 39486 11286 39516 11666
rect 39076 10627 39516 11286
rect 39076 10541 39169 10627
rect 39255 10541 39337 10627
rect 39423 10541 39516 10627
rect 39076 9115 39516 10541
rect 39076 9029 39169 9115
rect 39255 9029 39337 9115
rect 39423 9029 39516 9115
rect 39076 7666 39516 9029
rect 39076 7286 39106 7666
rect 39486 7286 39516 7666
rect 39076 6091 39516 7286
rect 39076 6005 39169 6091
rect 39255 6005 39337 6091
rect 39423 6005 39516 6091
rect 39076 4579 39516 6005
rect 39076 4493 39169 4579
rect 39255 4493 39337 4579
rect 39423 4493 39516 4579
rect 39076 3666 39516 4493
rect 39076 3286 39106 3666
rect 39486 3286 39516 3666
rect 39076 3067 39516 3286
rect 39076 2981 39169 3067
rect 39255 2981 39337 3067
rect 39423 2981 39516 3067
rect 39076 1555 39516 2981
rect 39076 1469 39169 1555
rect 39255 1469 39337 1555
rect 39423 1469 39516 1555
rect 39076 712 39516 1469
rect 40316 38599 40756 38682
rect 40316 38513 40409 38599
rect 40495 38513 40577 38599
rect 40663 38513 40756 38599
rect 40316 37087 40756 38513
rect 40316 37001 40409 37087
rect 40495 37001 40577 37087
rect 40663 37001 40756 37087
rect 40316 36906 40756 37001
rect 40316 36526 40346 36906
rect 40726 36526 40756 36906
rect 40316 35575 40756 36526
rect 40316 35489 40409 35575
rect 40495 35489 40577 35575
rect 40663 35489 40756 35575
rect 40316 34063 40756 35489
rect 40316 33977 40409 34063
rect 40495 33977 40577 34063
rect 40663 33977 40756 34063
rect 40316 32906 40756 33977
rect 40316 32526 40346 32906
rect 40726 32526 40756 32906
rect 40316 32465 40409 32526
rect 40495 32465 40577 32526
rect 40663 32465 40756 32526
rect 40316 31039 40756 32465
rect 40316 30953 40409 31039
rect 40495 30953 40577 31039
rect 40663 30953 40756 31039
rect 40316 29527 40756 30953
rect 40316 29441 40409 29527
rect 40495 29441 40577 29527
rect 40663 29441 40756 29527
rect 40316 28906 40756 29441
rect 40316 28526 40346 28906
rect 40726 28526 40756 28906
rect 40316 28015 40756 28526
rect 40316 27929 40409 28015
rect 40495 27929 40577 28015
rect 40663 27929 40756 28015
rect 40316 26503 40756 27929
rect 40316 26417 40409 26503
rect 40495 26417 40577 26503
rect 40663 26417 40756 26503
rect 40316 24991 40756 26417
rect 40316 24906 40409 24991
rect 40495 24906 40577 24991
rect 40663 24906 40756 24991
rect 40316 24526 40346 24906
rect 40726 24526 40756 24906
rect 40316 23479 40756 24526
rect 40316 23393 40409 23479
rect 40495 23393 40577 23479
rect 40663 23393 40756 23479
rect 40316 21967 40756 23393
rect 40316 21881 40409 21967
rect 40495 21881 40577 21967
rect 40663 21881 40756 21967
rect 40316 20906 40756 21881
rect 40316 20526 40346 20906
rect 40726 20526 40756 20906
rect 40316 20455 40756 20526
rect 40316 20369 40409 20455
rect 40495 20369 40577 20455
rect 40663 20369 40756 20455
rect 40316 18943 40756 20369
rect 40316 18857 40409 18943
rect 40495 18857 40577 18943
rect 40663 18857 40756 18943
rect 40316 17431 40756 18857
rect 40316 17345 40409 17431
rect 40495 17345 40577 17431
rect 40663 17345 40756 17431
rect 40316 16906 40756 17345
rect 40316 16526 40346 16906
rect 40726 16526 40756 16906
rect 40316 15919 40756 16526
rect 40316 15833 40409 15919
rect 40495 15833 40577 15919
rect 40663 15833 40756 15919
rect 40316 14407 40756 15833
rect 40316 14321 40409 14407
rect 40495 14321 40577 14407
rect 40663 14321 40756 14407
rect 40316 12906 40756 14321
rect 40316 12526 40346 12906
rect 40726 12526 40756 12906
rect 40316 11383 40756 12526
rect 40316 11297 40409 11383
rect 40495 11297 40577 11383
rect 40663 11297 40756 11383
rect 40316 9871 40756 11297
rect 40316 9785 40409 9871
rect 40495 9785 40577 9871
rect 40663 9785 40756 9871
rect 40316 8906 40756 9785
rect 40316 8526 40346 8906
rect 40726 8526 40756 8906
rect 40316 8359 40756 8526
rect 40316 8273 40409 8359
rect 40495 8273 40577 8359
rect 40663 8273 40756 8359
rect 40316 6847 40756 8273
rect 40316 6761 40409 6847
rect 40495 6761 40577 6847
rect 40663 6761 40756 6847
rect 40316 5335 40756 6761
rect 40316 5249 40409 5335
rect 40495 5249 40577 5335
rect 40663 5249 40756 5335
rect 40316 4906 40756 5249
rect 40316 4526 40346 4906
rect 40726 4526 40756 4906
rect 40316 3823 40756 4526
rect 40316 3737 40409 3823
rect 40495 3737 40577 3823
rect 40663 3737 40756 3823
rect 40316 2311 40756 3737
rect 40316 2225 40409 2311
rect 40495 2225 40577 2311
rect 40663 2225 40756 2311
rect 40316 799 40756 2225
rect 40316 713 40409 799
rect 40495 713 40577 799
rect 40663 713 40756 799
rect 40316 630 40756 713
rect 43076 37843 43516 38600
rect 43076 37757 43169 37843
rect 43255 37757 43337 37843
rect 43423 37757 43516 37843
rect 43076 36331 43516 37757
rect 43076 36245 43169 36331
rect 43255 36245 43337 36331
rect 43423 36245 43516 36331
rect 43076 35666 43516 36245
rect 43076 35286 43106 35666
rect 43486 35286 43516 35666
rect 43076 34819 43516 35286
rect 43076 34733 43169 34819
rect 43255 34733 43337 34819
rect 43423 34733 43516 34819
rect 43076 33307 43516 34733
rect 43076 33221 43169 33307
rect 43255 33221 43337 33307
rect 43423 33221 43516 33307
rect 43076 31795 43516 33221
rect 43076 31709 43169 31795
rect 43255 31709 43337 31795
rect 43423 31709 43516 31795
rect 43076 31666 43516 31709
rect 43076 31286 43106 31666
rect 43486 31286 43516 31666
rect 43076 30283 43516 31286
rect 43076 30197 43169 30283
rect 43255 30197 43337 30283
rect 43423 30197 43516 30283
rect 43076 28771 43516 30197
rect 43076 28685 43169 28771
rect 43255 28685 43337 28771
rect 43423 28685 43516 28771
rect 43076 27666 43516 28685
rect 43076 27286 43106 27666
rect 43486 27286 43516 27666
rect 43076 27259 43516 27286
rect 43076 27173 43169 27259
rect 43255 27173 43337 27259
rect 43423 27173 43516 27259
rect 43076 25747 43516 27173
rect 43076 25661 43169 25747
rect 43255 25661 43337 25747
rect 43423 25661 43516 25747
rect 43076 24235 43516 25661
rect 43076 24149 43169 24235
rect 43255 24149 43337 24235
rect 43423 24149 43516 24235
rect 43076 23666 43516 24149
rect 43076 23286 43106 23666
rect 43486 23286 43516 23666
rect 43076 22723 43516 23286
rect 43076 22637 43169 22723
rect 43255 22637 43337 22723
rect 43423 22637 43516 22723
rect 43076 21211 43516 22637
rect 43076 21125 43169 21211
rect 43255 21125 43337 21211
rect 43423 21125 43516 21211
rect 43076 19699 43516 21125
rect 43076 19666 43169 19699
rect 43255 19666 43337 19699
rect 43423 19666 43516 19699
rect 43076 19286 43106 19666
rect 43486 19286 43516 19666
rect 43076 18187 43516 19286
rect 43076 18101 43169 18187
rect 43255 18101 43337 18187
rect 43423 18101 43516 18187
rect 43076 16675 43516 18101
rect 43076 16589 43169 16675
rect 43255 16589 43337 16675
rect 43423 16589 43516 16675
rect 43076 15666 43516 16589
rect 43076 15286 43106 15666
rect 43486 15286 43516 15666
rect 43076 15163 43516 15286
rect 43076 15077 43169 15163
rect 43255 15077 43337 15163
rect 43423 15077 43516 15163
rect 43076 13651 43516 15077
rect 43076 13565 43169 13651
rect 43255 13565 43337 13651
rect 43423 13565 43516 13651
rect 43076 12139 43516 13565
rect 43076 12053 43169 12139
rect 43255 12053 43337 12139
rect 43423 12053 43516 12139
rect 43076 11666 43516 12053
rect 43076 11286 43106 11666
rect 43486 11286 43516 11666
rect 43076 10627 43516 11286
rect 43076 10541 43169 10627
rect 43255 10541 43337 10627
rect 43423 10541 43516 10627
rect 43076 9115 43516 10541
rect 43076 9029 43169 9115
rect 43255 9029 43337 9115
rect 43423 9029 43516 9115
rect 43076 7666 43516 9029
rect 43076 7286 43106 7666
rect 43486 7286 43516 7666
rect 43076 6091 43516 7286
rect 43076 6005 43169 6091
rect 43255 6005 43337 6091
rect 43423 6005 43516 6091
rect 43076 4579 43516 6005
rect 43076 4493 43169 4579
rect 43255 4493 43337 4579
rect 43423 4493 43516 4579
rect 43076 3666 43516 4493
rect 43076 3286 43106 3666
rect 43486 3286 43516 3666
rect 43076 3067 43516 3286
rect 43076 2981 43169 3067
rect 43255 2981 43337 3067
rect 43423 2981 43516 3067
rect 43076 1555 43516 2981
rect 43076 1469 43169 1555
rect 43255 1469 43337 1555
rect 43423 1469 43516 1555
rect 43076 712 43516 1469
rect 44316 38599 44756 38682
rect 44316 38513 44409 38599
rect 44495 38513 44577 38599
rect 44663 38513 44756 38599
rect 44316 37087 44756 38513
rect 44316 37001 44409 37087
rect 44495 37001 44577 37087
rect 44663 37001 44756 37087
rect 44316 36906 44756 37001
rect 44316 36526 44346 36906
rect 44726 36526 44756 36906
rect 44316 35575 44756 36526
rect 44316 35489 44409 35575
rect 44495 35489 44577 35575
rect 44663 35489 44756 35575
rect 44316 34063 44756 35489
rect 44316 33977 44409 34063
rect 44495 33977 44577 34063
rect 44663 33977 44756 34063
rect 44316 32906 44756 33977
rect 44316 32526 44346 32906
rect 44726 32526 44756 32906
rect 44316 32465 44409 32526
rect 44495 32465 44577 32526
rect 44663 32465 44756 32526
rect 44316 31039 44756 32465
rect 44316 30953 44409 31039
rect 44495 30953 44577 31039
rect 44663 30953 44756 31039
rect 44316 29527 44756 30953
rect 44316 29441 44409 29527
rect 44495 29441 44577 29527
rect 44663 29441 44756 29527
rect 44316 28906 44756 29441
rect 44316 28526 44346 28906
rect 44726 28526 44756 28906
rect 44316 28015 44756 28526
rect 44316 27929 44409 28015
rect 44495 27929 44577 28015
rect 44663 27929 44756 28015
rect 44316 26503 44756 27929
rect 44316 26417 44409 26503
rect 44495 26417 44577 26503
rect 44663 26417 44756 26503
rect 44316 24991 44756 26417
rect 44316 24906 44409 24991
rect 44495 24906 44577 24991
rect 44663 24906 44756 24991
rect 44316 24526 44346 24906
rect 44726 24526 44756 24906
rect 44316 23479 44756 24526
rect 44316 23393 44409 23479
rect 44495 23393 44577 23479
rect 44663 23393 44756 23479
rect 44316 21967 44756 23393
rect 44316 21881 44409 21967
rect 44495 21881 44577 21967
rect 44663 21881 44756 21967
rect 44316 20906 44756 21881
rect 44316 20526 44346 20906
rect 44726 20526 44756 20906
rect 44316 20455 44756 20526
rect 44316 20369 44409 20455
rect 44495 20369 44577 20455
rect 44663 20369 44756 20455
rect 44316 18943 44756 20369
rect 44316 18857 44409 18943
rect 44495 18857 44577 18943
rect 44663 18857 44756 18943
rect 44316 17431 44756 18857
rect 44316 17345 44409 17431
rect 44495 17345 44577 17431
rect 44663 17345 44756 17431
rect 44316 16906 44756 17345
rect 44316 16526 44346 16906
rect 44726 16526 44756 16906
rect 44316 15919 44756 16526
rect 44316 15833 44409 15919
rect 44495 15833 44577 15919
rect 44663 15833 44756 15919
rect 44316 14407 44756 15833
rect 44316 14321 44409 14407
rect 44495 14321 44577 14407
rect 44663 14321 44756 14407
rect 44316 12906 44756 14321
rect 44316 12526 44346 12906
rect 44726 12526 44756 12906
rect 44316 11383 44756 12526
rect 44316 11297 44409 11383
rect 44495 11297 44577 11383
rect 44663 11297 44756 11383
rect 44316 9871 44756 11297
rect 44316 9785 44409 9871
rect 44495 9785 44577 9871
rect 44663 9785 44756 9871
rect 44316 8906 44756 9785
rect 44316 8526 44346 8906
rect 44726 8526 44756 8906
rect 44316 8359 44756 8526
rect 44316 8273 44409 8359
rect 44495 8273 44577 8359
rect 44663 8273 44756 8359
rect 44316 6847 44756 8273
rect 44316 6761 44409 6847
rect 44495 6761 44577 6847
rect 44663 6761 44756 6847
rect 44316 5335 44756 6761
rect 44316 5249 44409 5335
rect 44495 5249 44577 5335
rect 44663 5249 44756 5335
rect 44316 4906 44756 5249
rect 44316 4526 44346 4906
rect 44726 4526 44756 4906
rect 44316 3823 44756 4526
rect 44316 3737 44409 3823
rect 44495 3737 44577 3823
rect 44663 3737 44756 3823
rect 44316 2311 44756 3737
rect 44316 2225 44409 2311
rect 44495 2225 44577 2311
rect 44663 2225 44756 2311
rect 44316 799 44756 2225
rect 44316 713 44409 799
rect 44495 713 44577 799
rect 44663 713 44756 799
rect 44316 630 44756 713
rect 47076 37843 47516 38600
rect 47076 37757 47169 37843
rect 47255 37757 47337 37843
rect 47423 37757 47516 37843
rect 47076 36331 47516 37757
rect 47076 36245 47169 36331
rect 47255 36245 47337 36331
rect 47423 36245 47516 36331
rect 47076 35666 47516 36245
rect 47076 35286 47106 35666
rect 47486 35286 47516 35666
rect 47076 34819 47516 35286
rect 47076 34733 47169 34819
rect 47255 34733 47337 34819
rect 47423 34733 47516 34819
rect 47076 33307 47516 34733
rect 47076 33221 47169 33307
rect 47255 33221 47337 33307
rect 47423 33221 47516 33307
rect 47076 31795 47516 33221
rect 47076 31709 47169 31795
rect 47255 31709 47337 31795
rect 47423 31709 47516 31795
rect 47076 31666 47516 31709
rect 47076 31286 47106 31666
rect 47486 31286 47516 31666
rect 47076 30283 47516 31286
rect 47076 30197 47169 30283
rect 47255 30197 47337 30283
rect 47423 30197 47516 30283
rect 47076 28771 47516 30197
rect 47076 28685 47169 28771
rect 47255 28685 47337 28771
rect 47423 28685 47516 28771
rect 47076 27666 47516 28685
rect 47076 27286 47106 27666
rect 47486 27286 47516 27666
rect 47076 27259 47516 27286
rect 47076 27173 47169 27259
rect 47255 27173 47337 27259
rect 47423 27173 47516 27259
rect 47076 25747 47516 27173
rect 47076 25661 47169 25747
rect 47255 25661 47337 25747
rect 47423 25661 47516 25747
rect 47076 24235 47516 25661
rect 47076 24149 47169 24235
rect 47255 24149 47337 24235
rect 47423 24149 47516 24235
rect 47076 23666 47516 24149
rect 47076 23286 47106 23666
rect 47486 23286 47516 23666
rect 47076 22723 47516 23286
rect 47076 22637 47169 22723
rect 47255 22637 47337 22723
rect 47423 22637 47516 22723
rect 47076 21211 47516 22637
rect 47076 21125 47169 21211
rect 47255 21125 47337 21211
rect 47423 21125 47516 21211
rect 47076 19699 47516 21125
rect 47076 19666 47169 19699
rect 47255 19666 47337 19699
rect 47423 19666 47516 19699
rect 47076 19286 47106 19666
rect 47486 19286 47516 19666
rect 47076 18187 47516 19286
rect 47076 18101 47169 18187
rect 47255 18101 47337 18187
rect 47423 18101 47516 18187
rect 47076 16675 47516 18101
rect 47076 16589 47169 16675
rect 47255 16589 47337 16675
rect 47423 16589 47516 16675
rect 47076 15666 47516 16589
rect 47076 15286 47106 15666
rect 47486 15286 47516 15666
rect 47076 15163 47516 15286
rect 47076 15077 47169 15163
rect 47255 15077 47337 15163
rect 47423 15077 47516 15163
rect 47076 13651 47516 15077
rect 47076 13565 47169 13651
rect 47255 13565 47337 13651
rect 47423 13565 47516 13651
rect 47076 12139 47516 13565
rect 47076 12053 47169 12139
rect 47255 12053 47337 12139
rect 47423 12053 47516 12139
rect 47076 11666 47516 12053
rect 47076 11286 47106 11666
rect 47486 11286 47516 11666
rect 47076 10627 47516 11286
rect 47076 10541 47169 10627
rect 47255 10541 47337 10627
rect 47423 10541 47516 10627
rect 47076 9115 47516 10541
rect 47076 9029 47169 9115
rect 47255 9029 47337 9115
rect 47423 9029 47516 9115
rect 47076 7666 47516 9029
rect 47076 7286 47106 7666
rect 47486 7286 47516 7666
rect 47076 6091 47516 7286
rect 47076 6005 47169 6091
rect 47255 6005 47337 6091
rect 47423 6005 47516 6091
rect 47076 4579 47516 6005
rect 47076 4493 47169 4579
rect 47255 4493 47337 4579
rect 47423 4493 47516 4579
rect 47076 3666 47516 4493
rect 47076 3286 47106 3666
rect 47486 3286 47516 3666
rect 47076 3067 47516 3286
rect 47076 2981 47169 3067
rect 47255 2981 47337 3067
rect 47423 2981 47516 3067
rect 47076 1555 47516 2981
rect 47076 1469 47169 1555
rect 47255 1469 47337 1555
rect 47423 1469 47516 1555
rect 47076 712 47516 1469
rect 48316 38599 48756 38682
rect 48316 38513 48409 38599
rect 48495 38513 48577 38599
rect 48663 38513 48756 38599
rect 48316 37087 48756 38513
rect 48316 37001 48409 37087
rect 48495 37001 48577 37087
rect 48663 37001 48756 37087
rect 48316 36906 48756 37001
rect 48316 36526 48346 36906
rect 48726 36526 48756 36906
rect 48316 35575 48756 36526
rect 48316 35489 48409 35575
rect 48495 35489 48577 35575
rect 48663 35489 48756 35575
rect 48316 34063 48756 35489
rect 48316 33977 48409 34063
rect 48495 33977 48577 34063
rect 48663 33977 48756 34063
rect 48316 32906 48756 33977
rect 48316 32526 48346 32906
rect 48726 32526 48756 32906
rect 48316 32465 48409 32526
rect 48495 32465 48577 32526
rect 48663 32465 48756 32526
rect 48316 31039 48756 32465
rect 48316 30953 48409 31039
rect 48495 30953 48577 31039
rect 48663 30953 48756 31039
rect 48316 29527 48756 30953
rect 48316 29441 48409 29527
rect 48495 29441 48577 29527
rect 48663 29441 48756 29527
rect 48316 28906 48756 29441
rect 48316 28526 48346 28906
rect 48726 28526 48756 28906
rect 48316 28015 48756 28526
rect 48316 27929 48409 28015
rect 48495 27929 48577 28015
rect 48663 27929 48756 28015
rect 48316 26503 48756 27929
rect 48316 26417 48409 26503
rect 48495 26417 48577 26503
rect 48663 26417 48756 26503
rect 48316 24991 48756 26417
rect 48316 24906 48409 24991
rect 48495 24906 48577 24991
rect 48663 24906 48756 24991
rect 48316 24526 48346 24906
rect 48726 24526 48756 24906
rect 48316 23479 48756 24526
rect 48316 23393 48409 23479
rect 48495 23393 48577 23479
rect 48663 23393 48756 23479
rect 48316 21967 48756 23393
rect 48316 21881 48409 21967
rect 48495 21881 48577 21967
rect 48663 21881 48756 21967
rect 48316 20906 48756 21881
rect 48316 20526 48346 20906
rect 48726 20526 48756 20906
rect 48316 20455 48756 20526
rect 48316 20369 48409 20455
rect 48495 20369 48577 20455
rect 48663 20369 48756 20455
rect 48316 18943 48756 20369
rect 48316 18857 48409 18943
rect 48495 18857 48577 18943
rect 48663 18857 48756 18943
rect 48316 17431 48756 18857
rect 48316 17345 48409 17431
rect 48495 17345 48577 17431
rect 48663 17345 48756 17431
rect 48316 16906 48756 17345
rect 48316 16526 48346 16906
rect 48726 16526 48756 16906
rect 48316 15919 48756 16526
rect 48316 15833 48409 15919
rect 48495 15833 48577 15919
rect 48663 15833 48756 15919
rect 48316 14407 48756 15833
rect 48316 14321 48409 14407
rect 48495 14321 48577 14407
rect 48663 14321 48756 14407
rect 48316 12906 48756 14321
rect 48316 12526 48346 12906
rect 48726 12526 48756 12906
rect 48316 11383 48756 12526
rect 48316 11297 48409 11383
rect 48495 11297 48577 11383
rect 48663 11297 48756 11383
rect 48316 9871 48756 11297
rect 48316 9785 48409 9871
rect 48495 9785 48577 9871
rect 48663 9785 48756 9871
rect 48316 8906 48756 9785
rect 48316 8526 48346 8906
rect 48726 8526 48756 8906
rect 48316 8359 48756 8526
rect 48316 8273 48409 8359
rect 48495 8273 48577 8359
rect 48663 8273 48756 8359
rect 48316 6847 48756 8273
rect 48316 6761 48409 6847
rect 48495 6761 48577 6847
rect 48663 6761 48756 6847
rect 48316 5335 48756 6761
rect 48316 5249 48409 5335
rect 48495 5249 48577 5335
rect 48663 5249 48756 5335
rect 48316 4906 48756 5249
rect 48316 4526 48346 4906
rect 48726 4526 48756 4906
rect 48316 3823 48756 4526
rect 48316 3737 48409 3823
rect 48495 3737 48577 3823
rect 48663 3737 48756 3823
rect 48316 2311 48756 3737
rect 48316 2225 48409 2311
rect 48495 2225 48577 2311
rect 48663 2225 48756 2311
rect 48316 799 48756 2225
rect 48316 713 48409 799
rect 48495 713 48577 799
rect 48663 713 48756 799
rect 48316 630 48756 713
rect 51076 37843 51516 38600
rect 51076 37757 51169 37843
rect 51255 37757 51337 37843
rect 51423 37757 51516 37843
rect 51076 36331 51516 37757
rect 51076 36245 51169 36331
rect 51255 36245 51337 36331
rect 51423 36245 51516 36331
rect 51076 35666 51516 36245
rect 51076 35286 51106 35666
rect 51486 35286 51516 35666
rect 51076 34819 51516 35286
rect 51076 34733 51169 34819
rect 51255 34733 51337 34819
rect 51423 34733 51516 34819
rect 51076 33307 51516 34733
rect 51076 33221 51169 33307
rect 51255 33221 51337 33307
rect 51423 33221 51516 33307
rect 51076 31795 51516 33221
rect 51076 31709 51169 31795
rect 51255 31709 51337 31795
rect 51423 31709 51516 31795
rect 51076 31666 51516 31709
rect 51076 31286 51106 31666
rect 51486 31286 51516 31666
rect 51076 30283 51516 31286
rect 51076 30197 51169 30283
rect 51255 30197 51337 30283
rect 51423 30197 51516 30283
rect 51076 28771 51516 30197
rect 51076 28685 51169 28771
rect 51255 28685 51337 28771
rect 51423 28685 51516 28771
rect 51076 27666 51516 28685
rect 51076 27286 51106 27666
rect 51486 27286 51516 27666
rect 51076 27259 51516 27286
rect 51076 27173 51169 27259
rect 51255 27173 51337 27259
rect 51423 27173 51516 27259
rect 51076 25747 51516 27173
rect 51076 25661 51169 25747
rect 51255 25661 51337 25747
rect 51423 25661 51516 25747
rect 51076 24235 51516 25661
rect 51076 24149 51169 24235
rect 51255 24149 51337 24235
rect 51423 24149 51516 24235
rect 51076 23666 51516 24149
rect 51076 23286 51106 23666
rect 51486 23286 51516 23666
rect 51076 22723 51516 23286
rect 51076 22637 51169 22723
rect 51255 22637 51337 22723
rect 51423 22637 51516 22723
rect 51076 21211 51516 22637
rect 51076 21125 51169 21211
rect 51255 21125 51337 21211
rect 51423 21125 51516 21211
rect 51076 19699 51516 21125
rect 51076 19666 51169 19699
rect 51255 19666 51337 19699
rect 51423 19666 51516 19699
rect 51076 19286 51106 19666
rect 51486 19286 51516 19666
rect 51076 18187 51516 19286
rect 51076 18101 51169 18187
rect 51255 18101 51337 18187
rect 51423 18101 51516 18187
rect 51076 16675 51516 18101
rect 51076 16589 51169 16675
rect 51255 16589 51337 16675
rect 51423 16589 51516 16675
rect 51076 15666 51516 16589
rect 51076 15286 51106 15666
rect 51486 15286 51516 15666
rect 51076 15163 51516 15286
rect 51076 15077 51169 15163
rect 51255 15077 51337 15163
rect 51423 15077 51516 15163
rect 51076 13651 51516 15077
rect 51076 13565 51169 13651
rect 51255 13565 51337 13651
rect 51423 13565 51516 13651
rect 51076 12139 51516 13565
rect 51076 12053 51169 12139
rect 51255 12053 51337 12139
rect 51423 12053 51516 12139
rect 51076 11666 51516 12053
rect 51076 11286 51106 11666
rect 51486 11286 51516 11666
rect 51076 10627 51516 11286
rect 51076 10541 51169 10627
rect 51255 10541 51337 10627
rect 51423 10541 51516 10627
rect 51076 9115 51516 10541
rect 51076 9029 51169 9115
rect 51255 9029 51337 9115
rect 51423 9029 51516 9115
rect 51076 7666 51516 9029
rect 51076 7286 51106 7666
rect 51486 7286 51516 7666
rect 51076 6091 51516 7286
rect 51076 6005 51169 6091
rect 51255 6005 51337 6091
rect 51423 6005 51516 6091
rect 51076 4579 51516 6005
rect 51076 4493 51169 4579
rect 51255 4493 51337 4579
rect 51423 4493 51516 4579
rect 51076 3666 51516 4493
rect 51076 3286 51106 3666
rect 51486 3286 51516 3666
rect 51076 3067 51516 3286
rect 51076 2981 51169 3067
rect 51255 2981 51337 3067
rect 51423 2981 51516 3067
rect 51076 1555 51516 2981
rect 51076 1469 51169 1555
rect 51255 1469 51337 1555
rect 51423 1469 51516 1555
rect 51076 712 51516 1469
rect 52316 38599 52756 38682
rect 52316 38513 52409 38599
rect 52495 38513 52577 38599
rect 52663 38513 52756 38599
rect 52316 37087 52756 38513
rect 52316 37001 52409 37087
rect 52495 37001 52577 37087
rect 52663 37001 52756 37087
rect 52316 36906 52756 37001
rect 52316 36526 52346 36906
rect 52726 36526 52756 36906
rect 52316 35575 52756 36526
rect 52316 35489 52409 35575
rect 52495 35489 52577 35575
rect 52663 35489 52756 35575
rect 52316 34063 52756 35489
rect 52316 33977 52409 34063
rect 52495 33977 52577 34063
rect 52663 33977 52756 34063
rect 52316 32906 52756 33977
rect 52316 32526 52346 32906
rect 52726 32526 52756 32906
rect 52316 32465 52409 32526
rect 52495 32465 52577 32526
rect 52663 32465 52756 32526
rect 52316 31039 52756 32465
rect 52316 30953 52409 31039
rect 52495 30953 52577 31039
rect 52663 30953 52756 31039
rect 52316 29527 52756 30953
rect 52316 29441 52409 29527
rect 52495 29441 52577 29527
rect 52663 29441 52756 29527
rect 52316 28906 52756 29441
rect 52316 28526 52346 28906
rect 52726 28526 52756 28906
rect 52316 28015 52756 28526
rect 52316 27929 52409 28015
rect 52495 27929 52577 28015
rect 52663 27929 52756 28015
rect 52316 26503 52756 27929
rect 52316 26417 52409 26503
rect 52495 26417 52577 26503
rect 52663 26417 52756 26503
rect 52316 24991 52756 26417
rect 52316 24906 52409 24991
rect 52495 24906 52577 24991
rect 52663 24906 52756 24991
rect 52316 24526 52346 24906
rect 52726 24526 52756 24906
rect 52316 23479 52756 24526
rect 52316 23393 52409 23479
rect 52495 23393 52577 23479
rect 52663 23393 52756 23479
rect 52316 21967 52756 23393
rect 52316 21881 52409 21967
rect 52495 21881 52577 21967
rect 52663 21881 52756 21967
rect 52316 20906 52756 21881
rect 52316 20526 52346 20906
rect 52726 20526 52756 20906
rect 52316 20455 52756 20526
rect 52316 20369 52409 20455
rect 52495 20369 52577 20455
rect 52663 20369 52756 20455
rect 52316 18943 52756 20369
rect 52316 18857 52409 18943
rect 52495 18857 52577 18943
rect 52663 18857 52756 18943
rect 52316 17431 52756 18857
rect 52316 17345 52409 17431
rect 52495 17345 52577 17431
rect 52663 17345 52756 17431
rect 52316 16906 52756 17345
rect 52316 16526 52346 16906
rect 52726 16526 52756 16906
rect 52316 15919 52756 16526
rect 52316 15833 52409 15919
rect 52495 15833 52577 15919
rect 52663 15833 52756 15919
rect 52316 14407 52756 15833
rect 52316 14321 52409 14407
rect 52495 14321 52577 14407
rect 52663 14321 52756 14407
rect 52316 12906 52756 14321
rect 52316 12526 52346 12906
rect 52726 12526 52756 12906
rect 52316 11383 52756 12526
rect 52316 11297 52409 11383
rect 52495 11297 52577 11383
rect 52663 11297 52756 11383
rect 52316 9871 52756 11297
rect 52316 9785 52409 9871
rect 52495 9785 52577 9871
rect 52663 9785 52756 9871
rect 52316 8906 52756 9785
rect 52316 8526 52346 8906
rect 52726 8526 52756 8906
rect 52316 8359 52756 8526
rect 52316 8273 52409 8359
rect 52495 8273 52577 8359
rect 52663 8273 52756 8359
rect 52316 6847 52756 8273
rect 52316 6761 52409 6847
rect 52495 6761 52577 6847
rect 52663 6761 52756 6847
rect 52316 5335 52756 6761
rect 52316 5249 52409 5335
rect 52495 5249 52577 5335
rect 52663 5249 52756 5335
rect 52316 4906 52756 5249
rect 52316 4526 52346 4906
rect 52726 4526 52756 4906
rect 52316 3823 52756 4526
rect 52316 3737 52409 3823
rect 52495 3737 52577 3823
rect 52663 3737 52756 3823
rect 52316 2311 52756 3737
rect 52316 2225 52409 2311
rect 52495 2225 52577 2311
rect 52663 2225 52756 2311
rect 52316 799 52756 2225
rect 52316 713 52409 799
rect 52495 713 52577 799
rect 52663 713 52756 799
rect 52316 630 52756 713
rect 55076 37843 55516 38600
rect 55076 37757 55169 37843
rect 55255 37757 55337 37843
rect 55423 37757 55516 37843
rect 55076 36331 55516 37757
rect 55076 36245 55169 36331
rect 55255 36245 55337 36331
rect 55423 36245 55516 36331
rect 55076 35666 55516 36245
rect 55076 35286 55106 35666
rect 55486 35286 55516 35666
rect 55076 34819 55516 35286
rect 55076 34733 55169 34819
rect 55255 34733 55337 34819
rect 55423 34733 55516 34819
rect 55076 33307 55516 34733
rect 55076 33221 55169 33307
rect 55255 33221 55337 33307
rect 55423 33221 55516 33307
rect 55076 31795 55516 33221
rect 55076 31709 55169 31795
rect 55255 31709 55337 31795
rect 55423 31709 55516 31795
rect 55076 31666 55516 31709
rect 55076 31286 55106 31666
rect 55486 31286 55516 31666
rect 55076 30283 55516 31286
rect 55076 30197 55169 30283
rect 55255 30197 55337 30283
rect 55423 30197 55516 30283
rect 55076 28771 55516 30197
rect 55076 28685 55169 28771
rect 55255 28685 55337 28771
rect 55423 28685 55516 28771
rect 55076 27666 55516 28685
rect 55076 27286 55106 27666
rect 55486 27286 55516 27666
rect 55076 27259 55516 27286
rect 55076 27173 55169 27259
rect 55255 27173 55337 27259
rect 55423 27173 55516 27259
rect 55076 25747 55516 27173
rect 55076 25661 55169 25747
rect 55255 25661 55337 25747
rect 55423 25661 55516 25747
rect 55076 24235 55516 25661
rect 55076 24149 55169 24235
rect 55255 24149 55337 24235
rect 55423 24149 55516 24235
rect 55076 23666 55516 24149
rect 55076 23286 55106 23666
rect 55486 23286 55516 23666
rect 55076 22723 55516 23286
rect 55076 22637 55169 22723
rect 55255 22637 55337 22723
rect 55423 22637 55516 22723
rect 55076 21211 55516 22637
rect 55076 21125 55169 21211
rect 55255 21125 55337 21211
rect 55423 21125 55516 21211
rect 55076 19699 55516 21125
rect 55076 19666 55169 19699
rect 55255 19666 55337 19699
rect 55423 19666 55516 19699
rect 55076 19286 55106 19666
rect 55486 19286 55516 19666
rect 55076 18187 55516 19286
rect 55076 18101 55169 18187
rect 55255 18101 55337 18187
rect 55423 18101 55516 18187
rect 55076 16675 55516 18101
rect 55076 16589 55169 16675
rect 55255 16589 55337 16675
rect 55423 16589 55516 16675
rect 55076 15666 55516 16589
rect 55076 15286 55106 15666
rect 55486 15286 55516 15666
rect 55076 15163 55516 15286
rect 55076 15077 55169 15163
rect 55255 15077 55337 15163
rect 55423 15077 55516 15163
rect 55076 13651 55516 15077
rect 55076 13565 55169 13651
rect 55255 13565 55337 13651
rect 55423 13565 55516 13651
rect 55076 12139 55516 13565
rect 55076 12053 55169 12139
rect 55255 12053 55337 12139
rect 55423 12053 55516 12139
rect 55076 11666 55516 12053
rect 55076 11286 55106 11666
rect 55486 11286 55516 11666
rect 55076 10627 55516 11286
rect 55076 10541 55169 10627
rect 55255 10541 55337 10627
rect 55423 10541 55516 10627
rect 55076 9115 55516 10541
rect 55076 9029 55169 9115
rect 55255 9029 55337 9115
rect 55423 9029 55516 9115
rect 55076 7666 55516 9029
rect 55076 7286 55106 7666
rect 55486 7286 55516 7666
rect 55076 6091 55516 7286
rect 55076 6005 55169 6091
rect 55255 6005 55337 6091
rect 55423 6005 55516 6091
rect 55076 4579 55516 6005
rect 55076 4493 55169 4579
rect 55255 4493 55337 4579
rect 55423 4493 55516 4579
rect 55076 3666 55516 4493
rect 55076 3286 55106 3666
rect 55486 3286 55516 3666
rect 55076 3067 55516 3286
rect 55076 2981 55169 3067
rect 55255 2981 55337 3067
rect 55423 2981 55516 3067
rect 55076 1555 55516 2981
rect 55076 1469 55169 1555
rect 55255 1469 55337 1555
rect 55423 1469 55516 1555
rect 55076 712 55516 1469
rect 56316 38599 56756 38682
rect 56316 38513 56409 38599
rect 56495 38513 56577 38599
rect 56663 38513 56756 38599
rect 56316 37087 56756 38513
rect 56316 37001 56409 37087
rect 56495 37001 56577 37087
rect 56663 37001 56756 37087
rect 56316 36906 56756 37001
rect 56316 36526 56346 36906
rect 56726 36526 56756 36906
rect 56316 35575 56756 36526
rect 56316 35489 56409 35575
rect 56495 35489 56577 35575
rect 56663 35489 56756 35575
rect 56316 34063 56756 35489
rect 56316 33977 56409 34063
rect 56495 33977 56577 34063
rect 56663 33977 56756 34063
rect 56316 32906 56756 33977
rect 56316 32526 56346 32906
rect 56726 32526 56756 32906
rect 56316 32465 56409 32526
rect 56495 32465 56577 32526
rect 56663 32465 56756 32526
rect 56316 31039 56756 32465
rect 56316 30953 56409 31039
rect 56495 30953 56577 31039
rect 56663 30953 56756 31039
rect 56316 29527 56756 30953
rect 56316 29441 56409 29527
rect 56495 29441 56577 29527
rect 56663 29441 56756 29527
rect 56316 28906 56756 29441
rect 56316 28526 56346 28906
rect 56726 28526 56756 28906
rect 56316 28015 56756 28526
rect 56316 27929 56409 28015
rect 56495 27929 56577 28015
rect 56663 27929 56756 28015
rect 56316 26503 56756 27929
rect 56316 26417 56409 26503
rect 56495 26417 56577 26503
rect 56663 26417 56756 26503
rect 56316 24991 56756 26417
rect 56316 24906 56409 24991
rect 56495 24906 56577 24991
rect 56663 24906 56756 24991
rect 56316 24526 56346 24906
rect 56726 24526 56756 24906
rect 56316 23479 56756 24526
rect 56316 23393 56409 23479
rect 56495 23393 56577 23479
rect 56663 23393 56756 23479
rect 56316 21967 56756 23393
rect 56316 21881 56409 21967
rect 56495 21881 56577 21967
rect 56663 21881 56756 21967
rect 56316 20906 56756 21881
rect 56316 20526 56346 20906
rect 56726 20526 56756 20906
rect 56316 20455 56756 20526
rect 56316 20369 56409 20455
rect 56495 20369 56577 20455
rect 56663 20369 56756 20455
rect 56316 18943 56756 20369
rect 56316 18857 56409 18943
rect 56495 18857 56577 18943
rect 56663 18857 56756 18943
rect 56316 17431 56756 18857
rect 56316 17345 56409 17431
rect 56495 17345 56577 17431
rect 56663 17345 56756 17431
rect 56316 16906 56756 17345
rect 56316 16526 56346 16906
rect 56726 16526 56756 16906
rect 56316 15919 56756 16526
rect 56316 15833 56409 15919
rect 56495 15833 56577 15919
rect 56663 15833 56756 15919
rect 56316 14407 56756 15833
rect 56316 14321 56409 14407
rect 56495 14321 56577 14407
rect 56663 14321 56756 14407
rect 56316 12906 56756 14321
rect 56316 12526 56346 12906
rect 56726 12526 56756 12906
rect 56316 11383 56756 12526
rect 56316 11297 56409 11383
rect 56495 11297 56577 11383
rect 56663 11297 56756 11383
rect 56316 9871 56756 11297
rect 56316 9785 56409 9871
rect 56495 9785 56577 9871
rect 56663 9785 56756 9871
rect 56316 8906 56756 9785
rect 56316 8526 56346 8906
rect 56726 8526 56756 8906
rect 56316 8359 56756 8526
rect 56316 8273 56409 8359
rect 56495 8273 56577 8359
rect 56663 8273 56756 8359
rect 56316 6847 56756 8273
rect 56316 6761 56409 6847
rect 56495 6761 56577 6847
rect 56663 6761 56756 6847
rect 56316 5335 56756 6761
rect 56316 5249 56409 5335
rect 56495 5249 56577 5335
rect 56663 5249 56756 5335
rect 56316 4906 56756 5249
rect 56316 4526 56346 4906
rect 56726 4526 56756 4906
rect 56316 3823 56756 4526
rect 56316 3737 56409 3823
rect 56495 3737 56577 3823
rect 56663 3737 56756 3823
rect 56316 2311 56756 3737
rect 56316 2225 56409 2311
rect 56495 2225 56577 2311
rect 56663 2225 56756 2311
rect 56316 799 56756 2225
rect 56316 713 56409 799
rect 56495 713 56577 799
rect 56663 713 56756 799
rect 56316 630 56756 713
rect 59076 37843 59516 38600
rect 59076 37757 59169 37843
rect 59255 37757 59337 37843
rect 59423 37757 59516 37843
rect 59076 36331 59516 37757
rect 59076 36245 59169 36331
rect 59255 36245 59337 36331
rect 59423 36245 59516 36331
rect 59076 35666 59516 36245
rect 59076 35286 59106 35666
rect 59486 35286 59516 35666
rect 59076 34819 59516 35286
rect 59076 34733 59169 34819
rect 59255 34733 59337 34819
rect 59423 34733 59516 34819
rect 59076 33307 59516 34733
rect 59076 33221 59169 33307
rect 59255 33221 59337 33307
rect 59423 33221 59516 33307
rect 59076 31795 59516 33221
rect 59076 31709 59169 31795
rect 59255 31709 59337 31795
rect 59423 31709 59516 31795
rect 59076 31666 59516 31709
rect 59076 31286 59106 31666
rect 59486 31286 59516 31666
rect 59076 30283 59516 31286
rect 59076 30197 59169 30283
rect 59255 30197 59337 30283
rect 59423 30197 59516 30283
rect 59076 28771 59516 30197
rect 59076 28685 59169 28771
rect 59255 28685 59337 28771
rect 59423 28685 59516 28771
rect 59076 27666 59516 28685
rect 59076 27286 59106 27666
rect 59486 27286 59516 27666
rect 59076 27259 59516 27286
rect 59076 27173 59169 27259
rect 59255 27173 59337 27259
rect 59423 27173 59516 27259
rect 59076 25747 59516 27173
rect 59076 25661 59169 25747
rect 59255 25661 59337 25747
rect 59423 25661 59516 25747
rect 59076 24235 59516 25661
rect 59076 24149 59169 24235
rect 59255 24149 59337 24235
rect 59423 24149 59516 24235
rect 59076 23666 59516 24149
rect 59076 23286 59106 23666
rect 59486 23286 59516 23666
rect 59076 22723 59516 23286
rect 59076 22637 59169 22723
rect 59255 22637 59337 22723
rect 59423 22637 59516 22723
rect 59076 21211 59516 22637
rect 59076 21125 59169 21211
rect 59255 21125 59337 21211
rect 59423 21125 59516 21211
rect 59076 19699 59516 21125
rect 59076 19666 59169 19699
rect 59255 19666 59337 19699
rect 59423 19666 59516 19699
rect 59076 19286 59106 19666
rect 59486 19286 59516 19666
rect 59076 18187 59516 19286
rect 59076 18101 59169 18187
rect 59255 18101 59337 18187
rect 59423 18101 59516 18187
rect 59076 16675 59516 18101
rect 59076 16589 59169 16675
rect 59255 16589 59337 16675
rect 59423 16589 59516 16675
rect 59076 15666 59516 16589
rect 59076 15286 59106 15666
rect 59486 15286 59516 15666
rect 59076 15163 59516 15286
rect 59076 15077 59169 15163
rect 59255 15077 59337 15163
rect 59423 15077 59516 15163
rect 59076 13651 59516 15077
rect 59076 13565 59169 13651
rect 59255 13565 59337 13651
rect 59423 13565 59516 13651
rect 59076 12139 59516 13565
rect 59076 12053 59169 12139
rect 59255 12053 59337 12139
rect 59423 12053 59516 12139
rect 59076 11666 59516 12053
rect 59076 11286 59106 11666
rect 59486 11286 59516 11666
rect 59076 10627 59516 11286
rect 59076 10541 59169 10627
rect 59255 10541 59337 10627
rect 59423 10541 59516 10627
rect 59076 9115 59516 10541
rect 59076 9029 59169 9115
rect 59255 9029 59337 9115
rect 59423 9029 59516 9115
rect 59076 7666 59516 9029
rect 59076 7286 59106 7666
rect 59486 7286 59516 7666
rect 59076 6091 59516 7286
rect 59076 6005 59169 6091
rect 59255 6005 59337 6091
rect 59423 6005 59516 6091
rect 59076 4579 59516 6005
rect 59076 4493 59169 4579
rect 59255 4493 59337 4579
rect 59423 4493 59516 4579
rect 59076 3666 59516 4493
rect 59076 3286 59106 3666
rect 59486 3286 59516 3666
rect 59076 3067 59516 3286
rect 59076 2981 59169 3067
rect 59255 2981 59337 3067
rect 59423 2981 59516 3067
rect 59076 1555 59516 2981
rect 59076 1469 59169 1555
rect 59255 1469 59337 1555
rect 59423 1469 59516 1555
rect 59076 712 59516 1469
rect 60316 38599 60756 38682
rect 60316 38513 60409 38599
rect 60495 38513 60577 38599
rect 60663 38513 60756 38599
rect 60316 37087 60756 38513
rect 60316 37001 60409 37087
rect 60495 37001 60577 37087
rect 60663 37001 60756 37087
rect 60316 36906 60756 37001
rect 60316 36526 60346 36906
rect 60726 36526 60756 36906
rect 60316 35575 60756 36526
rect 60316 35489 60409 35575
rect 60495 35489 60577 35575
rect 60663 35489 60756 35575
rect 60316 34063 60756 35489
rect 60316 33977 60409 34063
rect 60495 33977 60577 34063
rect 60663 33977 60756 34063
rect 60316 32906 60756 33977
rect 60316 32526 60346 32906
rect 60726 32526 60756 32906
rect 60316 32465 60409 32526
rect 60495 32465 60577 32526
rect 60663 32465 60756 32526
rect 60316 31039 60756 32465
rect 60316 30953 60409 31039
rect 60495 30953 60577 31039
rect 60663 30953 60756 31039
rect 60316 29527 60756 30953
rect 60316 29441 60409 29527
rect 60495 29441 60577 29527
rect 60663 29441 60756 29527
rect 60316 28906 60756 29441
rect 60316 28526 60346 28906
rect 60726 28526 60756 28906
rect 60316 28015 60756 28526
rect 60316 27929 60409 28015
rect 60495 27929 60577 28015
rect 60663 27929 60756 28015
rect 60316 26503 60756 27929
rect 60316 26417 60409 26503
rect 60495 26417 60577 26503
rect 60663 26417 60756 26503
rect 60316 24991 60756 26417
rect 60316 24906 60409 24991
rect 60495 24906 60577 24991
rect 60663 24906 60756 24991
rect 60316 24526 60346 24906
rect 60726 24526 60756 24906
rect 60316 23479 60756 24526
rect 60316 23393 60409 23479
rect 60495 23393 60577 23479
rect 60663 23393 60756 23479
rect 60316 21967 60756 23393
rect 60316 21881 60409 21967
rect 60495 21881 60577 21967
rect 60663 21881 60756 21967
rect 60316 20906 60756 21881
rect 60316 20526 60346 20906
rect 60726 20526 60756 20906
rect 60316 20455 60756 20526
rect 60316 20369 60409 20455
rect 60495 20369 60577 20455
rect 60663 20369 60756 20455
rect 60316 18943 60756 20369
rect 60316 18857 60409 18943
rect 60495 18857 60577 18943
rect 60663 18857 60756 18943
rect 60316 17431 60756 18857
rect 60316 17345 60409 17431
rect 60495 17345 60577 17431
rect 60663 17345 60756 17431
rect 60316 16906 60756 17345
rect 60316 16526 60346 16906
rect 60726 16526 60756 16906
rect 60316 15919 60756 16526
rect 60316 15833 60409 15919
rect 60495 15833 60577 15919
rect 60663 15833 60756 15919
rect 60316 14407 60756 15833
rect 60316 14321 60409 14407
rect 60495 14321 60577 14407
rect 60663 14321 60756 14407
rect 60316 12906 60756 14321
rect 60316 12526 60346 12906
rect 60726 12526 60756 12906
rect 60316 11383 60756 12526
rect 60316 11297 60409 11383
rect 60495 11297 60577 11383
rect 60663 11297 60756 11383
rect 60316 9871 60756 11297
rect 60316 9785 60409 9871
rect 60495 9785 60577 9871
rect 60663 9785 60756 9871
rect 60316 8906 60756 9785
rect 60316 8526 60346 8906
rect 60726 8526 60756 8906
rect 60316 8359 60756 8526
rect 60316 8273 60409 8359
rect 60495 8273 60577 8359
rect 60663 8273 60756 8359
rect 60316 6847 60756 8273
rect 60316 6761 60409 6847
rect 60495 6761 60577 6847
rect 60663 6761 60756 6847
rect 60316 5335 60756 6761
rect 60316 5249 60409 5335
rect 60495 5249 60577 5335
rect 60663 5249 60756 5335
rect 60316 4906 60756 5249
rect 60316 4526 60346 4906
rect 60726 4526 60756 4906
rect 60316 3823 60756 4526
rect 60316 3737 60409 3823
rect 60495 3737 60577 3823
rect 60663 3737 60756 3823
rect 60316 2311 60756 3737
rect 60316 2225 60409 2311
rect 60495 2225 60577 2311
rect 60663 2225 60756 2311
rect 60316 799 60756 2225
rect 60316 713 60409 799
rect 60495 713 60577 799
rect 60663 713 60756 799
rect 60316 630 60756 713
rect 63076 37843 63516 38600
rect 63076 37757 63169 37843
rect 63255 37757 63337 37843
rect 63423 37757 63516 37843
rect 63076 36331 63516 37757
rect 63076 36245 63169 36331
rect 63255 36245 63337 36331
rect 63423 36245 63516 36331
rect 63076 35666 63516 36245
rect 63076 35286 63106 35666
rect 63486 35286 63516 35666
rect 63076 34819 63516 35286
rect 63076 34733 63169 34819
rect 63255 34733 63337 34819
rect 63423 34733 63516 34819
rect 63076 33307 63516 34733
rect 63076 33221 63169 33307
rect 63255 33221 63337 33307
rect 63423 33221 63516 33307
rect 63076 31795 63516 33221
rect 63076 31709 63169 31795
rect 63255 31709 63337 31795
rect 63423 31709 63516 31795
rect 63076 31666 63516 31709
rect 63076 31286 63106 31666
rect 63486 31286 63516 31666
rect 63076 30283 63516 31286
rect 63076 30197 63169 30283
rect 63255 30197 63337 30283
rect 63423 30197 63516 30283
rect 63076 28771 63516 30197
rect 63076 28685 63169 28771
rect 63255 28685 63337 28771
rect 63423 28685 63516 28771
rect 63076 27666 63516 28685
rect 63076 27286 63106 27666
rect 63486 27286 63516 27666
rect 63076 27259 63516 27286
rect 63076 27173 63169 27259
rect 63255 27173 63337 27259
rect 63423 27173 63516 27259
rect 63076 25747 63516 27173
rect 63076 25661 63169 25747
rect 63255 25661 63337 25747
rect 63423 25661 63516 25747
rect 63076 24235 63516 25661
rect 63076 24149 63169 24235
rect 63255 24149 63337 24235
rect 63423 24149 63516 24235
rect 63076 23666 63516 24149
rect 63076 23286 63106 23666
rect 63486 23286 63516 23666
rect 63076 22723 63516 23286
rect 63076 22637 63169 22723
rect 63255 22637 63337 22723
rect 63423 22637 63516 22723
rect 63076 21211 63516 22637
rect 63076 21125 63169 21211
rect 63255 21125 63337 21211
rect 63423 21125 63516 21211
rect 63076 19699 63516 21125
rect 63076 19666 63169 19699
rect 63255 19666 63337 19699
rect 63423 19666 63516 19699
rect 63076 19286 63106 19666
rect 63486 19286 63516 19666
rect 63076 18187 63516 19286
rect 63076 18101 63169 18187
rect 63255 18101 63337 18187
rect 63423 18101 63516 18187
rect 63076 16675 63516 18101
rect 63076 16589 63169 16675
rect 63255 16589 63337 16675
rect 63423 16589 63516 16675
rect 63076 15666 63516 16589
rect 63076 15286 63106 15666
rect 63486 15286 63516 15666
rect 63076 15163 63516 15286
rect 63076 15077 63169 15163
rect 63255 15077 63337 15163
rect 63423 15077 63516 15163
rect 63076 13651 63516 15077
rect 63076 13565 63169 13651
rect 63255 13565 63337 13651
rect 63423 13565 63516 13651
rect 63076 12139 63516 13565
rect 63076 12053 63169 12139
rect 63255 12053 63337 12139
rect 63423 12053 63516 12139
rect 63076 11666 63516 12053
rect 63076 11286 63106 11666
rect 63486 11286 63516 11666
rect 63076 10627 63516 11286
rect 63076 10541 63169 10627
rect 63255 10541 63337 10627
rect 63423 10541 63516 10627
rect 63076 9115 63516 10541
rect 63076 9029 63169 9115
rect 63255 9029 63337 9115
rect 63423 9029 63516 9115
rect 63076 7666 63516 9029
rect 63076 7286 63106 7666
rect 63486 7286 63516 7666
rect 63076 6091 63516 7286
rect 63076 6005 63169 6091
rect 63255 6005 63337 6091
rect 63423 6005 63516 6091
rect 63076 4579 63516 6005
rect 63076 4493 63169 4579
rect 63255 4493 63337 4579
rect 63423 4493 63516 4579
rect 63076 3666 63516 4493
rect 63076 3286 63106 3666
rect 63486 3286 63516 3666
rect 63076 3067 63516 3286
rect 63076 2981 63169 3067
rect 63255 2981 63337 3067
rect 63423 2981 63516 3067
rect 63076 1555 63516 2981
rect 63076 1469 63169 1555
rect 63255 1469 63337 1555
rect 63423 1469 63516 1555
rect 63076 712 63516 1469
rect 64316 38599 64756 38682
rect 64316 38513 64409 38599
rect 64495 38513 64577 38599
rect 64663 38513 64756 38599
rect 64316 37087 64756 38513
rect 64316 37001 64409 37087
rect 64495 37001 64577 37087
rect 64663 37001 64756 37087
rect 64316 36906 64756 37001
rect 64316 36526 64346 36906
rect 64726 36526 64756 36906
rect 64316 35575 64756 36526
rect 64316 35489 64409 35575
rect 64495 35489 64577 35575
rect 64663 35489 64756 35575
rect 64316 34063 64756 35489
rect 64316 33977 64409 34063
rect 64495 33977 64577 34063
rect 64663 33977 64756 34063
rect 64316 32906 64756 33977
rect 64316 32526 64346 32906
rect 64726 32526 64756 32906
rect 64316 32465 64409 32526
rect 64495 32465 64577 32526
rect 64663 32465 64756 32526
rect 64316 31039 64756 32465
rect 64316 30953 64409 31039
rect 64495 30953 64577 31039
rect 64663 30953 64756 31039
rect 64316 29527 64756 30953
rect 64316 29441 64409 29527
rect 64495 29441 64577 29527
rect 64663 29441 64756 29527
rect 64316 28906 64756 29441
rect 64316 28526 64346 28906
rect 64726 28526 64756 28906
rect 64316 28015 64756 28526
rect 64316 27929 64409 28015
rect 64495 27929 64577 28015
rect 64663 27929 64756 28015
rect 64316 26503 64756 27929
rect 64316 26417 64409 26503
rect 64495 26417 64577 26503
rect 64663 26417 64756 26503
rect 64316 24991 64756 26417
rect 64316 24906 64409 24991
rect 64495 24906 64577 24991
rect 64663 24906 64756 24991
rect 64316 24526 64346 24906
rect 64726 24526 64756 24906
rect 64316 23479 64756 24526
rect 64316 23393 64409 23479
rect 64495 23393 64577 23479
rect 64663 23393 64756 23479
rect 64316 21967 64756 23393
rect 64316 21881 64409 21967
rect 64495 21881 64577 21967
rect 64663 21881 64756 21967
rect 64316 20906 64756 21881
rect 64316 20526 64346 20906
rect 64726 20526 64756 20906
rect 64316 20455 64756 20526
rect 64316 20369 64409 20455
rect 64495 20369 64577 20455
rect 64663 20369 64756 20455
rect 64316 18943 64756 20369
rect 64316 18857 64409 18943
rect 64495 18857 64577 18943
rect 64663 18857 64756 18943
rect 64316 17431 64756 18857
rect 64316 17345 64409 17431
rect 64495 17345 64577 17431
rect 64663 17345 64756 17431
rect 64316 16906 64756 17345
rect 64316 16526 64346 16906
rect 64726 16526 64756 16906
rect 64316 15919 64756 16526
rect 64316 15833 64409 15919
rect 64495 15833 64577 15919
rect 64663 15833 64756 15919
rect 64316 14407 64756 15833
rect 64316 14321 64409 14407
rect 64495 14321 64577 14407
rect 64663 14321 64756 14407
rect 64316 12906 64756 14321
rect 64316 12526 64346 12906
rect 64726 12526 64756 12906
rect 64316 11383 64756 12526
rect 64316 11297 64409 11383
rect 64495 11297 64577 11383
rect 64663 11297 64756 11383
rect 64316 9871 64756 11297
rect 64316 9785 64409 9871
rect 64495 9785 64577 9871
rect 64663 9785 64756 9871
rect 64316 8906 64756 9785
rect 64316 8526 64346 8906
rect 64726 8526 64756 8906
rect 64316 8359 64756 8526
rect 64316 8273 64409 8359
rect 64495 8273 64577 8359
rect 64663 8273 64756 8359
rect 64316 6847 64756 8273
rect 64316 6761 64409 6847
rect 64495 6761 64577 6847
rect 64663 6761 64756 6847
rect 64316 5335 64756 6761
rect 64316 5249 64409 5335
rect 64495 5249 64577 5335
rect 64663 5249 64756 5335
rect 64316 4906 64756 5249
rect 64316 4526 64346 4906
rect 64726 4526 64756 4906
rect 64316 3823 64756 4526
rect 64316 3737 64409 3823
rect 64495 3737 64577 3823
rect 64663 3737 64756 3823
rect 64316 2311 64756 3737
rect 64316 2225 64409 2311
rect 64495 2225 64577 2311
rect 64663 2225 64756 2311
rect 64316 799 64756 2225
rect 64316 713 64409 799
rect 64495 713 64577 799
rect 64663 713 64756 799
rect 64316 630 64756 713
rect 67076 37843 67516 38600
rect 67076 37757 67169 37843
rect 67255 37757 67337 37843
rect 67423 37757 67516 37843
rect 67076 36331 67516 37757
rect 67076 36245 67169 36331
rect 67255 36245 67337 36331
rect 67423 36245 67516 36331
rect 67076 35666 67516 36245
rect 67076 35286 67106 35666
rect 67486 35286 67516 35666
rect 67076 34819 67516 35286
rect 67076 34733 67169 34819
rect 67255 34733 67337 34819
rect 67423 34733 67516 34819
rect 67076 33307 67516 34733
rect 67076 33221 67169 33307
rect 67255 33221 67337 33307
rect 67423 33221 67516 33307
rect 67076 31795 67516 33221
rect 67076 31709 67169 31795
rect 67255 31709 67337 31795
rect 67423 31709 67516 31795
rect 67076 31666 67516 31709
rect 67076 31286 67106 31666
rect 67486 31286 67516 31666
rect 67076 30283 67516 31286
rect 67076 30197 67169 30283
rect 67255 30197 67337 30283
rect 67423 30197 67516 30283
rect 67076 28771 67516 30197
rect 67076 28685 67169 28771
rect 67255 28685 67337 28771
rect 67423 28685 67516 28771
rect 67076 27666 67516 28685
rect 67076 27286 67106 27666
rect 67486 27286 67516 27666
rect 67076 27259 67516 27286
rect 67076 27173 67169 27259
rect 67255 27173 67337 27259
rect 67423 27173 67516 27259
rect 67076 25747 67516 27173
rect 67076 25661 67169 25747
rect 67255 25661 67337 25747
rect 67423 25661 67516 25747
rect 67076 24235 67516 25661
rect 67076 24149 67169 24235
rect 67255 24149 67337 24235
rect 67423 24149 67516 24235
rect 67076 23666 67516 24149
rect 67076 23286 67106 23666
rect 67486 23286 67516 23666
rect 67076 22723 67516 23286
rect 67076 22637 67169 22723
rect 67255 22637 67337 22723
rect 67423 22637 67516 22723
rect 67076 21211 67516 22637
rect 67076 21125 67169 21211
rect 67255 21125 67337 21211
rect 67423 21125 67516 21211
rect 67076 19699 67516 21125
rect 67076 19666 67169 19699
rect 67255 19666 67337 19699
rect 67423 19666 67516 19699
rect 67076 19286 67106 19666
rect 67486 19286 67516 19666
rect 67076 18187 67516 19286
rect 67076 18101 67169 18187
rect 67255 18101 67337 18187
rect 67423 18101 67516 18187
rect 67076 16675 67516 18101
rect 67076 16589 67169 16675
rect 67255 16589 67337 16675
rect 67423 16589 67516 16675
rect 67076 15666 67516 16589
rect 67076 15286 67106 15666
rect 67486 15286 67516 15666
rect 67076 15163 67516 15286
rect 67076 15077 67169 15163
rect 67255 15077 67337 15163
rect 67423 15077 67516 15163
rect 67076 13651 67516 15077
rect 67076 13565 67169 13651
rect 67255 13565 67337 13651
rect 67423 13565 67516 13651
rect 67076 12139 67516 13565
rect 67076 12053 67169 12139
rect 67255 12053 67337 12139
rect 67423 12053 67516 12139
rect 67076 11666 67516 12053
rect 67076 11286 67106 11666
rect 67486 11286 67516 11666
rect 67076 10627 67516 11286
rect 67076 10541 67169 10627
rect 67255 10541 67337 10627
rect 67423 10541 67516 10627
rect 67076 9115 67516 10541
rect 67076 9029 67169 9115
rect 67255 9029 67337 9115
rect 67423 9029 67516 9115
rect 67076 7666 67516 9029
rect 67076 7286 67106 7666
rect 67486 7286 67516 7666
rect 67076 6091 67516 7286
rect 67076 6005 67169 6091
rect 67255 6005 67337 6091
rect 67423 6005 67516 6091
rect 67076 4579 67516 6005
rect 67076 4493 67169 4579
rect 67255 4493 67337 4579
rect 67423 4493 67516 4579
rect 67076 3666 67516 4493
rect 67076 3286 67106 3666
rect 67486 3286 67516 3666
rect 67076 3067 67516 3286
rect 67076 2981 67169 3067
rect 67255 2981 67337 3067
rect 67423 2981 67516 3067
rect 67076 1555 67516 2981
rect 67076 1469 67169 1555
rect 67255 1469 67337 1555
rect 67423 1469 67516 1555
rect 67076 712 67516 1469
rect 68316 38599 68756 38682
rect 68316 38513 68409 38599
rect 68495 38513 68577 38599
rect 68663 38513 68756 38599
rect 68316 37087 68756 38513
rect 68316 37001 68409 37087
rect 68495 37001 68577 37087
rect 68663 37001 68756 37087
rect 68316 36906 68756 37001
rect 68316 36526 68346 36906
rect 68726 36526 68756 36906
rect 68316 35575 68756 36526
rect 68316 35489 68409 35575
rect 68495 35489 68577 35575
rect 68663 35489 68756 35575
rect 68316 34063 68756 35489
rect 68316 33977 68409 34063
rect 68495 33977 68577 34063
rect 68663 33977 68756 34063
rect 68316 32906 68756 33977
rect 68316 32526 68346 32906
rect 68726 32526 68756 32906
rect 68316 32465 68409 32526
rect 68495 32465 68577 32526
rect 68663 32465 68756 32526
rect 68316 31039 68756 32465
rect 68316 30953 68409 31039
rect 68495 30953 68577 31039
rect 68663 30953 68756 31039
rect 68316 29527 68756 30953
rect 68316 29441 68409 29527
rect 68495 29441 68577 29527
rect 68663 29441 68756 29527
rect 68316 28906 68756 29441
rect 68316 28526 68346 28906
rect 68726 28526 68756 28906
rect 68316 28015 68756 28526
rect 68316 27929 68409 28015
rect 68495 27929 68577 28015
rect 68663 27929 68756 28015
rect 68316 26503 68756 27929
rect 68316 26417 68409 26503
rect 68495 26417 68577 26503
rect 68663 26417 68756 26503
rect 68316 24991 68756 26417
rect 68316 24906 68409 24991
rect 68495 24906 68577 24991
rect 68663 24906 68756 24991
rect 68316 24526 68346 24906
rect 68726 24526 68756 24906
rect 68316 23479 68756 24526
rect 68316 23393 68409 23479
rect 68495 23393 68577 23479
rect 68663 23393 68756 23479
rect 68316 21967 68756 23393
rect 68316 21881 68409 21967
rect 68495 21881 68577 21967
rect 68663 21881 68756 21967
rect 68316 20906 68756 21881
rect 68316 20526 68346 20906
rect 68726 20526 68756 20906
rect 68316 20455 68756 20526
rect 68316 20369 68409 20455
rect 68495 20369 68577 20455
rect 68663 20369 68756 20455
rect 68316 18943 68756 20369
rect 68316 18857 68409 18943
rect 68495 18857 68577 18943
rect 68663 18857 68756 18943
rect 68316 17431 68756 18857
rect 68316 17345 68409 17431
rect 68495 17345 68577 17431
rect 68663 17345 68756 17431
rect 68316 16906 68756 17345
rect 68316 16526 68346 16906
rect 68726 16526 68756 16906
rect 68316 15919 68756 16526
rect 68316 15833 68409 15919
rect 68495 15833 68577 15919
rect 68663 15833 68756 15919
rect 68316 14407 68756 15833
rect 68316 14321 68409 14407
rect 68495 14321 68577 14407
rect 68663 14321 68756 14407
rect 68316 12906 68756 14321
rect 68316 12526 68346 12906
rect 68726 12526 68756 12906
rect 68316 11383 68756 12526
rect 68316 11297 68409 11383
rect 68495 11297 68577 11383
rect 68663 11297 68756 11383
rect 68316 9871 68756 11297
rect 68316 9785 68409 9871
rect 68495 9785 68577 9871
rect 68663 9785 68756 9871
rect 68316 8906 68756 9785
rect 68316 8526 68346 8906
rect 68726 8526 68756 8906
rect 68316 8359 68756 8526
rect 68316 8273 68409 8359
rect 68495 8273 68577 8359
rect 68663 8273 68756 8359
rect 68316 6847 68756 8273
rect 68316 6761 68409 6847
rect 68495 6761 68577 6847
rect 68663 6761 68756 6847
rect 68316 5335 68756 6761
rect 68316 5249 68409 5335
rect 68495 5249 68577 5335
rect 68663 5249 68756 5335
rect 68316 4906 68756 5249
rect 68316 4526 68346 4906
rect 68726 4526 68756 4906
rect 68316 3823 68756 4526
rect 68316 3737 68409 3823
rect 68495 3737 68577 3823
rect 68663 3737 68756 3823
rect 68316 2311 68756 3737
rect 68316 2225 68409 2311
rect 68495 2225 68577 2311
rect 68663 2225 68756 2311
rect 68316 799 68756 2225
rect 68316 713 68409 799
rect 68495 713 68577 799
rect 68663 713 68756 799
rect 68316 630 68756 713
rect 71076 37843 71516 38600
rect 71076 37757 71169 37843
rect 71255 37757 71337 37843
rect 71423 37757 71516 37843
rect 71076 36331 71516 37757
rect 71076 36245 71169 36331
rect 71255 36245 71337 36331
rect 71423 36245 71516 36331
rect 71076 35666 71516 36245
rect 71076 35286 71106 35666
rect 71486 35286 71516 35666
rect 71076 34819 71516 35286
rect 71076 34733 71169 34819
rect 71255 34733 71337 34819
rect 71423 34733 71516 34819
rect 71076 31666 71516 34733
rect 71076 31286 71106 31666
rect 71486 31286 71516 31666
rect 71076 27666 71516 31286
rect 71076 27286 71106 27666
rect 71486 27286 71516 27666
rect 71076 23666 71516 27286
rect 71076 23286 71106 23666
rect 71486 23286 71516 23666
rect 71076 22723 71516 23286
rect 71076 22637 71169 22723
rect 71255 22637 71337 22723
rect 71423 22637 71516 22723
rect 71076 21211 71516 22637
rect 71076 21125 71169 21211
rect 71255 21125 71337 21211
rect 71423 21125 71516 21211
rect 71076 19699 71516 21125
rect 71076 19666 71169 19699
rect 71255 19666 71337 19699
rect 71423 19666 71516 19699
rect 71076 19286 71106 19666
rect 71486 19286 71516 19666
rect 71076 18187 71516 19286
rect 71076 18101 71169 18187
rect 71255 18101 71337 18187
rect 71423 18101 71516 18187
rect 71076 15666 71516 18101
rect 71076 15286 71106 15666
rect 71486 15286 71516 15666
rect 71076 11666 71516 15286
rect 71076 11286 71106 11666
rect 71486 11286 71516 11666
rect 71076 7666 71516 11286
rect 71076 7286 71106 7666
rect 71486 7286 71516 7666
rect 71076 6091 71516 7286
rect 71076 6005 71169 6091
rect 71255 6005 71337 6091
rect 71423 6005 71516 6091
rect 71076 4579 71516 6005
rect 71076 4493 71169 4579
rect 71255 4493 71337 4579
rect 71423 4493 71516 4579
rect 71076 3666 71516 4493
rect 71076 3286 71106 3666
rect 71486 3286 71516 3666
rect 71076 3067 71516 3286
rect 71076 2981 71169 3067
rect 71255 2981 71337 3067
rect 71423 2981 71516 3067
rect 71076 1555 71516 2981
rect 71076 1469 71169 1555
rect 71255 1469 71337 1555
rect 71423 1469 71516 1555
rect 71076 712 71516 1469
rect 72316 38599 72756 38682
rect 72316 38513 72409 38599
rect 72495 38513 72577 38599
rect 72663 38513 72756 38599
rect 72316 37087 72756 38513
rect 72316 37001 72409 37087
rect 72495 37001 72577 37087
rect 72663 37001 72756 37087
rect 72316 36906 72756 37001
rect 72316 36526 72346 36906
rect 72726 36526 72756 36906
rect 72316 35575 72756 36526
rect 72316 35489 72409 35575
rect 72495 35489 72577 35575
rect 72663 35489 72756 35575
rect 72316 34063 72756 35489
rect 72316 33977 72409 34063
rect 72495 33977 72577 34063
rect 72663 33977 72756 34063
rect 72316 32906 72756 33977
rect 72316 32526 72346 32906
rect 72726 32526 72756 32906
rect 72316 31122 72756 32526
rect 72316 31036 72409 31122
rect 72495 31036 72577 31122
rect 72663 31036 72756 31122
rect 72316 30954 72756 31036
rect 72316 30868 72409 30954
rect 72495 30868 72577 30954
rect 72663 30868 72756 30954
rect 72316 30786 72756 30868
rect 72316 30700 72409 30786
rect 72495 30700 72577 30786
rect 72663 30700 72756 30786
rect 72316 30618 72756 30700
rect 72316 30532 72409 30618
rect 72495 30532 72577 30618
rect 72663 30532 72756 30618
rect 72316 30450 72756 30532
rect 72316 30364 72409 30450
rect 72495 30364 72577 30450
rect 72663 30364 72756 30450
rect 72316 30282 72756 30364
rect 72316 30196 72409 30282
rect 72495 30196 72577 30282
rect 72663 30196 72756 30282
rect 72316 30114 72756 30196
rect 72316 30028 72409 30114
rect 72495 30028 72577 30114
rect 72663 30028 72756 30114
rect 72316 29946 72756 30028
rect 72316 29860 72409 29946
rect 72495 29860 72577 29946
rect 72663 29860 72756 29946
rect 72316 29778 72756 29860
rect 72316 29692 72409 29778
rect 72495 29692 72577 29778
rect 72663 29692 72756 29778
rect 72316 29610 72756 29692
rect 72316 29524 72409 29610
rect 72495 29524 72577 29610
rect 72663 29524 72756 29610
rect 72316 29442 72756 29524
rect 72316 29356 72409 29442
rect 72495 29356 72577 29442
rect 72663 29356 72756 29442
rect 72316 29274 72756 29356
rect 72316 29188 72409 29274
rect 72495 29188 72577 29274
rect 72663 29188 72756 29274
rect 72316 29106 72756 29188
rect 72316 29020 72409 29106
rect 72495 29020 72577 29106
rect 72663 29020 72756 29106
rect 72316 28906 72756 29020
rect 72316 28526 72346 28906
rect 72726 28526 72756 28906
rect 72316 24906 72756 28526
rect 72316 24526 72346 24906
rect 72726 24526 72756 24906
rect 72316 23479 72756 24526
rect 72316 23393 72409 23479
rect 72495 23393 72577 23479
rect 72663 23393 72756 23479
rect 72316 21967 72756 23393
rect 72316 21881 72409 21967
rect 72495 21881 72577 21967
rect 72663 21881 72756 21967
rect 72316 20906 72756 21881
rect 72316 20526 72346 20906
rect 72726 20526 72756 20906
rect 72316 20455 72756 20526
rect 72316 20369 72409 20455
rect 72495 20369 72577 20455
rect 72663 20369 72756 20455
rect 72316 18943 72756 20369
rect 72316 18857 72409 18943
rect 72495 18857 72577 18943
rect 72663 18857 72756 18943
rect 72316 17431 72756 18857
rect 72316 17345 72409 17431
rect 72495 17345 72577 17431
rect 72663 17345 72756 17431
rect 72316 16906 72756 17345
rect 72316 16526 72346 16906
rect 72726 16526 72756 16906
rect 72316 15122 72756 16526
rect 72316 15036 72409 15122
rect 72495 15036 72577 15122
rect 72663 15036 72756 15122
rect 72316 14954 72756 15036
rect 72316 14868 72409 14954
rect 72495 14868 72577 14954
rect 72663 14868 72756 14954
rect 72316 14786 72756 14868
rect 72316 14700 72409 14786
rect 72495 14700 72577 14786
rect 72663 14700 72756 14786
rect 72316 14618 72756 14700
rect 72316 14532 72409 14618
rect 72495 14532 72577 14618
rect 72663 14532 72756 14618
rect 72316 14450 72756 14532
rect 72316 14364 72409 14450
rect 72495 14364 72577 14450
rect 72663 14364 72756 14450
rect 72316 14282 72756 14364
rect 72316 14196 72409 14282
rect 72495 14196 72577 14282
rect 72663 14196 72756 14282
rect 72316 14114 72756 14196
rect 72316 14028 72409 14114
rect 72495 14028 72577 14114
rect 72663 14028 72756 14114
rect 72316 13946 72756 14028
rect 72316 13860 72409 13946
rect 72495 13860 72577 13946
rect 72663 13860 72756 13946
rect 72316 13778 72756 13860
rect 72316 13692 72409 13778
rect 72495 13692 72577 13778
rect 72663 13692 72756 13778
rect 72316 13610 72756 13692
rect 72316 13524 72409 13610
rect 72495 13524 72577 13610
rect 72663 13524 72756 13610
rect 72316 13442 72756 13524
rect 72316 13356 72409 13442
rect 72495 13356 72577 13442
rect 72663 13356 72756 13442
rect 72316 13274 72756 13356
rect 72316 13188 72409 13274
rect 72495 13188 72577 13274
rect 72663 13188 72756 13274
rect 72316 13106 72756 13188
rect 72316 13020 72409 13106
rect 72495 13020 72577 13106
rect 72663 13020 72756 13106
rect 72316 12906 72756 13020
rect 72316 12526 72346 12906
rect 72726 12526 72756 12906
rect 72316 8906 72756 12526
rect 72316 8526 72346 8906
rect 72726 8526 72756 8906
rect 72316 6847 72756 8526
rect 72316 6761 72409 6847
rect 72495 6761 72577 6847
rect 72663 6761 72756 6847
rect 72316 5335 72756 6761
rect 72316 5249 72409 5335
rect 72495 5249 72577 5335
rect 72663 5249 72756 5335
rect 72316 4906 72756 5249
rect 72316 4526 72346 4906
rect 72726 4526 72756 4906
rect 72316 3823 72756 4526
rect 72316 3737 72409 3823
rect 72495 3737 72577 3823
rect 72663 3737 72756 3823
rect 72316 2311 72756 3737
rect 72316 2225 72409 2311
rect 72495 2225 72577 2311
rect 72663 2225 72756 2311
rect 72316 799 72756 2225
rect 72316 713 72409 799
rect 72495 713 72577 799
rect 72663 713 72756 799
rect 72316 630 72756 713
rect 75076 37843 75516 38600
rect 75076 37757 75169 37843
rect 75255 37757 75337 37843
rect 75423 37757 75516 37843
rect 75076 36331 75516 37757
rect 75076 36245 75169 36331
rect 75255 36245 75337 36331
rect 75423 36245 75516 36331
rect 75076 35666 75516 36245
rect 75076 35286 75106 35666
rect 75486 35286 75516 35666
rect 75076 34819 75516 35286
rect 75076 34733 75169 34819
rect 75255 34733 75337 34819
rect 75423 34733 75516 34819
rect 75076 31666 75516 34733
rect 75076 31286 75106 31666
rect 75486 31286 75516 31666
rect 75076 28246 75516 31286
rect 75076 28160 75169 28246
rect 75255 28160 75337 28246
rect 75423 28160 75516 28246
rect 75076 28078 75516 28160
rect 75076 27992 75169 28078
rect 75255 27992 75337 28078
rect 75423 27992 75516 28078
rect 75076 27910 75516 27992
rect 75076 27824 75169 27910
rect 75255 27824 75337 27910
rect 75423 27824 75516 27910
rect 75076 27742 75516 27824
rect 75076 27666 75169 27742
rect 75255 27666 75337 27742
rect 75423 27666 75516 27742
rect 75076 27286 75106 27666
rect 75486 27286 75516 27666
rect 75076 27238 75516 27286
rect 75076 27152 75169 27238
rect 75255 27152 75337 27238
rect 75423 27152 75516 27238
rect 75076 27070 75516 27152
rect 75076 26984 75169 27070
rect 75255 26984 75337 27070
rect 75423 26984 75516 27070
rect 75076 26902 75516 26984
rect 75076 26816 75169 26902
rect 75255 26816 75337 26902
rect 75423 26816 75516 26902
rect 75076 26734 75516 26816
rect 75076 26648 75169 26734
rect 75255 26648 75337 26734
rect 75423 26648 75516 26734
rect 75076 26566 75516 26648
rect 75076 26480 75169 26566
rect 75255 26480 75337 26566
rect 75423 26480 75516 26566
rect 75076 26398 75516 26480
rect 75076 26312 75169 26398
rect 75255 26312 75337 26398
rect 75423 26312 75516 26398
rect 75076 26230 75516 26312
rect 75076 26144 75169 26230
rect 75255 26144 75337 26230
rect 75423 26144 75516 26230
rect 75076 23666 75516 26144
rect 75076 23286 75106 23666
rect 75486 23286 75516 23666
rect 75076 22723 75516 23286
rect 75076 22637 75169 22723
rect 75255 22637 75337 22723
rect 75423 22637 75516 22723
rect 75076 21211 75516 22637
rect 75076 21125 75169 21211
rect 75255 21125 75337 21211
rect 75423 21125 75516 21211
rect 75076 19699 75516 21125
rect 75076 19666 75169 19699
rect 75255 19666 75337 19699
rect 75423 19666 75516 19699
rect 75076 19286 75106 19666
rect 75486 19286 75516 19666
rect 75076 18187 75516 19286
rect 75076 18101 75169 18187
rect 75255 18101 75337 18187
rect 75423 18101 75516 18187
rect 75076 15666 75516 18101
rect 75076 15286 75106 15666
rect 75486 15286 75516 15666
rect 75076 12246 75516 15286
rect 75076 12160 75169 12246
rect 75255 12160 75337 12246
rect 75423 12160 75516 12246
rect 75076 12078 75516 12160
rect 75076 11992 75169 12078
rect 75255 11992 75337 12078
rect 75423 11992 75516 12078
rect 75076 11910 75516 11992
rect 75076 11824 75169 11910
rect 75255 11824 75337 11910
rect 75423 11824 75516 11910
rect 75076 11742 75516 11824
rect 75076 11666 75169 11742
rect 75255 11666 75337 11742
rect 75423 11666 75516 11742
rect 75076 11286 75106 11666
rect 75486 11286 75516 11666
rect 75076 11238 75516 11286
rect 75076 11152 75169 11238
rect 75255 11152 75337 11238
rect 75423 11152 75516 11238
rect 75076 11070 75516 11152
rect 75076 10984 75169 11070
rect 75255 10984 75337 11070
rect 75423 10984 75516 11070
rect 75076 10902 75516 10984
rect 75076 10816 75169 10902
rect 75255 10816 75337 10902
rect 75423 10816 75516 10902
rect 75076 10734 75516 10816
rect 75076 10648 75169 10734
rect 75255 10648 75337 10734
rect 75423 10648 75516 10734
rect 75076 10566 75516 10648
rect 75076 10480 75169 10566
rect 75255 10480 75337 10566
rect 75423 10480 75516 10566
rect 75076 10398 75516 10480
rect 75076 10312 75169 10398
rect 75255 10312 75337 10398
rect 75423 10312 75516 10398
rect 75076 10230 75516 10312
rect 75076 10144 75169 10230
rect 75255 10144 75337 10230
rect 75423 10144 75516 10230
rect 75076 7666 75516 10144
rect 75076 7286 75106 7666
rect 75486 7286 75516 7666
rect 75076 6091 75516 7286
rect 75076 6005 75169 6091
rect 75255 6005 75337 6091
rect 75423 6005 75516 6091
rect 75076 4579 75516 6005
rect 75076 4493 75169 4579
rect 75255 4493 75337 4579
rect 75423 4493 75516 4579
rect 75076 3666 75516 4493
rect 75076 3286 75106 3666
rect 75486 3286 75516 3666
rect 75076 3067 75516 3286
rect 75076 2981 75169 3067
rect 75255 2981 75337 3067
rect 75423 2981 75516 3067
rect 75076 1555 75516 2981
rect 75076 1469 75169 1555
rect 75255 1469 75337 1555
rect 75423 1469 75516 1555
rect 75076 712 75516 1469
rect 76316 38599 76756 38682
rect 76316 38513 76409 38599
rect 76495 38513 76577 38599
rect 76663 38513 76756 38599
rect 76316 37087 76756 38513
rect 76316 37001 76409 37087
rect 76495 37001 76577 37087
rect 76663 37001 76756 37087
rect 76316 36906 76756 37001
rect 76316 36526 76346 36906
rect 76726 36526 76756 36906
rect 76316 35575 76756 36526
rect 76316 35489 76409 35575
rect 76495 35489 76577 35575
rect 76663 35489 76756 35575
rect 76316 34063 76756 35489
rect 76316 33977 76409 34063
rect 76495 33977 76577 34063
rect 76663 33977 76756 34063
rect 76316 32906 76756 33977
rect 76316 32526 76346 32906
rect 76726 32526 76756 32906
rect 76316 31122 76756 32526
rect 76316 31036 76409 31122
rect 76495 31036 76577 31122
rect 76663 31036 76756 31122
rect 76316 30954 76756 31036
rect 76316 30868 76409 30954
rect 76495 30868 76577 30954
rect 76663 30868 76756 30954
rect 76316 30786 76756 30868
rect 76316 30700 76409 30786
rect 76495 30700 76577 30786
rect 76663 30700 76756 30786
rect 76316 30618 76756 30700
rect 76316 30532 76409 30618
rect 76495 30532 76577 30618
rect 76663 30532 76756 30618
rect 76316 30450 76756 30532
rect 76316 30364 76409 30450
rect 76495 30364 76577 30450
rect 76663 30364 76756 30450
rect 76316 30282 76756 30364
rect 76316 30196 76409 30282
rect 76495 30196 76577 30282
rect 76663 30196 76756 30282
rect 76316 30114 76756 30196
rect 76316 30028 76409 30114
rect 76495 30028 76577 30114
rect 76663 30028 76756 30114
rect 76316 29946 76756 30028
rect 76316 29860 76409 29946
rect 76495 29860 76577 29946
rect 76663 29860 76756 29946
rect 76316 29778 76756 29860
rect 76316 29692 76409 29778
rect 76495 29692 76577 29778
rect 76663 29692 76756 29778
rect 76316 29610 76756 29692
rect 76316 29524 76409 29610
rect 76495 29524 76577 29610
rect 76663 29524 76756 29610
rect 76316 29442 76756 29524
rect 76316 29356 76409 29442
rect 76495 29356 76577 29442
rect 76663 29356 76756 29442
rect 76316 29274 76756 29356
rect 76316 29188 76409 29274
rect 76495 29188 76577 29274
rect 76663 29188 76756 29274
rect 76316 29106 76756 29188
rect 76316 29020 76409 29106
rect 76495 29020 76577 29106
rect 76663 29020 76756 29106
rect 76316 28906 76756 29020
rect 76316 28526 76346 28906
rect 76726 28526 76756 28906
rect 76316 24906 76756 28526
rect 76316 24526 76346 24906
rect 76726 24526 76756 24906
rect 76316 23479 76756 24526
rect 76316 23393 76409 23479
rect 76495 23393 76577 23479
rect 76663 23393 76756 23479
rect 76316 21967 76756 23393
rect 76316 21881 76409 21967
rect 76495 21881 76577 21967
rect 76663 21881 76756 21967
rect 76316 20906 76756 21881
rect 76316 20526 76346 20906
rect 76726 20526 76756 20906
rect 76316 20455 76756 20526
rect 76316 20369 76409 20455
rect 76495 20369 76577 20455
rect 76663 20369 76756 20455
rect 76316 18943 76756 20369
rect 76316 18857 76409 18943
rect 76495 18857 76577 18943
rect 76663 18857 76756 18943
rect 76316 17431 76756 18857
rect 76316 17345 76409 17431
rect 76495 17345 76577 17431
rect 76663 17345 76756 17431
rect 76316 16906 76756 17345
rect 76316 16526 76346 16906
rect 76726 16526 76756 16906
rect 76316 15122 76756 16526
rect 76316 15036 76409 15122
rect 76495 15036 76577 15122
rect 76663 15036 76756 15122
rect 76316 14954 76756 15036
rect 76316 14868 76409 14954
rect 76495 14868 76577 14954
rect 76663 14868 76756 14954
rect 76316 14786 76756 14868
rect 76316 14700 76409 14786
rect 76495 14700 76577 14786
rect 76663 14700 76756 14786
rect 76316 14618 76756 14700
rect 76316 14532 76409 14618
rect 76495 14532 76577 14618
rect 76663 14532 76756 14618
rect 76316 14450 76756 14532
rect 76316 14364 76409 14450
rect 76495 14364 76577 14450
rect 76663 14364 76756 14450
rect 76316 14282 76756 14364
rect 76316 14196 76409 14282
rect 76495 14196 76577 14282
rect 76663 14196 76756 14282
rect 76316 14114 76756 14196
rect 76316 14028 76409 14114
rect 76495 14028 76577 14114
rect 76663 14028 76756 14114
rect 76316 13946 76756 14028
rect 76316 13860 76409 13946
rect 76495 13860 76577 13946
rect 76663 13860 76756 13946
rect 76316 13778 76756 13860
rect 76316 13692 76409 13778
rect 76495 13692 76577 13778
rect 76663 13692 76756 13778
rect 76316 13610 76756 13692
rect 76316 13524 76409 13610
rect 76495 13524 76577 13610
rect 76663 13524 76756 13610
rect 76316 13442 76756 13524
rect 76316 13356 76409 13442
rect 76495 13356 76577 13442
rect 76663 13356 76756 13442
rect 76316 13274 76756 13356
rect 76316 13188 76409 13274
rect 76495 13188 76577 13274
rect 76663 13188 76756 13274
rect 76316 13106 76756 13188
rect 76316 13020 76409 13106
rect 76495 13020 76577 13106
rect 76663 13020 76756 13106
rect 76316 12906 76756 13020
rect 76316 12526 76346 12906
rect 76726 12526 76756 12906
rect 76316 8906 76756 12526
rect 76316 8526 76346 8906
rect 76726 8526 76756 8906
rect 76316 6847 76756 8526
rect 76316 6761 76409 6847
rect 76495 6761 76577 6847
rect 76663 6761 76756 6847
rect 76316 5335 76756 6761
rect 76316 5249 76409 5335
rect 76495 5249 76577 5335
rect 76663 5249 76756 5335
rect 76316 4906 76756 5249
rect 76316 4526 76346 4906
rect 76726 4526 76756 4906
rect 76316 3823 76756 4526
rect 76316 3737 76409 3823
rect 76495 3737 76577 3823
rect 76663 3737 76756 3823
rect 76316 2311 76756 3737
rect 76316 2225 76409 2311
rect 76495 2225 76577 2311
rect 76663 2225 76756 2311
rect 76316 799 76756 2225
rect 76316 713 76409 799
rect 76495 713 76577 799
rect 76663 713 76756 799
rect 76316 630 76756 713
rect 79076 37843 79516 38600
rect 79076 37757 79169 37843
rect 79255 37757 79337 37843
rect 79423 37757 79516 37843
rect 79076 36331 79516 37757
rect 79076 36245 79169 36331
rect 79255 36245 79337 36331
rect 79423 36245 79516 36331
rect 79076 35666 79516 36245
rect 79076 35286 79106 35666
rect 79486 35286 79516 35666
rect 79076 34819 79516 35286
rect 79076 34733 79169 34819
rect 79255 34733 79337 34819
rect 79423 34733 79516 34819
rect 79076 31666 79516 34733
rect 79076 31286 79106 31666
rect 79486 31286 79516 31666
rect 79076 28246 79516 31286
rect 79076 28160 79169 28246
rect 79255 28160 79337 28246
rect 79423 28160 79516 28246
rect 79076 28078 79516 28160
rect 79076 27992 79169 28078
rect 79255 27992 79337 28078
rect 79423 27992 79516 28078
rect 79076 27910 79516 27992
rect 79076 27824 79169 27910
rect 79255 27824 79337 27910
rect 79423 27824 79516 27910
rect 79076 27742 79516 27824
rect 79076 27666 79169 27742
rect 79255 27666 79337 27742
rect 79423 27666 79516 27742
rect 79076 27286 79106 27666
rect 79486 27286 79516 27666
rect 79076 27238 79516 27286
rect 79076 27152 79169 27238
rect 79255 27152 79337 27238
rect 79423 27152 79516 27238
rect 79076 27070 79516 27152
rect 79076 26984 79169 27070
rect 79255 26984 79337 27070
rect 79423 26984 79516 27070
rect 79076 26902 79516 26984
rect 79076 26816 79169 26902
rect 79255 26816 79337 26902
rect 79423 26816 79516 26902
rect 79076 26734 79516 26816
rect 79076 26648 79169 26734
rect 79255 26648 79337 26734
rect 79423 26648 79516 26734
rect 79076 26566 79516 26648
rect 79076 26480 79169 26566
rect 79255 26480 79337 26566
rect 79423 26480 79516 26566
rect 79076 26398 79516 26480
rect 79076 26312 79169 26398
rect 79255 26312 79337 26398
rect 79423 26312 79516 26398
rect 79076 26230 79516 26312
rect 79076 26144 79169 26230
rect 79255 26144 79337 26230
rect 79423 26144 79516 26230
rect 79076 23666 79516 26144
rect 79076 23286 79106 23666
rect 79486 23286 79516 23666
rect 79076 22723 79516 23286
rect 79076 22637 79169 22723
rect 79255 22637 79337 22723
rect 79423 22637 79516 22723
rect 79076 21211 79516 22637
rect 79076 21125 79169 21211
rect 79255 21125 79337 21211
rect 79423 21125 79516 21211
rect 79076 19699 79516 21125
rect 79076 19666 79169 19699
rect 79255 19666 79337 19699
rect 79423 19666 79516 19699
rect 79076 19286 79106 19666
rect 79486 19286 79516 19666
rect 79076 18187 79516 19286
rect 79076 18101 79169 18187
rect 79255 18101 79337 18187
rect 79423 18101 79516 18187
rect 79076 15666 79516 18101
rect 79076 15286 79106 15666
rect 79486 15286 79516 15666
rect 79076 12246 79516 15286
rect 79076 12160 79169 12246
rect 79255 12160 79337 12246
rect 79423 12160 79516 12246
rect 79076 12078 79516 12160
rect 79076 11992 79169 12078
rect 79255 11992 79337 12078
rect 79423 11992 79516 12078
rect 79076 11910 79516 11992
rect 79076 11824 79169 11910
rect 79255 11824 79337 11910
rect 79423 11824 79516 11910
rect 79076 11742 79516 11824
rect 79076 11666 79169 11742
rect 79255 11666 79337 11742
rect 79423 11666 79516 11742
rect 79076 11286 79106 11666
rect 79486 11286 79516 11666
rect 79076 11238 79516 11286
rect 79076 11152 79169 11238
rect 79255 11152 79337 11238
rect 79423 11152 79516 11238
rect 79076 11070 79516 11152
rect 79076 10984 79169 11070
rect 79255 10984 79337 11070
rect 79423 10984 79516 11070
rect 79076 10902 79516 10984
rect 79076 10816 79169 10902
rect 79255 10816 79337 10902
rect 79423 10816 79516 10902
rect 79076 10734 79516 10816
rect 79076 10648 79169 10734
rect 79255 10648 79337 10734
rect 79423 10648 79516 10734
rect 79076 10566 79516 10648
rect 79076 10480 79169 10566
rect 79255 10480 79337 10566
rect 79423 10480 79516 10566
rect 79076 10398 79516 10480
rect 79076 10312 79169 10398
rect 79255 10312 79337 10398
rect 79423 10312 79516 10398
rect 79076 10230 79516 10312
rect 79076 10144 79169 10230
rect 79255 10144 79337 10230
rect 79423 10144 79516 10230
rect 79076 7666 79516 10144
rect 79076 7286 79106 7666
rect 79486 7286 79516 7666
rect 79076 6091 79516 7286
rect 79076 6005 79169 6091
rect 79255 6005 79337 6091
rect 79423 6005 79516 6091
rect 79076 4579 79516 6005
rect 79076 4493 79169 4579
rect 79255 4493 79337 4579
rect 79423 4493 79516 4579
rect 79076 3666 79516 4493
rect 79076 3286 79106 3666
rect 79486 3286 79516 3666
rect 79076 3067 79516 3286
rect 79076 2981 79169 3067
rect 79255 2981 79337 3067
rect 79423 2981 79516 3067
rect 79076 1555 79516 2981
rect 79076 1469 79169 1555
rect 79255 1469 79337 1555
rect 79423 1469 79516 1555
rect 79076 712 79516 1469
rect 80316 38599 80756 38682
rect 80316 38513 80409 38599
rect 80495 38513 80577 38599
rect 80663 38513 80756 38599
rect 80316 37087 80756 38513
rect 80316 37001 80409 37087
rect 80495 37001 80577 37087
rect 80663 37001 80756 37087
rect 80316 36906 80756 37001
rect 80316 36526 80346 36906
rect 80726 36526 80756 36906
rect 80316 35575 80756 36526
rect 80316 35489 80409 35575
rect 80495 35489 80577 35575
rect 80663 35489 80756 35575
rect 80316 34063 80756 35489
rect 80316 33977 80409 34063
rect 80495 33977 80577 34063
rect 80663 33977 80756 34063
rect 80316 32906 80756 33977
rect 80316 32526 80346 32906
rect 80726 32526 80756 32906
rect 80316 31122 80756 32526
rect 80316 31036 80409 31122
rect 80495 31036 80577 31122
rect 80663 31036 80756 31122
rect 80316 30954 80756 31036
rect 80316 30868 80409 30954
rect 80495 30868 80577 30954
rect 80663 30868 80756 30954
rect 80316 30786 80756 30868
rect 80316 30700 80409 30786
rect 80495 30700 80577 30786
rect 80663 30700 80756 30786
rect 80316 30618 80756 30700
rect 80316 30532 80409 30618
rect 80495 30532 80577 30618
rect 80663 30532 80756 30618
rect 80316 30450 80756 30532
rect 80316 30364 80409 30450
rect 80495 30364 80577 30450
rect 80663 30364 80756 30450
rect 80316 30282 80756 30364
rect 80316 30196 80409 30282
rect 80495 30196 80577 30282
rect 80663 30196 80756 30282
rect 80316 30114 80756 30196
rect 80316 30028 80409 30114
rect 80495 30028 80577 30114
rect 80663 30028 80756 30114
rect 80316 29946 80756 30028
rect 80316 29860 80409 29946
rect 80495 29860 80577 29946
rect 80663 29860 80756 29946
rect 80316 29778 80756 29860
rect 80316 29692 80409 29778
rect 80495 29692 80577 29778
rect 80663 29692 80756 29778
rect 80316 29610 80756 29692
rect 80316 29524 80409 29610
rect 80495 29524 80577 29610
rect 80663 29524 80756 29610
rect 80316 29442 80756 29524
rect 80316 29356 80409 29442
rect 80495 29356 80577 29442
rect 80663 29356 80756 29442
rect 80316 29274 80756 29356
rect 80316 29188 80409 29274
rect 80495 29188 80577 29274
rect 80663 29188 80756 29274
rect 80316 29106 80756 29188
rect 80316 29020 80409 29106
rect 80495 29020 80577 29106
rect 80663 29020 80756 29106
rect 80316 28906 80756 29020
rect 80316 28526 80346 28906
rect 80726 28526 80756 28906
rect 80316 24906 80756 28526
rect 80316 24526 80346 24906
rect 80726 24526 80756 24906
rect 80316 23479 80756 24526
rect 80316 23393 80409 23479
rect 80495 23393 80577 23479
rect 80663 23393 80756 23479
rect 80316 21967 80756 23393
rect 80316 21881 80409 21967
rect 80495 21881 80577 21967
rect 80663 21881 80756 21967
rect 80316 20906 80756 21881
rect 80316 20526 80346 20906
rect 80726 20526 80756 20906
rect 80316 20455 80756 20526
rect 80316 20369 80409 20455
rect 80495 20369 80577 20455
rect 80663 20369 80756 20455
rect 80316 18943 80756 20369
rect 80316 18857 80409 18943
rect 80495 18857 80577 18943
rect 80663 18857 80756 18943
rect 80316 17431 80756 18857
rect 80316 17345 80409 17431
rect 80495 17345 80577 17431
rect 80663 17345 80756 17431
rect 80316 16906 80756 17345
rect 80316 16526 80346 16906
rect 80726 16526 80756 16906
rect 80316 15122 80756 16526
rect 80316 15036 80409 15122
rect 80495 15036 80577 15122
rect 80663 15036 80756 15122
rect 80316 14954 80756 15036
rect 80316 14868 80409 14954
rect 80495 14868 80577 14954
rect 80663 14868 80756 14954
rect 80316 14786 80756 14868
rect 80316 14700 80409 14786
rect 80495 14700 80577 14786
rect 80663 14700 80756 14786
rect 80316 14618 80756 14700
rect 80316 14532 80409 14618
rect 80495 14532 80577 14618
rect 80663 14532 80756 14618
rect 80316 14450 80756 14532
rect 80316 14364 80409 14450
rect 80495 14364 80577 14450
rect 80663 14364 80756 14450
rect 80316 14282 80756 14364
rect 80316 14196 80409 14282
rect 80495 14196 80577 14282
rect 80663 14196 80756 14282
rect 80316 14114 80756 14196
rect 80316 14028 80409 14114
rect 80495 14028 80577 14114
rect 80663 14028 80756 14114
rect 80316 13946 80756 14028
rect 80316 13860 80409 13946
rect 80495 13860 80577 13946
rect 80663 13860 80756 13946
rect 80316 13778 80756 13860
rect 80316 13692 80409 13778
rect 80495 13692 80577 13778
rect 80663 13692 80756 13778
rect 80316 13610 80756 13692
rect 80316 13524 80409 13610
rect 80495 13524 80577 13610
rect 80663 13524 80756 13610
rect 80316 13442 80756 13524
rect 80316 13356 80409 13442
rect 80495 13356 80577 13442
rect 80663 13356 80756 13442
rect 80316 13274 80756 13356
rect 80316 13188 80409 13274
rect 80495 13188 80577 13274
rect 80663 13188 80756 13274
rect 80316 13106 80756 13188
rect 80316 13020 80409 13106
rect 80495 13020 80577 13106
rect 80663 13020 80756 13106
rect 80316 12906 80756 13020
rect 80316 12526 80346 12906
rect 80726 12526 80756 12906
rect 80316 8906 80756 12526
rect 80316 8526 80346 8906
rect 80726 8526 80756 8906
rect 80316 6847 80756 8526
rect 80316 6761 80409 6847
rect 80495 6761 80577 6847
rect 80663 6761 80756 6847
rect 80316 5335 80756 6761
rect 80316 5249 80409 5335
rect 80495 5249 80577 5335
rect 80663 5249 80756 5335
rect 80316 4906 80756 5249
rect 80316 4526 80346 4906
rect 80726 4526 80756 4906
rect 80316 3823 80756 4526
rect 80316 3737 80409 3823
rect 80495 3737 80577 3823
rect 80663 3737 80756 3823
rect 80316 2311 80756 3737
rect 80316 2225 80409 2311
rect 80495 2225 80577 2311
rect 80663 2225 80756 2311
rect 80316 799 80756 2225
rect 80316 713 80409 799
rect 80495 713 80577 799
rect 80663 713 80756 799
rect 80316 630 80756 713
rect 83076 37843 83516 38600
rect 83076 37757 83169 37843
rect 83255 37757 83337 37843
rect 83423 37757 83516 37843
rect 83076 36331 83516 37757
rect 83076 36245 83169 36331
rect 83255 36245 83337 36331
rect 83423 36245 83516 36331
rect 83076 35666 83516 36245
rect 83076 35286 83106 35666
rect 83486 35286 83516 35666
rect 83076 34819 83516 35286
rect 83076 34733 83169 34819
rect 83255 34733 83337 34819
rect 83423 34733 83516 34819
rect 83076 31666 83516 34733
rect 83076 31286 83106 31666
rect 83486 31286 83516 31666
rect 83076 28246 83516 31286
rect 83076 28160 83169 28246
rect 83255 28160 83337 28246
rect 83423 28160 83516 28246
rect 83076 28078 83516 28160
rect 83076 27992 83169 28078
rect 83255 27992 83337 28078
rect 83423 27992 83516 28078
rect 83076 27910 83516 27992
rect 83076 27824 83169 27910
rect 83255 27824 83337 27910
rect 83423 27824 83516 27910
rect 83076 27742 83516 27824
rect 83076 27666 83169 27742
rect 83255 27666 83337 27742
rect 83423 27666 83516 27742
rect 83076 27286 83106 27666
rect 83486 27286 83516 27666
rect 83076 27238 83516 27286
rect 83076 27152 83169 27238
rect 83255 27152 83337 27238
rect 83423 27152 83516 27238
rect 83076 27070 83516 27152
rect 83076 26984 83169 27070
rect 83255 26984 83337 27070
rect 83423 26984 83516 27070
rect 83076 26902 83516 26984
rect 83076 26816 83169 26902
rect 83255 26816 83337 26902
rect 83423 26816 83516 26902
rect 83076 26734 83516 26816
rect 83076 26648 83169 26734
rect 83255 26648 83337 26734
rect 83423 26648 83516 26734
rect 83076 26566 83516 26648
rect 83076 26480 83169 26566
rect 83255 26480 83337 26566
rect 83423 26480 83516 26566
rect 83076 26398 83516 26480
rect 83076 26312 83169 26398
rect 83255 26312 83337 26398
rect 83423 26312 83516 26398
rect 83076 26230 83516 26312
rect 83076 26144 83169 26230
rect 83255 26144 83337 26230
rect 83423 26144 83516 26230
rect 83076 23666 83516 26144
rect 83076 23286 83106 23666
rect 83486 23286 83516 23666
rect 83076 22723 83516 23286
rect 83076 22637 83169 22723
rect 83255 22637 83337 22723
rect 83423 22637 83516 22723
rect 83076 21211 83516 22637
rect 83076 21125 83169 21211
rect 83255 21125 83337 21211
rect 83423 21125 83516 21211
rect 83076 19699 83516 21125
rect 83076 19666 83169 19699
rect 83255 19666 83337 19699
rect 83423 19666 83516 19699
rect 83076 19286 83106 19666
rect 83486 19286 83516 19666
rect 83076 18187 83516 19286
rect 83076 18101 83169 18187
rect 83255 18101 83337 18187
rect 83423 18101 83516 18187
rect 83076 15666 83516 18101
rect 83076 15286 83106 15666
rect 83486 15286 83516 15666
rect 83076 12246 83516 15286
rect 83076 12160 83169 12246
rect 83255 12160 83337 12246
rect 83423 12160 83516 12246
rect 83076 12078 83516 12160
rect 83076 11992 83169 12078
rect 83255 11992 83337 12078
rect 83423 11992 83516 12078
rect 83076 11910 83516 11992
rect 83076 11824 83169 11910
rect 83255 11824 83337 11910
rect 83423 11824 83516 11910
rect 83076 11742 83516 11824
rect 83076 11666 83169 11742
rect 83255 11666 83337 11742
rect 83423 11666 83516 11742
rect 83076 11286 83106 11666
rect 83486 11286 83516 11666
rect 83076 11238 83516 11286
rect 83076 11152 83169 11238
rect 83255 11152 83337 11238
rect 83423 11152 83516 11238
rect 83076 11070 83516 11152
rect 83076 10984 83169 11070
rect 83255 10984 83337 11070
rect 83423 10984 83516 11070
rect 83076 10902 83516 10984
rect 83076 10816 83169 10902
rect 83255 10816 83337 10902
rect 83423 10816 83516 10902
rect 83076 10734 83516 10816
rect 83076 10648 83169 10734
rect 83255 10648 83337 10734
rect 83423 10648 83516 10734
rect 83076 10566 83516 10648
rect 83076 10480 83169 10566
rect 83255 10480 83337 10566
rect 83423 10480 83516 10566
rect 83076 10398 83516 10480
rect 83076 10312 83169 10398
rect 83255 10312 83337 10398
rect 83423 10312 83516 10398
rect 83076 10230 83516 10312
rect 83076 10144 83169 10230
rect 83255 10144 83337 10230
rect 83423 10144 83516 10230
rect 83076 7666 83516 10144
rect 83076 7286 83106 7666
rect 83486 7286 83516 7666
rect 83076 6091 83516 7286
rect 83076 6005 83169 6091
rect 83255 6005 83337 6091
rect 83423 6005 83516 6091
rect 83076 4579 83516 6005
rect 83076 4493 83169 4579
rect 83255 4493 83337 4579
rect 83423 4493 83516 4579
rect 83076 3666 83516 4493
rect 83076 3286 83106 3666
rect 83486 3286 83516 3666
rect 83076 3067 83516 3286
rect 83076 2981 83169 3067
rect 83255 2981 83337 3067
rect 83423 2981 83516 3067
rect 83076 1555 83516 2981
rect 83076 1469 83169 1555
rect 83255 1469 83337 1555
rect 83423 1469 83516 1555
rect 83076 712 83516 1469
rect 84316 38599 84756 38682
rect 84316 38513 84409 38599
rect 84495 38513 84577 38599
rect 84663 38513 84756 38599
rect 84316 37087 84756 38513
rect 84316 37001 84409 37087
rect 84495 37001 84577 37087
rect 84663 37001 84756 37087
rect 84316 36906 84756 37001
rect 84316 36526 84346 36906
rect 84726 36526 84756 36906
rect 84316 35575 84756 36526
rect 84316 35489 84409 35575
rect 84495 35489 84577 35575
rect 84663 35489 84756 35575
rect 84316 34063 84756 35489
rect 87076 37843 87516 38600
rect 87076 37757 87169 37843
rect 87255 37757 87337 37843
rect 87423 37757 87516 37843
rect 87076 36331 87516 37757
rect 87076 36245 87169 36331
rect 87255 36245 87337 36331
rect 87423 36245 87516 36331
rect 87076 35666 87516 36245
rect 87076 35286 87106 35666
rect 87486 35286 87516 35666
rect 84316 33977 84409 34063
rect 84495 33977 84577 34063
rect 84663 33977 84756 34063
rect 84316 32906 84756 33977
rect 84316 32526 84346 32906
rect 84726 32526 84756 32906
rect 84316 31122 84756 32526
rect 84316 31036 84409 31122
rect 84495 31036 84577 31122
rect 84663 31036 84756 31122
rect 84316 30954 84756 31036
rect 84316 30868 84409 30954
rect 84495 30868 84577 30954
rect 84663 30868 84756 30954
rect 84316 30786 84756 30868
rect 84316 30700 84409 30786
rect 84495 30700 84577 30786
rect 84663 30700 84756 30786
rect 84316 30618 84756 30700
rect 84316 30532 84409 30618
rect 84495 30532 84577 30618
rect 84663 30532 84756 30618
rect 84316 30450 84756 30532
rect 84316 30364 84409 30450
rect 84495 30364 84577 30450
rect 84663 30364 84756 30450
rect 84316 30282 84756 30364
rect 84316 30196 84409 30282
rect 84495 30196 84577 30282
rect 84663 30196 84756 30282
rect 84316 30114 84756 30196
rect 84316 30028 84409 30114
rect 84495 30028 84577 30114
rect 84663 30028 84756 30114
rect 84316 29946 84756 30028
rect 84316 29860 84409 29946
rect 84495 29860 84577 29946
rect 84663 29860 84756 29946
rect 84316 29778 84756 29860
rect 84316 29692 84409 29778
rect 84495 29692 84577 29778
rect 84663 29692 84756 29778
rect 84316 29610 84756 29692
rect 84316 29524 84409 29610
rect 84495 29524 84577 29610
rect 84663 29524 84756 29610
rect 84316 29442 84756 29524
rect 84316 29356 84409 29442
rect 84495 29356 84577 29442
rect 84663 29356 84756 29442
rect 84316 29274 84756 29356
rect 84316 29188 84409 29274
rect 84495 29188 84577 29274
rect 84663 29188 84756 29274
rect 84316 29106 84756 29188
rect 84316 29020 84409 29106
rect 84495 29020 84577 29106
rect 84663 29020 84756 29106
rect 84316 28906 84756 29020
rect 84316 28526 84346 28906
rect 84726 28526 84756 28906
rect 84316 24906 84756 28526
rect 84316 24526 84346 24906
rect 84726 24526 84756 24906
rect 84316 23479 84756 24526
rect 84316 23393 84409 23479
rect 84495 23393 84577 23479
rect 84663 23393 84756 23479
rect 84316 21967 84756 23393
rect 86348 34987 86676 35108
rect 86348 34901 86469 34987
rect 86555 34901 86676 34987
rect 86348 23143 86676 34901
rect 86348 23057 86469 23143
rect 86555 23057 86676 23143
rect 86348 22936 86676 23057
rect 87076 34819 87516 35286
rect 87076 34733 87169 34819
rect 87255 34733 87337 34819
rect 87423 34733 87516 34819
rect 87076 31666 87516 34733
rect 87076 31286 87106 31666
rect 87486 31286 87516 31666
rect 87076 28246 87516 31286
rect 87076 28160 87169 28246
rect 87255 28160 87337 28246
rect 87423 28160 87516 28246
rect 87076 28078 87516 28160
rect 87076 27992 87169 28078
rect 87255 27992 87337 28078
rect 87423 27992 87516 28078
rect 87076 27910 87516 27992
rect 87076 27824 87169 27910
rect 87255 27824 87337 27910
rect 87423 27824 87516 27910
rect 87076 27742 87516 27824
rect 87076 27666 87169 27742
rect 87255 27666 87337 27742
rect 87423 27666 87516 27742
rect 87076 27286 87106 27666
rect 87486 27286 87516 27666
rect 87076 27238 87516 27286
rect 87076 27152 87169 27238
rect 87255 27152 87337 27238
rect 87423 27152 87516 27238
rect 87076 27070 87516 27152
rect 87076 26984 87169 27070
rect 87255 26984 87337 27070
rect 87423 26984 87516 27070
rect 87076 26902 87516 26984
rect 87076 26816 87169 26902
rect 87255 26816 87337 26902
rect 87423 26816 87516 26902
rect 87076 26734 87516 26816
rect 87076 26648 87169 26734
rect 87255 26648 87337 26734
rect 87423 26648 87516 26734
rect 87076 26566 87516 26648
rect 87076 26480 87169 26566
rect 87255 26480 87337 26566
rect 87423 26480 87516 26566
rect 87076 26398 87516 26480
rect 87076 26312 87169 26398
rect 87255 26312 87337 26398
rect 87423 26312 87516 26398
rect 87076 26230 87516 26312
rect 87076 26144 87169 26230
rect 87255 26144 87337 26230
rect 87423 26144 87516 26230
rect 87076 23666 87516 26144
rect 87076 23286 87106 23666
rect 87486 23286 87516 23666
rect 84316 21881 84409 21967
rect 84495 21881 84577 21967
rect 84663 21881 84756 21967
rect 84316 20906 84756 21881
rect 84316 20526 84346 20906
rect 84726 20526 84756 20906
rect 84316 20455 84756 20526
rect 84316 20369 84409 20455
rect 84495 20369 84577 20455
rect 84663 20369 84756 20455
rect 84316 18943 84756 20369
rect 87076 22723 87516 23286
rect 87076 22637 87169 22723
rect 87255 22637 87337 22723
rect 87423 22637 87516 22723
rect 87076 21211 87516 22637
rect 87076 21125 87169 21211
rect 87255 21125 87337 21211
rect 87423 21125 87516 21211
rect 87076 19699 87516 21125
rect 87076 19666 87169 19699
rect 87255 19666 87337 19699
rect 87423 19666 87516 19699
rect 84316 18857 84409 18943
rect 84495 18857 84577 18943
rect 84663 18857 84756 18943
rect 84316 17431 84756 18857
rect 84316 17345 84409 17431
rect 84495 17345 84577 17431
rect 84663 17345 84756 17431
rect 84316 16906 84756 17345
rect 84316 16526 84346 16906
rect 84726 16526 84756 16906
rect 84316 15122 84756 16526
rect 84316 15036 84409 15122
rect 84495 15036 84577 15122
rect 84663 15036 84756 15122
rect 84316 14954 84756 15036
rect 84316 14868 84409 14954
rect 84495 14868 84577 14954
rect 84663 14868 84756 14954
rect 84316 14786 84756 14868
rect 84316 14700 84409 14786
rect 84495 14700 84577 14786
rect 84663 14700 84756 14786
rect 84316 14618 84756 14700
rect 84316 14532 84409 14618
rect 84495 14532 84577 14618
rect 84663 14532 84756 14618
rect 84316 14450 84756 14532
rect 84316 14364 84409 14450
rect 84495 14364 84577 14450
rect 84663 14364 84756 14450
rect 84316 14282 84756 14364
rect 84316 14196 84409 14282
rect 84495 14196 84577 14282
rect 84663 14196 84756 14282
rect 84316 14114 84756 14196
rect 84316 14028 84409 14114
rect 84495 14028 84577 14114
rect 84663 14028 84756 14114
rect 84316 13946 84756 14028
rect 84316 13860 84409 13946
rect 84495 13860 84577 13946
rect 84663 13860 84756 13946
rect 84316 13778 84756 13860
rect 84316 13692 84409 13778
rect 84495 13692 84577 13778
rect 84663 13692 84756 13778
rect 84316 13610 84756 13692
rect 84316 13524 84409 13610
rect 84495 13524 84577 13610
rect 84663 13524 84756 13610
rect 84316 13442 84756 13524
rect 84316 13356 84409 13442
rect 84495 13356 84577 13442
rect 84663 13356 84756 13442
rect 84316 13274 84756 13356
rect 84316 13188 84409 13274
rect 84495 13188 84577 13274
rect 84663 13188 84756 13274
rect 84316 13106 84756 13188
rect 84316 13020 84409 13106
rect 84495 13020 84577 13106
rect 84663 13020 84756 13106
rect 84316 12906 84756 13020
rect 84316 12526 84346 12906
rect 84726 12526 84756 12906
rect 84316 8906 84756 12526
rect 84316 8526 84346 8906
rect 84726 8526 84756 8906
rect 84316 6847 84756 8526
rect 86348 19363 86676 19484
rect 86348 19277 86469 19363
rect 86555 19277 86676 19363
rect 86348 7435 86676 19277
rect 86348 7349 86469 7435
rect 86555 7349 86676 7435
rect 86348 7228 86676 7349
rect 87076 19286 87106 19666
rect 87486 19286 87516 19666
rect 87076 18187 87516 19286
rect 87076 18101 87169 18187
rect 87255 18101 87337 18187
rect 87423 18101 87516 18187
rect 87076 15666 87516 18101
rect 87076 15286 87106 15666
rect 87486 15286 87516 15666
rect 87076 12246 87516 15286
rect 87076 12160 87169 12246
rect 87255 12160 87337 12246
rect 87423 12160 87516 12246
rect 87076 12078 87516 12160
rect 87076 11992 87169 12078
rect 87255 11992 87337 12078
rect 87423 11992 87516 12078
rect 87076 11910 87516 11992
rect 87076 11824 87169 11910
rect 87255 11824 87337 11910
rect 87423 11824 87516 11910
rect 87076 11742 87516 11824
rect 87076 11666 87169 11742
rect 87255 11666 87337 11742
rect 87423 11666 87516 11742
rect 87076 11286 87106 11666
rect 87486 11286 87516 11666
rect 87076 11238 87516 11286
rect 87076 11152 87169 11238
rect 87255 11152 87337 11238
rect 87423 11152 87516 11238
rect 87076 11070 87516 11152
rect 87076 10984 87169 11070
rect 87255 10984 87337 11070
rect 87423 10984 87516 11070
rect 87076 10902 87516 10984
rect 87076 10816 87169 10902
rect 87255 10816 87337 10902
rect 87423 10816 87516 10902
rect 87076 10734 87516 10816
rect 87076 10648 87169 10734
rect 87255 10648 87337 10734
rect 87423 10648 87516 10734
rect 87076 10566 87516 10648
rect 87076 10480 87169 10566
rect 87255 10480 87337 10566
rect 87423 10480 87516 10566
rect 87076 10398 87516 10480
rect 87076 10312 87169 10398
rect 87255 10312 87337 10398
rect 87423 10312 87516 10398
rect 87076 10230 87516 10312
rect 87076 10144 87169 10230
rect 87255 10144 87337 10230
rect 87423 10144 87516 10230
rect 87076 7666 87516 10144
rect 87076 7286 87106 7666
rect 87486 7286 87516 7666
rect 84316 6761 84409 6847
rect 84495 6761 84577 6847
rect 84663 6761 84756 6847
rect 84316 5335 84756 6761
rect 84316 5249 84409 5335
rect 84495 5249 84577 5335
rect 84663 5249 84756 5335
rect 84316 4906 84756 5249
rect 84316 4526 84346 4906
rect 84726 4526 84756 4906
rect 84316 3823 84756 4526
rect 84316 3737 84409 3823
rect 84495 3737 84577 3823
rect 84663 3737 84756 3823
rect 84316 2311 84756 3737
rect 84316 2225 84409 2311
rect 84495 2225 84577 2311
rect 84663 2225 84756 2311
rect 84316 799 84756 2225
rect 84316 713 84409 799
rect 84495 713 84577 799
rect 84663 713 84756 799
rect 84316 630 84756 713
rect 87076 6091 87516 7286
rect 87076 6005 87169 6091
rect 87255 6005 87337 6091
rect 87423 6005 87516 6091
rect 87076 4579 87516 6005
rect 87076 4493 87169 4579
rect 87255 4493 87337 4579
rect 87423 4493 87516 4579
rect 87076 3666 87516 4493
rect 87076 3286 87106 3666
rect 87486 3286 87516 3666
rect 87076 3067 87516 3286
rect 87076 2981 87169 3067
rect 87255 2981 87337 3067
rect 87423 2981 87516 3067
rect 87076 1555 87516 2981
rect 87076 1469 87169 1555
rect 87255 1469 87337 1555
rect 87423 1469 87516 1555
rect 87076 712 87516 1469
rect 88316 38599 88756 38682
rect 88316 38513 88409 38599
rect 88495 38513 88577 38599
rect 88663 38513 88756 38599
rect 88316 37087 88756 38513
rect 88316 37001 88409 37087
rect 88495 37001 88577 37087
rect 88663 37001 88756 37087
rect 88316 36906 88756 37001
rect 88316 36526 88346 36906
rect 88726 36526 88756 36906
rect 88316 35575 88756 36526
rect 88316 35489 88409 35575
rect 88495 35489 88577 35575
rect 88663 35489 88756 35575
rect 88316 34063 88756 35489
rect 88316 33977 88409 34063
rect 88495 33977 88577 34063
rect 88663 33977 88756 34063
rect 88316 32906 88756 33977
rect 88316 32526 88346 32906
rect 88726 32526 88756 32906
rect 88316 31122 88756 32526
rect 88316 31036 88409 31122
rect 88495 31036 88577 31122
rect 88663 31036 88756 31122
rect 88316 30954 88756 31036
rect 88316 30868 88409 30954
rect 88495 30868 88577 30954
rect 88663 30868 88756 30954
rect 88316 30786 88756 30868
rect 88316 30700 88409 30786
rect 88495 30700 88577 30786
rect 88663 30700 88756 30786
rect 88316 30618 88756 30700
rect 88316 30532 88409 30618
rect 88495 30532 88577 30618
rect 88663 30532 88756 30618
rect 88316 30450 88756 30532
rect 88316 30364 88409 30450
rect 88495 30364 88577 30450
rect 88663 30364 88756 30450
rect 88316 30282 88756 30364
rect 88316 30196 88409 30282
rect 88495 30196 88577 30282
rect 88663 30196 88756 30282
rect 88316 30114 88756 30196
rect 88316 30028 88409 30114
rect 88495 30028 88577 30114
rect 88663 30028 88756 30114
rect 88316 29946 88756 30028
rect 88316 29860 88409 29946
rect 88495 29860 88577 29946
rect 88663 29860 88756 29946
rect 88316 29778 88756 29860
rect 88316 29692 88409 29778
rect 88495 29692 88577 29778
rect 88663 29692 88756 29778
rect 88316 29610 88756 29692
rect 88316 29524 88409 29610
rect 88495 29524 88577 29610
rect 88663 29524 88756 29610
rect 88316 29442 88756 29524
rect 88316 29356 88409 29442
rect 88495 29356 88577 29442
rect 88663 29356 88756 29442
rect 88316 29274 88756 29356
rect 88316 29188 88409 29274
rect 88495 29188 88577 29274
rect 88663 29188 88756 29274
rect 88316 29106 88756 29188
rect 88316 29020 88409 29106
rect 88495 29020 88577 29106
rect 88663 29020 88756 29106
rect 88316 28906 88756 29020
rect 88316 28526 88346 28906
rect 88726 28526 88756 28906
rect 88316 24906 88756 28526
rect 88316 24526 88346 24906
rect 88726 24526 88756 24906
rect 88316 23479 88756 24526
rect 88316 23393 88409 23479
rect 88495 23393 88577 23479
rect 88663 23393 88756 23479
rect 88316 21967 88756 23393
rect 88316 21881 88409 21967
rect 88495 21881 88577 21967
rect 88663 21881 88756 21967
rect 88316 20906 88756 21881
rect 88316 20526 88346 20906
rect 88726 20526 88756 20906
rect 88316 20455 88756 20526
rect 88316 20369 88409 20455
rect 88495 20369 88577 20455
rect 88663 20369 88756 20455
rect 88316 18943 88756 20369
rect 88316 18857 88409 18943
rect 88495 18857 88577 18943
rect 88663 18857 88756 18943
rect 88316 17431 88756 18857
rect 88316 17345 88409 17431
rect 88495 17345 88577 17431
rect 88663 17345 88756 17431
rect 88316 16906 88756 17345
rect 88316 16526 88346 16906
rect 88726 16526 88756 16906
rect 88316 15122 88756 16526
rect 88316 15036 88409 15122
rect 88495 15036 88577 15122
rect 88663 15036 88756 15122
rect 88316 14954 88756 15036
rect 88316 14868 88409 14954
rect 88495 14868 88577 14954
rect 88663 14868 88756 14954
rect 88316 14786 88756 14868
rect 88316 14700 88409 14786
rect 88495 14700 88577 14786
rect 88663 14700 88756 14786
rect 88316 14618 88756 14700
rect 88316 14532 88409 14618
rect 88495 14532 88577 14618
rect 88663 14532 88756 14618
rect 88316 14450 88756 14532
rect 88316 14364 88409 14450
rect 88495 14364 88577 14450
rect 88663 14364 88756 14450
rect 88316 14282 88756 14364
rect 88316 14196 88409 14282
rect 88495 14196 88577 14282
rect 88663 14196 88756 14282
rect 88316 14114 88756 14196
rect 88316 14028 88409 14114
rect 88495 14028 88577 14114
rect 88663 14028 88756 14114
rect 88316 13946 88756 14028
rect 88316 13860 88409 13946
rect 88495 13860 88577 13946
rect 88663 13860 88756 13946
rect 88316 13778 88756 13860
rect 88316 13692 88409 13778
rect 88495 13692 88577 13778
rect 88663 13692 88756 13778
rect 88316 13610 88756 13692
rect 88316 13524 88409 13610
rect 88495 13524 88577 13610
rect 88663 13524 88756 13610
rect 88316 13442 88756 13524
rect 88316 13356 88409 13442
rect 88495 13356 88577 13442
rect 88663 13356 88756 13442
rect 88316 13274 88756 13356
rect 88316 13188 88409 13274
rect 88495 13188 88577 13274
rect 88663 13188 88756 13274
rect 88316 13106 88756 13188
rect 88316 13020 88409 13106
rect 88495 13020 88577 13106
rect 88663 13020 88756 13106
rect 88316 12906 88756 13020
rect 88316 12526 88346 12906
rect 88726 12526 88756 12906
rect 88316 8906 88756 12526
rect 88316 8526 88346 8906
rect 88726 8526 88756 8906
rect 88316 6847 88756 8526
rect 88316 6761 88409 6847
rect 88495 6761 88577 6847
rect 88663 6761 88756 6847
rect 88316 5335 88756 6761
rect 88316 5249 88409 5335
rect 88495 5249 88577 5335
rect 88663 5249 88756 5335
rect 88316 4906 88756 5249
rect 88316 4526 88346 4906
rect 88726 4526 88756 4906
rect 88316 3823 88756 4526
rect 88316 3737 88409 3823
rect 88495 3737 88577 3823
rect 88663 3737 88756 3823
rect 88316 2311 88756 3737
rect 88316 2225 88409 2311
rect 88495 2225 88577 2311
rect 88663 2225 88756 2311
rect 88316 799 88756 2225
rect 88316 713 88409 799
rect 88495 713 88577 799
rect 88663 713 88756 799
rect 88316 630 88756 713
rect 91076 37843 91516 38600
rect 91076 37757 91169 37843
rect 91255 37757 91337 37843
rect 91423 37757 91516 37843
rect 91076 36331 91516 37757
rect 91076 36245 91169 36331
rect 91255 36245 91337 36331
rect 91423 36245 91516 36331
rect 91076 35666 91516 36245
rect 91076 35286 91106 35666
rect 91486 35286 91516 35666
rect 91076 34819 91516 35286
rect 91076 34733 91169 34819
rect 91255 34733 91337 34819
rect 91423 34733 91516 34819
rect 91076 31666 91516 34733
rect 91076 31286 91106 31666
rect 91486 31286 91516 31666
rect 91076 28246 91516 31286
rect 91076 28160 91169 28246
rect 91255 28160 91337 28246
rect 91423 28160 91516 28246
rect 91076 28078 91516 28160
rect 91076 27992 91169 28078
rect 91255 27992 91337 28078
rect 91423 27992 91516 28078
rect 91076 27910 91516 27992
rect 91076 27824 91169 27910
rect 91255 27824 91337 27910
rect 91423 27824 91516 27910
rect 91076 27742 91516 27824
rect 91076 27666 91169 27742
rect 91255 27666 91337 27742
rect 91423 27666 91516 27742
rect 91076 27286 91106 27666
rect 91486 27286 91516 27666
rect 91076 27238 91516 27286
rect 91076 27152 91169 27238
rect 91255 27152 91337 27238
rect 91423 27152 91516 27238
rect 91076 27070 91516 27152
rect 91076 26984 91169 27070
rect 91255 26984 91337 27070
rect 91423 26984 91516 27070
rect 91076 26902 91516 26984
rect 91076 26816 91169 26902
rect 91255 26816 91337 26902
rect 91423 26816 91516 26902
rect 91076 26734 91516 26816
rect 91076 26648 91169 26734
rect 91255 26648 91337 26734
rect 91423 26648 91516 26734
rect 91076 26566 91516 26648
rect 91076 26480 91169 26566
rect 91255 26480 91337 26566
rect 91423 26480 91516 26566
rect 91076 26398 91516 26480
rect 91076 26312 91169 26398
rect 91255 26312 91337 26398
rect 91423 26312 91516 26398
rect 91076 26230 91516 26312
rect 91076 26144 91169 26230
rect 91255 26144 91337 26230
rect 91423 26144 91516 26230
rect 91076 23666 91516 26144
rect 91076 23286 91106 23666
rect 91486 23286 91516 23666
rect 91076 22723 91516 23286
rect 91076 22637 91169 22723
rect 91255 22637 91337 22723
rect 91423 22637 91516 22723
rect 91076 21211 91516 22637
rect 91076 21125 91169 21211
rect 91255 21125 91337 21211
rect 91423 21125 91516 21211
rect 91076 19699 91516 21125
rect 91076 19666 91169 19699
rect 91255 19666 91337 19699
rect 91423 19666 91516 19699
rect 91076 19286 91106 19666
rect 91486 19286 91516 19666
rect 91076 18187 91516 19286
rect 91076 18101 91169 18187
rect 91255 18101 91337 18187
rect 91423 18101 91516 18187
rect 91076 15666 91516 18101
rect 91076 15286 91106 15666
rect 91486 15286 91516 15666
rect 91076 12246 91516 15286
rect 91076 12160 91169 12246
rect 91255 12160 91337 12246
rect 91423 12160 91516 12246
rect 91076 12078 91516 12160
rect 91076 11992 91169 12078
rect 91255 11992 91337 12078
rect 91423 11992 91516 12078
rect 91076 11910 91516 11992
rect 91076 11824 91169 11910
rect 91255 11824 91337 11910
rect 91423 11824 91516 11910
rect 91076 11742 91516 11824
rect 91076 11666 91169 11742
rect 91255 11666 91337 11742
rect 91423 11666 91516 11742
rect 91076 11286 91106 11666
rect 91486 11286 91516 11666
rect 91076 11238 91516 11286
rect 91076 11152 91169 11238
rect 91255 11152 91337 11238
rect 91423 11152 91516 11238
rect 91076 11070 91516 11152
rect 91076 10984 91169 11070
rect 91255 10984 91337 11070
rect 91423 10984 91516 11070
rect 91076 10902 91516 10984
rect 91076 10816 91169 10902
rect 91255 10816 91337 10902
rect 91423 10816 91516 10902
rect 91076 10734 91516 10816
rect 91076 10648 91169 10734
rect 91255 10648 91337 10734
rect 91423 10648 91516 10734
rect 91076 10566 91516 10648
rect 91076 10480 91169 10566
rect 91255 10480 91337 10566
rect 91423 10480 91516 10566
rect 91076 10398 91516 10480
rect 91076 10312 91169 10398
rect 91255 10312 91337 10398
rect 91423 10312 91516 10398
rect 91076 10230 91516 10312
rect 91076 10144 91169 10230
rect 91255 10144 91337 10230
rect 91423 10144 91516 10230
rect 91076 7666 91516 10144
rect 91076 7286 91106 7666
rect 91486 7286 91516 7666
rect 91076 6091 91516 7286
rect 91076 6005 91169 6091
rect 91255 6005 91337 6091
rect 91423 6005 91516 6091
rect 91076 4579 91516 6005
rect 91076 4493 91169 4579
rect 91255 4493 91337 4579
rect 91423 4493 91516 4579
rect 91076 3666 91516 4493
rect 91076 3286 91106 3666
rect 91486 3286 91516 3666
rect 91076 3067 91516 3286
rect 91076 2981 91169 3067
rect 91255 2981 91337 3067
rect 91423 2981 91516 3067
rect 91076 1555 91516 2981
rect 91076 1469 91169 1555
rect 91255 1469 91337 1555
rect 91423 1469 91516 1555
rect 91076 712 91516 1469
rect 92316 38599 92756 38682
rect 92316 38513 92409 38599
rect 92495 38513 92577 38599
rect 92663 38513 92756 38599
rect 92316 37087 92756 38513
rect 92316 37001 92409 37087
rect 92495 37001 92577 37087
rect 92663 37001 92756 37087
rect 92316 36906 92756 37001
rect 92316 36526 92346 36906
rect 92726 36526 92756 36906
rect 92316 35575 92756 36526
rect 92316 35489 92409 35575
rect 92495 35489 92577 35575
rect 92663 35489 92756 35575
rect 92316 34063 92756 35489
rect 92316 33977 92409 34063
rect 92495 33977 92577 34063
rect 92663 33977 92756 34063
rect 92316 32906 92756 33977
rect 92316 32526 92346 32906
rect 92726 32526 92756 32906
rect 92316 31122 92756 32526
rect 92316 31036 92409 31122
rect 92495 31036 92577 31122
rect 92663 31036 92756 31122
rect 92316 30954 92756 31036
rect 92316 30868 92409 30954
rect 92495 30868 92577 30954
rect 92663 30868 92756 30954
rect 92316 30786 92756 30868
rect 92316 30700 92409 30786
rect 92495 30700 92577 30786
rect 92663 30700 92756 30786
rect 92316 30618 92756 30700
rect 92316 30532 92409 30618
rect 92495 30532 92577 30618
rect 92663 30532 92756 30618
rect 92316 30450 92756 30532
rect 92316 30364 92409 30450
rect 92495 30364 92577 30450
rect 92663 30364 92756 30450
rect 92316 30282 92756 30364
rect 92316 30196 92409 30282
rect 92495 30196 92577 30282
rect 92663 30196 92756 30282
rect 92316 30114 92756 30196
rect 92316 30028 92409 30114
rect 92495 30028 92577 30114
rect 92663 30028 92756 30114
rect 92316 29946 92756 30028
rect 92316 29860 92409 29946
rect 92495 29860 92577 29946
rect 92663 29860 92756 29946
rect 92316 29778 92756 29860
rect 92316 29692 92409 29778
rect 92495 29692 92577 29778
rect 92663 29692 92756 29778
rect 92316 29610 92756 29692
rect 92316 29524 92409 29610
rect 92495 29524 92577 29610
rect 92663 29524 92756 29610
rect 92316 29442 92756 29524
rect 92316 29356 92409 29442
rect 92495 29356 92577 29442
rect 92663 29356 92756 29442
rect 92316 29274 92756 29356
rect 92316 29188 92409 29274
rect 92495 29188 92577 29274
rect 92663 29188 92756 29274
rect 92316 29106 92756 29188
rect 92316 29020 92409 29106
rect 92495 29020 92577 29106
rect 92663 29020 92756 29106
rect 92316 28906 92756 29020
rect 92316 28526 92346 28906
rect 92726 28526 92756 28906
rect 92316 24906 92756 28526
rect 92316 24526 92346 24906
rect 92726 24526 92756 24906
rect 92316 23479 92756 24526
rect 92316 23393 92409 23479
rect 92495 23393 92577 23479
rect 92663 23393 92756 23479
rect 92316 21967 92756 23393
rect 92316 21881 92409 21967
rect 92495 21881 92577 21967
rect 92663 21881 92756 21967
rect 92316 20906 92756 21881
rect 92316 20526 92346 20906
rect 92726 20526 92756 20906
rect 92316 20455 92756 20526
rect 92316 20369 92409 20455
rect 92495 20369 92577 20455
rect 92663 20369 92756 20455
rect 92316 18943 92756 20369
rect 92316 18857 92409 18943
rect 92495 18857 92577 18943
rect 92663 18857 92756 18943
rect 92316 17431 92756 18857
rect 92316 17345 92409 17431
rect 92495 17345 92577 17431
rect 92663 17345 92756 17431
rect 92316 16906 92756 17345
rect 92316 16526 92346 16906
rect 92726 16526 92756 16906
rect 92316 15122 92756 16526
rect 92316 15036 92409 15122
rect 92495 15036 92577 15122
rect 92663 15036 92756 15122
rect 92316 14954 92756 15036
rect 92316 14868 92409 14954
rect 92495 14868 92577 14954
rect 92663 14868 92756 14954
rect 92316 14786 92756 14868
rect 92316 14700 92409 14786
rect 92495 14700 92577 14786
rect 92663 14700 92756 14786
rect 92316 14618 92756 14700
rect 92316 14532 92409 14618
rect 92495 14532 92577 14618
rect 92663 14532 92756 14618
rect 92316 14450 92756 14532
rect 92316 14364 92409 14450
rect 92495 14364 92577 14450
rect 92663 14364 92756 14450
rect 92316 14282 92756 14364
rect 92316 14196 92409 14282
rect 92495 14196 92577 14282
rect 92663 14196 92756 14282
rect 92316 14114 92756 14196
rect 92316 14028 92409 14114
rect 92495 14028 92577 14114
rect 92663 14028 92756 14114
rect 92316 13946 92756 14028
rect 92316 13860 92409 13946
rect 92495 13860 92577 13946
rect 92663 13860 92756 13946
rect 92316 13778 92756 13860
rect 92316 13692 92409 13778
rect 92495 13692 92577 13778
rect 92663 13692 92756 13778
rect 92316 13610 92756 13692
rect 92316 13524 92409 13610
rect 92495 13524 92577 13610
rect 92663 13524 92756 13610
rect 92316 13442 92756 13524
rect 92316 13356 92409 13442
rect 92495 13356 92577 13442
rect 92663 13356 92756 13442
rect 92316 13274 92756 13356
rect 92316 13188 92409 13274
rect 92495 13188 92577 13274
rect 92663 13188 92756 13274
rect 92316 13106 92756 13188
rect 92316 13020 92409 13106
rect 92495 13020 92577 13106
rect 92663 13020 92756 13106
rect 92316 12906 92756 13020
rect 92316 12526 92346 12906
rect 92726 12526 92756 12906
rect 92316 8906 92756 12526
rect 92316 8526 92346 8906
rect 92726 8526 92756 8906
rect 92316 6847 92756 8526
rect 92316 6761 92409 6847
rect 92495 6761 92577 6847
rect 92663 6761 92756 6847
rect 92316 5335 92756 6761
rect 92316 5249 92409 5335
rect 92495 5249 92577 5335
rect 92663 5249 92756 5335
rect 92316 4906 92756 5249
rect 92316 4526 92346 4906
rect 92726 4526 92756 4906
rect 92316 3823 92756 4526
rect 92316 3737 92409 3823
rect 92495 3737 92577 3823
rect 92663 3737 92756 3823
rect 92316 2311 92756 3737
rect 92316 2225 92409 2311
rect 92495 2225 92577 2311
rect 92663 2225 92756 2311
rect 92316 799 92756 2225
rect 92316 713 92409 799
rect 92495 713 92577 799
rect 92663 713 92756 799
rect 92316 630 92756 713
rect 95076 37843 95516 38600
rect 95076 37757 95169 37843
rect 95255 37757 95337 37843
rect 95423 37757 95516 37843
rect 95076 36331 95516 37757
rect 95076 36245 95169 36331
rect 95255 36245 95337 36331
rect 95423 36245 95516 36331
rect 95076 35666 95516 36245
rect 95076 35286 95106 35666
rect 95486 35286 95516 35666
rect 95076 34819 95516 35286
rect 95076 34733 95169 34819
rect 95255 34733 95337 34819
rect 95423 34733 95516 34819
rect 95076 31666 95516 34733
rect 95076 31286 95106 31666
rect 95486 31286 95516 31666
rect 95076 28246 95516 31286
rect 95076 28160 95169 28246
rect 95255 28160 95337 28246
rect 95423 28160 95516 28246
rect 95076 28078 95516 28160
rect 95076 27992 95169 28078
rect 95255 27992 95337 28078
rect 95423 27992 95516 28078
rect 95076 27910 95516 27992
rect 95076 27824 95169 27910
rect 95255 27824 95337 27910
rect 95423 27824 95516 27910
rect 95076 27742 95516 27824
rect 95076 27666 95169 27742
rect 95255 27666 95337 27742
rect 95423 27666 95516 27742
rect 95076 27286 95106 27666
rect 95486 27286 95516 27666
rect 95076 27238 95516 27286
rect 95076 27152 95169 27238
rect 95255 27152 95337 27238
rect 95423 27152 95516 27238
rect 95076 27070 95516 27152
rect 95076 26984 95169 27070
rect 95255 26984 95337 27070
rect 95423 26984 95516 27070
rect 95076 26902 95516 26984
rect 95076 26816 95169 26902
rect 95255 26816 95337 26902
rect 95423 26816 95516 26902
rect 95076 26734 95516 26816
rect 95076 26648 95169 26734
rect 95255 26648 95337 26734
rect 95423 26648 95516 26734
rect 95076 26566 95516 26648
rect 95076 26480 95169 26566
rect 95255 26480 95337 26566
rect 95423 26480 95516 26566
rect 95076 26398 95516 26480
rect 95076 26312 95169 26398
rect 95255 26312 95337 26398
rect 95423 26312 95516 26398
rect 95076 26230 95516 26312
rect 95076 26144 95169 26230
rect 95255 26144 95337 26230
rect 95423 26144 95516 26230
rect 95076 23666 95516 26144
rect 95076 23286 95106 23666
rect 95486 23286 95516 23666
rect 95076 22723 95516 23286
rect 95076 22637 95169 22723
rect 95255 22637 95337 22723
rect 95423 22637 95516 22723
rect 95076 21211 95516 22637
rect 95076 21125 95169 21211
rect 95255 21125 95337 21211
rect 95423 21125 95516 21211
rect 95076 19699 95516 21125
rect 95076 19666 95169 19699
rect 95255 19666 95337 19699
rect 95423 19666 95516 19699
rect 95076 19286 95106 19666
rect 95486 19286 95516 19666
rect 95076 18187 95516 19286
rect 95076 18101 95169 18187
rect 95255 18101 95337 18187
rect 95423 18101 95516 18187
rect 95076 15666 95516 18101
rect 95076 15286 95106 15666
rect 95486 15286 95516 15666
rect 95076 12246 95516 15286
rect 95076 12160 95169 12246
rect 95255 12160 95337 12246
rect 95423 12160 95516 12246
rect 95076 12078 95516 12160
rect 95076 11992 95169 12078
rect 95255 11992 95337 12078
rect 95423 11992 95516 12078
rect 95076 11910 95516 11992
rect 95076 11824 95169 11910
rect 95255 11824 95337 11910
rect 95423 11824 95516 11910
rect 95076 11742 95516 11824
rect 95076 11666 95169 11742
rect 95255 11666 95337 11742
rect 95423 11666 95516 11742
rect 95076 11286 95106 11666
rect 95486 11286 95516 11666
rect 95076 11238 95516 11286
rect 95076 11152 95169 11238
rect 95255 11152 95337 11238
rect 95423 11152 95516 11238
rect 95076 11070 95516 11152
rect 95076 10984 95169 11070
rect 95255 10984 95337 11070
rect 95423 10984 95516 11070
rect 95076 10902 95516 10984
rect 95076 10816 95169 10902
rect 95255 10816 95337 10902
rect 95423 10816 95516 10902
rect 95076 10734 95516 10816
rect 95076 10648 95169 10734
rect 95255 10648 95337 10734
rect 95423 10648 95516 10734
rect 95076 10566 95516 10648
rect 95076 10480 95169 10566
rect 95255 10480 95337 10566
rect 95423 10480 95516 10566
rect 95076 10398 95516 10480
rect 95076 10312 95169 10398
rect 95255 10312 95337 10398
rect 95423 10312 95516 10398
rect 95076 10230 95516 10312
rect 95076 10144 95169 10230
rect 95255 10144 95337 10230
rect 95423 10144 95516 10230
rect 95076 7666 95516 10144
rect 95076 7286 95106 7666
rect 95486 7286 95516 7666
rect 95076 6091 95516 7286
rect 95076 6005 95169 6091
rect 95255 6005 95337 6091
rect 95423 6005 95516 6091
rect 95076 4579 95516 6005
rect 95076 4493 95169 4579
rect 95255 4493 95337 4579
rect 95423 4493 95516 4579
rect 95076 3666 95516 4493
rect 95076 3286 95106 3666
rect 95486 3286 95516 3666
rect 95076 3067 95516 3286
rect 95076 2981 95169 3067
rect 95255 2981 95337 3067
rect 95423 2981 95516 3067
rect 95076 1555 95516 2981
rect 95076 1469 95169 1555
rect 95255 1469 95337 1555
rect 95423 1469 95516 1555
rect 95076 712 95516 1469
rect 96316 38599 96756 38682
rect 96316 38513 96409 38599
rect 96495 38513 96577 38599
rect 96663 38513 96756 38599
rect 96316 37087 96756 38513
rect 96316 37001 96409 37087
rect 96495 37001 96577 37087
rect 96663 37001 96756 37087
rect 96316 36906 96756 37001
rect 96316 36526 96346 36906
rect 96726 36526 96756 36906
rect 96316 35575 96756 36526
rect 96316 35489 96409 35575
rect 96495 35489 96577 35575
rect 96663 35489 96756 35575
rect 96316 34063 96756 35489
rect 96316 33977 96409 34063
rect 96495 33977 96577 34063
rect 96663 33977 96756 34063
rect 96316 32906 96756 33977
rect 96316 32526 96346 32906
rect 96726 32526 96756 32906
rect 96316 31122 96756 32526
rect 96316 31036 96409 31122
rect 96495 31036 96577 31122
rect 96663 31036 96756 31122
rect 96316 30954 96756 31036
rect 96316 30868 96409 30954
rect 96495 30868 96577 30954
rect 96663 30868 96756 30954
rect 96316 30786 96756 30868
rect 96316 30700 96409 30786
rect 96495 30700 96577 30786
rect 96663 30700 96756 30786
rect 96316 30618 96756 30700
rect 96316 30532 96409 30618
rect 96495 30532 96577 30618
rect 96663 30532 96756 30618
rect 96316 30450 96756 30532
rect 96316 30364 96409 30450
rect 96495 30364 96577 30450
rect 96663 30364 96756 30450
rect 96316 30282 96756 30364
rect 96316 30196 96409 30282
rect 96495 30196 96577 30282
rect 96663 30196 96756 30282
rect 96316 30114 96756 30196
rect 96316 30028 96409 30114
rect 96495 30028 96577 30114
rect 96663 30028 96756 30114
rect 96316 29946 96756 30028
rect 96316 29860 96409 29946
rect 96495 29860 96577 29946
rect 96663 29860 96756 29946
rect 96316 29778 96756 29860
rect 96316 29692 96409 29778
rect 96495 29692 96577 29778
rect 96663 29692 96756 29778
rect 96316 29610 96756 29692
rect 96316 29524 96409 29610
rect 96495 29524 96577 29610
rect 96663 29524 96756 29610
rect 96316 29442 96756 29524
rect 96316 29356 96409 29442
rect 96495 29356 96577 29442
rect 96663 29356 96756 29442
rect 96316 29274 96756 29356
rect 96316 29188 96409 29274
rect 96495 29188 96577 29274
rect 96663 29188 96756 29274
rect 96316 29106 96756 29188
rect 96316 29020 96409 29106
rect 96495 29020 96577 29106
rect 96663 29020 96756 29106
rect 96316 28906 96756 29020
rect 96316 28526 96346 28906
rect 96726 28526 96756 28906
rect 96316 24906 96756 28526
rect 96316 24526 96346 24906
rect 96726 24526 96756 24906
rect 96316 23479 96756 24526
rect 96316 23393 96409 23479
rect 96495 23393 96577 23479
rect 96663 23393 96756 23479
rect 96316 21967 96756 23393
rect 96316 21881 96409 21967
rect 96495 21881 96577 21967
rect 96663 21881 96756 21967
rect 96316 20906 96756 21881
rect 96316 20526 96346 20906
rect 96726 20526 96756 20906
rect 96316 20455 96756 20526
rect 96316 20369 96409 20455
rect 96495 20369 96577 20455
rect 96663 20369 96756 20455
rect 96316 18943 96756 20369
rect 96316 18857 96409 18943
rect 96495 18857 96577 18943
rect 96663 18857 96756 18943
rect 96316 17431 96756 18857
rect 96316 17345 96409 17431
rect 96495 17345 96577 17431
rect 96663 17345 96756 17431
rect 96316 16906 96756 17345
rect 96316 16526 96346 16906
rect 96726 16526 96756 16906
rect 96316 15122 96756 16526
rect 96316 15036 96409 15122
rect 96495 15036 96577 15122
rect 96663 15036 96756 15122
rect 96316 14954 96756 15036
rect 96316 14868 96409 14954
rect 96495 14868 96577 14954
rect 96663 14868 96756 14954
rect 96316 14786 96756 14868
rect 96316 14700 96409 14786
rect 96495 14700 96577 14786
rect 96663 14700 96756 14786
rect 96316 14618 96756 14700
rect 96316 14532 96409 14618
rect 96495 14532 96577 14618
rect 96663 14532 96756 14618
rect 96316 14450 96756 14532
rect 96316 14364 96409 14450
rect 96495 14364 96577 14450
rect 96663 14364 96756 14450
rect 96316 14282 96756 14364
rect 96316 14196 96409 14282
rect 96495 14196 96577 14282
rect 96663 14196 96756 14282
rect 96316 14114 96756 14196
rect 96316 14028 96409 14114
rect 96495 14028 96577 14114
rect 96663 14028 96756 14114
rect 96316 13946 96756 14028
rect 96316 13860 96409 13946
rect 96495 13860 96577 13946
rect 96663 13860 96756 13946
rect 96316 13778 96756 13860
rect 96316 13692 96409 13778
rect 96495 13692 96577 13778
rect 96663 13692 96756 13778
rect 96316 13610 96756 13692
rect 96316 13524 96409 13610
rect 96495 13524 96577 13610
rect 96663 13524 96756 13610
rect 96316 13442 96756 13524
rect 96316 13356 96409 13442
rect 96495 13356 96577 13442
rect 96663 13356 96756 13442
rect 96316 13274 96756 13356
rect 96316 13188 96409 13274
rect 96495 13188 96577 13274
rect 96663 13188 96756 13274
rect 96316 13106 96756 13188
rect 96316 13020 96409 13106
rect 96495 13020 96577 13106
rect 96663 13020 96756 13106
rect 96316 12906 96756 13020
rect 96316 12526 96346 12906
rect 96726 12526 96756 12906
rect 96316 8906 96756 12526
rect 96316 8526 96346 8906
rect 96726 8526 96756 8906
rect 96316 6847 96756 8526
rect 96316 6761 96409 6847
rect 96495 6761 96577 6847
rect 96663 6761 96756 6847
rect 96316 5335 96756 6761
rect 96316 5249 96409 5335
rect 96495 5249 96577 5335
rect 96663 5249 96756 5335
rect 96316 4906 96756 5249
rect 96316 4526 96346 4906
rect 96726 4526 96756 4906
rect 96316 3823 96756 4526
rect 96316 3737 96409 3823
rect 96495 3737 96577 3823
rect 96663 3737 96756 3823
rect 96316 2311 96756 3737
rect 96316 2225 96409 2311
rect 96495 2225 96577 2311
rect 96663 2225 96756 2311
rect 96316 799 96756 2225
rect 96316 713 96409 799
rect 96495 713 96577 799
rect 96663 713 96756 799
rect 96316 630 96756 713
rect 99076 37843 99516 38600
rect 99076 37757 99169 37843
rect 99255 37757 99337 37843
rect 99423 37757 99516 37843
rect 99076 36331 99516 37757
rect 99076 36245 99169 36331
rect 99255 36245 99337 36331
rect 99423 36245 99516 36331
rect 99076 35666 99516 36245
rect 99076 35286 99106 35666
rect 99486 35286 99516 35666
rect 99076 34819 99516 35286
rect 99076 34733 99169 34819
rect 99255 34733 99337 34819
rect 99423 34733 99516 34819
rect 99076 31666 99516 34733
rect 99076 31286 99106 31666
rect 99486 31286 99516 31666
rect 99076 27666 99516 31286
rect 99076 27286 99106 27666
rect 99486 27286 99516 27666
rect 99076 23666 99516 27286
rect 99076 23286 99106 23666
rect 99486 23286 99516 23666
rect 99076 22723 99516 23286
rect 99076 22637 99169 22723
rect 99255 22637 99337 22723
rect 99423 22637 99516 22723
rect 99076 21211 99516 22637
rect 99076 21125 99169 21211
rect 99255 21125 99337 21211
rect 99423 21125 99516 21211
rect 99076 19699 99516 21125
rect 99076 19666 99169 19699
rect 99255 19666 99337 19699
rect 99423 19666 99516 19699
rect 99076 19286 99106 19666
rect 99486 19286 99516 19666
rect 99076 18187 99516 19286
rect 99076 18101 99169 18187
rect 99255 18101 99337 18187
rect 99423 18101 99516 18187
rect 99076 15666 99516 18101
rect 99076 15286 99106 15666
rect 99486 15286 99516 15666
rect 99076 11666 99516 15286
rect 99076 11286 99106 11666
rect 99486 11286 99516 11666
rect 99076 7666 99516 11286
rect 99076 7286 99106 7666
rect 99486 7286 99516 7666
rect 99076 6091 99516 7286
rect 99076 6005 99169 6091
rect 99255 6005 99337 6091
rect 99423 6005 99516 6091
rect 99076 4579 99516 6005
rect 99076 4493 99169 4579
rect 99255 4493 99337 4579
rect 99423 4493 99516 4579
rect 99076 3666 99516 4493
rect 99076 3286 99106 3666
rect 99486 3286 99516 3666
rect 99076 3067 99516 3286
rect 99076 2981 99169 3067
rect 99255 2981 99337 3067
rect 99423 2981 99516 3067
rect 99076 1555 99516 2981
rect 99076 1469 99169 1555
rect 99255 1469 99337 1555
rect 99423 1469 99516 1555
rect 99076 712 99516 1469
<< via6 >>
rect 3106 35286 3486 35666
rect 3106 31286 3486 31666
rect 3106 27286 3486 27666
rect 3106 23286 3486 23666
rect 3106 19613 3169 19666
rect 3169 19613 3255 19666
rect 3255 19613 3337 19666
rect 3337 19613 3423 19666
rect 3423 19613 3486 19666
rect 3106 19286 3486 19613
rect 3106 15286 3486 15666
rect 3106 11286 3486 11666
rect 3106 7603 3486 7666
rect 3106 7517 3169 7603
rect 3169 7517 3255 7603
rect 3255 7517 3337 7603
rect 3337 7517 3423 7603
rect 3423 7517 3486 7603
rect 3106 7286 3486 7517
rect 3106 3286 3486 3666
rect 4346 36526 4726 36906
rect 4346 32551 4726 32906
rect 4346 32526 4409 32551
rect 4409 32526 4495 32551
rect 4495 32526 4577 32551
rect 4577 32526 4663 32551
rect 4663 32526 4726 32551
rect 4346 28526 4726 28906
rect 4346 24905 4409 24906
rect 4409 24905 4495 24906
rect 4495 24905 4577 24906
rect 4577 24905 4663 24906
rect 4663 24905 4726 24906
rect 4346 24526 4726 24905
rect 4346 20526 4726 20906
rect 4346 16526 4726 16906
rect 4346 12895 4726 12906
rect 4346 12809 4409 12895
rect 4409 12809 4495 12895
rect 4495 12809 4577 12895
rect 4577 12809 4663 12895
rect 4663 12809 4726 12895
rect 4346 12526 4726 12809
rect 4346 8526 4726 8906
rect 4346 4526 4726 4906
rect 7106 35286 7486 35666
rect 7106 31286 7486 31666
rect 7106 27286 7486 27666
rect 7106 23286 7486 23666
rect 7106 19613 7169 19666
rect 7169 19613 7255 19666
rect 7255 19613 7337 19666
rect 7337 19613 7423 19666
rect 7423 19613 7486 19666
rect 7106 19286 7486 19613
rect 7106 15286 7486 15666
rect 7106 11286 7486 11666
rect 7106 7603 7486 7666
rect 7106 7517 7169 7603
rect 7169 7517 7255 7603
rect 7255 7517 7337 7603
rect 7337 7517 7423 7603
rect 7423 7517 7486 7603
rect 7106 7286 7486 7517
rect 7106 3286 7486 3666
rect 8346 36526 8726 36906
rect 8346 32551 8726 32906
rect 8346 32526 8409 32551
rect 8409 32526 8495 32551
rect 8495 32526 8577 32551
rect 8577 32526 8663 32551
rect 8663 32526 8726 32551
rect 8346 28526 8726 28906
rect 8346 24905 8409 24906
rect 8409 24905 8495 24906
rect 8495 24905 8577 24906
rect 8577 24905 8663 24906
rect 8663 24905 8726 24906
rect 8346 24526 8726 24905
rect 8346 20526 8726 20906
rect 8346 16526 8726 16906
rect 8346 12895 8726 12906
rect 8346 12809 8409 12895
rect 8409 12809 8495 12895
rect 8495 12809 8577 12895
rect 8577 12809 8663 12895
rect 8663 12809 8726 12895
rect 8346 12526 8726 12809
rect 8346 8526 8726 8906
rect 8346 4526 8726 4906
rect 11106 35286 11486 35666
rect 11106 31286 11486 31666
rect 11106 27286 11486 27666
rect 11106 23286 11486 23666
rect 11106 19613 11169 19666
rect 11169 19613 11255 19666
rect 11255 19613 11337 19666
rect 11337 19613 11423 19666
rect 11423 19613 11486 19666
rect 11106 19286 11486 19613
rect 11106 15286 11486 15666
rect 11106 11286 11486 11666
rect 11106 7603 11486 7666
rect 11106 7517 11169 7603
rect 11169 7517 11255 7603
rect 11255 7517 11337 7603
rect 11337 7517 11423 7603
rect 11423 7517 11486 7603
rect 11106 7286 11486 7517
rect 11106 3286 11486 3666
rect 12346 36526 12726 36906
rect 12346 32551 12726 32906
rect 12346 32526 12409 32551
rect 12409 32526 12495 32551
rect 12495 32526 12577 32551
rect 12577 32526 12663 32551
rect 12663 32526 12726 32551
rect 12346 28526 12726 28906
rect 12346 24905 12409 24906
rect 12409 24905 12495 24906
rect 12495 24905 12577 24906
rect 12577 24905 12663 24906
rect 12663 24905 12726 24906
rect 12346 24526 12726 24905
rect 12346 20526 12726 20906
rect 12346 16526 12726 16906
rect 12346 12895 12726 12906
rect 12346 12809 12409 12895
rect 12409 12809 12495 12895
rect 12495 12809 12577 12895
rect 12577 12809 12663 12895
rect 12663 12809 12726 12895
rect 12346 12526 12726 12809
rect 12346 8526 12726 8906
rect 12346 4526 12726 4906
rect 15106 35286 15486 35666
rect 15106 31286 15486 31666
rect 15106 27286 15486 27666
rect 15106 23286 15486 23666
rect 15106 19613 15169 19666
rect 15169 19613 15255 19666
rect 15255 19613 15337 19666
rect 15337 19613 15423 19666
rect 15423 19613 15486 19666
rect 15106 19286 15486 19613
rect 15106 15286 15486 15666
rect 15106 11286 15486 11666
rect 15106 7603 15486 7666
rect 15106 7517 15169 7603
rect 15169 7517 15255 7603
rect 15255 7517 15337 7603
rect 15337 7517 15423 7603
rect 15423 7517 15486 7603
rect 15106 7286 15486 7517
rect 15106 3286 15486 3666
rect 16346 36526 16726 36906
rect 16346 32551 16726 32906
rect 16346 32526 16409 32551
rect 16409 32526 16495 32551
rect 16495 32526 16577 32551
rect 16577 32526 16663 32551
rect 16663 32526 16726 32551
rect 16346 28526 16726 28906
rect 16346 24905 16409 24906
rect 16409 24905 16495 24906
rect 16495 24905 16577 24906
rect 16577 24905 16663 24906
rect 16663 24905 16726 24906
rect 16346 24526 16726 24905
rect 16346 20526 16726 20906
rect 16346 16526 16726 16906
rect 16346 12895 16726 12906
rect 16346 12809 16409 12895
rect 16409 12809 16495 12895
rect 16495 12809 16577 12895
rect 16577 12809 16663 12895
rect 16663 12809 16726 12895
rect 16346 12526 16726 12809
rect 16346 8526 16726 8906
rect 16346 4526 16726 4906
rect 19106 35286 19486 35666
rect 19106 31286 19486 31666
rect 19106 27286 19486 27666
rect 19106 23286 19486 23666
rect 19106 19613 19169 19666
rect 19169 19613 19255 19666
rect 19255 19613 19337 19666
rect 19337 19613 19423 19666
rect 19423 19613 19486 19666
rect 19106 19286 19486 19613
rect 19106 15286 19486 15666
rect 19106 11286 19486 11666
rect 19106 7603 19486 7666
rect 19106 7517 19169 7603
rect 19169 7517 19255 7603
rect 19255 7517 19337 7603
rect 19337 7517 19423 7603
rect 19423 7517 19486 7603
rect 19106 7286 19486 7517
rect 19106 3286 19486 3666
rect 20346 36526 20726 36906
rect 20346 32551 20726 32906
rect 20346 32526 20409 32551
rect 20409 32526 20495 32551
rect 20495 32526 20577 32551
rect 20577 32526 20663 32551
rect 20663 32526 20726 32551
rect 20346 28526 20726 28906
rect 20346 24905 20409 24906
rect 20409 24905 20495 24906
rect 20495 24905 20577 24906
rect 20577 24905 20663 24906
rect 20663 24905 20726 24906
rect 20346 24526 20726 24905
rect 20346 20526 20726 20906
rect 20346 16526 20726 16906
rect 20346 12895 20726 12906
rect 20346 12809 20409 12895
rect 20409 12809 20495 12895
rect 20495 12809 20577 12895
rect 20577 12809 20663 12895
rect 20663 12809 20726 12895
rect 20346 12526 20726 12809
rect 20346 8526 20726 8906
rect 20346 4526 20726 4906
rect 23106 35286 23486 35666
rect 23106 31286 23486 31666
rect 23106 27286 23486 27666
rect 23106 23286 23486 23666
rect 23106 19613 23169 19666
rect 23169 19613 23255 19666
rect 23255 19613 23337 19666
rect 23337 19613 23423 19666
rect 23423 19613 23486 19666
rect 23106 19286 23486 19613
rect 23106 15286 23486 15666
rect 23106 11286 23486 11666
rect 23106 7603 23486 7666
rect 23106 7517 23169 7603
rect 23169 7517 23255 7603
rect 23255 7517 23337 7603
rect 23337 7517 23423 7603
rect 23423 7517 23486 7603
rect 23106 7286 23486 7517
rect 23106 3286 23486 3666
rect 24346 36526 24726 36906
rect 24346 32551 24726 32906
rect 24346 32526 24409 32551
rect 24409 32526 24495 32551
rect 24495 32526 24577 32551
rect 24577 32526 24663 32551
rect 24663 32526 24726 32551
rect 24346 28526 24726 28906
rect 24346 24905 24409 24906
rect 24409 24905 24495 24906
rect 24495 24905 24577 24906
rect 24577 24905 24663 24906
rect 24663 24905 24726 24906
rect 24346 24526 24726 24905
rect 24346 20526 24726 20906
rect 24346 16526 24726 16906
rect 24346 12895 24726 12906
rect 24346 12809 24409 12895
rect 24409 12809 24495 12895
rect 24495 12809 24577 12895
rect 24577 12809 24663 12895
rect 24663 12809 24726 12895
rect 24346 12526 24726 12809
rect 24346 8526 24726 8906
rect 24346 4526 24726 4906
rect 27106 35286 27486 35666
rect 27106 31286 27486 31666
rect 27106 27286 27486 27666
rect 27106 23286 27486 23666
rect 27106 19613 27169 19666
rect 27169 19613 27255 19666
rect 27255 19613 27337 19666
rect 27337 19613 27423 19666
rect 27423 19613 27486 19666
rect 27106 19286 27486 19613
rect 27106 15286 27486 15666
rect 27106 11286 27486 11666
rect 27106 7603 27486 7666
rect 27106 7517 27169 7603
rect 27169 7517 27255 7603
rect 27255 7517 27337 7603
rect 27337 7517 27423 7603
rect 27423 7517 27486 7603
rect 27106 7286 27486 7517
rect 27106 3286 27486 3666
rect 28346 36526 28726 36906
rect 28346 32551 28726 32906
rect 28346 32526 28409 32551
rect 28409 32526 28495 32551
rect 28495 32526 28577 32551
rect 28577 32526 28663 32551
rect 28663 32526 28726 32551
rect 28346 28526 28726 28906
rect 28346 24905 28409 24906
rect 28409 24905 28495 24906
rect 28495 24905 28577 24906
rect 28577 24905 28663 24906
rect 28663 24905 28726 24906
rect 28346 24526 28726 24905
rect 28346 20526 28726 20906
rect 28346 16526 28726 16906
rect 28346 12895 28726 12906
rect 28346 12809 28409 12895
rect 28409 12809 28495 12895
rect 28495 12809 28577 12895
rect 28577 12809 28663 12895
rect 28663 12809 28726 12895
rect 28346 12526 28726 12809
rect 28346 8526 28726 8906
rect 28346 4526 28726 4906
rect 31106 35286 31486 35666
rect 31106 31286 31486 31666
rect 31106 27286 31486 27666
rect 31106 23286 31486 23666
rect 31106 19613 31169 19666
rect 31169 19613 31255 19666
rect 31255 19613 31337 19666
rect 31337 19613 31423 19666
rect 31423 19613 31486 19666
rect 31106 19286 31486 19613
rect 31106 15286 31486 15666
rect 31106 11286 31486 11666
rect 31106 7603 31486 7666
rect 31106 7517 31169 7603
rect 31169 7517 31255 7603
rect 31255 7517 31337 7603
rect 31337 7517 31423 7603
rect 31423 7517 31486 7603
rect 31106 7286 31486 7517
rect 31106 3286 31486 3666
rect 32346 36526 32726 36906
rect 32346 32551 32726 32906
rect 32346 32526 32409 32551
rect 32409 32526 32495 32551
rect 32495 32526 32577 32551
rect 32577 32526 32663 32551
rect 32663 32526 32726 32551
rect 32346 28526 32726 28906
rect 32346 24905 32409 24906
rect 32409 24905 32495 24906
rect 32495 24905 32577 24906
rect 32577 24905 32663 24906
rect 32663 24905 32726 24906
rect 32346 24526 32726 24905
rect 32346 20526 32726 20906
rect 32346 16526 32726 16906
rect 32346 12895 32726 12906
rect 32346 12809 32409 12895
rect 32409 12809 32495 12895
rect 32495 12809 32577 12895
rect 32577 12809 32663 12895
rect 32663 12809 32726 12895
rect 32346 12526 32726 12809
rect 32346 8526 32726 8906
rect 32346 4526 32726 4906
rect 35106 35286 35486 35666
rect 35106 31286 35486 31666
rect 35106 27286 35486 27666
rect 35106 23286 35486 23666
rect 35106 19613 35169 19666
rect 35169 19613 35255 19666
rect 35255 19613 35337 19666
rect 35337 19613 35423 19666
rect 35423 19613 35486 19666
rect 35106 19286 35486 19613
rect 35106 15286 35486 15666
rect 35106 11286 35486 11666
rect 35106 7603 35486 7666
rect 35106 7517 35169 7603
rect 35169 7517 35255 7603
rect 35255 7517 35337 7603
rect 35337 7517 35423 7603
rect 35423 7517 35486 7603
rect 35106 7286 35486 7517
rect 35106 3286 35486 3666
rect 36346 36526 36726 36906
rect 36346 32551 36726 32906
rect 36346 32526 36409 32551
rect 36409 32526 36495 32551
rect 36495 32526 36577 32551
rect 36577 32526 36663 32551
rect 36663 32526 36726 32551
rect 36346 28526 36726 28906
rect 36346 24905 36409 24906
rect 36409 24905 36495 24906
rect 36495 24905 36577 24906
rect 36577 24905 36663 24906
rect 36663 24905 36726 24906
rect 36346 24526 36726 24905
rect 36346 20526 36726 20906
rect 36346 16526 36726 16906
rect 36346 12895 36726 12906
rect 36346 12809 36409 12895
rect 36409 12809 36495 12895
rect 36495 12809 36577 12895
rect 36577 12809 36663 12895
rect 36663 12809 36726 12895
rect 36346 12526 36726 12809
rect 36346 8526 36726 8906
rect 36346 4526 36726 4906
rect 39106 35286 39486 35666
rect 39106 31286 39486 31666
rect 39106 27286 39486 27666
rect 39106 23286 39486 23666
rect 39106 19613 39169 19666
rect 39169 19613 39255 19666
rect 39255 19613 39337 19666
rect 39337 19613 39423 19666
rect 39423 19613 39486 19666
rect 39106 19286 39486 19613
rect 39106 15286 39486 15666
rect 39106 11286 39486 11666
rect 39106 7603 39486 7666
rect 39106 7517 39169 7603
rect 39169 7517 39255 7603
rect 39255 7517 39337 7603
rect 39337 7517 39423 7603
rect 39423 7517 39486 7603
rect 39106 7286 39486 7517
rect 39106 3286 39486 3666
rect 40346 36526 40726 36906
rect 40346 32551 40726 32906
rect 40346 32526 40409 32551
rect 40409 32526 40495 32551
rect 40495 32526 40577 32551
rect 40577 32526 40663 32551
rect 40663 32526 40726 32551
rect 40346 28526 40726 28906
rect 40346 24905 40409 24906
rect 40409 24905 40495 24906
rect 40495 24905 40577 24906
rect 40577 24905 40663 24906
rect 40663 24905 40726 24906
rect 40346 24526 40726 24905
rect 40346 20526 40726 20906
rect 40346 16526 40726 16906
rect 40346 12895 40726 12906
rect 40346 12809 40409 12895
rect 40409 12809 40495 12895
rect 40495 12809 40577 12895
rect 40577 12809 40663 12895
rect 40663 12809 40726 12895
rect 40346 12526 40726 12809
rect 40346 8526 40726 8906
rect 40346 4526 40726 4906
rect 43106 35286 43486 35666
rect 43106 31286 43486 31666
rect 43106 27286 43486 27666
rect 43106 23286 43486 23666
rect 43106 19613 43169 19666
rect 43169 19613 43255 19666
rect 43255 19613 43337 19666
rect 43337 19613 43423 19666
rect 43423 19613 43486 19666
rect 43106 19286 43486 19613
rect 43106 15286 43486 15666
rect 43106 11286 43486 11666
rect 43106 7603 43486 7666
rect 43106 7517 43169 7603
rect 43169 7517 43255 7603
rect 43255 7517 43337 7603
rect 43337 7517 43423 7603
rect 43423 7517 43486 7603
rect 43106 7286 43486 7517
rect 43106 3286 43486 3666
rect 44346 36526 44726 36906
rect 44346 32551 44726 32906
rect 44346 32526 44409 32551
rect 44409 32526 44495 32551
rect 44495 32526 44577 32551
rect 44577 32526 44663 32551
rect 44663 32526 44726 32551
rect 44346 28526 44726 28906
rect 44346 24905 44409 24906
rect 44409 24905 44495 24906
rect 44495 24905 44577 24906
rect 44577 24905 44663 24906
rect 44663 24905 44726 24906
rect 44346 24526 44726 24905
rect 44346 20526 44726 20906
rect 44346 16526 44726 16906
rect 44346 12895 44726 12906
rect 44346 12809 44409 12895
rect 44409 12809 44495 12895
rect 44495 12809 44577 12895
rect 44577 12809 44663 12895
rect 44663 12809 44726 12895
rect 44346 12526 44726 12809
rect 44346 8526 44726 8906
rect 44346 4526 44726 4906
rect 47106 35286 47486 35666
rect 47106 31286 47486 31666
rect 47106 27286 47486 27666
rect 47106 23286 47486 23666
rect 47106 19613 47169 19666
rect 47169 19613 47255 19666
rect 47255 19613 47337 19666
rect 47337 19613 47423 19666
rect 47423 19613 47486 19666
rect 47106 19286 47486 19613
rect 47106 15286 47486 15666
rect 47106 11286 47486 11666
rect 47106 7603 47486 7666
rect 47106 7517 47169 7603
rect 47169 7517 47255 7603
rect 47255 7517 47337 7603
rect 47337 7517 47423 7603
rect 47423 7517 47486 7603
rect 47106 7286 47486 7517
rect 47106 3286 47486 3666
rect 48346 36526 48726 36906
rect 48346 32551 48726 32906
rect 48346 32526 48409 32551
rect 48409 32526 48495 32551
rect 48495 32526 48577 32551
rect 48577 32526 48663 32551
rect 48663 32526 48726 32551
rect 48346 28526 48726 28906
rect 48346 24905 48409 24906
rect 48409 24905 48495 24906
rect 48495 24905 48577 24906
rect 48577 24905 48663 24906
rect 48663 24905 48726 24906
rect 48346 24526 48726 24905
rect 48346 20526 48726 20906
rect 48346 16526 48726 16906
rect 48346 12895 48726 12906
rect 48346 12809 48409 12895
rect 48409 12809 48495 12895
rect 48495 12809 48577 12895
rect 48577 12809 48663 12895
rect 48663 12809 48726 12895
rect 48346 12526 48726 12809
rect 48346 8526 48726 8906
rect 48346 4526 48726 4906
rect 51106 35286 51486 35666
rect 51106 31286 51486 31666
rect 51106 27286 51486 27666
rect 51106 23286 51486 23666
rect 51106 19613 51169 19666
rect 51169 19613 51255 19666
rect 51255 19613 51337 19666
rect 51337 19613 51423 19666
rect 51423 19613 51486 19666
rect 51106 19286 51486 19613
rect 51106 15286 51486 15666
rect 51106 11286 51486 11666
rect 51106 7603 51486 7666
rect 51106 7517 51169 7603
rect 51169 7517 51255 7603
rect 51255 7517 51337 7603
rect 51337 7517 51423 7603
rect 51423 7517 51486 7603
rect 51106 7286 51486 7517
rect 51106 3286 51486 3666
rect 52346 36526 52726 36906
rect 52346 32551 52726 32906
rect 52346 32526 52409 32551
rect 52409 32526 52495 32551
rect 52495 32526 52577 32551
rect 52577 32526 52663 32551
rect 52663 32526 52726 32551
rect 52346 28526 52726 28906
rect 52346 24905 52409 24906
rect 52409 24905 52495 24906
rect 52495 24905 52577 24906
rect 52577 24905 52663 24906
rect 52663 24905 52726 24906
rect 52346 24526 52726 24905
rect 52346 20526 52726 20906
rect 52346 16526 52726 16906
rect 52346 12895 52726 12906
rect 52346 12809 52409 12895
rect 52409 12809 52495 12895
rect 52495 12809 52577 12895
rect 52577 12809 52663 12895
rect 52663 12809 52726 12895
rect 52346 12526 52726 12809
rect 52346 8526 52726 8906
rect 52346 4526 52726 4906
rect 55106 35286 55486 35666
rect 55106 31286 55486 31666
rect 55106 27286 55486 27666
rect 55106 23286 55486 23666
rect 55106 19613 55169 19666
rect 55169 19613 55255 19666
rect 55255 19613 55337 19666
rect 55337 19613 55423 19666
rect 55423 19613 55486 19666
rect 55106 19286 55486 19613
rect 55106 15286 55486 15666
rect 55106 11286 55486 11666
rect 55106 7603 55486 7666
rect 55106 7517 55169 7603
rect 55169 7517 55255 7603
rect 55255 7517 55337 7603
rect 55337 7517 55423 7603
rect 55423 7517 55486 7603
rect 55106 7286 55486 7517
rect 55106 3286 55486 3666
rect 56346 36526 56726 36906
rect 56346 32551 56726 32906
rect 56346 32526 56409 32551
rect 56409 32526 56495 32551
rect 56495 32526 56577 32551
rect 56577 32526 56663 32551
rect 56663 32526 56726 32551
rect 56346 28526 56726 28906
rect 56346 24905 56409 24906
rect 56409 24905 56495 24906
rect 56495 24905 56577 24906
rect 56577 24905 56663 24906
rect 56663 24905 56726 24906
rect 56346 24526 56726 24905
rect 56346 20526 56726 20906
rect 56346 16526 56726 16906
rect 56346 12895 56726 12906
rect 56346 12809 56409 12895
rect 56409 12809 56495 12895
rect 56495 12809 56577 12895
rect 56577 12809 56663 12895
rect 56663 12809 56726 12895
rect 56346 12526 56726 12809
rect 56346 8526 56726 8906
rect 56346 4526 56726 4906
rect 59106 35286 59486 35666
rect 59106 31286 59486 31666
rect 59106 27286 59486 27666
rect 59106 23286 59486 23666
rect 59106 19613 59169 19666
rect 59169 19613 59255 19666
rect 59255 19613 59337 19666
rect 59337 19613 59423 19666
rect 59423 19613 59486 19666
rect 59106 19286 59486 19613
rect 59106 15286 59486 15666
rect 59106 11286 59486 11666
rect 59106 7603 59486 7666
rect 59106 7517 59169 7603
rect 59169 7517 59255 7603
rect 59255 7517 59337 7603
rect 59337 7517 59423 7603
rect 59423 7517 59486 7603
rect 59106 7286 59486 7517
rect 59106 3286 59486 3666
rect 60346 36526 60726 36906
rect 60346 32551 60726 32906
rect 60346 32526 60409 32551
rect 60409 32526 60495 32551
rect 60495 32526 60577 32551
rect 60577 32526 60663 32551
rect 60663 32526 60726 32551
rect 60346 28526 60726 28906
rect 60346 24905 60409 24906
rect 60409 24905 60495 24906
rect 60495 24905 60577 24906
rect 60577 24905 60663 24906
rect 60663 24905 60726 24906
rect 60346 24526 60726 24905
rect 60346 20526 60726 20906
rect 60346 16526 60726 16906
rect 60346 12895 60726 12906
rect 60346 12809 60409 12895
rect 60409 12809 60495 12895
rect 60495 12809 60577 12895
rect 60577 12809 60663 12895
rect 60663 12809 60726 12895
rect 60346 12526 60726 12809
rect 60346 8526 60726 8906
rect 60346 4526 60726 4906
rect 63106 35286 63486 35666
rect 63106 31286 63486 31666
rect 63106 27286 63486 27666
rect 63106 23286 63486 23666
rect 63106 19613 63169 19666
rect 63169 19613 63255 19666
rect 63255 19613 63337 19666
rect 63337 19613 63423 19666
rect 63423 19613 63486 19666
rect 63106 19286 63486 19613
rect 63106 15286 63486 15666
rect 63106 11286 63486 11666
rect 63106 7603 63486 7666
rect 63106 7517 63169 7603
rect 63169 7517 63255 7603
rect 63255 7517 63337 7603
rect 63337 7517 63423 7603
rect 63423 7517 63486 7603
rect 63106 7286 63486 7517
rect 63106 3286 63486 3666
rect 64346 36526 64726 36906
rect 64346 32551 64726 32906
rect 64346 32526 64409 32551
rect 64409 32526 64495 32551
rect 64495 32526 64577 32551
rect 64577 32526 64663 32551
rect 64663 32526 64726 32551
rect 64346 28526 64726 28906
rect 64346 24905 64409 24906
rect 64409 24905 64495 24906
rect 64495 24905 64577 24906
rect 64577 24905 64663 24906
rect 64663 24905 64726 24906
rect 64346 24526 64726 24905
rect 64346 20526 64726 20906
rect 64346 16526 64726 16906
rect 64346 12895 64726 12906
rect 64346 12809 64409 12895
rect 64409 12809 64495 12895
rect 64495 12809 64577 12895
rect 64577 12809 64663 12895
rect 64663 12809 64726 12895
rect 64346 12526 64726 12809
rect 64346 8526 64726 8906
rect 64346 4526 64726 4906
rect 67106 35286 67486 35666
rect 67106 31286 67486 31666
rect 67106 27286 67486 27666
rect 67106 23286 67486 23666
rect 67106 19613 67169 19666
rect 67169 19613 67255 19666
rect 67255 19613 67337 19666
rect 67337 19613 67423 19666
rect 67423 19613 67486 19666
rect 67106 19286 67486 19613
rect 67106 15286 67486 15666
rect 67106 11286 67486 11666
rect 67106 7603 67486 7666
rect 67106 7517 67169 7603
rect 67169 7517 67255 7603
rect 67255 7517 67337 7603
rect 67337 7517 67423 7603
rect 67423 7517 67486 7603
rect 67106 7286 67486 7517
rect 67106 3286 67486 3666
rect 68346 36526 68726 36906
rect 68346 32551 68726 32906
rect 68346 32526 68409 32551
rect 68409 32526 68495 32551
rect 68495 32526 68577 32551
rect 68577 32526 68663 32551
rect 68663 32526 68726 32551
rect 68346 28526 68726 28906
rect 68346 24905 68409 24906
rect 68409 24905 68495 24906
rect 68495 24905 68577 24906
rect 68577 24905 68663 24906
rect 68663 24905 68726 24906
rect 68346 24526 68726 24905
rect 68346 20526 68726 20906
rect 68346 16526 68726 16906
rect 68346 12895 68726 12906
rect 68346 12809 68409 12895
rect 68409 12809 68495 12895
rect 68495 12809 68577 12895
rect 68577 12809 68663 12895
rect 68663 12809 68726 12895
rect 68346 12526 68726 12809
rect 68346 8526 68726 8906
rect 68346 4526 68726 4906
rect 71106 35286 71486 35666
rect 71106 31286 71486 31666
rect 71106 27286 71486 27666
rect 71106 23286 71486 23666
rect 71106 19613 71169 19666
rect 71169 19613 71255 19666
rect 71255 19613 71337 19666
rect 71337 19613 71423 19666
rect 71423 19613 71486 19666
rect 71106 19286 71486 19613
rect 71106 15286 71486 15666
rect 71106 11286 71486 11666
rect 71106 7603 71486 7666
rect 71106 7517 71169 7603
rect 71169 7517 71255 7603
rect 71255 7517 71337 7603
rect 71337 7517 71423 7603
rect 71423 7517 71486 7603
rect 71106 7286 71486 7517
rect 71106 3286 71486 3666
rect 72346 36526 72726 36906
rect 72346 32526 72726 32906
rect 72346 28526 72726 28906
rect 72346 24526 72726 24906
rect 72346 20526 72726 20906
rect 72346 16526 72726 16906
rect 72346 12526 72726 12906
rect 72346 8526 72726 8906
rect 72346 4526 72726 4906
rect 75106 35286 75486 35666
rect 75106 31286 75486 31666
rect 75106 27656 75169 27666
rect 75169 27656 75255 27666
rect 75255 27656 75337 27666
rect 75337 27656 75423 27666
rect 75423 27656 75486 27666
rect 75106 27574 75486 27656
rect 75106 27488 75169 27574
rect 75169 27488 75255 27574
rect 75255 27488 75337 27574
rect 75337 27488 75423 27574
rect 75423 27488 75486 27574
rect 75106 27406 75486 27488
rect 75106 27320 75169 27406
rect 75169 27320 75255 27406
rect 75255 27320 75337 27406
rect 75337 27320 75423 27406
rect 75423 27320 75486 27406
rect 75106 27286 75486 27320
rect 75106 23286 75486 23666
rect 75106 19613 75169 19666
rect 75169 19613 75255 19666
rect 75255 19613 75337 19666
rect 75337 19613 75423 19666
rect 75423 19613 75486 19666
rect 75106 19286 75486 19613
rect 75106 15286 75486 15666
rect 75106 11656 75169 11666
rect 75169 11656 75255 11666
rect 75255 11656 75337 11666
rect 75337 11656 75423 11666
rect 75423 11656 75486 11666
rect 75106 11574 75486 11656
rect 75106 11488 75169 11574
rect 75169 11488 75255 11574
rect 75255 11488 75337 11574
rect 75337 11488 75423 11574
rect 75423 11488 75486 11574
rect 75106 11406 75486 11488
rect 75106 11320 75169 11406
rect 75169 11320 75255 11406
rect 75255 11320 75337 11406
rect 75337 11320 75423 11406
rect 75423 11320 75486 11406
rect 75106 11286 75486 11320
rect 75106 7603 75486 7666
rect 75106 7517 75169 7603
rect 75169 7517 75255 7603
rect 75255 7517 75337 7603
rect 75337 7517 75423 7603
rect 75423 7517 75486 7603
rect 75106 7286 75486 7517
rect 75106 3286 75486 3666
rect 76346 36526 76726 36906
rect 76346 32526 76726 32906
rect 76346 28526 76726 28906
rect 76346 24526 76726 24906
rect 76346 20526 76726 20906
rect 76346 16526 76726 16906
rect 76346 12526 76726 12906
rect 76346 8526 76726 8906
rect 76346 4526 76726 4906
rect 79106 35286 79486 35666
rect 79106 31286 79486 31666
rect 79106 27656 79169 27666
rect 79169 27656 79255 27666
rect 79255 27656 79337 27666
rect 79337 27656 79423 27666
rect 79423 27656 79486 27666
rect 79106 27574 79486 27656
rect 79106 27488 79169 27574
rect 79169 27488 79255 27574
rect 79255 27488 79337 27574
rect 79337 27488 79423 27574
rect 79423 27488 79486 27574
rect 79106 27406 79486 27488
rect 79106 27320 79169 27406
rect 79169 27320 79255 27406
rect 79255 27320 79337 27406
rect 79337 27320 79423 27406
rect 79423 27320 79486 27406
rect 79106 27286 79486 27320
rect 79106 23286 79486 23666
rect 79106 19613 79169 19666
rect 79169 19613 79255 19666
rect 79255 19613 79337 19666
rect 79337 19613 79423 19666
rect 79423 19613 79486 19666
rect 79106 19286 79486 19613
rect 79106 15286 79486 15666
rect 79106 11656 79169 11666
rect 79169 11656 79255 11666
rect 79255 11656 79337 11666
rect 79337 11656 79423 11666
rect 79423 11656 79486 11666
rect 79106 11574 79486 11656
rect 79106 11488 79169 11574
rect 79169 11488 79255 11574
rect 79255 11488 79337 11574
rect 79337 11488 79423 11574
rect 79423 11488 79486 11574
rect 79106 11406 79486 11488
rect 79106 11320 79169 11406
rect 79169 11320 79255 11406
rect 79255 11320 79337 11406
rect 79337 11320 79423 11406
rect 79423 11320 79486 11406
rect 79106 11286 79486 11320
rect 79106 7603 79486 7666
rect 79106 7517 79169 7603
rect 79169 7517 79255 7603
rect 79255 7517 79337 7603
rect 79337 7517 79423 7603
rect 79423 7517 79486 7603
rect 79106 7286 79486 7517
rect 79106 3286 79486 3666
rect 80346 36526 80726 36906
rect 80346 32526 80726 32906
rect 80346 28526 80726 28906
rect 80346 24526 80726 24906
rect 80346 20526 80726 20906
rect 80346 16526 80726 16906
rect 80346 12526 80726 12906
rect 80346 8526 80726 8906
rect 80346 4526 80726 4906
rect 83106 35286 83486 35666
rect 83106 31286 83486 31666
rect 83106 27656 83169 27666
rect 83169 27656 83255 27666
rect 83255 27656 83337 27666
rect 83337 27656 83423 27666
rect 83423 27656 83486 27666
rect 83106 27574 83486 27656
rect 83106 27488 83169 27574
rect 83169 27488 83255 27574
rect 83255 27488 83337 27574
rect 83337 27488 83423 27574
rect 83423 27488 83486 27574
rect 83106 27406 83486 27488
rect 83106 27320 83169 27406
rect 83169 27320 83255 27406
rect 83255 27320 83337 27406
rect 83337 27320 83423 27406
rect 83423 27320 83486 27406
rect 83106 27286 83486 27320
rect 83106 23286 83486 23666
rect 83106 19613 83169 19666
rect 83169 19613 83255 19666
rect 83255 19613 83337 19666
rect 83337 19613 83423 19666
rect 83423 19613 83486 19666
rect 83106 19286 83486 19613
rect 83106 15286 83486 15666
rect 83106 11656 83169 11666
rect 83169 11656 83255 11666
rect 83255 11656 83337 11666
rect 83337 11656 83423 11666
rect 83423 11656 83486 11666
rect 83106 11574 83486 11656
rect 83106 11488 83169 11574
rect 83169 11488 83255 11574
rect 83255 11488 83337 11574
rect 83337 11488 83423 11574
rect 83423 11488 83486 11574
rect 83106 11406 83486 11488
rect 83106 11320 83169 11406
rect 83169 11320 83255 11406
rect 83255 11320 83337 11406
rect 83337 11320 83423 11406
rect 83423 11320 83486 11406
rect 83106 11286 83486 11320
rect 83106 7603 83486 7666
rect 83106 7517 83169 7603
rect 83169 7517 83255 7603
rect 83255 7517 83337 7603
rect 83337 7517 83423 7603
rect 83423 7517 83486 7603
rect 83106 7286 83486 7517
rect 83106 3286 83486 3666
rect 84346 36526 84726 36906
rect 87106 35286 87486 35666
rect 84346 32526 84726 32906
rect 84346 28526 84726 28906
rect 84346 24526 84726 24906
rect 87106 31286 87486 31666
rect 87106 27656 87169 27666
rect 87169 27656 87255 27666
rect 87255 27656 87337 27666
rect 87337 27656 87423 27666
rect 87423 27656 87486 27666
rect 87106 27574 87486 27656
rect 87106 27488 87169 27574
rect 87169 27488 87255 27574
rect 87255 27488 87337 27574
rect 87337 27488 87423 27574
rect 87423 27488 87486 27574
rect 87106 27406 87486 27488
rect 87106 27320 87169 27406
rect 87169 27320 87255 27406
rect 87255 27320 87337 27406
rect 87337 27320 87423 27406
rect 87423 27320 87486 27406
rect 87106 27286 87486 27320
rect 87106 23286 87486 23666
rect 84346 20526 84726 20906
rect 84346 16526 84726 16906
rect 84346 12526 84726 12906
rect 84346 8526 84726 8906
rect 87106 19613 87169 19666
rect 87169 19613 87255 19666
rect 87255 19613 87337 19666
rect 87337 19613 87423 19666
rect 87423 19613 87486 19666
rect 87106 19286 87486 19613
rect 87106 15286 87486 15666
rect 87106 11656 87169 11666
rect 87169 11656 87255 11666
rect 87255 11656 87337 11666
rect 87337 11656 87423 11666
rect 87423 11656 87486 11666
rect 87106 11574 87486 11656
rect 87106 11488 87169 11574
rect 87169 11488 87255 11574
rect 87255 11488 87337 11574
rect 87337 11488 87423 11574
rect 87423 11488 87486 11574
rect 87106 11406 87486 11488
rect 87106 11320 87169 11406
rect 87169 11320 87255 11406
rect 87255 11320 87337 11406
rect 87337 11320 87423 11406
rect 87423 11320 87486 11406
rect 87106 11286 87486 11320
rect 87106 7603 87486 7666
rect 87106 7517 87169 7603
rect 87169 7517 87255 7603
rect 87255 7517 87337 7603
rect 87337 7517 87423 7603
rect 87423 7517 87486 7603
rect 87106 7286 87486 7517
rect 84346 4526 84726 4906
rect 87106 3286 87486 3666
rect 88346 36526 88726 36906
rect 88346 32526 88726 32906
rect 88346 28526 88726 28906
rect 88346 24526 88726 24906
rect 88346 20526 88726 20906
rect 88346 16526 88726 16906
rect 88346 12526 88726 12906
rect 88346 8526 88726 8906
rect 88346 4526 88726 4906
rect 91106 35286 91486 35666
rect 91106 31286 91486 31666
rect 91106 27656 91169 27666
rect 91169 27656 91255 27666
rect 91255 27656 91337 27666
rect 91337 27656 91423 27666
rect 91423 27656 91486 27666
rect 91106 27574 91486 27656
rect 91106 27488 91169 27574
rect 91169 27488 91255 27574
rect 91255 27488 91337 27574
rect 91337 27488 91423 27574
rect 91423 27488 91486 27574
rect 91106 27406 91486 27488
rect 91106 27320 91169 27406
rect 91169 27320 91255 27406
rect 91255 27320 91337 27406
rect 91337 27320 91423 27406
rect 91423 27320 91486 27406
rect 91106 27286 91486 27320
rect 91106 23286 91486 23666
rect 91106 19613 91169 19666
rect 91169 19613 91255 19666
rect 91255 19613 91337 19666
rect 91337 19613 91423 19666
rect 91423 19613 91486 19666
rect 91106 19286 91486 19613
rect 91106 15286 91486 15666
rect 91106 11656 91169 11666
rect 91169 11656 91255 11666
rect 91255 11656 91337 11666
rect 91337 11656 91423 11666
rect 91423 11656 91486 11666
rect 91106 11574 91486 11656
rect 91106 11488 91169 11574
rect 91169 11488 91255 11574
rect 91255 11488 91337 11574
rect 91337 11488 91423 11574
rect 91423 11488 91486 11574
rect 91106 11406 91486 11488
rect 91106 11320 91169 11406
rect 91169 11320 91255 11406
rect 91255 11320 91337 11406
rect 91337 11320 91423 11406
rect 91423 11320 91486 11406
rect 91106 11286 91486 11320
rect 91106 7603 91486 7666
rect 91106 7517 91169 7603
rect 91169 7517 91255 7603
rect 91255 7517 91337 7603
rect 91337 7517 91423 7603
rect 91423 7517 91486 7603
rect 91106 7286 91486 7517
rect 91106 3286 91486 3666
rect 92346 36526 92726 36906
rect 92346 32526 92726 32906
rect 92346 28526 92726 28906
rect 92346 24526 92726 24906
rect 92346 20526 92726 20906
rect 92346 16526 92726 16906
rect 92346 12526 92726 12906
rect 92346 8526 92726 8906
rect 92346 4526 92726 4906
rect 95106 35286 95486 35666
rect 95106 31286 95486 31666
rect 95106 27656 95169 27666
rect 95169 27656 95255 27666
rect 95255 27656 95337 27666
rect 95337 27656 95423 27666
rect 95423 27656 95486 27666
rect 95106 27574 95486 27656
rect 95106 27488 95169 27574
rect 95169 27488 95255 27574
rect 95255 27488 95337 27574
rect 95337 27488 95423 27574
rect 95423 27488 95486 27574
rect 95106 27406 95486 27488
rect 95106 27320 95169 27406
rect 95169 27320 95255 27406
rect 95255 27320 95337 27406
rect 95337 27320 95423 27406
rect 95423 27320 95486 27406
rect 95106 27286 95486 27320
rect 95106 23286 95486 23666
rect 95106 19613 95169 19666
rect 95169 19613 95255 19666
rect 95255 19613 95337 19666
rect 95337 19613 95423 19666
rect 95423 19613 95486 19666
rect 95106 19286 95486 19613
rect 95106 15286 95486 15666
rect 95106 11656 95169 11666
rect 95169 11656 95255 11666
rect 95255 11656 95337 11666
rect 95337 11656 95423 11666
rect 95423 11656 95486 11666
rect 95106 11574 95486 11656
rect 95106 11488 95169 11574
rect 95169 11488 95255 11574
rect 95255 11488 95337 11574
rect 95337 11488 95423 11574
rect 95423 11488 95486 11574
rect 95106 11406 95486 11488
rect 95106 11320 95169 11406
rect 95169 11320 95255 11406
rect 95255 11320 95337 11406
rect 95337 11320 95423 11406
rect 95423 11320 95486 11406
rect 95106 11286 95486 11320
rect 95106 7603 95486 7666
rect 95106 7517 95169 7603
rect 95169 7517 95255 7603
rect 95255 7517 95337 7603
rect 95337 7517 95423 7603
rect 95423 7517 95486 7603
rect 95106 7286 95486 7517
rect 95106 3286 95486 3666
rect 96346 36526 96726 36906
rect 96346 32526 96726 32906
rect 96346 28526 96726 28906
rect 96346 24526 96726 24906
rect 96346 20526 96726 20906
rect 96346 16526 96726 16906
rect 96346 12526 96726 12906
rect 96346 8526 96726 8906
rect 96346 4526 96726 4906
rect 99106 35286 99486 35666
rect 99106 31286 99486 31666
rect 99106 27286 99486 27666
rect 99106 23286 99486 23666
rect 99106 19613 99169 19666
rect 99169 19613 99255 19666
rect 99255 19613 99337 19666
rect 99337 19613 99423 19666
rect 99423 19613 99486 19666
rect 99106 19286 99486 19613
rect 99106 15286 99486 15666
rect 99106 11286 99486 11666
rect 99106 7603 99486 7666
rect 99106 7517 99169 7603
rect 99169 7517 99255 7603
rect 99255 7517 99337 7603
rect 99337 7517 99423 7603
rect 99423 7517 99486 7603
rect 99106 7286 99486 7517
rect 99106 3286 99486 3666
<< metal7 >>
rect 532 36906 99404 36936
rect 532 36526 4346 36906
rect 4726 36526 8346 36906
rect 8726 36526 12346 36906
rect 12726 36526 16346 36906
rect 16726 36526 20346 36906
rect 20726 36526 24346 36906
rect 24726 36526 28346 36906
rect 28726 36526 32346 36906
rect 32726 36526 36346 36906
rect 36726 36526 40346 36906
rect 40726 36526 44346 36906
rect 44726 36526 48346 36906
rect 48726 36526 52346 36906
rect 52726 36526 56346 36906
rect 56726 36526 60346 36906
rect 60726 36526 64346 36906
rect 64726 36526 68346 36906
rect 68726 36526 72346 36906
rect 72726 36526 76346 36906
rect 76726 36526 80346 36906
rect 80726 36526 84346 36906
rect 84726 36526 88346 36906
rect 88726 36526 92346 36906
rect 92726 36526 96346 36906
rect 96726 36526 99404 36906
rect 532 36496 99404 36526
rect 532 35666 99516 35696
rect 532 35286 3106 35666
rect 3486 35286 7106 35666
rect 7486 35286 11106 35666
rect 11486 35286 15106 35666
rect 15486 35286 19106 35666
rect 19486 35286 23106 35666
rect 23486 35286 27106 35666
rect 27486 35286 31106 35666
rect 31486 35286 35106 35666
rect 35486 35286 39106 35666
rect 39486 35286 43106 35666
rect 43486 35286 47106 35666
rect 47486 35286 51106 35666
rect 51486 35286 55106 35666
rect 55486 35286 59106 35666
rect 59486 35286 63106 35666
rect 63486 35286 67106 35666
rect 67486 35286 71106 35666
rect 71486 35286 75106 35666
rect 75486 35286 79106 35666
rect 79486 35286 83106 35666
rect 83486 35286 87106 35666
rect 87486 35286 91106 35666
rect 91486 35286 95106 35666
rect 95486 35286 99106 35666
rect 99486 35286 99516 35666
rect 532 35256 99516 35286
rect 532 32906 99404 32936
rect 532 32526 4346 32906
rect 4726 32526 8346 32906
rect 8726 32526 12346 32906
rect 12726 32526 16346 32906
rect 16726 32526 20346 32906
rect 20726 32526 24346 32906
rect 24726 32526 28346 32906
rect 28726 32526 32346 32906
rect 32726 32526 36346 32906
rect 36726 32526 40346 32906
rect 40726 32526 44346 32906
rect 44726 32526 48346 32906
rect 48726 32526 52346 32906
rect 52726 32526 56346 32906
rect 56726 32526 60346 32906
rect 60726 32526 64346 32906
rect 64726 32526 68346 32906
rect 68726 32526 72346 32906
rect 72726 32526 76346 32906
rect 76726 32526 80346 32906
rect 80726 32526 84346 32906
rect 84726 32526 88346 32906
rect 88726 32526 92346 32906
rect 92726 32526 96346 32906
rect 96726 32526 99404 32906
rect 532 32496 99404 32526
rect 532 31666 99516 31696
rect 532 31286 3106 31666
rect 3486 31286 7106 31666
rect 7486 31286 11106 31666
rect 11486 31286 15106 31666
rect 15486 31286 19106 31666
rect 19486 31286 23106 31666
rect 23486 31286 27106 31666
rect 27486 31286 31106 31666
rect 31486 31286 35106 31666
rect 35486 31286 39106 31666
rect 39486 31286 43106 31666
rect 43486 31286 47106 31666
rect 47486 31286 51106 31666
rect 51486 31286 55106 31666
rect 55486 31286 59106 31666
rect 59486 31286 63106 31666
rect 63486 31286 67106 31666
rect 67486 31286 71106 31666
rect 71486 31286 75106 31666
rect 75486 31286 79106 31666
rect 79486 31286 83106 31666
rect 83486 31286 87106 31666
rect 87486 31286 91106 31666
rect 91486 31286 95106 31666
rect 95486 31286 99106 31666
rect 99486 31286 99516 31666
rect 532 31256 99516 31286
rect 532 28906 99404 28936
rect 532 28526 4346 28906
rect 4726 28526 8346 28906
rect 8726 28526 12346 28906
rect 12726 28526 16346 28906
rect 16726 28526 20346 28906
rect 20726 28526 24346 28906
rect 24726 28526 28346 28906
rect 28726 28526 32346 28906
rect 32726 28526 36346 28906
rect 36726 28526 40346 28906
rect 40726 28526 44346 28906
rect 44726 28526 48346 28906
rect 48726 28526 52346 28906
rect 52726 28526 56346 28906
rect 56726 28526 60346 28906
rect 60726 28526 64346 28906
rect 64726 28526 68346 28906
rect 68726 28526 72346 28906
rect 72726 28526 76346 28906
rect 76726 28526 80346 28906
rect 80726 28526 84346 28906
rect 84726 28526 88346 28906
rect 88726 28526 92346 28906
rect 92726 28526 96346 28906
rect 96726 28526 99404 28906
rect 532 28496 99404 28526
rect 532 27666 99516 27696
rect 532 27286 3106 27666
rect 3486 27286 7106 27666
rect 7486 27286 11106 27666
rect 11486 27286 15106 27666
rect 15486 27286 19106 27666
rect 19486 27286 23106 27666
rect 23486 27286 27106 27666
rect 27486 27286 31106 27666
rect 31486 27286 35106 27666
rect 35486 27286 39106 27666
rect 39486 27286 43106 27666
rect 43486 27286 47106 27666
rect 47486 27286 51106 27666
rect 51486 27286 55106 27666
rect 55486 27286 59106 27666
rect 59486 27286 63106 27666
rect 63486 27286 67106 27666
rect 67486 27286 71106 27666
rect 71486 27286 75106 27666
rect 75486 27286 79106 27666
rect 79486 27286 83106 27666
rect 83486 27286 87106 27666
rect 87486 27286 91106 27666
rect 91486 27286 95106 27666
rect 95486 27286 99106 27666
rect 99486 27286 99516 27666
rect 532 27256 99516 27286
rect 532 24906 99404 24936
rect 532 24526 4346 24906
rect 4726 24526 8346 24906
rect 8726 24526 12346 24906
rect 12726 24526 16346 24906
rect 16726 24526 20346 24906
rect 20726 24526 24346 24906
rect 24726 24526 28346 24906
rect 28726 24526 32346 24906
rect 32726 24526 36346 24906
rect 36726 24526 40346 24906
rect 40726 24526 44346 24906
rect 44726 24526 48346 24906
rect 48726 24526 52346 24906
rect 52726 24526 56346 24906
rect 56726 24526 60346 24906
rect 60726 24526 64346 24906
rect 64726 24526 68346 24906
rect 68726 24526 72346 24906
rect 72726 24526 76346 24906
rect 76726 24526 80346 24906
rect 80726 24526 84346 24906
rect 84726 24526 88346 24906
rect 88726 24526 92346 24906
rect 92726 24526 96346 24906
rect 96726 24526 99404 24906
rect 532 24496 99404 24526
rect 532 23666 99516 23696
rect 532 23286 3106 23666
rect 3486 23286 7106 23666
rect 7486 23286 11106 23666
rect 11486 23286 15106 23666
rect 15486 23286 19106 23666
rect 19486 23286 23106 23666
rect 23486 23286 27106 23666
rect 27486 23286 31106 23666
rect 31486 23286 35106 23666
rect 35486 23286 39106 23666
rect 39486 23286 43106 23666
rect 43486 23286 47106 23666
rect 47486 23286 51106 23666
rect 51486 23286 55106 23666
rect 55486 23286 59106 23666
rect 59486 23286 63106 23666
rect 63486 23286 67106 23666
rect 67486 23286 71106 23666
rect 71486 23286 75106 23666
rect 75486 23286 79106 23666
rect 79486 23286 83106 23666
rect 83486 23286 87106 23666
rect 87486 23286 91106 23666
rect 91486 23286 95106 23666
rect 95486 23286 99106 23666
rect 99486 23286 99516 23666
rect 532 23256 99516 23286
rect 532 20906 99404 20936
rect 532 20526 4346 20906
rect 4726 20526 8346 20906
rect 8726 20526 12346 20906
rect 12726 20526 16346 20906
rect 16726 20526 20346 20906
rect 20726 20526 24346 20906
rect 24726 20526 28346 20906
rect 28726 20526 32346 20906
rect 32726 20526 36346 20906
rect 36726 20526 40346 20906
rect 40726 20526 44346 20906
rect 44726 20526 48346 20906
rect 48726 20526 52346 20906
rect 52726 20526 56346 20906
rect 56726 20526 60346 20906
rect 60726 20526 64346 20906
rect 64726 20526 68346 20906
rect 68726 20526 72346 20906
rect 72726 20526 76346 20906
rect 76726 20526 80346 20906
rect 80726 20526 84346 20906
rect 84726 20526 88346 20906
rect 88726 20526 92346 20906
rect 92726 20526 96346 20906
rect 96726 20526 99404 20906
rect 532 20496 99404 20526
rect 532 19666 99516 19696
rect 532 19286 3106 19666
rect 3486 19286 7106 19666
rect 7486 19286 11106 19666
rect 11486 19286 15106 19666
rect 15486 19286 19106 19666
rect 19486 19286 23106 19666
rect 23486 19286 27106 19666
rect 27486 19286 31106 19666
rect 31486 19286 35106 19666
rect 35486 19286 39106 19666
rect 39486 19286 43106 19666
rect 43486 19286 47106 19666
rect 47486 19286 51106 19666
rect 51486 19286 55106 19666
rect 55486 19286 59106 19666
rect 59486 19286 63106 19666
rect 63486 19286 67106 19666
rect 67486 19286 71106 19666
rect 71486 19286 75106 19666
rect 75486 19286 79106 19666
rect 79486 19286 83106 19666
rect 83486 19286 87106 19666
rect 87486 19286 91106 19666
rect 91486 19286 95106 19666
rect 95486 19286 99106 19666
rect 99486 19286 99516 19666
rect 532 19256 99516 19286
rect 532 16906 99404 16936
rect 532 16526 4346 16906
rect 4726 16526 8346 16906
rect 8726 16526 12346 16906
rect 12726 16526 16346 16906
rect 16726 16526 20346 16906
rect 20726 16526 24346 16906
rect 24726 16526 28346 16906
rect 28726 16526 32346 16906
rect 32726 16526 36346 16906
rect 36726 16526 40346 16906
rect 40726 16526 44346 16906
rect 44726 16526 48346 16906
rect 48726 16526 52346 16906
rect 52726 16526 56346 16906
rect 56726 16526 60346 16906
rect 60726 16526 64346 16906
rect 64726 16526 68346 16906
rect 68726 16526 72346 16906
rect 72726 16526 76346 16906
rect 76726 16526 80346 16906
rect 80726 16526 84346 16906
rect 84726 16526 88346 16906
rect 88726 16526 92346 16906
rect 92726 16526 96346 16906
rect 96726 16526 99404 16906
rect 532 16496 99404 16526
rect 532 15666 99516 15696
rect 532 15286 3106 15666
rect 3486 15286 7106 15666
rect 7486 15286 11106 15666
rect 11486 15286 15106 15666
rect 15486 15286 19106 15666
rect 19486 15286 23106 15666
rect 23486 15286 27106 15666
rect 27486 15286 31106 15666
rect 31486 15286 35106 15666
rect 35486 15286 39106 15666
rect 39486 15286 43106 15666
rect 43486 15286 47106 15666
rect 47486 15286 51106 15666
rect 51486 15286 55106 15666
rect 55486 15286 59106 15666
rect 59486 15286 63106 15666
rect 63486 15286 67106 15666
rect 67486 15286 71106 15666
rect 71486 15286 75106 15666
rect 75486 15286 79106 15666
rect 79486 15286 83106 15666
rect 83486 15286 87106 15666
rect 87486 15286 91106 15666
rect 91486 15286 95106 15666
rect 95486 15286 99106 15666
rect 99486 15286 99516 15666
rect 532 15256 99516 15286
rect 532 12906 99404 12936
rect 532 12526 4346 12906
rect 4726 12526 8346 12906
rect 8726 12526 12346 12906
rect 12726 12526 16346 12906
rect 16726 12526 20346 12906
rect 20726 12526 24346 12906
rect 24726 12526 28346 12906
rect 28726 12526 32346 12906
rect 32726 12526 36346 12906
rect 36726 12526 40346 12906
rect 40726 12526 44346 12906
rect 44726 12526 48346 12906
rect 48726 12526 52346 12906
rect 52726 12526 56346 12906
rect 56726 12526 60346 12906
rect 60726 12526 64346 12906
rect 64726 12526 68346 12906
rect 68726 12526 72346 12906
rect 72726 12526 76346 12906
rect 76726 12526 80346 12906
rect 80726 12526 84346 12906
rect 84726 12526 88346 12906
rect 88726 12526 92346 12906
rect 92726 12526 96346 12906
rect 96726 12526 99404 12906
rect 532 12496 99404 12526
rect 532 11666 99516 11696
rect 532 11286 3106 11666
rect 3486 11286 7106 11666
rect 7486 11286 11106 11666
rect 11486 11286 15106 11666
rect 15486 11286 19106 11666
rect 19486 11286 23106 11666
rect 23486 11286 27106 11666
rect 27486 11286 31106 11666
rect 31486 11286 35106 11666
rect 35486 11286 39106 11666
rect 39486 11286 43106 11666
rect 43486 11286 47106 11666
rect 47486 11286 51106 11666
rect 51486 11286 55106 11666
rect 55486 11286 59106 11666
rect 59486 11286 63106 11666
rect 63486 11286 67106 11666
rect 67486 11286 71106 11666
rect 71486 11286 75106 11666
rect 75486 11286 79106 11666
rect 79486 11286 83106 11666
rect 83486 11286 87106 11666
rect 87486 11286 91106 11666
rect 91486 11286 95106 11666
rect 95486 11286 99106 11666
rect 99486 11286 99516 11666
rect 532 11256 99516 11286
rect 532 8906 99404 8936
rect 532 8526 4346 8906
rect 4726 8526 8346 8906
rect 8726 8526 12346 8906
rect 12726 8526 16346 8906
rect 16726 8526 20346 8906
rect 20726 8526 24346 8906
rect 24726 8526 28346 8906
rect 28726 8526 32346 8906
rect 32726 8526 36346 8906
rect 36726 8526 40346 8906
rect 40726 8526 44346 8906
rect 44726 8526 48346 8906
rect 48726 8526 52346 8906
rect 52726 8526 56346 8906
rect 56726 8526 60346 8906
rect 60726 8526 64346 8906
rect 64726 8526 68346 8906
rect 68726 8526 72346 8906
rect 72726 8526 76346 8906
rect 76726 8526 80346 8906
rect 80726 8526 84346 8906
rect 84726 8526 88346 8906
rect 88726 8526 92346 8906
rect 92726 8526 96346 8906
rect 96726 8526 99404 8906
rect 532 8496 99404 8526
rect 532 7666 99516 7696
rect 532 7286 3106 7666
rect 3486 7286 7106 7666
rect 7486 7286 11106 7666
rect 11486 7286 15106 7666
rect 15486 7286 19106 7666
rect 19486 7286 23106 7666
rect 23486 7286 27106 7666
rect 27486 7286 31106 7666
rect 31486 7286 35106 7666
rect 35486 7286 39106 7666
rect 39486 7286 43106 7666
rect 43486 7286 47106 7666
rect 47486 7286 51106 7666
rect 51486 7286 55106 7666
rect 55486 7286 59106 7666
rect 59486 7286 63106 7666
rect 63486 7286 67106 7666
rect 67486 7286 71106 7666
rect 71486 7286 75106 7666
rect 75486 7286 79106 7666
rect 79486 7286 83106 7666
rect 83486 7286 87106 7666
rect 87486 7286 91106 7666
rect 91486 7286 95106 7666
rect 95486 7286 99106 7666
rect 99486 7286 99516 7666
rect 532 7256 99516 7286
rect 532 4906 99404 4936
rect 532 4526 4346 4906
rect 4726 4526 8346 4906
rect 8726 4526 12346 4906
rect 12726 4526 16346 4906
rect 16726 4526 20346 4906
rect 20726 4526 24346 4906
rect 24726 4526 28346 4906
rect 28726 4526 32346 4906
rect 32726 4526 36346 4906
rect 36726 4526 40346 4906
rect 40726 4526 44346 4906
rect 44726 4526 48346 4906
rect 48726 4526 52346 4906
rect 52726 4526 56346 4906
rect 56726 4526 60346 4906
rect 60726 4526 64346 4906
rect 64726 4526 68346 4906
rect 68726 4526 72346 4906
rect 72726 4526 76346 4906
rect 76726 4526 80346 4906
rect 80726 4526 84346 4906
rect 84726 4526 88346 4906
rect 88726 4526 92346 4906
rect 92726 4526 96346 4906
rect 96726 4526 99404 4906
rect 532 4496 99404 4526
rect 532 3666 99516 3696
rect 532 3286 3106 3666
rect 3486 3286 7106 3666
rect 7486 3286 11106 3666
rect 11486 3286 15106 3666
rect 15486 3286 19106 3666
rect 19486 3286 23106 3666
rect 23486 3286 27106 3666
rect 27486 3286 31106 3666
rect 31486 3286 35106 3666
rect 35486 3286 39106 3666
rect 39486 3286 43106 3666
rect 43486 3286 47106 3666
rect 47486 3286 51106 3666
rect 51486 3286 55106 3666
rect 55486 3286 59106 3666
rect 59486 3286 63106 3666
rect 63486 3286 67106 3666
rect 67486 3286 71106 3666
rect 71486 3286 75106 3666
rect 75486 3286 79106 3666
rect 79486 3286 83106 3666
rect 83486 3286 87106 3666
rect 87486 3286 91106 3666
rect 91486 3286 95106 3666
rect 95486 3286 99106 3666
rect 99486 3286 99516 3666
rect 532 3256 99516 3286
use sg13g2_buf_1  _08_
timestamp 1676381911
transform -1 0 1920 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _09_
timestamp 1676381911
transform -1 0 2304 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _10_
timestamp 1676381911
transform -1 0 2016 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _11_
timestamp 1676381911
transform -1 0 1632 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _12_
timestamp 1676381911
transform -1 0 2016 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _13_
timestamp 1676381911
transform -1 0 2304 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _14_
timestamp 1676381911
transform -1 0 1536 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _15_
timestamp 1676381911
transform -1 0 1920 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _16_
timestamp 1676381911
transform -1 0 1728 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _17_
timestamp 1676381911
transform -1 0 2112 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _18_
timestamp 1676381911
transform -1 0 1632 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _19_
timestamp 1676381911
transform -1 0 1824 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _20_
timestamp 1676381911
transform -1 0 1728 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _21_
timestamp 1676381911
transform -1 0 1632 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _22_
timestamp 1676381911
transform -1 0 1632 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _23_
timestamp 1676381911
transform -1 0 1728 0 -1 11340
box -48 -56 432 834
use dac128module  dacH
timestamp 0
transform 1 0 72000 0 1 26014
box 0 0 1 1
use dac128module  dacL
timestamp 0
transform 1 0 72000 0 1 10014
box 0 0 1 1
use sg13g2_buf_1  digitalenH.g\[0\].u.buff
timestamp 1676381911
transform 1 0 69312 0 -1 26460
box -48 -56 432 834
use sg13g2_inv_1  digitalenH.g\[0\].u.inv
timestamp 1676382929
transform 1 0 69024 0 -1 26460
box -48 -56 336 834
use sg13g2_buf_1  digitalenH.g\[1\].u.buff
timestamp 1676381911
transform -1 0 98784 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalenH.g\[1\].u.inv
timestamp 1676382929
transform -1 0 99072 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalenH.g\[2\].u.buff
timestamp 1676381911
transform -1 0 98784 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalenH.g\[2\].u.inv
timestamp 1676382929
transform 1 0 99072 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalenH.g\[3\].u.buff
timestamp 1676381911
transform 1 0 69312 0 1 30996
box -48 -56 432 834
use sg13g2_inv_1  digitalenH.g\[3\].u.inv
timestamp 1676382929
transform 1 0 69504 0 -1 30996
box -48 -56 336 834
use sg13g2_buf_1  digitalenL.g\[0\].u.buff
timestamp 1676381911
transform 1 0 69312 0 -1 9828
box -48 -56 432 834
use sg13g2_inv_1  digitalenL.g\[0\].u.inv
timestamp 1676382929
transform 1 0 69696 0 -1 9828
box -48 -56 336 834
use sg13g2_buf_1  digitalenL.g\[1\].u.buff
timestamp 1676381911
transform -1 0 98784 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalenL.g\[1\].u.inv
timestamp 1676382929
transform 1 0 98592 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalenL.g\[2\].u.buff
timestamp 1676381911
transform 1 0 96864 0 -1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalenL.g\[2\].u.inv
timestamp 1676382929
transform -1 0 98496 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalenL.g\[3\].u.buff
timestamp 1676381911
transform 1 0 69120 0 -1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalenL.g\[3\].u.inv
timestamp 1676382929
transform 1 0 68928 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[0\].u.buff
timestamp 1676381911
transform 1 0 68736 0 -1 27972
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[0\].u.inv
timestamp 1676382929
transform -1 0 68736 0 -1 26460
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[1\].u.buff
timestamp 1676381911
transform 1 0 69600 0 1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[1\].u.inv
timestamp 1676382929
transform 1 0 68736 0 -1 26460
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[2\].u.buff
timestamp 1676381911
transform 1 0 69408 0 1 26460
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[2\].u.inv
timestamp 1676382929
transform 1 0 73248 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[3\].u.buff
timestamp 1676381911
transform 1 0 67680 0 -1 26460
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[3\].u.inv
timestamp 1676382929
transform 1 0 69696 0 -1 26460
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[4\].u.buff
timestamp 1676381911
transform 1 0 68544 0 1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[4\].u.inv
timestamp 1676382929
transform 1 0 73728 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[5\].u.buff
timestamp 1676381911
transform -1 0 74880 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[5\].u.inv
timestamp 1676382929
transform 1 0 72960 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[6\].u.buff
timestamp 1676381911
transform 1 0 74688 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[6\].u.inv
timestamp 1676382929
transform -1 0 67680 0 -1 26460
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[7\].u.buff
timestamp 1676381911
transform -1 0 75840 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[7\].u.inv
timestamp 1676382929
transform -1 0 74304 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[8\].u.buff
timestamp 1676381911
transform -1 0 76224 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[8\].u.inv
timestamp 1676382929
transform 1 0 75648 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[9\].u.buff
timestamp 1676381911
transform 1 0 76032 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[9\].u.inv
timestamp 1676382929
transform 1 0 75744 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[10\].u.buff
timestamp 1676381911
transform 1 0 76512 0 -1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[10\].u.inv
timestamp 1676382929
transform 1 0 76512 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[11\].u.buff
timestamp 1676381911
transform 1 0 76800 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[11\].u.inv
timestamp 1676382929
transform 1 0 77088 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[12\].u.buff
timestamp 1676381911
transform 1 0 77184 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[12\].u.inv
timestamp 1676382929
transform 1 0 77472 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[13\].u.buff
timestamp 1676381911
transform 1 0 77664 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[13\].u.inv
timestamp 1676382929
transform -1 0 78240 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[14\].u.buff
timestamp 1676381911
transform 1 0 78048 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[14\].u.inv
timestamp 1676382929
transform -1 0 79392 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[15\].u.buff
timestamp 1676381911
transform 1 0 78336 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[15\].u.inv
timestamp 1676382929
transform 1 0 78720 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[16\].u.buff
timestamp 1676381911
transform 1 0 78816 0 -1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[16\].u.inv
timestamp 1676382929
transform -1 0 79680 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[17\].u.buff
timestamp 1676381911
transform 1 0 79200 0 -1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[17\].u.inv
timestamp 1676382929
transform 1 0 79680 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[18\].u.buff
timestamp 1676381911
transform 1 0 79488 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[18\].u.inv
timestamp 1676382929
transform -1 0 81120 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[19\].u.buff
timestamp 1676381911
transform 1 0 79872 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[19\].u.inv
timestamp 1676382929
transform -1 0 81408 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[20\].u.buff
timestamp 1676381911
transform 1 0 80352 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[20\].u.inv
timestamp 1676382929
transform -1 0 81024 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[21\].u.buff
timestamp 1676381911
transform 1 0 80736 0 -1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[21\].u.inv
timestamp 1676382929
transform -1 0 81696 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[22\].u.buff
timestamp 1676381911
transform 1 0 81216 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[22\].u.inv
timestamp 1676382929
transform -1 0 81984 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[23\].u.buff
timestamp 1676381911
transform 1 0 81600 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[23\].u.inv
timestamp 1676382929
transform -1 0 82272 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[24\].u.buff
timestamp 1676381911
transform 1 0 82080 0 -1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[24\].u.inv
timestamp 1676382929
transform -1 0 82752 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[25\].u.buff
timestamp 1676381911
transform 1 0 82368 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[25\].u.inv
timestamp 1676382929
transform 1 0 82752 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[26\].u.buff
timestamp 1676381911
transform -1 0 83328 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[26\].u.inv
timestamp 1676382929
transform -1 0 84192 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[27\].u.buff
timestamp 1676381911
transform 1 0 83328 0 -1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[27\].u.inv
timestamp 1676382929
transform 1 0 83424 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[28\].u.buff
timestamp 1676381911
transform 1 0 83712 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[28\].u.inv
timestamp 1676382929
transform -1 0 84384 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[29\].u.buff
timestamp 1676381911
transform 1 0 84096 0 -1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[29\].u.inv
timestamp 1676382929
transform 1 0 84288 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[30\].u.buff
timestamp 1676381911
transform 1 0 84480 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[30\].u.inv
timestamp 1676382929
transform 1 0 84672 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[31\].u.buff
timestamp 1676381911
transform 1 0 84864 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[31\].u.inv
timestamp 1676382929
transform 1 0 85056 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[32\].u.buff
timestamp 1676381911
transform -1 0 85728 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[32\].u.inv
timestamp 1676382929
transform 1 0 85344 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[33\].u.buff
timestamp 1676381911
transform 1 0 85728 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[33\].u.inv
timestamp 1676382929
transform 1 0 85824 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[34\].u.buff
timestamp 1676381911
transform 1 0 86016 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[34\].u.inv
timestamp 1676382929
transform -1 0 86592 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[35\].u.buff
timestamp 1676381911
transform 1 0 86496 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[35\].u.inv
timestamp 1676382929
transform 1 0 86688 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[36\].u.buff
timestamp 1676381911
transform 1 0 86880 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[36\].u.inv
timestamp 1676382929
transform -1 0 87936 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[37\].u.buff
timestamp 1676381911
transform 1 0 87168 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[37\].u.inv
timestamp 1676382929
transform 1 0 86880 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[38\].u.buff
timestamp 1676381911
transform 1 0 87552 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[38\].u.inv
timestamp 1676382929
transform -1 0 88224 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[39\].u.buff
timestamp 1676381911
transform 1 0 87936 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[39\].u.inv
timestamp 1676382929
transform -1 0 88608 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[40\].u.buff
timestamp 1676381911
transform 1 0 88320 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[40\].u.inv
timestamp 1676382929
transform 1 0 88704 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[41\].u.buff
timestamp 1676381911
transform 1 0 88800 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[41\].u.inv
timestamp 1676382929
transform -1 0 89280 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[42\].u.buff
timestamp 1676381911
transform 1 0 89280 0 -1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[42\].u.inv
timestamp 1676382929
transform -1 0 89568 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[43\].u.buff
timestamp 1676381911
transform 1 0 89664 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[43\].u.inv
timestamp 1676382929
transform -1 0 90720 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[44\].u.buff
timestamp 1676381911
transform -1 0 90528 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[44\].u.inv
timestamp 1676382929
transform -1 0 91008 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[45\].u.buff
timestamp 1676381911
transform 1 0 90528 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[45\].u.inv
timestamp 1676382929
transform -1 0 91296 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[46\].u.buff
timestamp 1676381911
transform -1 0 91968 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[46\].u.inv
timestamp 1676382929
transform 1 0 91008 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[47\].u.buff
timestamp 1676381911
transform 1 0 91200 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[47\].u.inv
timestamp 1676382929
transform 1 0 90912 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[48\].u.buff
timestamp 1676381911
transform -1 0 92352 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[48\].u.inv
timestamp 1676382929
transform 1 0 91296 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[49\].u.buff
timestamp 1676381911
transform -1 0 92736 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[49\].u.inv
timestamp 1676382929
transform -1 0 93888 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[50\].u.buff
timestamp 1676381911
transform -1 0 93120 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[50\].u.inv
timestamp 1676382929
transform 1 0 92640 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[51\].u.buff
timestamp 1676381911
transform 1 0 92832 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[51\].u.inv
timestamp 1676382929
transform -1 0 93504 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[52\].u.buff
timestamp 1676381911
transform 1 0 93216 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[52\].u.inv
timestamp 1676382929
transform -1 0 94176 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[53\].u.buff
timestamp 1676381911
transform 1 0 93696 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[53\].u.inv
timestamp 1676382929
transform 1 0 93408 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[54\].u.buff
timestamp 1676381911
transform 1 0 94080 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[54\].u.inv
timestamp 1676382929
transform 1 0 94464 0 1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[55\].u.buff
timestamp 1676381911
transform 1 0 94368 0 -1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[55\].u.inv
timestamp 1676382929
transform -1 0 95040 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[56\].u.buff
timestamp 1676381911
transform 1 0 94848 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[56\].u.inv
timestamp 1676382929
transform -1 0 95424 0 -1 21924
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[57\].u.buff
timestamp 1676381911
transform 1 0 95232 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[57\].u.inv
timestamp 1676382929
transform 1 0 95232 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[58\].u.buff
timestamp 1676381911
transform 1 0 95616 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[58\].u.inv
timestamp 1676382929
transform -1 0 96672 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[59\].u.buff
timestamp 1676381911
transform 1 0 96000 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[59\].u.inv
timestamp 1676382929
transform -1 0 96960 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[60\].u.buff
timestamp 1676381911
transform 1 0 96480 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[60\].u.inv
timestamp 1676382929
transform -1 0 97248 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[61\].u.buff
timestamp 1676381911
transform -1 0 97344 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[61\].u.inv
timestamp 1676382929
transform -1 0 97536 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[62\].u.buff
timestamp 1676381911
transform -1 0 97920 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[62\].u.inv
timestamp 1676382929
transform -1 0 97920 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[63\].u.buff
timestamp 1676381911
transform -1 0 98304 0 1 21924
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[63\].u.inv
timestamp 1676382929
transform -1 0 98304 0 -1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[64\].u.buff
timestamp 1676381911
transform 1 0 97728 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[64\].u.inv
timestamp 1676382929
transform 1 0 98784 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[65\].u.buff
timestamp 1676381911
transform 1 0 97440 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[65\].u.inv
timestamp 1676382929
transform -1 0 98400 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[66\].u.buff
timestamp 1676381911
transform 1 0 96960 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[66\].u.inv
timestamp 1676382929
transform 1 0 96672 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[67\].u.buff
timestamp 1676381911
transform 1 0 96480 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[67\].u.inv
timestamp 1676382929
transform 1 0 97824 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[68\].u.buff
timestamp 1676381911
transform 1 0 96096 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[68\].u.inv
timestamp 1676382929
transform -1 0 97152 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[69\].u.buff
timestamp 1676381911
transform 1 0 95712 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[69\].u.inv
timestamp 1676382929
transform -1 0 95328 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[70\].u.buff
timestamp 1676381911
transform 1 0 95328 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[70\].u.inv
timestamp 1676382929
transform -1 0 95712 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[71\].u.buff
timestamp 1676381911
transform 1 0 94944 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[71\].u.inv
timestamp 1676382929
transform 1 0 94848 0 1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[72\].u.buff
timestamp 1676381911
transform 1 0 94560 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[72\].u.inv
timestamp 1676382929
transform -1 0 94944 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[73\].u.buff
timestamp 1676381911
transform -1 0 94656 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[73\].u.inv
timestamp 1676382929
transform 1 0 94176 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[74\].u.buff
timestamp 1676381911
transform 1 0 93792 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[74\].u.inv
timestamp 1676382929
transform -1 0 94080 0 1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[75\].u.buff
timestamp 1676381911
transform 1 0 93312 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[75\].u.inv
timestamp 1676382929
transform 1 0 93024 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[76\].u.buff
timestamp 1676381911
transform 1 0 93024 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[76\].u.inv
timestamp 1676382929
transform -1 0 93696 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[77\].u.buff
timestamp 1676381911
transform 1 0 92544 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[77\].u.inv
timestamp 1676382929
transform -1 0 92160 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[78\].u.buff
timestamp 1676381911
transform 1 0 92160 0 1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[78\].u.inv
timestamp 1676382929
transform 1 0 92160 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[79\].u.buff
timestamp 1676381911
transform 1 0 91680 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[79\].u.inv
timestamp 1676382929
transform 1 0 91392 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[80\].u.buff
timestamp 1676381911
transform 1 0 90624 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[80\].u.inv
timestamp 1676382929
transform -1 0 91872 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[81\].u.buff
timestamp 1676381911
transform 1 0 91008 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[81\].u.inv
timestamp 1676382929
transform -1 0 91584 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[82\].u.buff
timestamp 1676381911
transform 1 0 90432 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[82\].u.inv
timestamp 1676382929
transform 1 0 90144 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[83\].u.buff
timestamp 1676381911
transform 1 0 90144 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[83\].u.inv
timestamp 1676382929
transform 1 0 90144 0 1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[84\].u.buff
timestamp 1676381911
transform 1 0 89760 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[84\].u.inv
timestamp 1676382929
transform 1 0 89760 0 1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[85\].u.buff
timestamp 1676381911
transform 1 0 89376 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[85\].u.inv
timestamp 1676382929
transform -1 0 90048 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[86\].u.buff
timestamp 1676381911
transform 1 0 88992 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[86\].u.inv
timestamp 1676382929
transform -1 0 89760 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[87\].u.buff
timestamp 1676381911
transform 1 0 88608 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[87\].u.inv
timestamp 1676382929
transform 1 0 88608 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[88\].u.buff
timestamp 1676381911
transform 1 0 88224 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[88\].u.inv
timestamp 1676382929
transform -1 0 87840 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[89\].u.buff
timestamp 1676381911
transform 1 0 87744 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[89\].u.inv
timestamp 1676382929
transform 1 0 87744 0 1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[90\].u.buff
timestamp 1676381911
transform -1 0 88608 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[90\].u.inv
timestamp 1676382929
transform 1 0 87264 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[91\].u.buff
timestamp 1676381911
transform -1 0 87552 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[91\].u.inv
timestamp 1676382929
transform 1 0 86976 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[92\].u.buff
timestamp 1676381911
transform -1 0 87168 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[92\].u.inv
timestamp 1676382929
transform 1 0 86496 0 1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[93\].u.buff
timestamp 1676381911
transform 1 0 86016 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[93\].u.inv
timestamp 1676382929
transform -1 0 86976 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[94\].u.buff
timestamp 1676381911
transform 1 0 85728 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[94\].u.inv
timestamp 1676382929
transform 1 0 85728 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[95\].u.buff
timestamp 1676381911
transform 1 0 85344 0 1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[95\].u.inv
timestamp 1676382929
transform 1 0 85344 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[96\].u.buff
timestamp 1676381911
transform 1 0 84960 0 1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[96\].u.inv
timestamp 1676382929
transform 1 0 84960 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[97\].u.buff
timestamp 1676381911
transform 1 0 84576 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[97\].u.inv
timestamp 1676382929
transform -1 0 84576 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[98\].u.buff
timestamp 1676381911
transform 1 0 84192 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[98\].u.inv
timestamp 1676382929
transform 1 0 84576 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[99\].u.buff
timestamp 1676381911
transform 1 0 83808 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[99\].u.inv
timestamp 1676382929
transform -1 0 84288 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[100\].u.buff
timestamp 1676381911
transform 1 0 83424 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[100\].u.inv
timestamp 1676382929
transform -1 0 84000 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[101\].u.buff
timestamp 1676381911
transform -1 0 83424 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[101\].u.inv
timestamp 1676382929
transform -1 0 83712 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[102\].u.buff
timestamp 1676381911
transform 1 0 82560 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[102\].u.inv
timestamp 1676382929
transform 1 0 82272 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[103\].u.buff
timestamp 1676381911
transform 1 0 82176 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[103\].u.inv
timestamp 1676382929
transform 1 0 82560 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[104\].u.buff
timestamp 1676381911
transform 1 0 81696 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[104\].u.inv
timestamp 1676382929
transform 1 0 81120 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[105\].u.buff
timestamp 1676381911
transform 1 0 81312 0 1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[105\].u.inv
timestamp 1676382929
transform -1 0 81696 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[106\].u.buff
timestamp 1676381911
transform 1 0 80832 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[106\].u.inv
timestamp 1676382929
transform 1 0 80544 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[107\].u.buff
timestamp 1676381911
transform 1 0 80352 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[107\].u.inv
timestamp 1676382929
transform 1 0 80064 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[108\].u.buff
timestamp 1676381911
transform 1 0 80064 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[108\].u.inv
timestamp 1676382929
transform 1 0 80160 0 1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[109\].u.buff
timestamp 1676381911
transform 1 0 79680 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[109\].u.inv
timestamp 1676382929
transform 1 0 79680 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[110\].u.buff
timestamp 1676381911
transform 1 0 79296 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[110\].u.inv
timestamp 1676382929
transform 1 0 79296 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[111\].u.buff
timestamp 1676381911
transform -1 0 79488 0 1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[111\].u.inv
timestamp 1676382929
transform 1 0 78816 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[112\].u.buff
timestamp 1676381911
transform 1 0 78528 0 1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[112\].u.inv
timestamp 1676382929
transform 1 0 78432 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[113\].u.buff
timestamp 1676381911
transform 1 0 78144 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[113\].u.inv
timestamp 1676382929
transform -1 0 78816 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[114\].u.buff
timestamp 1676381911
transform 1 0 77760 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[114\].u.inv
timestamp 1676382929
transform 1 0 77472 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[115\].u.buff
timestamp 1676381911
transform 1 0 77376 0 1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[115\].u.inv
timestamp 1676382929
transform 1 0 76608 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[116\].u.buff
timestamp 1676381911
transform 1 0 76896 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[116\].u.inv
timestamp 1676382929
transform -1 0 77664 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[117\].u.buff
timestamp 1676381911
transform 1 0 76512 0 1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[117\].u.inv
timestamp 1676382929
transform 1 0 76608 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[118\].u.buff
timestamp 1676381911
transform 1 0 76128 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[118\].u.inv
timestamp 1676382929
transform 1 0 75840 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[119\].u.buff
timestamp 1676381911
transform 1 0 75552 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[119\].u.inv
timestamp 1676382929
transform -1 0 76224 0 -1 35532
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[120\].u.buff
timestamp 1676381911
transform 1 0 75072 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[120\].u.inv
timestamp 1676382929
transform -1 0 75744 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[121\].u.buff
timestamp 1676381911
transform 1 0 74784 0 1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[121\].u.inv
timestamp 1676382929
transform 1 0 74784 0 1 34020
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[122\].u.buff
timestamp 1676381911
transform 1 0 74016 0 -1 35532
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[122\].u.inv
timestamp 1676382929
transform 1 0 69696 0 -1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[123\].u.buff
timestamp 1676381911
transform 1 0 73824 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[123\].u.inv
timestamp 1676382929
transform 1 0 68448 0 -1 30996
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[124\].u.buff
timestamp 1676381911
transform 1 0 73344 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[124\].u.inv
timestamp 1676382929
transform -1 0 67392 0 1 30996
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[125\].u.buff
timestamp 1676381911
transform 1 0 67296 0 -1 30996
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[125\].u.inv
timestamp 1676382929
transform 1 0 69696 0 1 30996
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[126\].u.buff
timestamp 1676381911
transform 1 0 68544 0 1 30996
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[126\].u.inv
timestamp 1676382929
transform 1 0 69216 0 -1 30996
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[127\].u.buff
timestamp 1676381911
transform 1 0 68928 0 1 30996
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[127\].u.inv
timestamp 1676382929
transform 1 0 68928 0 -1 30996
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[0\].u.buff
timestamp 1676381911
transform 1 0 68928 0 -1 9828
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[0\].u.inv
timestamp 1676382929
transform -1 0 68448 0 1 9828
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[1\].u.buff
timestamp 1676381911
transform 1 0 68928 0 1 9828
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[1\].u.inv
timestamp 1676382929
transform 1 0 69600 0 1 9828
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[2\].u.buff
timestamp 1676381911
transform 1 0 67392 0 1 9828
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[2\].u.inv
timestamp 1676382929
transform 1 0 69312 0 1 9828
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[3\].u.buff
timestamp 1676381911
transform 1 0 69216 0 -1 11340
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[3\].u.inv
timestamp 1676382929
transform 1 0 73248 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[4\].u.buff
timestamp 1676381911
transform 1 0 73536 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[4\].u.inv
timestamp 1676382929
transform 1 0 69696 0 -1 11340
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[5\].u.buff
timestamp 1676381911
transform -1 0 75552 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[5\].u.inv
timestamp 1676382929
transform 1 0 74016 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[6\].u.buff
timestamp 1676381911
transform 1 0 74688 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[6\].u.inv
timestamp 1676382929
transform 1 0 75072 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[7\].u.buff
timestamp 1676381911
transform 1 0 75072 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[7\].u.inv
timestamp 1676382929
transform 1 0 75360 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[8\].u.buff
timestamp 1676381911
transform 1 0 75648 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[8\].u.inv
timestamp 1676382929
transform 1 0 75648 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[9\].u.buff
timestamp 1676381911
transform 1 0 76032 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[9\].u.inv
timestamp 1676382929
transform 1 0 76224 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[10\].u.buff
timestamp 1676381911
transform 1 0 76416 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[10\].u.inv
timestamp 1676382929
transform 1 0 76608 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[11\].u.buff
timestamp 1676381911
transform 1 0 76896 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[11\].u.inv
timestamp 1676382929
transform -1 0 76800 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[12\].u.buff
timestamp 1676381911
transform 1 0 76800 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[12\].u.inv
timestamp 1676382929
transform -1 0 78240 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[13\].u.buff
timestamp 1676381911
transform 1 0 77664 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[13\].u.inv
timestamp 1676382929
transform -1 0 78528 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[14\].u.buff
timestamp 1676381911
transform 1 0 78048 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[14\].u.inv
timestamp 1676382929
transform 1 0 78144 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[15\].u.buff
timestamp 1676381911
transform 1 0 78528 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[15\].u.inv
timestamp 1676382929
transform 1 0 78624 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[16\].u.buff
timestamp 1676381911
transform 1 0 78816 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[16\].u.inv
timestamp 1676382929
transform 1 0 79008 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[17\].u.buff
timestamp 1676381911
transform -1 0 79680 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[17\].u.inv
timestamp 1676382929
transform 1 0 79296 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[18\].u.buff
timestamp 1676381911
transform 1 0 79584 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[18\].u.inv
timestamp 1676382929
transform 1 0 79872 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[19\].u.buff
timestamp 1676381911
transform 1 0 79872 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[19\].u.inv
timestamp 1676382929
transform -1 0 80544 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[20\].u.buff
timestamp 1676381911
transform 1 0 80352 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[20\].u.inv
timestamp 1676382929
transform -1 0 81888 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[21\].u.buff
timestamp 1676381911
transform 1 0 80832 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[21\].u.inv
timestamp 1676382929
transform 1 0 81024 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[22\].u.buff
timestamp 1676381911
transform 1 0 81216 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[22\].u.inv
timestamp 1676382929
transform 1 0 81888 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[23\].u.buff
timestamp 1676381911
transform 1 0 81600 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[23\].u.inv
timestamp 1676382929
transform 1 0 81312 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[24\].u.buff
timestamp 1676381911
transform 1 0 81984 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[24\].u.inv
timestamp 1676382929
transform 1 0 82176 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[25\].u.buff
timestamp 1676381911
transform 1 0 82368 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[25\].u.inv
timestamp 1676382929
transform -1 0 83232 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[26\].u.buff
timestamp 1676381911
transform 1 0 82656 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[26\].u.inv
timestamp 1676382929
transform 1 0 83232 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[27\].u.buff
timestamp 1676381911
transform 1 0 83136 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[27\].u.inv
timestamp 1676382929
transform 1 0 83424 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[28\].u.buff
timestamp 1676381911
transform 1 0 83616 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[28\].u.inv
timestamp 1676382929
transform 1 0 83712 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[29\].u.buff
timestamp 1676381911
transform 1 0 84096 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[29\].u.inv
timestamp 1676382929
transform 1 0 85536 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[30\].u.buff
timestamp 1676381911
transform 1 0 84480 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[30\].u.inv
timestamp 1676382929
transform 1 0 84480 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[31\].u.buff
timestamp 1676381911
transform 1 0 84768 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[31\].u.inv
timestamp 1676382929
transform -1 0 85152 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[32\].u.buff
timestamp 1676381911
transform 1 0 85152 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[32\].u.inv
timestamp 1676382929
transform 1 0 85344 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[33\].u.buff
timestamp 1676381911
transform 1 0 85536 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[33\].u.inv
timestamp 1676382929
transform 1 0 86784 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[34\].u.buff
timestamp 1676381911
transform 1 0 86016 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[34\].u.inv
timestamp 1676382929
transform -1 0 87360 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[35\].u.buff
timestamp 1676381911
transform 1 0 86496 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[35\].u.inv
timestamp 1676382929
transform -1 0 87648 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[36\].u.buff
timestamp 1676381911
transform 1 0 86784 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[36\].u.inv
timestamp 1676382929
transform -1 0 87936 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[37\].u.buff
timestamp 1676381911
transform 1 0 87264 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[37\].u.inv
timestamp 1676382929
transform 1 0 87456 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[38\].u.buff
timestamp 1676381911
transform 1 0 87648 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[38\].u.inv
timestamp 1676382929
transform -1 0 89184 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[39\].u.buff
timestamp 1676381911
transform 1 0 88032 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[39\].u.inv
timestamp 1676382929
transform -1 0 88704 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[40\].u.buff
timestamp 1676381911
transform 1 0 88512 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[40\].u.inv
timestamp 1676382929
transform -1 0 88992 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[41\].u.buff
timestamp 1676381911
transform 1 0 88800 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[41\].u.inv
timestamp 1676382929
transform 1 0 89088 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[42\].u.buff
timestamp 1676381911
transform -1 0 89760 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[42\].u.inv
timestamp 1676382929
transform 1 0 89472 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[43\].u.buff
timestamp 1676381911
transform 1 0 89376 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[43\].u.inv
timestamp 1676382929
transform -1 0 90816 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[44\].u.buff
timestamp 1676381911
transform -1 0 90528 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[44\].u.inv
timestamp 1676382929
transform 1 0 90240 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[45\].u.buff
timestamp 1676381911
transform 1 0 90336 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[45\].u.inv
timestamp 1676382929
transform 1 0 91680 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[46\].u.buff
timestamp 1676381911
transform 1 0 90816 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[46\].u.inv
timestamp 1676382929
transform -1 0 91488 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[47\].u.buff
timestamp 1676381911
transform 1 0 90912 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[47\].u.inv
timestamp 1676382929
transform 1 0 91488 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[48\].u.buff
timestamp 1676381911
transform 1 0 91584 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[48\].u.inv
timestamp 1676382929
transform 1 0 92448 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[49\].u.buff
timestamp 1676381911
transform 1 0 92064 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[49\].u.inv
timestamp 1676382929
transform -1 0 93504 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[50\].u.buff
timestamp 1676381911
transform -1 0 93216 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[50\].u.inv
timestamp 1676382929
transform -1 0 93024 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[51\].u.buff
timestamp 1676381911
transform 1 0 92928 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[51\].u.inv
timestamp 1676382929
transform -1 0 93408 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[52\].u.buff
timestamp 1676381911
transform 1 0 93312 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[52\].u.inv
timestamp 1676382929
transform -1 0 93792 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[53\].u.buff
timestamp 1676381911
transform 1 0 93792 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[53\].u.inv
timestamp 1676382929
transform 1 0 93792 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[54\].u.buff
timestamp 1676381911
transform -1 0 94560 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[54\].u.inv
timestamp 1676382929
transform 1 0 93600 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[55\].u.buff
timestamp 1676381911
transform -1 0 95040 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[55\].u.inv
timestamp 1676382929
transform 1 0 94656 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[56\].u.buff
timestamp 1676381911
transform -1 0 95424 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[56\].u.inv
timestamp 1676382929
transform 1 0 95808 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[57\].u.buff
timestamp 1676381911
transform 1 0 95040 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[57\].u.inv
timestamp 1676382929
transform -1 0 95808 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[58\].u.buff
timestamp 1676381911
transform 1 0 95424 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[58\].u.inv
timestamp 1676382929
transform 1 0 95808 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[59\].u.buff
timestamp 1676381911
transform 1 0 95616 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[59\].u.inv
timestamp 1676382929
transform -1 0 97056 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[60\].u.buff
timestamp 1676381911
transform 1 0 96288 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[60\].u.inv
timestamp 1676382929
transform -1 0 97344 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[61\].u.buff
timestamp 1676381911
transform 1 0 96864 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[61\].u.inv
timestamp 1676382929
transform 1 0 97248 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[62\].u.buff
timestamp 1676381911
transform -1 0 97728 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[62\].u.inv
timestamp 1676382929
transform -1 0 97920 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[63\].u.buff
timestamp 1676381911
transform -1 0 98304 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[63\].u.inv
timestamp 1676382929
transform 1 0 97920 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[64\].u.buff
timestamp 1676381911
transform -1 0 98592 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[64\].u.inv
timestamp 1676382929
transform 1 0 98592 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[65\].u.buff
timestamp 1676381911
transform -1 0 98016 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[65\].u.inv
timestamp 1676382929
transform -1 0 97728 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[66\].u.buff
timestamp 1676381911
transform 1 0 96960 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[66\].u.inv
timestamp 1676382929
transform -1 0 97056 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[67\].u.buff
timestamp 1676381911
transform 1 0 96576 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[67\].u.inv
timestamp 1676382929
transform 1 0 97344 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[68\].u.buff
timestamp 1676381911
transform 1 0 96192 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[68\].u.inv
timestamp 1676382929
transform -1 0 96480 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[69\].u.buff
timestamp 1676381911
transform 1 0 95808 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[69\].u.inv
timestamp 1676382929
transform -1 0 96096 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[70\].u.buff
timestamp 1676381911
transform 1 0 95424 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[70\].u.inv
timestamp 1676382929
transform 1 0 95328 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[71\].u.buff
timestamp 1676381911
transform 1 0 94944 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[71\].u.inv
timestamp 1676382929
transform 1 0 94656 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[72\].u.buff
timestamp 1676381911
transform -1 0 95040 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[72\].u.inv
timestamp 1676382929
transform 1 0 95040 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[73\].u.buff
timestamp 1676381911
transform 1 0 94176 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[73\].u.inv
timestamp 1676382929
transform 1 0 94176 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[74\].u.buff
timestamp 1676381911
transform 1 0 93792 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[74\].u.inv
timestamp 1676382929
transform -1 0 94176 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[75\].u.buff
timestamp 1676381911
transform -1 0 93888 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[75\].u.inv
timestamp 1676382929
transform 1 0 92736 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[76\].u.buff
timestamp 1676381911
transform 1 0 93024 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[76\].u.inv
timestamp 1676382929
transform -1 0 93312 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[77\].u.buff
timestamp 1676381911
transform 1 0 92448 0 1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[77\].u.inv
timestamp 1676382929
transform -1 0 93024 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[78\].u.buff
timestamp 1676381911
transform -1 0 92736 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[78\].u.inv
timestamp 1676382929
transform 1 0 92160 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[79\].u.buff
timestamp 1676381911
transform -1 0 92352 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[79\].u.inv
timestamp 1676382929
transform 1 0 91776 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[80\].u.buff
timestamp 1676381911
transform 1 0 91200 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[80\].u.inv
timestamp 1676382929
transform 1 0 91296 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[81\].u.buff
timestamp 1676381911
transform -1 0 91968 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[81\].u.inv
timestamp 1676382929
transform 1 0 90912 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[82\].u.buff
timestamp 1676381911
transform 1 0 90528 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[82\].u.inv
timestamp 1676382929
transform 1 0 90528 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[83\].u.buff
timestamp 1676381911
transform 1 0 90048 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[83\].u.inv
timestamp 1676382929
transform 1 0 90144 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[84\].u.buff
timestamp 1676381911
transform 1 0 89664 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[84\].u.inv
timestamp 1676382929
transform 1 0 89376 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[85\].u.buff
timestamp 1676381911
transform 1 0 89376 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[85\].u.inv
timestamp 1676382929
transform -1 0 90048 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[86\].u.buff
timestamp 1676381911
transform 1 0 88896 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[86\].u.inv
timestamp 1676382929
transform 1 0 88992 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[87\].u.buff
timestamp 1676381911
transform 1 0 88512 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[87\].u.inv
timestamp 1676382929
transform 1 0 88512 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[88\].u.buff
timestamp 1676381911
transform 1 0 88128 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[88\].u.inv
timestamp 1676382929
transform 1 0 88128 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[89\].u.buff
timestamp 1676381911
transform 1 0 87648 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[89\].u.inv
timestamp 1676382929
transform -1 0 88608 0 1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[90\].u.buff
timestamp 1676381911
transform 1 0 87360 0 1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[90\].u.inv
timestamp 1676382929
transform 1 0 87360 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[91\].u.buff
timestamp 1676381911
transform 1 0 86976 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[91\].u.inv
timestamp 1676382929
transform 1 0 86976 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[92\].u.buff
timestamp 1676381911
transform 1 0 86496 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[92\].u.inv
timestamp 1676382929
transform 1 0 86496 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[93\].u.buff
timestamp 1676381911
transform 1 0 86112 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[93\].u.inv
timestamp 1676382929
transform 1 0 86208 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[94\].u.buff
timestamp 1676381911
transform 1 0 85824 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[94\].u.inv
timestamp 1676382929
transform 1 0 85728 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[95\].u.buff
timestamp 1676381911
transform 1 0 85440 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[95\].u.inv
timestamp 1676382929
transform 1 0 85344 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[96\].u.buff
timestamp 1676381911
transform 1 0 84864 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[96\].u.inv
timestamp 1676382929
transform -1 0 84864 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[97\].u.buff
timestamp 1676381911
transform 1 0 84576 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[97\].u.inv
timestamp 1676382929
transform 1 0 84960 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[98\].u.buff
timestamp 1676381911
transform 1 0 84192 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[98\].u.inv
timestamp 1676382929
transform 1 0 84096 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[99\].u.buff
timestamp 1676381911
transform 1 0 83712 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[99\].u.inv
timestamp 1676382929
transform 1 0 83712 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[100\].u.buff
timestamp 1676381911
transform 1 0 83328 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[100\].u.inv
timestamp 1676382929
transform 1 0 83328 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[101\].u.buff
timestamp 1676381911
transform 1 0 82944 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[101\].u.inv
timestamp 1676382929
transform 1 0 82944 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[102\].u.buff
timestamp 1676381911
transform 1 0 82560 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[102\].u.inv
timestamp 1676382929
transform 1 0 82560 0 1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[103\].u.buff
timestamp 1676381911
transform 1 0 82176 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[103\].u.inv
timestamp 1676382929
transform 1 0 82176 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[104\].u.buff
timestamp 1676381911
transform 1 0 81696 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[104\].u.inv
timestamp 1676382929
transform -1 0 82080 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[105\].u.buff
timestamp 1676381911
transform 1 0 81312 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[105\].u.inv
timestamp 1676382929
transform 1 0 81408 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[106\].u.buff
timestamp 1676381911
transform 1 0 80928 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[106\].u.inv
timestamp 1676382929
transform -1 0 81408 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[107\].u.buff
timestamp 1676381911
transform 1 0 80448 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[107\].u.inv
timestamp 1676382929
transform -1 0 81120 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[108\].u.buff
timestamp 1676381911
transform 1 0 80064 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[108\].u.inv
timestamp 1676382929
transform 1 0 79968 0 1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[109\].u.buff
timestamp 1676381911
transform 1 0 79776 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[109\].u.inv
timestamp 1676382929
transform 1 0 79776 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[110\].u.buff
timestamp 1676381911
transform 1 0 79296 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[110\].u.inv
timestamp 1676382929
transform 1 0 79392 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[111\].u.buff
timestamp 1676381911
transform 1 0 78336 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[111\].u.inv
timestamp 1676382929
transform -1 0 79296 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[112\].u.buff
timestamp 1676381911
transform 1 0 78624 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[112\].u.inv
timestamp 1676382929
transform 1 0 78528 0 1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[113\].u.buff
timestamp 1676381911
transform 1 0 78144 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[113\].u.inv
timestamp 1676382929
transform 1 0 78048 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[114\].u.buff
timestamp 1676381911
transform 1 0 77568 0 1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[114\].u.inv
timestamp 1676382929
transform 1 0 77664 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[115\].u.buff
timestamp 1676381911
transform 1 0 77280 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[115\].u.inv
timestamp 1676382929
transform 1 0 77376 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[116\].u.buff
timestamp 1676381911
transform 1 0 76896 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[116\].u.inv
timestamp 1676382929
transform 1 0 76992 0 1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[117\].u.buff
timestamp 1676381911
transform 1 0 76512 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[117\].u.inv
timestamp 1676382929
transform 1 0 76416 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[118\].u.buff
timestamp 1676381911
transform 1 0 76128 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[118\].u.inv
timestamp 1676382929
transform 1 0 76512 0 1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[119\].u.buff
timestamp 1676381911
transform 1 0 75744 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[119\].u.inv
timestamp 1676382929
transform 1 0 75552 0 1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[120\].u.buff
timestamp 1676381911
transform 1 0 75264 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[120\].u.inv
timestamp 1676382929
transform 1 0 74976 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[121\].u.buff
timestamp 1676381911
transform 1 0 74496 0 -1 18900
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[121\].u.inv
timestamp 1676382929
transform -1 0 75936 0 1 17388
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[122\].u.buff
timestamp 1676381911
transform 1 0 74400 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[122\].u.inv
timestamp 1676382929
transform -1 0 74400 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[123\].u.buff
timestamp 1676381911
transform 1 0 74016 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[123\].u.inv
timestamp 1676382929
transform 1 0 69696 0 -1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[124\].u.buff
timestamp 1676381911
transform 1 0 73632 0 1 17388
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[124\].u.inv
timestamp 1676382929
transform 1 0 68544 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[125\].u.buff
timestamp 1676381911
transform 1 0 69600 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[125\].u.inv
timestamp 1676382929
transform 1 0 72864 0 -1 18900
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[126\].u.buff
timestamp 1676381911
transform 1 0 67104 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[126\].u.inv
timestamp 1676382929
transform 1 0 69312 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[127\].u.buff
timestamp 1676381911
transform 1 0 69024 0 1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[127\].u.inv
timestamp 1676382929
transform -1 0 68256 0 1 14364
box -48 -56 336 834
use sg13g2_buf_2  fanout21
timestamp 1676381867
transform 1 0 69120 0 1 24948
box -48 -56 528 834
use sg13g2_buf_1  fanout22
timestamp 1676381911
transform -1 0 68064 0 1 26460
box -48 -56 432 834
use sg13g2_buf_2  fanout23
timestamp 1676381867
transform 1 0 67392 0 1 30996
box -48 -56 528 834
use sg13g2_buf_1  fanout24
timestamp 1676381911
transform -1 0 68448 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  fanout25
timestamp 1676381911
transform -1 0 75456 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout26
timestamp 1676381911
transform -1 0 77952 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout27
timestamp 1676381911
transform 1 0 78720 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout28
timestamp 1676381911
transform 1 0 74304 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout29
timestamp 1676381911
transform -1 0 75360 0 1 21924
box -48 -56 432 834
use sg13g2_buf_2  fanout30
timestamp 1676381867
transform -1 0 80448 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_1  fanout31
timestamp 1676381911
transform -1 0 80832 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_2  fanout32
timestamp 1676381867
transform 1 0 83040 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_1  fanout33
timestamp 1676381911
transform -1 0 83904 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout34
timestamp 1676381911
transform -1 0 75744 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout35
timestamp 1676381911
transform 1 0 73632 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout36
timestamp 1676381911
transform 1 0 76992 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout37
timestamp 1676381911
transform 1 0 78912 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout38
timestamp 1676381911
transform -1 0 74784 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout39
timestamp 1676381911
transform -1 0 74784 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout40
timestamp 1676381911
transform -1 0 81120 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout41
timestamp 1676381911
transform 1 0 81408 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout42
timestamp 1676381911
transform 1 0 83040 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout43
timestamp 1676381911
transform 1 0 84960 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout44
timestamp 1676381911
transform -1 0 82176 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout45
timestamp 1676381911
transform 1 0 85632 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout46
timestamp 1676381911
transform -1 0 87648 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_2  fanout47
timestamp 1676381867
transform -1 0 90048 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_1  fanout48
timestamp 1676381911
transform -1 0 90432 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout49
timestamp 1676381911
transform -1 0 86496 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  fanout50
timestamp 1676381911
transform 1 0 92352 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout51
timestamp 1676381911
transform 1 0 91968 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_2  fanout52
timestamp 1676381867
transform 1 0 95520 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_1  fanout53
timestamp 1676381911
transform 1 0 96000 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout54
timestamp 1676381911
transform 1 0 91584 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout55
timestamp 1676381911
transform -1 0 86688 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout56
timestamp 1676381911
transform 1 0 87840 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout57
timestamp 1676381911
transform -1 0 89472 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout58
timestamp 1676381911
transform 1 0 90912 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout59
timestamp 1676381911
transform -1 0 86784 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout60
timestamp 1676381911
transform 1 0 92160 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout61
timestamp 1676381911
transform -1 0 94272 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  fanout62
timestamp 1676381911
transform -1 0 96192 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout63
timestamp 1676381911
transform 1 0 96192 0 1 34020
box -48 -56 432 834
use sg13g2_buf_2  fanout64
timestamp 1676381867
transform -1 0 93024 0 1 34020
box -48 -56 528 834
use sg13g2_buf_2  fanout65
timestamp 1676381867
transform -1 0 86880 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_1  fanout66
timestamp 1676381911
transform 1 0 76224 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  fanout67
timestamp 1676381911
transform -1 0 2112 0 1 8316
box -48 -56 432 834
use sg13g2_buf_2  fanout68
timestamp 1676381867
transform -1 0 68928 0 1 9828
box -48 -56 528 834
use sg13g2_buf_2  fanout69
timestamp 1676381867
transform 1 0 68064 0 -1 15876
box -48 -56 528 834
use sg13g2_buf_1  fanout70
timestamp 1676381911
transform -1 0 67872 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout71
timestamp 1676381911
transform 1 0 74304 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout72
timestamp 1676381911
transform -1 0 75168 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout73
timestamp 1676381911
transform -1 0 77952 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout74
timestamp 1676381911
transform -1 0 80352 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout75
timestamp 1676381911
transform -1 0 77568 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout76
timestamp 1676381911
transform -1 0 74400 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout77
timestamp 1676381911
transform -1 0 81216 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout78
timestamp 1676381911
transform -1 0 82944 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout79
timestamp 1676381911
transform -1 0 84384 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout80
timestamp 1676381911
transform 1 0 85152 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout81
timestamp 1676381911
transform 1 0 80448 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout82
timestamp 1676381911
transform -1 0 74784 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout83
timestamp 1676381911
transform -1 0 75264 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout84
timestamp 1676381911
transform 1 0 74688 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout85
timestamp 1676381911
transform -1 0 78336 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout86
timestamp 1676381911
transform -1 0 79104 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_2  fanout87
timestamp 1676381867
transform 1 0 75072 0 1 18900
box -48 -56 528 834
use sg13g2_buf_1  fanout88
timestamp 1676381911
transform -1 0 80640 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout89
timestamp 1676381911
transform -1 0 82176 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout90
timestamp 1676381911
transform -1 0 84192 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout91
timestamp 1676381911
transform 1 0 85536 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout92
timestamp 1676381911
transform -1 0 80736 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout93
timestamp 1676381911
transform 1 0 86016 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout94
timestamp 1676381911
transform 1 0 87936 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout95
timestamp 1676381911
transform -1 0 90144 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout96
timestamp 1676381911
transform 1 0 91296 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout97
timestamp 1676381911
transform -1 0 86784 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout98
timestamp 1676381911
transform 1 0 92064 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout99
timestamp 1676381911
transform -1 0 94272 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout100
timestamp 1676381911
transform -1 0 96384 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout101
timestamp 1676381911
transform 1 0 96384 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout102
timestamp 1676381911
transform -1 0 92832 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout103
timestamp 1676381911
transform 1 0 94272 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout104
timestamp 1676381911
transform -1 0 86688 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout105
timestamp 1676381911
transform -1 0 88320 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout106
timestamp 1676381911
transform -1 0 89856 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout107
timestamp 1676381911
transform 1 0 91296 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout108
timestamp 1676381911
transform 1 0 89856 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout109
timestamp 1676381911
transform -1 0 93216 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout110
timestamp 1676381911
transform -1 0 94272 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout111
timestamp 1676381911
transform -1 0 95904 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout112
timestamp 1676381911
transform 1 0 97056 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout113
timestamp 1676381911
transform -1 0 93312 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout114
timestamp 1676381911
transform 1 0 86688 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  fanout115
timestamp 1676381911
transform 1 0 86784 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout116
timestamp 1676381911
transform 1 0 75456 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  fanout117
timestamp 1676381911
transform -1 0 2112 0 -1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679581782
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679581782
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679581782
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679581782
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679581782
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679581782
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679581782
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679581782
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679581782
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679581782
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679581782
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679581782
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679581782
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679581782
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679581782
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679581782
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679581782
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679581782
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679581782
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679581782
transform 1 0 55008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679581782
transform 1 0 55680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679581782
transform 1 0 56352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679581782
transform 1 0 57024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679581782
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679581782
transform 1 0 58368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679581782
transform 1 0 59040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679581782
transform 1 0 59712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679581782
transform 1 0 60384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679581782
transform 1 0 61056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679581782
transform 1 0 61728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679581782
transform 1 0 62400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679581782
transform 1 0 63072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679581782
transform 1 0 63744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679581782
transform 1 0 64416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679581782
transform 1 0 65088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679581782
transform 1 0 65760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679581782
transform 1 0 66432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679581782
transform 1 0 67104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679581782
transform 1 0 67776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679581782
transform 1 0 68448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679581782
transform 1 0 69120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679581782
transform 1 0 69792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679581782
transform 1 0 70464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679581782
transform 1 0 71136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679581782
transform 1 0 71808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_749
timestamp 1679581782
transform 1 0 72480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_756
timestamp 1679581782
transform 1 0 73152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_763
timestamp 1679581782
transform 1 0 73824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_770
timestamp 1679581782
transform 1 0 74496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_777
timestamp 1679581782
transform 1 0 75168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_784
timestamp 1679581782
transform 1 0 75840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_791
timestamp 1679581782
transform 1 0 76512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_798
timestamp 1679581782
transform 1 0 77184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_805
timestamp 1679581782
transform 1 0 77856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_812
timestamp 1679581782
transform 1 0 78528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_819
timestamp 1679581782
transform 1 0 79200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_826
timestamp 1679581782
transform 1 0 79872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_833
timestamp 1679581782
transform 1 0 80544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_840
timestamp 1679581782
transform 1 0 81216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_847
timestamp 1679581782
transform 1 0 81888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_854
timestamp 1679581782
transform 1 0 82560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_861
timestamp 1679581782
transform 1 0 83232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_868
timestamp 1679581782
transform 1 0 83904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_875
timestamp 1679581782
transform 1 0 84576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_882
timestamp 1679581782
transform 1 0 85248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_889
timestamp 1679581782
transform 1 0 85920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_896
timestamp 1679581782
transform 1 0 86592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_903
timestamp 1679581782
transform 1 0 87264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_910
timestamp 1679581782
transform 1 0 87936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_917
timestamp 1679581782
transform 1 0 88608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_924
timestamp 1679581782
transform 1 0 89280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_931
timestamp 1679581782
transform 1 0 89952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_938
timestamp 1679581782
transform 1 0 90624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_945
timestamp 1679581782
transform 1 0 91296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_952
timestamp 1679581782
transform 1 0 91968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_959
timestamp 1679581782
transform 1 0 92640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_966
timestamp 1679581782
transform 1 0 93312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_973
timestamp 1679581782
transform 1 0 93984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_980
timestamp 1679581782
transform 1 0 94656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_987
timestamp 1679581782
transform 1 0 95328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_994
timestamp 1679581782
transform 1 0 96000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1001
timestamp 1679581782
transform 1 0 96672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1008
timestamp 1679581782
transform 1 0 97344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1015
timestamp 1679581782
transform 1 0 98016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1022
timestamp 1679581782
transform 1 0 98688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679581782
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679581782
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679581782
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679581782
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679581782
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679581782
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679581782
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679581782
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679581782
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679581782
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679581782
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679581782
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679581782
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679581782
transform 1 0 30816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679581782
transform 1 0 31488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679581782
transform 1 0 32160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679581782
transform 1 0 32832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679581782
transform 1 0 33504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679581782
transform 1 0 34176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679581782
transform 1 0 34848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679581782
transform 1 0 35520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679581782
transform 1 0 36192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679581782
transform 1 0 36864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679581782
transform 1 0 37536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679581782
transform 1 0 38208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679581782
transform 1 0 38880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 39552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 40896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 41568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 42912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 43584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 44256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 44928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 45600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 46272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 46944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679581782
transform 1 0 48288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679581782
transform 1 0 48960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679581782
transform 1 0 49632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679581782
transform 1 0 50304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679581782
transform 1 0 52992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679581782
transform 1 0 53664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679581782
transform 1 0 54336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679581782
transform 1 0 55008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679581782
transform 1 0 55680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679581782
transform 1 0 56352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679581782
transform 1 0 57024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_595
timestamp 1679581782
transform 1 0 57696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_602
timestamp 1679581782
transform 1 0 58368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679581782
transform 1 0 59040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_616
timestamp 1679581782
transform 1 0 59712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_623
timestamp 1679581782
transform 1 0 60384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_630
timestamp 1679581782
transform 1 0 61056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_637
timestamp 1679581782
transform 1 0 61728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_644
timestamp 1679581782
transform 1 0 62400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_651
timestamp 1679581782
transform 1 0 63072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_658
timestamp 1679581782
transform 1 0 63744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_665
timestamp 1679581782
transform 1 0 64416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_672
timestamp 1679581782
transform 1 0 65088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_679
timestamp 1679581782
transform 1 0 65760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_686
timestamp 1679581782
transform 1 0 66432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_693
timestamp 1679581782
transform 1 0 67104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_700
timestamp 1679581782
transform 1 0 67776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_707
timestamp 1679581782
transform 1 0 68448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_714
timestamp 1679581782
transform 1 0 69120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_721
timestamp 1679581782
transform 1 0 69792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_728
timestamp 1679581782
transform 1 0 70464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_735
timestamp 1679581782
transform 1 0 71136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_742
timestamp 1679581782
transform 1 0 71808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_749
timestamp 1679581782
transform 1 0 72480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_756
timestamp 1679581782
transform 1 0 73152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_763
timestamp 1679581782
transform 1 0 73824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_770
timestamp 1679581782
transform 1 0 74496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_777
timestamp 1679581782
transform 1 0 75168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_784
timestamp 1679581782
transform 1 0 75840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_791
timestamp 1679581782
transform 1 0 76512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_798
timestamp 1679581782
transform 1 0 77184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_805
timestamp 1679581782
transform 1 0 77856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_812
timestamp 1679581782
transform 1 0 78528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_819
timestamp 1679581782
transform 1 0 79200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_826
timestamp 1679581782
transform 1 0 79872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_833
timestamp 1679581782
transform 1 0 80544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_840
timestamp 1679581782
transform 1 0 81216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_847
timestamp 1679581782
transform 1 0 81888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_854
timestamp 1679581782
transform 1 0 82560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_861
timestamp 1679581782
transform 1 0 83232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_868
timestamp 1679581782
transform 1 0 83904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_875
timestamp 1679581782
transform 1 0 84576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_882
timestamp 1679581782
transform 1 0 85248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_889
timestamp 1679581782
transform 1 0 85920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_896
timestamp 1679581782
transform 1 0 86592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_903
timestamp 1679581782
transform 1 0 87264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_910
timestamp 1679581782
transform 1 0 87936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_917
timestamp 1679581782
transform 1 0 88608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_924
timestamp 1679581782
transform 1 0 89280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_931
timestamp 1679581782
transform 1 0 89952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_938
timestamp 1679581782
transform 1 0 90624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_945
timestamp 1679581782
transform 1 0 91296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_952
timestamp 1679581782
transform 1 0 91968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_959
timestamp 1679581782
transform 1 0 92640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_966
timestamp 1679581782
transform 1 0 93312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_973
timestamp 1679581782
transform 1 0 93984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_980
timestamp 1679581782
transform 1 0 94656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_987
timestamp 1679581782
transform 1 0 95328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_994
timestamp 1679581782
transform 1 0 96000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1001
timestamp 1679581782
transform 1 0 96672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1008
timestamp 1679581782
transform 1 0 97344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1015
timestamp 1679581782
transform 1 0 98016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1022
timestamp 1679581782
transform 1 0 98688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679581782
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679581782
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_67
timestamp 1679581782
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_74
timestamp 1679581782
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679581782
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679581782
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679581782
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679581782
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679581782
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_116
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_123
timestamp 1679581782
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_130
timestamp 1679581782
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_137
timestamp 1679581782
transform 1 0 13728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 15744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_165
timestamp 1679581782
transform 1 0 16416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_172
timestamp 1679581782
transform 1 0 17088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1679581782
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_200
timestamp 1679581782
transform 1 0 19776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_207
timestamp 1679581782
transform 1 0 20448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_214
timestamp 1679581782
transform 1 0 21120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_221
timestamp 1679581782
transform 1 0 21792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_228
timestamp 1679581782
transform 1 0 22464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_235
timestamp 1679581782
transform 1 0 23136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_242
timestamp 1679581782
transform 1 0 23808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_249
timestamp 1679581782
transform 1 0 24480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_256
timestamp 1679581782
transform 1 0 25152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_263
timestamp 1679581782
transform 1 0 25824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_270
timestamp 1679581782
transform 1 0 26496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_277
timestamp 1679581782
transform 1 0 27168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_284
timestamp 1679581782
transform 1 0 27840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_291
timestamp 1679581782
transform 1 0 28512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_298
timestamp 1679581782
transform 1 0 29184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_305
timestamp 1679581782
transform 1 0 29856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_312
timestamp 1679581782
transform 1 0 30528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_319
timestamp 1679581782
transform 1 0 31200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_326
timestamp 1679581782
transform 1 0 31872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_333
timestamp 1679581782
transform 1 0 32544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_340
timestamp 1679581782
transform 1 0 33216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_347
timestamp 1679581782
transform 1 0 33888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_354
timestamp 1679581782
transform 1 0 34560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_361
timestamp 1679581782
transform 1 0 35232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_368
timestamp 1679581782
transform 1 0 35904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_375
timestamp 1679581782
transform 1 0 36576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_382
timestamp 1679581782
transform 1 0 37248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_389
timestamp 1679581782
transform 1 0 37920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_396
timestamp 1679581782
transform 1 0 38592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_403
timestamp 1679581782
transform 1 0 39264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_410
timestamp 1679581782
transform 1 0 39936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_417
timestamp 1679581782
transform 1 0 40608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_424
timestamp 1679581782
transform 1 0 41280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_431
timestamp 1679581782
transform 1 0 41952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_438
timestamp 1679581782
transform 1 0 42624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_445
timestamp 1679581782
transform 1 0 43296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_452
timestamp 1679581782
transform 1 0 43968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_459
timestamp 1679581782
transform 1 0 44640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_466
timestamp 1679581782
transform 1 0 45312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_473
timestamp 1679581782
transform 1 0 45984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_480
timestamp 1679581782
transform 1 0 46656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_487
timestamp 1679581782
transform 1 0 47328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_494
timestamp 1679581782
transform 1 0 48000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_501
timestamp 1679581782
transform 1 0 48672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_508
timestamp 1679581782
transform 1 0 49344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_515
timestamp 1679581782
transform 1 0 50016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_522
timestamp 1679581782
transform 1 0 50688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_529
timestamp 1679581782
transform 1 0 51360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_536
timestamp 1679581782
transform 1 0 52032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_543
timestamp 1679581782
transform 1 0 52704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_550
timestamp 1679581782
transform 1 0 53376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_557
timestamp 1679581782
transform 1 0 54048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_564
timestamp 1679581782
transform 1 0 54720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_571
timestamp 1679581782
transform 1 0 55392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_578
timestamp 1679581782
transform 1 0 56064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_585
timestamp 1679581782
transform 1 0 56736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_592
timestamp 1679581782
transform 1 0 57408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_599
timestamp 1679581782
transform 1 0 58080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_606
timestamp 1679581782
transform 1 0 58752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_613
timestamp 1679581782
transform 1 0 59424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_620
timestamp 1679581782
transform 1 0 60096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_627
timestamp 1679581782
transform 1 0 60768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_634
timestamp 1679581782
transform 1 0 61440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_641
timestamp 1679581782
transform 1 0 62112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_648
timestamp 1679581782
transform 1 0 62784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_655
timestamp 1679581782
transform 1 0 63456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_662
timestamp 1679581782
transform 1 0 64128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_669
timestamp 1679581782
transform 1 0 64800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_676
timestamp 1679581782
transform 1 0 65472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_683
timestamp 1679581782
transform 1 0 66144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_690
timestamp 1679581782
transform 1 0 66816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_697
timestamp 1679581782
transform 1 0 67488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_704
timestamp 1679581782
transform 1 0 68160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_711
timestamp 1679581782
transform 1 0 68832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_718
timestamp 1679581782
transform 1 0 69504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_725
timestamp 1679581782
transform 1 0 70176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_732
timestamp 1679581782
transform 1 0 70848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_739
timestamp 1679581782
transform 1 0 71520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_746
timestamp 1679581782
transform 1 0 72192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_753
timestamp 1679581782
transform 1 0 72864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_760
timestamp 1679581782
transform 1 0 73536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_767
timestamp 1679581782
transform 1 0 74208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_774
timestamp 1679581782
transform 1 0 74880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_781
timestamp 1679581782
transform 1 0 75552 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_788
timestamp 1679581782
transform 1 0 76224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_795
timestamp 1679581782
transform 1 0 76896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_802
timestamp 1679581782
transform 1 0 77568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_809
timestamp 1679581782
transform 1 0 78240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_816
timestamp 1679581782
transform 1 0 78912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_823
timestamp 1679581782
transform 1 0 79584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_830
timestamp 1679581782
transform 1 0 80256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_837
timestamp 1679581782
transform 1 0 80928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_844
timestamp 1679581782
transform 1 0 81600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_851
timestamp 1679581782
transform 1 0 82272 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_858
timestamp 1679581782
transform 1 0 82944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_865
timestamp 1679581782
transform 1 0 83616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_872
timestamp 1679581782
transform 1 0 84288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_879
timestamp 1679581782
transform 1 0 84960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_886
timestamp 1679581782
transform 1 0 85632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_893
timestamp 1679581782
transform 1 0 86304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_900
timestamp 1679581782
transform 1 0 86976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_907
timestamp 1679581782
transform 1 0 87648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_914
timestamp 1679581782
transform 1 0 88320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_921
timestamp 1679581782
transform 1 0 88992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_928
timestamp 1679581782
transform 1 0 89664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_935
timestamp 1679581782
transform 1 0 90336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_942
timestamp 1679581782
transform 1 0 91008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_949
timestamp 1679581782
transform 1 0 91680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_956
timestamp 1679581782
transform 1 0 92352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_963
timestamp 1679581782
transform 1 0 93024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_970
timestamp 1679581782
transform 1 0 93696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_977
timestamp 1679581782
transform 1 0 94368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_984
timestamp 1679581782
transform 1 0 95040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_991
timestamp 1679581782
transform 1 0 95712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_998
timestamp 1679581782
transform 1 0 96384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1005
timestamp 1679581782
transform 1 0 97056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1012
timestamp 1679581782
transform 1 0 97728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1019
timestamp 1679581782
transform 1 0 98400 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_1026
timestamp 1677580104
transform 1 0 99072 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_1028
timestamp 1677579658
transform 1 0 99264 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 4992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 5664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 7680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679581782
transform 1 0 9024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 9696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679581782
transform 1 0 11040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 11712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679581782
transform 1 0 12384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_130
timestamp 1679581782
transform 1 0 13056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_137
timestamp 1679581782
transform 1 0 13728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_144
timestamp 1679581782
transform 1 0 14400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_151
timestamp 1679581782
transform 1 0 15072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_158
timestamp 1679581782
transform 1 0 15744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_165
timestamp 1679581782
transform 1 0 16416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_172
timestamp 1679581782
transform 1 0 17088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_179
timestamp 1679581782
transform 1 0 17760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_186
timestamp 1679581782
transform 1 0 18432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_193
timestamp 1679581782
transform 1 0 19104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_200
timestamp 1679581782
transform 1 0 19776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_207
timestamp 1679581782
transform 1 0 20448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_214
timestamp 1679581782
transform 1 0 21120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_221
timestamp 1679581782
transform 1 0 21792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_228
timestamp 1679581782
transform 1 0 22464 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_235
timestamp 1679581782
transform 1 0 23136 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_242
timestamp 1679581782
transform 1 0 23808 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_249
timestamp 1679581782
transform 1 0 24480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_256
timestamp 1679581782
transform 1 0 25152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_263
timestamp 1679581782
transform 1 0 25824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_270
timestamp 1679581782
transform 1 0 26496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_277
timestamp 1679581782
transform 1 0 27168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_284
timestamp 1679581782
transform 1 0 27840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_291
timestamp 1679581782
transform 1 0 28512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_298
timestamp 1679581782
transform 1 0 29184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_305
timestamp 1679581782
transform 1 0 29856 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_312
timestamp 1679581782
transform 1 0 30528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_319
timestamp 1679581782
transform 1 0 31200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_326
timestamp 1679581782
transform 1 0 31872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_333
timestamp 1679581782
transform 1 0 32544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_340
timestamp 1679581782
transform 1 0 33216 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_347
timestamp 1679581782
transform 1 0 33888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_354
timestamp 1679581782
transform 1 0 34560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_361
timestamp 1679581782
transform 1 0 35232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_368
timestamp 1679581782
transform 1 0 35904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_375
timestamp 1679581782
transform 1 0 36576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_382
timestamp 1679581782
transform 1 0 37248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_389
timestamp 1679581782
transform 1 0 37920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_396
timestamp 1679581782
transform 1 0 38592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_403
timestamp 1679581782
transform 1 0 39264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_410
timestamp 1679581782
transform 1 0 39936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_417
timestamp 1679581782
transform 1 0 40608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_424
timestamp 1679581782
transform 1 0 41280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_431
timestamp 1679581782
transform 1 0 41952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_438
timestamp 1679581782
transform 1 0 42624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_445
timestamp 1679581782
transform 1 0 43296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_452
timestamp 1679581782
transform 1 0 43968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_459
timestamp 1679581782
transform 1 0 44640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_466
timestamp 1679581782
transform 1 0 45312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_473
timestamp 1679581782
transform 1 0 45984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_480
timestamp 1679581782
transform 1 0 46656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_487
timestamp 1679581782
transform 1 0 47328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_494
timestamp 1679581782
transform 1 0 48000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_501
timestamp 1679581782
transform 1 0 48672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_508
timestamp 1679581782
transform 1 0 49344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_515
timestamp 1679581782
transform 1 0 50016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_522
timestamp 1679581782
transform 1 0 50688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_529
timestamp 1679581782
transform 1 0 51360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_536
timestamp 1679581782
transform 1 0 52032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_543
timestamp 1679581782
transform 1 0 52704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_550
timestamp 1679581782
transform 1 0 53376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_557
timestamp 1679581782
transform 1 0 54048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_564
timestamp 1679581782
transform 1 0 54720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_571
timestamp 1679581782
transform 1 0 55392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_578
timestamp 1679581782
transform 1 0 56064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_585
timestamp 1679581782
transform 1 0 56736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_592
timestamp 1679581782
transform 1 0 57408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_599
timestamp 1679581782
transform 1 0 58080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_606
timestamp 1679581782
transform 1 0 58752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_613
timestamp 1679581782
transform 1 0 59424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_620
timestamp 1679581782
transform 1 0 60096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_627
timestamp 1679581782
transform 1 0 60768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_634
timestamp 1679581782
transform 1 0 61440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_641
timestamp 1679581782
transform 1 0 62112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_648
timestamp 1679581782
transform 1 0 62784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_655
timestamp 1679581782
transform 1 0 63456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_662
timestamp 1679581782
transform 1 0 64128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_669
timestamp 1679581782
transform 1 0 64800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_676
timestamp 1679581782
transform 1 0 65472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_683
timestamp 1679581782
transform 1 0 66144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_690
timestamp 1679581782
transform 1 0 66816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_697
timestamp 1679581782
transform 1 0 67488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_704
timestamp 1679581782
transform 1 0 68160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_711
timestamp 1679581782
transform 1 0 68832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_718
timestamp 1679581782
transform 1 0 69504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_725
timestamp 1679581782
transform 1 0 70176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_732
timestamp 1679581782
transform 1 0 70848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_739
timestamp 1679581782
transform 1 0 71520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_746
timestamp 1679581782
transform 1 0 72192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_753
timestamp 1679581782
transform 1 0 72864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_760
timestamp 1679581782
transform 1 0 73536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_767
timestamp 1679581782
transform 1 0 74208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_774
timestamp 1679581782
transform 1 0 74880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_781
timestamp 1679581782
transform 1 0 75552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_788
timestamp 1679581782
transform 1 0 76224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_795
timestamp 1679581782
transform 1 0 76896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_802
timestamp 1679581782
transform 1 0 77568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_809
timestamp 1679581782
transform 1 0 78240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_816
timestamp 1679581782
transform 1 0 78912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_823
timestamp 1679581782
transform 1 0 79584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_830
timestamp 1679581782
transform 1 0 80256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_837
timestamp 1679581782
transform 1 0 80928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_844
timestamp 1679581782
transform 1 0 81600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_851
timestamp 1679581782
transform 1 0 82272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_858
timestamp 1679581782
transform 1 0 82944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_865
timestamp 1679581782
transform 1 0 83616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_872
timestamp 1679581782
transform 1 0 84288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_879
timestamp 1679581782
transform 1 0 84960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_886
timestamp 1679581782
transform 1 0 85632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_893
timestamp 1679581782
transform 1 0 86304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_900
timestamp 1679581782
transform 1 0 86976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_907
timestamp 1679581782
transform 1 0 87648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_914
timestamp 1679581782
transform 1 0 88320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_921
timestamp 1679581782
transform 1 0 88992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_928
timestamp 1679581782
transform 1 0 89664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_935
timestamp 1679581782
transform 1 0 90336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_942
timestamp 1679581782
transform 1 0 91008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_949
timestamp 1679581782
transform 1 0 91680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_956
timestamp 1679581782
transform 1 0 92352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_963
timestamp 1679581782
transform 1 0 93024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_970
timestamp 1679581782
transform 1 0 93696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_977
timestamp 1679581782
transform 1 0 94368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_984
timestamp 1679581782
transform 1 0 95040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_991
timestamp 1679581782
transform 1 0 95712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_998
timestamp 1679581782
transform 1 0 96384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1005
timestamp 1679581782
transform 1 0 97056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1012
timestamp 1679581782
transform 1 0 97728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1019
timestamp 1679581782
transform 1 0 98400 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_1026
timestamp 1677580104
transform 1 0 99072 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_1028
timestamp 1677579658
transform 1 0 99264 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_4
timestamp 1679581782
transform 1 0 960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_11
timestamp 1679581782
transform 1 0 1632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_18
timestamp 1679581782
transform 1 0 2304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_25
timestamp 1679581782
transform 1 0 2976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_32
timestamp 1679581782
transform 1 0 3648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_39
timestamp 1679581782
transform 1 0 4320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_46
timestamp 1679581782
transform 1 0 4992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_53
timestamp 1679581782
transform 1 0 5664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_60
timestamp 1679581782
transform 1 0 6336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_67
timestamp 1679581782
transform 1 0 7008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_74
timestamp 1679581782
transform 1 0 7680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_81
timestamp 1679581782
transform 1 0 8352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_88
timestamp 1679581782
transform 1 0 9024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_95
timestamp 1679581782
transform 1 0 9696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_102
timestamp 1679581782
transform 1 0 10368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_109
timestamp 1679581782
transform 1 0 11040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_116
timestamp 1679581782
transform 1 0 11712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_123
timestamp 1679581782
transform 1 0 12384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_130
timestamp 1679581782
transform 1 0 13056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_137
timestamp 1679581782
transform 1 0 13728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_144
timestamp 1679581782
transform 1 0 14400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_151
timestamp 1679581782
transform 1 0 15072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_158
timestamp 1679581782
transform 1 0 15744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_165
timestamp 1679581782
transform 1 0 16416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_172
timestamp 1679581782
transform 1 0 17088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_179
timestamp 1679581782
transform 1 0 17760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_186
timestamp 1679581782
transform 1 0 18432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_193
timestamp 1679581782
transform 1 0 19104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_200
timestamp 1679581782
transform 1 0 19776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_207
timestamp 1679581782
transform 1 0 20448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_214
timestamp 1679581782
transform 1 0 21120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_221
timestamp 1679581782
transform 1 0 21792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_228
timestamp 1679581782
transform 1 0 22464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_235
timestamp 1679581782
transform 1 0 23136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_242
timestamp 1679581782
transform 1 0 23808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_249
timestamp 1679581782
transform 1 0 24480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_256
timestamp 1679581782
transform 1 0 25152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_263
timestamp 1679581782
transform 1 0 25824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_270
timestamp 1679581782
transform 1 0 26496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_277
timestamp 1679581782
transform 1 0 27168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_284
timestamp 1679581782
transform 1 0 27840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_291
timestamp 1679581782
transform 1 0 28512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_298
timestamp 1679581782
transform 1 0 29184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_305
timestamp 1679581782
transform 1 0 29856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_312
timestamp 1679581782
transform 1 0 30528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_319
timestamp 1679581782
transform 1 0 31200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_326
timestamp 1679581782
transform 1 0 31872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_333
timestamp 1679581782
transform 1 0 32544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_340
timestamp 1679581782
transform 1 0 33216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_347
timestamp 1679581782
transform 1 0 33888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_354
timestamp 1679581782
transform 1 0 34560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_361
timestamp 1679581782
transform 1 0 35232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_368
timestamp 1679581782
transform 1 0 35904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_375
timestamp 1679581782
transform 1 0 36576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_382
timestamp 1679581782
transform 1 0 37248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_389
timestamp 1679581782
transform 1 0 37920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_396
timestamp 1679581782
transform 1 0 38592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_403
timestamp 1679581782
transform 1 0 39264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_410
timestamp 1679581782
transform 1 0 39936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_417
timestamp 1679581782
transform 1 0 40608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_424
timestamp 1679581782
transform 1 0 41280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_431
timestamp 1679581782
transform 1 0 41952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_438
timestamp 1679581782
transform 1 0 42624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_445
timestamp 1679581782
transform 1 0 43296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_452
timestamp 1679581782
transform 1 0 43968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_459
timestamp 1679581782
transform 1 0 44640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_466
timestamp 1679581782
transform 1 0 45312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_473
timestamp 1679581782
transform 1 0 45984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_480
timestamp 1679581782
transform 1 0 46656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_487
timestamp 1679581782
transform 1 0 47328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_494
timestamp 1679581782
transform 1 0 48000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_501
timestamp 1679581782
transform 1 0 48672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_508
timestamp 1679581782
transform 1 0 49344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_515
timestamp 1679581782
transform 1 0 50016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_522
timestamp 1679581782
transform 1 0 50688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_529
timestamp 1679581782
transform 1 0 51360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_536
timestamp 1679581782
transform 1 0 52032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_543
timestamp 1679581782
transform 1 0 52704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_550
timestamp 1679581782
transform 1 0 53376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_557
timestamp 1679581782
transform 1 0 54048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_564
timestamp 1679581782
transform 1 0 54720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_571
timestamp 1679581782
transform 1 0 55392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_578
timestamp 1679581782
transform 1 0 56064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_585
timestamp 1679581782
transform 1 0 56736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_592
timestamp 1679581782
transform 1 0 57408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_599
timestamp 1679581782
transform 1 0 58080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_606
timestamp 1679581782
transform 1 0 58752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_613
timestamp 1679581782
transform 1 0 59424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_620
timestamp 1679581782
transform 1 0 60096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_627
timestamp 1679581782
transform 1 0 60768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_634
timestamp 1679581782
transform 1 0 61440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_641
timestamp 1679581782
transform 1 0 62112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_648
timestamp 1679581782
transform 1 0 62784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_655
timestamp 1679581782
transform 1 0 63456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_662
timestamp 1679581782
transform 1 0 64128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_669
timestamp 1679581782
transform 1 0 64800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_676
timestamp 1679581782
transform 1 0 65472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_683
timestamp 1679581782
transform 1 0 66144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_690
timestamp 1679581782
transform 1 0 66816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_697
timestamp 1679581782
transform 1 0 67488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_704
timestamp 1679581782
transform 1 0 68160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_711
timestamp 1679581782
transform 1 0 68832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_718
timestamp 1679581782
transform 1 0 69504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_725
timestamp 1679581782
transform 1 0 70176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_732
timestamp 1679581782
transform 1 0 70848 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_739
timestamp 1679581782
transform 1 0 71520 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_746
timestamp 1679581782
transform 1 0 72192 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_753
timestamp 1679581782
transform 1 0 72864 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_760
timestamp 1679581782
transform 1 0 73536 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_767
timestamp 1679581782
transform 1 0 74208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_774
timestamp 1679581782
transform 1 0 74880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_781
timestamp 1679581782
transform 1 0 75552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_788
timestamp 1679581782
transform 1 0 76224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_795
timestamp 1679581782
transform 1 0 76896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_802
timestamp 1679581782
transform 1 0 77568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_809
timestamp 1679581782
transform 1 0 78240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_816
timestamp 1679581782
transform 1 0 78912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_823
timestamp 1679581782
transform 1 0 79584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_830
timestamp 1679581782
transform 1 0 80256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_837
timestamp 1679581782
transform 1 0 80928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_844
timestamp 1679581782
transform 1 0 81600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_851
timestamp 1679581782
transform 1 0 82272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_858
timestamp 1679581782
transform 1 0 82944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_865
timestamp 1679581782
transform 1 0 83616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_872
timestamp 1679581782
transform 1 0 84288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_879
timestamp 1679581782
transform 1 0 84960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_886
timestamp 1679581782
transform 1 0 85632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_893
timestamp 1679581782
transform 1 0 86304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_900
timestamp 1679581782
transform 1 0 86976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_907
timestamp 1679581782
transform 1 0 87648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_914
timestamp 1679581782
transform 1 0 88320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_921
timestamp 1679581782
transform 1 0 88992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_928
timestamp 1679581782
transform 1 0 89664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_935
timestamp 1679581782
transform 1 0 90336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_942
timestamp 1679581782
transform 1 0 91008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_949
timestamp 1679581782
transform 1 0 91680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_956
timestamp 1679581782
transform 1 0 92352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_963
timestamp 1679581782
transform 1 0 93024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_970
timestamp 1679581782
transform 1 0 93696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_977
timestamp 1679581782
transform 1 0 94368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_984
timestamp 1679581782
transform 1 0 95040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_991
timestamp 1679581782
transform 1 0 95712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_998
timestamp 1679581782
transform 1 0 96384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1005
timestamp 1679581782
transform 1 0 97056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1012
timestamp 1679581782
transform 1 0 97728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1019
timestamp 1679581782
transform 1 0 98400 0 1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_1026
timestamp 1677580104
transform 1 0 99072 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_1028
timestamp 1677579658
transform 1 0 99264 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_4
timestamp 1677580104
transform 1 0 960 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_32
timestamp 1679581782
transform 1 0 3648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679581782
transform 1 0 4320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_46
timestamp 1679581782
transform 1 0 4992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_53
timestamp 1679581782
transform 1 0 5664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1679581782
transform 1 0 6336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_67
timestamp 1679581782
transform 1 0 7008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_74
timestamp 1679581782
transform 1 0 7680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679581782
transform 1 0 8352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679581782
transform 1 0 9024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679581782
transform 1 0 9696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679581782
transform 1 0 10368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_109
timestamp 1679581782
transform 1 0 11040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_116
timestamp 1679581782
transform 1 0 11712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_123
timestamp 1679581782
transform 1 0 12384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_130
timestamp 1679581782
transform 1 0 13056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_137
timestamp 1679581782
transform 1 0 13728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_144
timestamp 1679581782
transform 1 0 14400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_151
timestamp 1679581782
transform 1 0 15072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_158
timestamp 1679581782
transform 1 0 15744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_165
timestamp 1679581782
transform 1 0 16416 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_172
timestamp 1679581782
transform 1 0 17088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_179
timestamp 1679581782
transform 1 0 17760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_186
timestamp 1679581782
transform 1 0 18432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_193
timestamp 1679581782
transform 1 0 19104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_200
timestamp 1679581782
transform 1 0 19776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_207
timestamp 1679581782
transform 1 0 20448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_214
timestamp 1679581782
transform 1 0 21120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_221
timestamp 1679581782
transform 1 0 21792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_228
timestamp 1679581782
transform 1 0 22464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_235
timestamp 1679581782
transform 1 0 23136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_242
timestamp 1679581782
transform 1 0 23808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_249
timestamp 1679581782
transform 1 0 24480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_256
timestamp 1679581782
transform 1 0 25152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_263
timestamp 1679581782
transform 1 0 25824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_270
timestamp 1679581782
transform 1 0 26496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_277
timestamp 1679581782
transform 1 0 27168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_284
timestamp 1679581782
transform 1 0 27840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_291
timestamp 1679581782
transform 1 0 28512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_298
timestamp 1679581782
transform 1 0 29184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_305
timestamp 1679581782
transform 1 0 29856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_312
timestamp 1679581782
transform 1 0 30528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_319
timestamp 1679581782
transform 1 0 31200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_326
timestamp 1679581782
transform 1 0 31872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_333
timestamp 1679581782
transform 1 0 32544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_340
timestamp 1679581782
transform 1 0 33216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_347
timestamp 1679581782
transform 1 0 33888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_354
timestamp 1679581782
transform 1 0 34560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_361
timestamp 1679581782
transform 1 0 35232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_368
timestamp 1679581782
transform 1 0 35904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_375
timestamp 1679581782
transform 1 0 36576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_382
timestamp 1679581782
transform 1 0 37248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_389
timestamp 1679581782
transform 1 0 37920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_396
timestamp 1679581782
transform 1 0 38592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_403
timestamp 1679581782
transform 1 0 39264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_410
timestamp 1679581782
transform 1 0 39936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_417
timestamp 1679581782
transform 1 0 40608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_424
timestamp 1679581782
transform 1 0 41280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_431
timestamp 1679581782
transform 1 0 41952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_438
timestamp 1679581782
transform 1 0 42624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_445
timestamp 1679581782
transform 1 0 43296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_452
timestamp 1679581782
transform 1 0 43968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_459
timestamp 1679581782
transform 1 0 44640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_466
timestamp 1679581782
transform 1 0 45312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_473
timestamp 1679581782
transform 1 0 45984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_480
timestamp 1679581782
transform 1 0 46656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_487
timestamp 1679581782
transform 1 0 47328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_494
timestamp 1679581782
transform 1 0 48000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_501
timestamp 1679581782
transform 1 0 48672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_508
timestamp 1679581782
transform 1 0 49344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_515
timestamp 1679581782
transform 1 0 50016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_522
timestamp 1679581782
transform 1 0 50688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_529
timestamp 1679581782
transform 1 0 51360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_536
timestamp 1679581782
transform 1 0 52032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_543
timestamp 1679581782
transform 1 0 52704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_550
timestamp 1679581782
transform 1 0 53376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_557
timestamp 1679581782
transform 1 0 54048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_564
timestamp 1679581782
transform 1 0 54720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_571
timestamp 1679581782
transform 1 0 55392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_578
timestamp 1679581782
transform 1 0 56064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_585
timestamp 1679581782
transform 1 0 56736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_592
timestamp 1679581782
transform 1 0 57408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_599
timestamp 1679581782
transform 1 0 58080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_606
timestamp 1679581782
transform 1 0 58752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_613
timestamp 1679581782
transform 1 0 59424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_620
timestamp 1679581782
transform 1 0 60096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_627
timestamp 1679581782
transform 1 0 60768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_634
timestamp 1679581782
transform 1 0 61440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_641
timestamp 1679581782
transform 1 0 62112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_648
timestamp 1679581782
transform 1 0 62784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_655
timestamp 1679581782
transform 1 0 63456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_662
timestamp 1679581782
transform 1 0 64128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_669
timestamp 1679581782
transform 1 0 64800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_676
timestamp 1679581782
transform 1 0 65472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_683
timestamp 1679581782
transform 1 0 66144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_690
timestamp 1679581782
transform 1 0 66816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_697
timestamp 1679581782
transform 1 0 67488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_704
timestamp 1679581782
transform 1 0 68160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_711
timestamp 1679581782
transform 1 0 68832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_718
timestamp 1679581782
transform 1 0 69504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_725
timestamp 1679581782
transform 1 0 70176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_732
timestamp 1679581782
transform 1 0 70848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_739
timestamp 1679581782
transform 1 0 71520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_746
timestamp 1679581782
transform 1 0 72192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_753
timestamp 1679581782
transform 1 0 72864 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_760
timestamp 1679581782
transform 1 0 73536 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_767
timestamp 1679581782
transform 1 0 74208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_774
timestamp 1679581782
transform 1 0 74880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_781
timestamp 1679581782
transform 1 0 75552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_788
timestamp 1679581782
transform 1 0 76224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_795
timestamp 1679581782
transform 1 0 76896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_802
timestamp 1679581782
transform 1 0 77568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_809
timestamp 1679581782
transform 1 0 78240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_816
timestamp 1679581782
transform 1 0 78912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_823
timestamp 1679581782
transform 1 0 79584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_830
timestamp 1679581782
transform 1 0 80256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_837
timestamp 1679581782
transform 1 0 80928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_844
timestamp 1679581782
transform 1 0 81600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_851
timestamp 1679581782
transform 1 0 82272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_858
timestamp 1679581782
transform 1 0 82944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_865
timestamp 1679581782
transform 1 0 83616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_872
timestamp 1679581782
transform 1 0 84288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_879
timestamp 1679581782
transform 1 0 84960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_886
timestamp 1679581782
transform 1 0 85632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_893
timestamp 1679581782
transform 1 0 86304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_900
timestamp 1679581782
transform 1 0 86976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_907
timestamp 1679581782
transform 1 0 87648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_914
timestamp 1679581782
transform 1 0 88320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_921
timestamp 1679581782
transform 1 0 88992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_928
timestamp 1679581782
transform 1 0 89664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_935
timestamp 1679581782
transform 1 0 90336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_942
timestamp 1679581782
transform 1 0 91008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_949
timestamp 1679581782
transform 1 0 91680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_956
timestamp 1679581782
transform 1 0 92352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_963
timestamp 1679581782
transform 1 0 93024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_970
timestamp 1679581782
transform 1 0 93696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_977
timestamp 1679581782
transform 1 0 94368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_984
timestamp 1679581782
transform 1 0 95040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_991
timestamp 1679581782
transform 1 0 95712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_998
timestamp 1679577901
transform 1 0 96384 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_1002
timestamp 1677579658
transform 1 0 96768 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_1007
timestamp 1679581782
transform 1 0 97248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1014
timestamp 1679581782
transform 1 0 97920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1021
timestamp 1679581782
transform 1 0 98592 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_1028
timestamp 1677579658
transform 1 0 99264 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_4
timestamp 1679577901
transform 1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_16
timestamp 1679581782
transform 1 0 2112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_23
timestamp 1679581782
transform 1 0 2784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_30
timestamp 1679581782
transform 1 0 3456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_37
timestamp 1679581782
transform 1 0 4128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_44
timestamp 1679581782
transform 1 0 4800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_51
timestamp 1679581782
transform 1 0 5472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_58
timestamp 1679581782
transform 1 0 6144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_65
timestamp 1679581782
transform 1 0 6816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_72
timestamp 1679581782
transform 1 0 7488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_79
timestamp 1679581782
transform 1 0 8160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_86
timestamp 1679581782
transform 1 0 8832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_93
timestamp 1679581782
transform 1 0 9504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_100
timestamp 1679581782
transform 1 0 10176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_107
timestamp 1679581782
transform 1 0 10848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_114
timestamp 1679581782
transform 1 0 11520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_121
timestamp 1679581782
transform 1 0 12192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_128
timestamp 1679581782
transform 1 0 12864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_135
timestamp 1679581782
transform 1 0 13536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_142
timestamp 1679581782
transform 1 0 14208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_149
timestamp 1679581782
transform 1 0 14880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_156
timestamp 1679581782
transform 1 0 15552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_163
timestamp 1679581782
transform 1 0 16224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_170
timestamp 1679581782
transform 1 0 16896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_177
timestamp 1679581782
transform 1 0 17568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_184
timestamp 1679581782
transform 1 0 18240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_191
timestamp 1679581782
transform 1 0 18912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_198
timestamp 1679581782
transform 1 0 19584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_205
timestamp 1679581782
transform 1 0 20256 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_212
timestamp 1679581782
transform 1 0 20928 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_219
timestamp 1679581782
transform 1 0 21600 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_226
timestamp 1679581782
transform 1 0 22272 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_233
timestamp 1679581782
transform 1 0 22944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_240
timestamp 1679581782
transform 1 0 23616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_247
timestamp 1679581782
transform 1 0 24288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_254
timestamp 1679581782
transform 1 0 24960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_261
timestamp 1679581782
transform 1 0 25632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_268
timestamp 1679581782
transform 1 0 26304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_275
timestamp 1679581782
transform 1 0 26976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_282
timestamp 1679581782
transform 1 0 27648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_289
timestamp 1679581782
transform 1 0 28320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_296
timestamp 1679581782
transform 1 0 28992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_303
timestamp 1679581782
transform 1 0 29664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_310
timestamp 1679581782
transform 1 0 30336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_317
timestamp 1679581782
transform 1 0 31008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_324
timestamp 1679581782
transform 1 0 31680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_331
timestamp 1679581782
transform 1 0 32352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_338
timestamp 1679581782
transform 1 0 33024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_345
timestamp 1679581782
transform 1 0 33696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_352
timestamp 1679581782
transform 1 0 34368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_359
timestamp 1679581782
transform 1 0 35040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_366
timestamp 1679581782
transform 1 0 35712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_373
timestamp 1679581782
transform 1 0 36384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_380
timestamp 1679581782
transform 1 0 37056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_387
timestamp 1679581782
transform 1 0 37728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_394
timestamp 1679581782
transform 1 0 38400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_401
timestamp 1679581782
transform 1 0 39072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_408
timestamp 1679581782
transform 1 0 39744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_415
timestamp 1679581782
transform 1 0 40416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_422
timestamp 1679581782
transform 1 0 41088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_429
timestamp 1679581782
transform 1 0 41760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_436
timestamp 1679581782
transform 1 0 42432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_443
timestamp 1679581782
transform 1 0 43104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_450
timestamp 1679581782
transform 1 0 43776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_457
timestamp 1679581782
transform 1 0 44448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_464
timestamp 1679581782
transform 1 0 45120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_471
timestamp 1679581782
transform 1 0 45792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_478
timestamp 1679581782
transform 1 0 46464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_485
timestamp 1679581782
transform 1 0 47136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_492
timestamp 1679581782
transform 1 0 47808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_499
timestamp 1679581782
transform 1 0 48480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_506
timestamp 1679581782
transform 1 0 49152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_513
timestamp 1679581782
transform 1 0 49824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_520
timestamp 1679581782
transform 1 0 50496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_527
timestamp 1679581782
transform 1 0 51168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_534
timestamp 1679581782
transform 1 0 51840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_541
timestamp 1679581782
transform 1 0 52512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_548
timestamp 1679581782
transform 1 0 53184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_555
timestamp 1679581782
transform 1 0 53856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_562
timestamp 1679581782
transform 1 0 54528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_569
timestamp 1679581782
transform 1 0 55200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_576
timestamp 1679581782
transform 1 0 55872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_583
timestamp 1679581782
transform 1 0 56544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_590
timestamp 1679581782
transform 1 0 57216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_597
timestamp 1679581782
transform 1 0 57888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_604
timestamp 1679581782
transform 1 0 58560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_611
timestamp 1679581782
transform 1 0 59232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_618
timestamp 1679581782
transform 1 0 59904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_625
timestamp 1679581782
transform 1 0 60576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_632
timestamp 1679581782
transform 1 0 61248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_639
timestamp 1679581782
transform 1 0 61920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_646
timestamp 1679581782
transform 1 0 62592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_653
timestamp 1679581782
transform 1 0 63264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_660
timestamp 1679581782
transform 1 0 63936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_667
timestamp 1679581782
transform 1 0 64608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_674
timestamp 1679581782
transform 1 0 65280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_681
timestamp 1679581782
transform 1 0 65952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_688
timestamp 1679581782
transform 1 0 66624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_695
timestamp 1679581782
transform 1 0 67296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_702
timestamp 1679581782
transform 1 0 67968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_709
timestamp 1679581782
transform 1 0 68640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_716
timestamp 1679581782
transform 1 0 69312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_723
timestamp 1679581782
transform 1 0 69984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_730
timestamp 1679581782
transform 1 0 70656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_737
timestamp 1679581782
transform 1 0 71328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_744
timestamp 1679581782
transform 1 0 72000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_751
timestamp 1679581782
transform 1 0 72672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_758
timestamp 1679581782
transform 1 0 73344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_765
timestamp 1679581782
transform 1 0 74016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_772
timestamp 1679577901
transform 1 0 74688 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_780
timestamp 1679581782
transform 1 0 75456 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_787
timestamp 1677580104
transform 1 0 76128 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_789
timestamp 1677579658
transform 1 0 76320 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_794
timestamp 1679581782
transform 1 0 76800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_801
timestamp 1679581782
transform 1 0 77472 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_811
timestamp 1677579658
transform 1 0 78432 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_816
timestamp 1679581782
transform 1 0 78912 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_823
timestamp 1677580104
transform 1 0 79584 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_825
timestamp 1677579658
transform 1 0 79776 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_833
timestamp 1679577901
transform 1 0 80544 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_837
timestamp 1677579658
transform 1 0 80928 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_841
timestamp 1679581782
transform 1 0 81312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_848
timestamp 1679577901
transform 1 0 81984 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_856
timestamp 1679581782
transform 1 0 82752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_866
timestamp 1679581782
transform 1 0 83712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_873
timestamp 1679581782
transform 1 0 84384 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_880
timestamp 1677580104
transform 1 0 85056 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_882
timestamp 1677579658
transform 1 0 85248 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_886
timestamp 1679581782
transform 1 0 85632 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_893
timestamp 1677580104
transform 1 0 86304 0 1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_899
timestamp 1679577901
transform 1 0 86880 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_903
timestamp 1677580104
transform 1 0 87264 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_908
timestamp 1679581782
transform 1 0 87744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_915
timestamp 1679577901
transform 1 0 88416 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_923
timestamp 1677580104
transform 1 0 89184 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_925
timestamp 1677579658
transform 1 0 89376 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_929
timestamp 1679577901
transform 1 0 89760 0 1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_6_937
timestamp 1679581782
transform 1 0 90528 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_944
timestamp 1677580104
transform 1 0 91200 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_946
timestamp 1677579658
transform 1 0 91392 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_950
timestamp 1679581782
transform 1 0 91776 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_957
timestamp 1677580104
transform 1 0 92448 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_959
timestamp 1677579658
transform 1 0 92640 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_963
timestamp 1677579658
transform 1 0 93024 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_967
timestamp 1677579658
transform 1 0 93408 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_974
timestamp 1679581782
transform 1 0 94080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_981
timestamp 1679581782
transform 1 0 94752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_995
timestamp 1679581782
transform 1 0 96096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1002
timestamp 1679581782
transform 1 0 96768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1009
timestamp 1679581782
transform 1 0 97440 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_1016
timestamp 1677579658
transform 1 0 98112 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_1020
timestamp 1677579658
transform 1 0 98496 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_1024
timestamp 1679577901
transform 1 0 98880 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_1028
timestamp 1677579658
transform 1 0 99264 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_11
timestamp 1679581782
transform 1 0 1632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_18
timestamp 1679581782
transform 1 0 2304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_25
timestamp 1679581782
transform 1 0 2976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_32
timestamp 1679581782
transform 1 0 3648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_39
timestamp 1679581782
transform 1 0 4320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_46
timestamp 1679581782
transform 1 0 4992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_53
timestamp 1679581782
transform 1 0 5664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_60
timestamp 1679581782
transform 1 0 6336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_67
timestamp 1679581782
transform 1 0 7008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_74
timestamp 1679581782
transform 1 0 7680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_81
timestamp 1679581782
transform 1 0 8352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_88
timestamp 1679581782
transform 1 0 9024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_95
timestamp 1679581782
transform 1 0 9696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_102
timestamp 1679581782
transform 1 0 10368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_109
timestamp 1679581782
transform 1 0 11040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_116
timestamp 1679581782
transform 1 0 11712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_123
timestamp 1679581782
transform 1 0 12384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_130
timestamp 1679581782
transform 1 0 13056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_137
timestamp 1679581782
transform 1 0 13728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_144
timestamp 1679581782
transform 1 0 14400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_151
timestamp 1679581782
transform 1 0 15072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_158
timestamp 1679581782
transform 1 0 15744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_165
timestamp 1679581782
transform 1 0 16416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_172
timestamp 1679581782
transform 1 0 17088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_179
timestamp 1679581782
transform 1 0 17760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_186
timestamp 1679581782
transform 1 0 18432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_193
timestamp 1679581782
transform 1 0 19104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_200
timestamp 1679581782
transform 1 0 19776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_207
timestamp 1679581782
transform 1 0 20448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_214
timestamp 1679581782
transform 1 0 21120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_221
timestamp 1679581782
transform 1 0 21792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_228
timestamp 1679581782
transform 1 0 22464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_235
timestamp 1679581782
transform 1 0 23136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_242
timestamp 1679581782
transform 1 0 23808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_249
timestamp 1679581782
transform 1 0 24480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_256
timestamp 1679581782
transform 1 0 25152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_263
timestamp 1679581782
transform 1 0 25824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_270
timestamp 1679581782
transform 1 0 26496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_277
timestamp 1679581782
transform 1 0 27168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_284
timestamp 1679581782
transform 1 0 27840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_291
timestamp 1679581782
transform 1 0 28512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_298
timestamp 1679581782
transform 1 0 29184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_305
timestamp 1679581782
transform 1 0 29856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_312
timestamp 1679581782
transform 1 0 30528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_319
timestamp 1679581782
transform 1 0 31200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_326
timestamp 1679581782
transform 1 0 31872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_333
timestamp 1679581782
transform 1 0 32544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_340
timestamp 1679581782
transform 1 0 33216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_347
timestamp 1679581782
transform 1 0 33888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_354
timestamp 1679581782
transform 1 0 34560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_361
timestamp 1679581782
transform 1 0 35232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_368
timestamp 1679581782
transform 1 0 35904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_375
timestamp 1679581782
transform 1 0 36576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_382
timestamp 1679581782
transform 1 0 37248 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_389
timestamp 1679581782
transform 1 0 37920 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_396
timestamp 1679581782
transform 1 0 38592 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_403
timestamp 1679581782
transform 1 0 39264 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_410
timestamp 1679581782
transform 1 0 39936 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_417
timestamp 1679581782
transform 1 0 40608 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_424
timestamp 1679581782
transform 1 0 41280 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_431
timestamp 1679581782
transform 1 0 41952 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_438
timestamp 1679581782
transform 1 0 42624 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_445
timestamp 1679581782
transform 1 0 43296 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_452
timestamp 1679581782
transform 1 0 43968 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_459
timestamp 1679581782
transform 1 0 44640 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_466
timestamp 1679581782
transform 1 0 45312 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_473
timestamp 1679581782
transform 1 0 45984 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_480
timestamp 1679581782
transform 1 0 46656 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_487
timestamp 1679581782
transform 1 0 47328 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_494
timestamp 1679581782
transform 1 0 48000 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_501
timestamp 1679581782
transform 1 0 48672 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_508
timestamp 1679581782
transform 1 0 49344 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_515
timestamp 1679581782
transform 1 0 50016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_522
timestamp 1679581782
transform 1 0 50688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_529
timestamp 1679581782
transform 1 0 51360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_536
timestamp 1679581782
transform 1 0 52032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_543
timestamp 1679581782
transform 1 0 52704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_550
timestamp 1679581782
transform 1 0 53376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_557
timestamp 1679581782
transform 1 0 54048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_564
timestamp 1679581782
transform 1 0 54720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_571
timestamp 1679581782
transform 1 0 55392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_578
timestamp 1679581782
transform 1 0 56064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_585
timestamp 1679581782
transform 1 0 56736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_592
timestamp 1679581782
transform 1 0 57408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_599
timestamp 1679581782
transform 1 0 58080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_606
timestamp 1679581782
transform 1 0 58752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_613
timestamp 1679581782
transform 1 0 59424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_620
timestamp 1679581782
transform 1 0 60096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_627
timestamp 1679581782
transform 1 0 60768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_634
timestamp 1679581782
transform 1 0 61440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_641
timestamp 1679581782
transform 1 0 62112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_648
timestamp 1679581782
transform 1 0 62784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_655
timestamp 1679581782
transform 1 0 63456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_662
timestamp 1679581782
transform 1 0 64128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_669
timestamp 1679581782
transform 1 0 64800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_676
timestamp 1679581782
transform 1 0 65472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_683
timestamp 1679581782
transform 1 0 66144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_690
timestamp 1679581782
transform 1 0 66816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_697
timestamp 1679581782
transform 1 0 67488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_704
timestamp 1679581782
transform 1 0 68160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_711
timestamp 1679581782
transform 1 0 68832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_718
timestamp 1679581782
transform 1 0 69504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_725
timestamp 1679581782
transform 1 0 70176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_732
timestamp 1679581782
transform 1 0 70848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_739
timestamp 1679581782
transform 1 0 71520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_746
timestamp 1679581782
transform 1 0 72192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_753
timestamp 1679581782
transform 1 0 72864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_760
timestamp 1679577901
transform 1 0 73536 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_764
timestamp 1677579658
transform 1 0 73920 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_785
timestamp 1677580104
transform 1 0 75936 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_787
timestamp 1677579658
transform 1 0 76128 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_791
timestamp 1677579658
transform 1 0 76512 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_799
timestamp 1679577901
transform 1 0 77280 0 -1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_7_811
timestamp 1679577901
transform 1 0 78432 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_819
timestamp 1677579658
transform 1 0 79200 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_824
timestamp 1677580104
transform 1 0 79680 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_829
timestamp 1677580104
transform 1 0 80160 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_835
timestamp 1677579658
transform 1 0 80736 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_840
timestamp 1677579658
transform 1 0 81216 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_852
timestamp 1677580104
transform 1 0 82368 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_854
timestamp 1677579658
transform 1 0 82560 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_859
timestamp 1677579658
transform 1 0 83040 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_864
timestamp 1677579658
transform 1 0 83520 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_869
timestamp 1677579658
transform 1 0 84000 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_889
timestamp 1677579658
transform 1 0 85920 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_894
timestamp 1679577901
transform 1 0 86400 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_902
timestamp 1677579658
transform 1 0 87168 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_921
timestamp 1677579658
transform 1 0 88992 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_929
timestamp 1679577901
transform 1 0 89760 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_933
timestamp 1677580104
transform 1 0 90144 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_939
timestamp 1677579658
transform 1 0 90720 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_947
timestamp 1677579658
transform 1 0 91488 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_952
timestamp 1677579658
transform 1 0 91968 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_960
timestamp 1677580104
transform 1 0 92736 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_970
timestamp 1677579658
transform 1 0 93696 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_979
timestamp 1677579658
transform 1 0 94560 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_983
timestamp 1677579658
transform 1 0 94944 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_988
timestamp 1677579658
transform 1 0 95424 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_995
timestamp 1677580104
transform 1 0 96096 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_1001
timestamp 1677580104
transform 1 0 96672 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_1010
timestamp 1677579658
transform 1 0 97536 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_1017
timestamp 1679581782
transform 1 0 98208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_1024
timestamp 1679577901
transform 1 0 98880 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_1028
timestamp 1677579658
transform 1 0 99264 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_4
timestamp 1679581782
transform 1 0 960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_11
timestamp 1679581782
transform 1 0 1632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_18
timestamp 1679581782
transform 1 0 2304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_25
timestamp 1679581782
transform 1 0 2976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_32
timestamp 1679581782
transform 1 0 3648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_39
timestamp 1679581782
transform 1 0 4320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_46
timestamp 1679581782
transform 1 0 4992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_53
timestamp 1679581782
transform 1 0 5664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_60
timestamp 1679581782
transform 1 0 6336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_67
timestamp 1679581782
transform 1 0 7008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_74
timestamp 1679581782
transform 1 0 7680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_81
timestamp 1679581782
transform 1 0 8352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_88
timestamp 1679581782
transform 1 0 9024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_95
timestamp 1679581782
transform 1 0 9696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_102
timestamp 1679581782
transform 1 0 10368 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_109
timestamp 1679581782
transform 1 0 11040 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_116
timestamp 1679581782
transform 1 0 11712 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_123
timestamp 1679581782
transform 1 0 12384 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_130
timestamp 1679581782
transform 1 0 13056 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_137
timestamp 1679581782
transform 1 0 13728 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_144
timestamp 1679581782
transform 1 0 14400 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_151
timestamp 1679581782
transform 1 0 15072 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_158
timestamp 1679581782
transform 1 0 15744 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_165
timestamp 1679581782
transform 1 0 16416 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_172
timestamp 1679581782
transform 1 0 17088 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_179
timestamp 1679581782
transform 1 0 17760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_186
timestamp 1679581782
transform 1 0 18432 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_193
timestamp 1679581782
transform 1 0 19104 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_200
timestamp 1679581782
transform 1 0 19776 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_207
timestamp 1679581782
transform 1 0 20448 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_214
timestamp 1679581782
transform 1 0 21120 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_221
timestamp 1679581782
transform 1 0 21792 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_228
timestamp 1679581782
transform 1 0 22464 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_235
timestamp 1679581782
transform 1 0 23136 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_242
timestamp 1679581782
transform 1 0 23808 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_249
timestamp 1679581782
transform 1 0 24480 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_256
timestamp 1679581782
transform 1 0 25152 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_263
timestamp 1679581782
transform 1 0 25824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_270
timestamp 1679581782
transform 1 0 26496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_277
timestamp 1679581782
transform 1 0 27168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_284
timestamp 1679581782
transform 1 0 27840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_291
timestamp 1679581782
transform 1 0 28512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_298
timestamp 1679581782
transform 1 0 29184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_305
timestamp 1679581782
transform 1 0 29856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_312
timestamp 1679581782
transform 1 0 30528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_319
timestamp 1679581782
transform 1 0 31200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_326
timestamp 1679581782
transform 1 0 31872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_333
timestamp 1679581782
transform 1 0 32544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_340
timestamp 1679581782
transform 1 0 33216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_347
timestamp 1679581782
transform 1 0 33888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_354
timestamp 1679581782
transform 1 0 34560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_361
timestamp 1679581782
transform 1 0 35232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_368
timestamp 1679581782
transform 1 0 35904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_375
timestamp 1679581782
transform 1 0 36576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_382
timestamp 1679581782
transform 1 0 37248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_389
timestamp 1679581782
transform 1 0 37920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_396
timestamp 1679581782
transform 1 0 38592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_403
timestamp 1679581782
transform 1 0 39264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_410
timestamp 1679581782
transform 1 0 39936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_417
timestamp 1679581782
transform 1 0 40608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_424
timestamp 1679581782
transform 1 0 41280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_431
timestamp 1679581782
transform 1 0 41952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_438
timestamp 1679581782
transform 1 0 42624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_445
timestamp 1679581782
transform 1 0 43296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_452
timestamp 1679581782
transform 1 0 43968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_459
timestamp 1679581782
transform 1 0 44640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_466
timestamp 1679581782
transform 1 0 45312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_473
timestamp 1679581782
transform 1 0 45984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_480
timestamp 1679581782
transform 1 0 46656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_487
timestamp 1679581782
transform 1 0 47328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_494
timestamp 1679581782
transform 1 0 48000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_501
timestamp 1679581782
transform 1 0 48672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_508
timestamp 1679581782
transform 1 0 49344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_515
timestamp 1679581782
transform 1 0 50016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_522
timestamp 1679581782
transform 1 0 50688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_529
timestamp 1679581782
transform 1 0 51360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_536
timestamp 1679581782
transform 1 0 52032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_543
timestamp 1679581782
transform 1 0 52704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_550
timestamp 1679581782
transform 1 0 53376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_557
timestamp 1679581782
transform 1 0 54048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_564
timestamp 1679581782
transform 1 0 54720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_571
timestamp 1679581782
transform 1 0 55392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_578
timestamp 1679581782
transform 1 0 56064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_585
timestamp 1679581782
transform 1 0 56736 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_592
timestamp 1679581782
transform 1 0 57408 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_599
timestamp 1679581782
transform 1 0 58080 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_606
timestamp 1679581782
transform 1 0 58752 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_613
timestamp 1679581782
transform 1 0 59424 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_620
timestamp 1679581782
transform 1 0 60096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_627
timestamp 1679581782
transform 1 0 60768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_634
timestamp 1679581782
transform 1 0 61440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_641
timestamp 1679581782
transform 1 0 62112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_648
timestamp 1679581782
transform 1 0 62784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_655
timestamp 1679581782
transform 1 0 63456 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_662
timestamp 1679581782
transform 1 0 64128 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_669
timestamp 1679581782
transform 1 0 64800 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_676
timestamp 1679581782
transform 1 0 65472 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_683
timestamp 1679581782
transform 1 0 66144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_690
timestamp 1679581782
transform 1 0 66816 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_697
timestamp 1679581782
transform 1 0 67488 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_704
timestamp 1679581782
transform 1 0 68160 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_711
timestamp 1679581782
transform 1 0 68832 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_718
timestamp 1679581782
transform 1 0 69504 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_725
timestamp 1679581782
transform 1 0 70176 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_732
timestamp 1679581782
transform 1 0 70848 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_739
timestamp 1679581782
transform 1 0 71520 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_746
timestamp 1679581782
transform 1 0 72192 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_753
timestamp 1679577901
transform 1 0 72864 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_764
timestamp 1677579658
transform 1 0 73920 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_781
timestamp 1677579658
transform 1 0 75552 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_790
timestamp 1677579658
transform 1 0 76416 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_812
timestamp 1677579658
transform 1 0 78528 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_816
timestamp 1677579658
transform 1 0 78912 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_831
timestamp 1677579658
transform 1 0 80352 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_853
timestamp 1677579658
transform 1 0 82464 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_864
timestamp 1677580104
transform 1 0 83520 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_873
timestamp 1677579658
transform 1 0 84384 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_888
timestamp 1677580104
transform 1 0 85824 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_914
timestamp 1677580104
transform 1 0 88320 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_923
timestamp 1677580104
transform 1 0 89184 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_933
timestamp 1677579658
transform 1 0 90144 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_940
timestamp 1677579658
transform 1 0 90816 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_952
timestamp 1677579658
transform 1 0 91968 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_968
timestamp 1677579658
transform 1 0 93504 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_988
timestamp 1677580104
transform 1 0 95424 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_1012
timestamp 1677580104
transform 1 0 97728 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_1018
timestamp 1677579658
transform 1 0 98304 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_1023
timestamp 1679577901
transform 1 0 98784 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_1027
timestamp 1677580104
transform 1 0 99168 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_4
timestamp 1679577901
transform 1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_8
timestamp 1677579658
transform 1 0 1344 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_13
timestamp 1679581782
transform 1 0 1824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_20
timestamp 1679581782
transform 1 0 2496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_27
timestamp 1679581782
transform 1 0 3168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_34
timestamp 1679581782
transform 1 0 3840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_41
timestamp 1679581782
transform 1 0 4512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_48
timestamp 1679581782
transform 1 0 5184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_55
timestamp 1679581782
transform 1 0 5856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_62
timestamp 1679581782
transform 1 0 6528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_69
timestamp 1679581782
transform 1 0 7200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_76
timestamp 1679581782
transform 1 0 7872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_83
timestamp 1679581782
transform 1 0 8544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_90
timestamp 1679581782
transform 1 0 9216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_97
timestamp 1679581782
transform 1 0 9888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_104
timestamp 1679581782
transform 1 0 10560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_111
timestamp 1679581782
transform 1 0 11232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_118
timestamp 1679581782
transform 1 0 11904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_125
timestamp 1679581782
transform 1 0 12576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_132
timestamp 1679581782
transform 1 0 13248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_139
timestamp 1679581782
transform 1 0 13920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_146
timestamp 1679581782
transform 1 0 14592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_153
timestamp 1679581782
transform 1 0 15264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_160
timestamp 1679581782
transform 1 0 15936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_167
timestamp 1679581782
transform 1 0 16608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_174
timestamp 1679581782
transform 1 0 17280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_181
timestamp 1679581782
transform 1 0 17952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_188
timestamp 1679581782
transform 1 0 18624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_195
timestamp 1679581782
transform 1 0 19296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_202
timestamp 1679581782
transform 1 0 19968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_209
timestamp 1679581782
transform 1 0 20640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_216
timestamp 1679581782
transform 1 0 21312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_223
timestamp 1679581782
transform 1 0 21984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_230
timestamp 1679581782
transform 1 0 22656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_237
timestamp 1679581782
transform 1 0 23328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_244
timestamp 1679581782
transform 1 0 24000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_251
timestamp 1679581782
transform 1 0 24672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_258
timestamp 1679581782
transform 1 0 25344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_265
timestamp 1679581782
transform 1 0 26016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_272
timestamp 1679581782
transform 1 0 26688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_279
timestamp 1679581782
transform 1 0 27360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_286
timestamp 1679581782
transform 1 0 28032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_293
timestamp 1679581782
transform 1 0 28704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_300
timestamp 1679581782
transform 1 0 29376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_307
timestamp 1679581782
transform 1 0 30048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_314
timestamp 1679581782
transform 1 0 30720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_321
timestamp 1679581782
transform 1 0 31392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_328
timestamp 1679581782
transform 1 0 32064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_335
timestamp 1679581782
transform 1 0 32736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_342
timestamp 1679581782
transform 1 0 33408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_349
timestamp 1679581782
transform 1 0 34080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_356
timestamp 1679581782
transform 1 0 34752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_363
timestamp 1679581782
transform 1 0 35424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_370
timestamp 1679581782
transform 1 0 36096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_377
timestamp 1679581782
transform 1 0 36768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_384
timestamp 1679581782
transform 1 0 37440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_391
timestamp 1679581782
transform 1 0 38112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_398
timestamp 1679581782
transform 1 0 38784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_405
timestamp 1679581782
transform 1 0 39456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_412
timestamp 1679581782
transform 1 0 40128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_419
timestamp 1679581782
transform 1 0 40800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_426
timestamp 1679581782
transform 1 0 41472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_433
timestamp 1679581782
transform 1 0 42144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_440
timestamp 1679581782
transform 1 0 42816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_447
timestamp 1679581782
transform 1 0 43488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_454
timestamp 1679581782
transform 1 0 44160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_461
timestamp 1679581782
transform 1 0 44832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_468
timestamp 1679581782
transform 1 0 45504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_475
timestamp 1679581782
transform 1 0 46176 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_482
timestamp 1679581782
transform 1 0 46848 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_489
timestamp 1679581782
transform 1 0 47520 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_496
timestamp 1679581782
transform 1 0 48192 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_503
timestamp 1679581782
transform 1 0 48864 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_510
timestamp 1679581782
transform 1 0 49536 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_517
timestamp 1679581782
transform 1 0 50208 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_524
timestamp 1679581782
transform 1 0 50880 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_531
timestamp 1679581782
transform 1 0 51552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_538
timestamp 1679581782
transform 1 0 52224 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_545
timestamp 1679581782
transform 1 0 52896 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_552
timestamp 1679581782
transform 1 0 53568 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_559
timestamp 1679581782
transform 1 0 54240 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_566
timestamp 1679581782
transform 1 0 54912 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_573
timestamp 1679581782
transform 1 0 55584 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_580
timestamp 1679581782
transform 1 0 56256 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_587
timestamp 1679581782
transform 1 0 56928 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_594
timestamp 1679581782
transform 1 0 57600 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_601
timestamp 1679581782
transform 1 0 58272 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_608
timestamp 1679581782
transform 1 0 58944 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_615
timestamp 1679581782
transform 1 0 59616 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_622
timestamp 1679581782
transform 1 0 60288 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_629
timestamp 1679581782
transform 1 0 60960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_636
timestamp 1679581782
transform 1 0 61632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_643
timestamp 1679581782
transform 1 0 62304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_650
timestamp 1679581782
transform 1 0 62976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_657
timestamp 1679581782
transform 1 0 63648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_664
timestamp 1679581782
transform 1 0 64320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_671
timestamp 1679581782
transform 1 0 64992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_678
timestamp 1679581782
transform 1 0 65664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_685
timestamp 1679581782
transform 1 0 66336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_692
timestamp 1679581782
transform 1 0 67008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_699
timestamp 1679581782
transform 1 0 67680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_706
timestamp 1679581782
transform 1 0 68352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_713
timestamp 1679581782
transform 1 0 69024 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_720
timestamp 1677580104
transform 1 0 69696 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_722
timestamp 1677579658
transform 1 0 69888 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_4
timestamp 1679577901
transform 1 0 960 0 1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_16
timestamp 1679581782
transform 1 0 2112 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_23
timestamp 1679581782
transform 1 0 2784 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_30
timestamp 1679581782
transform 1 0 3456 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_37
timestamp 1679581782
transform 1 0 4128 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_44
timestamp 1679581782
transform 1 0 4800 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_51
timestamp 1679581782
transform 1 0 5472 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_58
timestamp 1679581782
transform 1 0 6144 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_65
timestamp 1679581782
transform 1 0 6816 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_72
timestamp 1679581782
transform 1 0 7488 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_79
timestamp 1679581782
transform 1 0 8160 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_86
timestamp 1679581782
transform 1 0 8832 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_93
timestamp 1679581782
transform 1 0 9504 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_100
timestamp 1679581782
transform 1 0 10176 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_107
timestamp 1679581782
transform 1 0 10848 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_114
timestamp 1679581782
transform 1 0 11520 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_121
timestamp 1679581782
transform 1 0 12192 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_128
timestamp 1679581782
transform 1 0 12864 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_135
timestamp 1679581782
transform 1 0 13536 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_142
timestamp 1679581782
transform 1 0 14208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_149
timestamp 1679581782
transform 1 0 14880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_156
timestamp 1679581782
transform 1 0 15552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_163
timestamp 1679581782
transform 1 0 16224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_170
timestamp 1679581782
transform 1 0 16896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_177
timestamp 1679581782
transform 1 0 17568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_184
timestamp 1679581782
transform 1 0 18240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_191
timestamp 1679581782
transform 1 0 18912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_198
timestamp 1679581782
transform 1 0 19584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_205
timestamp 1679581782
transform 1 0 20256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_212
timestamp 1679581782
transform 1 0 20928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_219
timestamp 1679581782
transform 1 0 21600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_226
timestamp 1679581782
transform 1 0 22272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_233
timestamp 1679581782
transform 1 0 22944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_240
timestamp 1679581782
transform 1 0 23616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_247
timestamp 1679581782
transform 1 0 24288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_254
timestamp 1679581782
transform 1 0 24960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_261
timestamp 1679581782
transform 1 0 25632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_268
timestamp 1679581782
transform 1 0 26304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_275
timestamp 1679581782
transform 1 0 26976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_282
timestamp 1679581782
transform 1 0 27648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_289
timestamp 1679581782
transform 1 0 28320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_296
timestamp 1679581782
transform 1 0 28992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_303
timestamp 1679581782
transform 1 0 29664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_310
timestamp 1679581782
transform 1 0 30336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_317
timestamp 1679581782
transform 1 0 31008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_324
timestamp 1679581782
transform 1 0 31680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_331
timestamp 1679581782
transform 1 0 32352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_338
timestamp 1679581782
transform 1 0 33024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_345
timestamp 1679581782
transform 1 0 33696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_352
timestamp 1679581782
transform 1 0 34368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_359
timestamp 1679581782
transform 1 0 35040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_366
timestamp 1679581782
transform 1 0 35712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_373
timestamp 1679581782
transform 1 0 36384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_380
timestamp 1679581782
transform 1 0 37056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_387
timestamp 1679581782
transform 1 0 37728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_394
timestamp 1679581782
transform 1 0 38400 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_401
timestamp 1679581782
transform 1 0 39072 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_408
timestamp 1679581782
transform 1 0 39744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_415
timestamp 1679581782
transform 1 0 40416 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_422
timestamp 1679581782
transform 1 0 41088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_429
timestamp 1679581782
transform 1 0 41760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_436
timestamp 1679581782
transform 1 0 42432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_443
timestamp 1679581782
transform 1 0 43104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_450
timestamp 1679581782
transform 1 0 43776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_457
timestamp 1679581782
transform 1 0 44448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_464
timestamp 1679581782
transform 1 0 45120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_471
timestamp 1679581782
transform 1 0 45792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_478
timestamp 1679581782
transform 1 0 46464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_485
timestamp 1679581782
transform 1 0 47136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_492
timestamp 1679581782
transform 1 0 47808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_499
timestamp 1679581782
transform 1 0 48480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_506
timestamp 1679581782
transform 1 0 49152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_513
timestamp 1679581782
transform 1 0 49824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_520
timestamp 1679581782
transform 1 0 50496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_527
timestamp 1679581782
transform 1 0 51168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_534
timestamp 1679581782
transform 1 0 51840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_541
timestamp 1679581782
transform 1 0 52512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_548
timestamp 1679581782
transform 1 0 53184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_555
timestamp 1679581782
transform 1 0 53856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_562
timestamp 1679581782
transform 1 0 54528 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_569
timestamp 1679581782
transform 1 0 55200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_576
timestamp 1679581782
transform 1 0 55872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_583
timestamp 1679581782
transform 1 0 56544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_590
timestamp 1679581782
transform 1 0 57216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_597
timestamp 1679581782
transform 1 0 57888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_604
timestamp 1679581782
transform 1 0 58560 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_611
timestamp 1679581782
transform 1 0 59232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_618
timestamp 1679581782
transform 1 0 59904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_625
timestamp 1679581782
transform 1 0 60576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_632
timestamp 1679581782
transform 1 0 61248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_639
timestamp 1679581782
transform 1 0 61920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_646
timestamp 1679581782
transform 1 0 62592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_653
timestamp 1679581782
transform 1 0 63264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_660
timestamp 1679581782
transform 1 0 63936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_667
timestamp 1679581782
transform 1 0 64608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_674
timestamp 1679581782
transform 1 0 65280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_681
timestamp 1679581782
transform 1 0 65952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_688
timestamp 1679581782
transform 1 0 66624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_695
timestamp 1679581782
transform 1 0 67296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_702
timestamp 1679581782
transform 1 0 67968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_709
timestamp 1679581782
transform 1 0 68640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_716
timestamp 1679581782
transform 1 0 69312 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_4
timestamp 1677580104
transform 1 0 960 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_6
timestamp 1677579658
transform 1 0 1152 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_11
timestamp 1679581782
transform 1 0 1632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_18
timestamp 1679581782
transform 1 0 2304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_25
timestamp 1679581782
transform 1 0 2976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_32
timestamp 1679581782
transform 1 0 3648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_39
timestamp 1679581782
transform 1 0 4320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_46
timestamp 1679581782
transform 1 0 4992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_53
timestamp 1679581782
transform 1 0 5664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_60
timestamp 1679581782
transform 1 0 6336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_67
timestamp 1679581782
transform 1 0 7008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_74
timestamp 1679581782
transform 1 0 7680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_81
timestamp 1679581782
transform 1 0 8352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_88
timestamp 1679581782
transform 1 0 9024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_95
timestamp 1679581782
transform 1 0 9696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_102
timestamp 1679581782
transform 1 0 10368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_109
timestamp 1679581782
transform 1 0 11040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_116
timestamp 1679581782
transform 1 0 11712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_123
timestamp 1679581782
transform 1 0 12384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_130
timestamp 1679581782
transform 1 0 13056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_137
timestamp 1679581782
transform 1 0 13728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_144
timestamp 1679581782
transform 1 0 14400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_151
timestamp 1679581782
transform 1 0 15072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_158
timestamp 1679581782
transform 1 0 15744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_165
timestamp 1679581782
transform 1 0 16416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_172
timestamp 1679581782
transform 1 0 17088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_179
timestamp 1679581782
transform 1 0 17760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_186
timestamp 1679581782
transform 1 0 18432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_193
timestamp 1679581782
transform 1 0 19104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_200
timestamp 1679581782
transform 1 0 19776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_207
timestamp 1679581782
transform 1 0 20448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_214
timestamp 1679581782
transform 1 0 21120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_221
timestamp 1679581782
transform 1 0 21792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_228
timestamp 1679581782
transform 1 0 22464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_235
timestamp 1679581782
transform 1 0 23136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_242
timestamp 1679581782
transform 1 0 23808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_249
timestamp 1679581782
transform 1 0 24480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_256
timestamp 1679581782
transform 1 0 25152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_263
timestamp 1679581782
transform 1 0 25824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_270
timestamp 1679581782
transform 1 0 26496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_277
timestamp 1679581782
transform 1 0 27168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_284
timestamp 1679581782
transform 1 0 27840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_291
timestamp 1679581782
transform 1 0 28512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_298
timestamp 1679581782
transform 1 0 29184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_305
timestamp 1679581782
transform 1 0 29856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_312
timestamp 1679581782
transform 1 0 30528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_319
timestamp 1679581782
transform 1 0 31200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_326
timestamp 1679581782
transform 1 0 31872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_333
timestamp 1679581782
transform 1 0 32544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_340
timestamp 1679581782
transform 1 0 33216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_347
timestamp 1679581782
transform 1 0 33888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_354
timestamp 1679581782
transform 1 0 34560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_361
timestamp 1679581782
transform 1 0 35232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_368
timestamp 1679581782
transform 1 0 35904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_375
timestamp 1679581782
transform 1 0 36576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_382
timestamp 1679581782
transform 1 0 37248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_389
timestamp 1679581782
transform 1 0 37920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_396
timestamp 1679581782
transform 1 0 38592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_403
timestamp 1679581782
transform 1 0 39264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_410
timestamp 1679581782
transform 1 0 39936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_417
timestamp 1679581782
transform 1 0 40608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_424
timestamp 1679581782
transform 1 0 41280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_431
timestamp 1679581782
transform 1 0 41952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_438
timestamp 1679581782
transform 1 0 42624 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_445
timestamp 1679581782
transform 1 0 43296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_452
timestamp 1679581782
transform 1 0 43968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_459
timestamp 1679581782
transform 1 0 44640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_466
timestamp 1679581782
transform 1 0 45312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_473
timestamp 1679581782
transform 1 0 45984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_480
timestamp 1679581782
transform 1 0 46656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_487
timestamp 1679581782
transform 1 0 47328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_494
timestamp 1679581782
transform 1 0 48000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_501
timestamp 1679581782
transform 1 0 48672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_508
timestamp 1679581782
transform 1 0 49344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_515
timestamp 1679581782
transform 1 0 50016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_522
timestamp 1679581782
transform 1 0 50688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_529
timestamp 1679581782
transform 1 0 51360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_536
timestamp 1679581782
transform 1 0 52032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_543
timestamp 1679581782
transform 1 0 52704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_550
timestamp 1679581782
transform 1 0 53376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_557
timestamp 1679581782
transform 1 0 54048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_564
timestamp 1679581782
transform 1 0 54720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_571
timestamp 1679581782
transform 1 0 55392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_578
timestamp 1679581782
transform 1 0 56064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_585
timestamp 1679581782
transform 1 0 56736 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_592
timestamp 1679581782
transform 1 0 57408 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_599
timestamp 1679581782
transform 1 0 58080 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_606
timestamp 1679581782
transform 1 0 58752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_613
timestamp 1679581782
transform 1 0 59424 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_620
timestamp 1679581782
transform 1 0 60096 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_627
timestamp 1679581782
transform 1 0 60768 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_634
timestamp 1679581782
transform 1 0 61440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_641
timestamp 1679581782
transform 1 0 62112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_648
timestamp 1679581782
transform 1 0 62784 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_655
timestamp 1679581782
transform 1 0 63456 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_662
timestamp 1679581782
transform 1 0 64128 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_669
timestamp 1679581782
transform 1 0 64800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_676
timestamp 1679581782
transform 1 0 65472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_683
timestamp 1679581782
transform 1 0 66144 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_690
timestamp 1679581782
transform 1 0 66816 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_697
timestamp 1679581782
transform 1 0 67488 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_704
timestamp 1679581782
transform 1 0 68160 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_711
timestamp 1677579658
transform 1 0 68832 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_4
timestamp 1677580104
transform 1 0 960 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_6
timestamp 1677579658
transform 1 0 1152 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_11
timestamp 1679581782
transform 1 0 1632 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_18
timestamp 1679581782
transform 1 0 2304 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_25
timestamp 1679581782
transform 1 0 2976 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_32
timestamp 1679581782
transform 1 0 3648 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_39
timestamp 1679581782
transform 1 0 4320 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_46
timestamp 1679581782
transform 1 0 4992 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_53
timestamp 1679581782
transform 1 0 5664 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_60
timestamp 1679581782
transform 1 0 6336 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_67
timestamp 1679581782
transform 1 0 7008 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_74
timestamp 1679581782
transform 1 0 7680 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_81
timestamp 1679581782
transform 1 0 8352 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_88
timestamp 1679581782
transform 1 0 9024 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_95
timestamp 1679581782
transform 1 0 9696 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_102
timestamp 1679581782
transform 1 0 10368 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_109
timestamp 1679581782
transform 1 0 11040 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_116
timestamp 1679581782
transform 1 0 11712 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_123
timestamp 1679581782
transform 1 0 12384 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_130
timestamp 1679581782
transform 1 0 13056 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_137
timestamp 1679581782
transform 1 0 13728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_144
timestamp 1679581782
transform 1 0 14400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_151
timestamp 1679581782
transform 1 0 15072 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_158
timestamp 1679581782
transform 1 0 15744 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_165
timestamp 1679581782
transform 1 0 16416 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_172
timestamp 1679581782
transform 1 0 17088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_179
timestamp 1679581782
transform 1 0 17760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_186
timestamp 1679581782
transform 1 0 18432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_193
timestamp 1679581782
transform 1 0 19104 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_200
timestamp 1679581782
transform 1 0 19776 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_207
timestamp 1679581782
transform 1 0 20448 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_214
timestamp 1679581782
transform 1 0 21120 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_221
timestamp 1679581782
transform 1 0 21792 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_228
timestamp 1679581782
transform 1 0 22464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_235
timestamp 1679581782
transform 1 0 23136 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_242
timestamp 1679581782
transform 1 0 23808 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_249
timestamp 1679581782
transform 1 0 24480 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_256
timestamp 1679581782
transform 1 0 25152 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_263
timestamp 1679581782
transform 1 0 25824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_270
timestamp 1679581782
transform 1 0 26496 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_277
timestamp 1679581782
transform 1 0 27168 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_284
timestamp 1679581782
transform 1 0 27840 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_291
timestamp 1679581782
transform 1 0 28512 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_298
timestamp 1679581782
transform 1 0 29184 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_305
timestamp 1679581782
transform 1 0 29856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_312
timestamp 1679581782
transform 1 0 30528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_319
timestamp 1679581782
transform 1 0 31200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_326
timestamp 1679581782
transform 1 0 31872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_333
timestamp 1679581782
transform 1 0 32544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_340
timestamp 1679581782
transform 1 0 33216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_347
timestamp 1679581782
transform 1 0 33888 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_354
timestamp 1679581782
transform 1 0 34560 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_361
timestamp 1679581782
transform 1 0 35232 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_368
timestamp 1679581782
transform 1 0 35904 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_375
timestamp 1679581782
transform 1 0 36576 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_382
timestamp 1679581782
transform 1 0 37248 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_389
timestamp 1679581782
transform 1 0 37920 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_396
timestamp 1679581782
transform 1 0 38592 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_403
timestamp 1679581782
transform 1 0 39264 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_410
timestamp 1679581782
transform 1 0 39936 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_417
timestamp 1679581782
transform 1 0 40608 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_424
timestamp 1679581782
transform 1 0 41280 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_431
timestamp 1679581782
transform 1 0 41952 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_438
timestamp 1679581782
transform 1 0 42624 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_445
timestamp 1679581782
transform 1 0 43296 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_452
timestamp 1679581782
transform 1 0 43968 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_459
timestamp 1679581782
transform 1 0 44640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_466
timestamp 1679581782
transform 1 0 45312 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_473
timestamp 1679581782
transform 1 0 45984 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_480
timestamp 1679581782
transform 1 0 46656 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_487
timestamp 1679581782
transform 1 0 47328 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_494
timestamp 1679581782
transform 1 0 48000 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_501
timestamp 1679581782
transform 1 0 48672 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_508
timestamp 1679581782
transform 1 0 49344 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_515
timestamp 1679581782
transform 1 0 50016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_522
timestamp 1679581782
transform 1 0 50688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_529
timestamp 1679581782
transform 1 0 51360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_536
timestamp 1679581782
transform 1 0 52032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_543
timestamp 1679581782
transform 1 0 52704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_550
timestamp 1679581782
transform 1 0 53376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_557
timestamp 1679581782
transform 1 0 54048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_564
timestamp 1679581782
transform 1 0 54720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_571
timestamp 1679581782
transform 1 0 55392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_578
timestamp 1679581782
transform 1 0 56064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_585
timestamp 1679581782
transform 1 0 56736 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_592
timestamp 1679581782
transform 1 0 57408 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_599
timestamp 1679581782
transform 1 0 58080 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_606
timestamp 1679581782
transform 1 0 58752 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_613
timestamp 1679581782
transform 1 0 59424 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_620
timestamp 1679581782
transform 1 0 60096 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_627
timestamp 1679581782
transform 1 0 60768 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_634
timestamp 1679581782
transform 1 0 61440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_641
timestamp 1679581782
transform 1 0 62112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_648
timestamp 1679581782
transform 1 0 62784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_655
timestamp 1679581782
transform 1 0 63456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_662
timestamp 1679581782
transform 1 0 64128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_669
timestamp 1679581782
transform 1 0 64800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_676
timestamp 1679581782
transform 1 0 65472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_683
timestamp 1679581782
transform 1 0 66144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_690
timestamp 1679577901
transform 1 0 66816 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_694
timestamp 1677580104
transform 1 0 67200 0 1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_12_700
timestamp 1679577901
transform 1 0 67776 0 1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_12_722
timestamp 1677579658
transform 1 0 69888 0 1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_13_4
timestamp 1679577901
transform 1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_13_12
timestamp 1679581782
transform 1 0 1728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_19
timestamp 1679581782
transform 1 0 2400 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_26
timestamp 1679581782
transform 1 0 3072 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_33
timestamp 1679581782
transform 1 0 3744 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_40
timestamp 1679581782
transform 1 0 4416 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_47
timestamp 1679581782
transform 1 0 5088 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_54
timestamp 1679581782
transform 1 0 5760 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_61
timestamp 1679581782
transform 1 0 6432 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_68
timestamp 1679581782
transform 1 0 7104 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_75
timestamp 1679581782
transform 1 0 7776 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_82
timestamp 1679581782
transform 1 0 8448 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_89
timestamp 1679581782
transform 1 0 9120 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_96
timestamp 1679581782
transform 1 0 9792 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_103
timestamp 1679581782
transform 1 0 10464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_110
timestamp 1679581782
transform 1 0 11136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_117
timestamp 1679581782
transform 1 0 11808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_124
timestamp 1679581782
transform 1 0 12480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_131
timestamp 1679581782
transform 1 0 13152 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_138
timestamp 1679581782
transform 1 0 13824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_145
timestamp 1679581782
transform 1 0 14496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_152
timestamp 1679581782
transform 1 0 15168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_159
timestamp 1679581782
transform 1 0 15840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_166
timestamp 1679581782
transform 1 0 16512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_173
timestamp 1679581782
transform 1 0 17184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_180
timestamp 1679581782
transform 1 0 17856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_187
timestamp 1679581782
transform 1 0 18528 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_194
timestamp 1679581782
transform 1 0 19200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_201
timestamp 1679581782
transform 1 0 19872 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_208
timestamp 1679581782
transform 1 0 20544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_215
timestamp 1679581782
transform 1 0 21216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_222
timestamp 1679581782
transform 1 0 21888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_229
timestamp 1679581782
transform 1 0 22560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_236
timestamp 1679581782
transform 1 0 23232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_243
timestamp 1679581782
transform 1 0 23904 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_250
timestamp 1679581782
transform 1 0 24576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_257
timestamp 1679581782
transform 1 0 25248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_264
timestamp 1679581782
transform 1 0 25920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_271
timestamp 1679581782
transform 1 0 26592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_278
timestamp 1679581782
transform 1 0 27264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_285
timestamp 1679581782
transform 1 0 27936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_292
timestamp 1679581782
transform 1 0 28608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_299
timestamp 1679581782
transform 1 0 29280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_306
timestamp 1679581782
transform 1 0 29952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_313
timestamp 1679581782
transform 1 0 30624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_320
timestamp 1679581782
transform 1 0 31296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_327
timestamp 1679581782
transform 1 0 31968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_334
timestamp 1679581782
transform 1 0 32640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_341
timestamp 1679581782
transform 1 0 33312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_348
timestamp 1679581782
transform 1 0 33984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_355
timestamp 1679581782
transform 1 0 34656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_362
timestamp 1679581782
transform 1 0 35328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_369
timestamp 1679581782
transform 1 0 36000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_376
timestamp 1679581782
transform 1 0 36672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_383
timestamp 1679581782
transform 1 0 37344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_390
timestamp 1679581782
transform 1 0 38016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_397
timestamp 1679581782
transform 1 0 38688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_404
timestamp 1679581782
transform 1 0 39360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_411
timestamp 1679581782
transform 1 0 40032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_418
timestamp 1679581782
transform 1 0 40704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_425
timestamp 1679581782
transform 1 0 41376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_432
timestamp 1679581782
transform 1 0 42048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_439
timestamp 1679581782
transform 1 0 42720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_446
timestamp 1679581782
transform 1 0 43392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_453
timestamp 1679581782
transform 1 0 44064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_460
timestamp 1679581782
transform 1 0 44736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_467
timestamp 1679581782
transform 1 0 45408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_474
timestamp 1679581782
transform 1 0 46080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_481
timestamp 1679581782
transform 1 0 46752 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_488
timestamp 1679581782
transform 1 0 47424 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_495
timestamp 1679581782
transform 1 0 48096 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_502
timestamp 1679581782
transform 1 0 48768 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_509
timestamp 1679581782
transform 1 0 49440 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_516
timestamp 1679581782
transform 1 0 50112 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_523
timestamp 1679581782
transform 1 0 50784 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_530
timestamp 1679581782
transform 1 0 51456 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_537
timestamp 1679581782
transform 1 0 52128 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_544
timestamp 1679581782
transform 1 0 52800 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_551
timestamp 1679581782
transform 1 0 53472 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_558
timestamp 1679581782
transform 1 0 54144 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_565
timestamp 1679581782
transform 1 0 54816 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_572
timestamp 1679581782
transform 1 0 55488 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_579
timestamp 1679581782
transform 1 0 56160 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_586
timestamp 1679581782
transform 1 0 56832 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_593
timestamp 1679581782
transform 1 0 57504 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_600
timestamp 1679581782
transform 1 0 58176 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_607
timestamp 1679581782
transform 1 0 58848 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_614
timestamp 1679581782
transform 1 0 59520 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_621
timestamp 1679581782
transform 1 0 60192 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_628
timestamp 1679581782
transform 1 0 60864 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_635
timestamp 1679581782
transform 1 0 61536 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_642
timestamp 1679581782
transform 1 0 62208 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_649
timestamp 1679581782
transform 1 0 62880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_656
timestamp 1679581782
transform 1 0 63552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_663
timestamp 1679581782
transform 1 0 64224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_670
timestamp 1679581782
transform 1 0 64896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_677
timestamp 1679581782
transform 1 0 65568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_684
timestamp 1679581782
transform 1 0 66240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_691
timestamp 1679581782
transform 1 0 66912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_698
timestamp 1679581782
transform 1 0 67584 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_705
timestamp 1679581782
transform 1 0 68256 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_712
timestamp 1677580104
transform 1 0 68928 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_714
timestamp 1677579658
transform 1 0 69120 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_719
timestamp 1677579658
transform 1 0 69600 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679581782
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_11
timestamp 1677580104
transform 1 0 1632 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_13
timestamp 1677579658
transform 1 0 1824 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_18
timestamp 1679581782
transform 1 0 2304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_25
timestamp 1679581782
transform 1 0 2976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_32
timestamp 1679581782
transform 1 0 3648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_39
timestamp 1679581782
transform 1 0 4320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_46
timestamp 1679581782
transform 1 0 4992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_53
timestamp 1679581782
transform 1 0 5664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_60
timestamp 1679581782
transform 1 0 6336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_67
timestamp 1679581782
transform 1 0 7008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_74
timestamp 1679581782
transform 1 0 7680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_81
timestamp 1679581782
transform 1 0 8352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_88
timestamp 1679581782
transform 1 0 9024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_95
timestamp 1679581782
transform 1 0 9696 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_102
timestamp 1679581782
transform 1 0 10368 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_109
timestamp 1679581782
transform 1 0 11040 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_116
timestamp 1679581782
transform 1 0 11712 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_123
timestamp 1679581782
transform 1 0 12384 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_130
timestamp 1679581782
transform 1 0 13056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_137
timestamp 1679581782
transform 1 0 13728 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_144
timestamp 1679581782
transform 1 0 14400 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_151
timestamp 1679581782
transform 1 0 15072 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_158
timestamp 1679581782
transform 1 0 15744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_165
timestamp 1679581782
transform 1 0 16416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_172
timestamp 1679581782
transform 1 0 17088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_179
timestamp 1679581782
transform 1 0 17760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_186
timestamp 1679581782
transform 1 0 18432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_193
timestamp 1679581782
transform 1 0 19104 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_200
timestamp 1679581782
transform 1 0 19776 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_207
timestamp 1679581782
transform 1 0 20448 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_214
timestamp 1679581782
transform 1 0 21120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_221
timestamp 1679581782
transform 1 0 21792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_228
timestamp 1679581782
transform 1 0 22464 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_235
timestamp 1679581782
transform 1 0 23136 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_242
timestamp 1679581782
transform 1 0 23808 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_249
timestamp 1679581782
transform 1 0 24480 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_256
timestamp 1679581782
transform 1 0 25152 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_263
timestamp 1679581782
transform 1 0 25824 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_270
timestamp 1679581782
transform 1 0 26496 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_277
timestamp 1679581782
transform 1 0 27168 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_284
timestamp 1679581782
transform 1 0 27840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_291
timestamp 1679581782
transform 1 0 28512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_298
timestamp 1679581782
transform 1 0 29184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_305
timestamp 1679581782
transform 1 0 29856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_312
timestamp 1679581782
transform 1 0 30528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_319
timestamp 1679581782
transform 1 0 31200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_326
timestamp 1679581782
transform 1 0 31872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_333
timestamp 1679581782
transform 1 0 32544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_340
timestamp 1679581782
transform 1 0 33216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_347
timestamp 1679581782
transform 1 0 33888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_354
timestamp 1679581782
transform 1 0 34560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_361
timestamp 1679581782
transform 1 0 35232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_368
timestamp 1679581782
transform 1 0 35904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_375
timestamp 1679581782
transform 1 0 36576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_382
timestamp 1679581782
transform 1 0 37248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_389
timestamp 1679581782
transform 1 0 37920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_396
timestamp 1679581782
transform 1 0 38592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_403
timestamp 1679581782
transform 1 0 39264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_410
timestamp 1679581782
transform 1 0 39936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_417
timestamp 1679581782
transform 1 0 40608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_424
timestamp 1679581782
transform 1 0 41280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_431
timestamp 1679581782
transform 1 0 41952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_438
timestamp 1679581782
transform 1 0 42624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_445
timestamp 1679581782
transform 1 0 43296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_452
timestamp 1679581782
transform 1 0 43968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_459
timestamp 1679581782
transform 1 0 44640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_466
timestamp 1679581782
transform 1 0 45312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_473
timestamp 1679581782
transform 1 0 45984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_480
timestamp 1679581782
transform 1 0 46656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_487
timestamp 1679581782
transform 1 0 47328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_494
timestamp 1679581782
transform 1 0 48000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_501
timestamp 1679581782
transform 1 0 48672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_508
timestamp 1679581782
transform 1 0 49344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_515
timestamp 1679581782
transform 1 0 50016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_522
timestamp 1679581782
transform 1 0 50688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_529
timestamp 1679581782
transform 1 0 51360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_536
timestamp 1679581782
transform 1 0 52032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_543
timestamp 1679581782
transform 1 0 52704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_550
timestamp 1679581782
transform 1 0 53376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_557
timestamp 1679581782
transform 1 0 54048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_564
timestamp 1679581782
transform 1 0 54720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_571
timestamp 1679581782
transform 1 0 55392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_578
timestamp 1679581782
transform 1 0 56064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_585
timestamp 1679581782
transform 1 0 56736 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_592
timestamp 1679581782
transform 1 0 57408 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_599
timestamp 1679581782
transform 1 0 58080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_606
timestamp 1679581782
transform 1 0 58752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_613
timestamp 1679581782
transform 1 0 59424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_620
timestamp 1679581782
transform 1 0 60096 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_627
timestamp 1679581782
transform 1 0 60768 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_634
timestamp 1679581782
transform 1 0 61440 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_641
timestamp 1679581782
transform 1 0 62112 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_648
timestamp 1679581782
transform 1 0 62784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_655
timestamp 1679581782
transform 1 0 63456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_662
timestamp 1679581782
transform 1 0 64128 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_669
timestamp 1679581782
transform 1 0 64800 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_676
timestamp 1679581782
transform 1 0 65472 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_683
timestamp 1679581782
transform 1 0 66144 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_690
timestamp 1679581782
transform 1 0 66816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_697
timestamp 1679581782
transform 1 0 67488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_704
timestamp 1679581782
transform 1 0 68160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_711
timestamp 1679581782
transform 1 0 68832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_14_718
timestamp 1679577901
transform 1 0 69504 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_722
timestamp 1677579658
transform 1 0 69888 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_4
timestamp 1679577901
transform 1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_8
timestamp 1677580104
transform 1 0 1344 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_14
timestamp 1679581782
transform 1 0 1920 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_21
timestamp 1679581782
transform 1 0 2592 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_28
timestamp 1679581782
transform 1 0 3264 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_35
timestamp 1679581782
transform 1 0 3936 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_42
timestamp 1679581782
transform 1 0 4608 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_49
timestamp 1679581782
transform 1 0 5280 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_56
timestamp 1679581782
transform 1 0 5952 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_63
timestamp 1679581782
transform 1 0 6624 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_70
timestamp 1679581782
transform 1 0 7296 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_77
timestamp 1679581782
transform 1 0 7968 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_84
timestamp 1679581782
transform 1 0 8640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_91
timestamp 1679581782
transform 1 0 9312 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_98
timestamp 1679581782
transform 1 0 9984 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_105
timestamp 1679581782
transform 1 0 10656 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_112
timestamp 1679581782
transform 1 0 11328 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_119
timestamp 1679581782
transform 1 0 12000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_126
timestamp 1679581782
transform 1 0 12672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_133
timestamp 1679581782
transform 1 0 13344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_140
timestamp 1679581782
transform 1 0 14016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_147
timestamp 1679581782
transform 1 0 14688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_154
timestamp 1679581782
transform 1 0 15360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_161
timestamp 1679581782
transform 1 0 16032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_168
timestamp 1679581782
transform 1 0 16704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_175
timestamp 1679581782
transform 1 0 17376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_182
timestamp 1679581782
transform 1 0 18048 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_189
timestamp 1679581782
transform 1 0 18720 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_196
timestamp 1679581782
transform 1 0 19392 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_203
timestamp 1679581782
transform 1 0 20064 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_210
timestamp 1679581782
transform 1 0 20736 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_217
timestamp 1679581782
transform 1 0 21408 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_224
timestamp 1679581782
transform 1 0 22080 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_231
timestamp 1679581782
transform 1 0 22752 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_238
timestamp 1679581782
transform 1 0 23424 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_245
timestamp 1679581782
transform 1 0 24096 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_252
timestamp 1679581782
transform 1 0 24768 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_259
timestamp 1679581782
transform 1 0 25440 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_266
timestamp 1679581782
transform 1 0 26112 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_273
timestamp 1679581782
transform 1 0 26784 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_280
timestamp 1679581782
transform 1 0 27456 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_287
timestamp 1679581782
transform 1 0 28128 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_294
timestamp 1679581782
transform 1 0 28800 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_301
timestamp 1679581782
transform 1 0 29472 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_308
timestamp 1679581782
transform 1 0 30144 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_315
timestamp 1679581782
transform 1 0 30816 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_322
timestamp 1679581782
transform 1 0 31488 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_329
timestamp 1679581782
transform 1 0 32160 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_336
timestamp 1679581782
transform 1 0 32832 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_343
timestamp 1679581782
transform 1 0 33504 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_350
timestamp 1679581782
transform 1 0 34176 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_357
timestamp 1679581782
transform 1 0 34848 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_364
timestamp 1679581782
transform 1 0 35520 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_371
timestamp 1679581782
transform 1 0 36192 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_378
timestamp 1679581782
transform 1 0 36864 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_385
timestamp 1679581782
transform 1 0 37536 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_392
timestamp 1679581782
transform 1 0 38208 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_399
timestamp 1679581782
transform 1 0 38880 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_406
timestamp 1679581782
transform 1 0 39552 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_413
timestamp 1679581782
transform 1 0 40224 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_420
timestamp 1679581782
transform 1 0 40896 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_427
timestamp 1679581782
transform 1 0 41568 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_434
timestamp 1679581782
transform 1 0 42240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_441
timestamp 1679581782
transform 1 0 42912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_448
timestamp 1679581782
transform 1 0 43584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_455
timestamp 1679581782
transform 1 0 44256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_462
timestamp 1679581782
transform 1 0 44928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_469
timestamp 1679581782
transform 1 0 45600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_476
timestamp 1679581782
transform 1 0 46272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_483
timestamp 1679581782
transform 1 0 46944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_490
timestamp 1679581782
transform 1 0 47616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_497
timestamp 1679581782
transform 1 0 48288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_504
timestamp 1679581782
transform 1 0 48960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_511
timestamp 1679581782
transform 1 0 49632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_518
timestamp 1679581782
transform 1 0 50304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_525
timestamp 1679581782
transform 1 0 50976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_532
timestamp 1679581782
transform 1 0 51648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_539
timestamp 1679581782
transform 1 0 52320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_546
timestamp 1679581782
transform 1 0 52992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_553
timestamp 1679581782
transform 1 0 53664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_560
timestamp 1679581782
transform 1 0 54336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_567
timestamp 1679581782
transform 1 0 55008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_574
timestamp 1679581782
transform 1 0 55680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_581
timestamp 1679581782
transform 1 0 56352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_588
timestamp 1679581782
transform 1 0 57024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_595
timestamp 1679581782
transform 1 0 57696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_602
timestamp 1679581782
transform 1 0 58368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_609
timestamp 1679581782
transform 1 0 59040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_616
timestamp 1679581782
transform 1 0 59712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_623
timestamp 1679581782
transform 1 0 60384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_630
timestamp 1679581782
transform 1 0 61056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_637
timestamp 1679581782
transform 1 0 61728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_644
timestamp 1679581782
transform 1 0 62400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_651
timestamp 1679581782
transform 1 0 63072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_658
timestamp 1679581782
transform 1 0 63744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_665
timestamp 1679581782
transform 1 0 64416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_672
timestamp 1679581782
transform 1 0 65088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_679
timestamp 1679581782
transform 1 0 65760 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_686
timestamp 1679581782
transform 1 0 66432 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_693
timestamp 1679581782
transform 1 0 67104 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_700
timestamp 1679581782
transform 1 0 67776 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_707
timestamp 1679581782
transform 1 0 68448 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_714
timestamp 1679581782
transform 1 0 69120 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_721
timestamp 1677580104
transform 1 0 69792 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_4
timestamp 1679581782
transform 1 0 960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_15
timestamp 1679581782
transform 1 0 2016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_22
timestamp 1679581782
transform 1 0 2688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_29
timestamp 1679581782
transform 1 0 3360 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_36
timestamp 1679581782
transform 1 0 4032 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_43
timestamp 1679581782
transform 1 0 4704 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_50
timestamp 1679581782
transform 1 0 5376 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_57
timestamp 1679581782
transform 1 0 6048 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_64
timestamp 1679581782
transform 1 0 6720 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_71
timestamp 1679581782
transform 1 0 7392 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_78
timestamp 1679581782
transform 1 0 8064 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_85
timestamp 1679581782
transform 1 0 8736 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_92
timestamp 1679581782
transform 1 0 9408 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_99
timestamp 1679581782
transform 1 0 10080 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_106
timestamp 1679581782
transform 1 0 10752 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_113
timestamp 1679581782
transform 1 0 11424 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_120
timestamp 1679581782
transform 1 0 12096 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_127
timestamp 1679581782
transform 1 0 12768 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_134
timestamp 1679581782
transform 1 0 13440 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_141
timestamp 1679581782
transform 1 0 14112 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_148
timestamp 1679581782
transform 1 0 14784 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_155
timestamp 1679581782
transform 1 0 15456 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_162
timestamp 1679581782
transform 1 0 16128 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_169
timestamp 1679581782
transform 1 0 16800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_176
timestamp 1679581782
transform 1 0 17472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_183
timestamp 1679581782
transform 1 0 18144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_190
timestamp 1679581782
transform 1 0 18816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_197
timestamp 1679581782
transform 1 0 19488 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_204
timestamp 1679581782
transform 1 0 20160 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_211
timestamp 1679581782
transform 1 0 20832 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_218
timestamp 1679581782
transform 1 0 21504 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_225
timestamp 1679581782
transform 1 0 22176 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_232
timestamp 1679581782
transform 1 0 22848 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_239
timestamp 1679581782
transform 1 0 23520 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_246
timestamp 1679581782
transform 1 0 24192 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_253
timestamp 1679581782
transform 1 0 24864 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_260
timestamp 1679581782
transform 1 0 25536 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_267
timestamp 1679581782
transform 1 0 26208 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_274
timestamp 1679581782
transform 1 0 26880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_281
timestamp 1679581782
transform 1 0 27552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_288
timestamp 1679581782
transform 1 0 28224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_295
timestamp 1679581782
transform 1 0 28896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_302
timestamp 1679581782
transform 1 0 29568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_309
timestamp 1679581782
transform 1 0 30240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_316
timestamp 1679581782
transform 1 0 30912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_323
timestamp 1679581782
transform 1 0 31584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_330
timestamp 1679581782
transform 1 0 32256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_337
timestamp 1679581782
transform 1 0 32928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_344
timestamp 1679581782
transform 1 0 33600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_351
timestamp 1679581782
transform 1 0 34272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_358
timestamp 1679581782
transform 1 0 34944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_365
timestamp 1679581782
transform 1 0 35616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_372
timestamp 1679581782
transform 1 0 36288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_379
timestamp 1679581782
transform 1 0 36960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_386
timestamp 1679581782
transform 1 0 37632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_393
timestamp 1679581782
transform 1 0 38304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_400
timestamp 1679581782
transform 1 0 38976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_407
timestamp 1679581782
transform 1 0 39648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_414
timestamp 1679581782
transform 1 0 40320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_421
timestamp 1679581782
transform 1 0 40992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_428
timestamp 1679581782
transform 1 0 41664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_435
timestamp 1679581782
transform 1 0 42336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_442
timestamp 1679581782
transform 1 0 43008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_449
timestamp 1679581782
transform 1 0 43680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_456
timestamp 1679581782
transform 1 0 44352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_463
timestamp 1679581782
transform 1 0 45024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_470
timestamp 1679581782
transform 1 0 45696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_477
timestamp 1679581782
transform 1 0 46368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_484
timestamp 1679581782
transform 1 0 47040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_491
timestamp 1679581782
transform 1 0 47712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_498
timestamp 1679581782
transform 1 0 48384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_505
timestamp 1679581782
transform 1 0 49056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_512
timestamp 1679581782
transform 1 0 49728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_519
timestamp 1679581782
transform 1 0 50400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_526
timestamp 1679581782
transform 1 0 51072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_533
timestamp 1679581782
transform 1 0 51744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_540
timestamp 1679581782
transform 1 0 52416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_547
timestamp 1679581782
transform 1 0 53088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_554
timestamp 1679581782
transform 1 0 53760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_561
timestamp 1679581782
transform 1 0 54432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_568
timestamp 1679581782
transform 1 0 55104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_575
timestamp 1679581782
transform 1 0 55776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_582
timestamp 1679581782
transform 1 0 56448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_589
timestamp 1679581782
transform 1 0 57120 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_596
timestamp 1679581782
transform 1 0 57792 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_603
timestamp 1679581782
transform 1 0 58464 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_610
timestamp 1679581782
transform 1 0 59136 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_617
timestamp 1679581782
transform 1 0 59808 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_624
timestamp 1679581782
transform 1 0 60480 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_631
timestamp 1679581782
transform 1 0 61152 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_638
timestamp 1679581782
transform 1 0 61824 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_645
timestamp 1679581782
transform 1 0 62496 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_652
timestamp 1679581782
transform 1 0 63168 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_659
timestamp 1679581782
transform 1 0 63840 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_666
timestamp 1679581782
transform 1 0 64512 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_673
timestamp 1679581782
transform 1 0 65184 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_680
timestamp 1679581782
transform 1 0 65856 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_687
timestamp 1679581782
transform 1 0 66528 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_694
timestamp 1679581782
transform 1 0 67200 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_701
timestamp 1679581782
transform 1 0 67872 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_708
timestamp 1679581782
transform 1 0 68544 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_715
timestamp 1679581782
transform 1 0 69216 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_722
timestamp 1677579658
transform 1 0 69888 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679581782
transform 1 0 576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_11
timestamp 1679581782
transform 1 0 1632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_18
timestamp 1679581782
transform 1 0 2304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_25
timestamp 1679581782
transform 1 0 2976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_32
timestamp 1679581782
transform 1 0 3648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_39
timestamp 1679581782
transform 1 0 4320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_46
timestamp 1679581782
transform 1 0 4992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_53
timestamp 1679581782
transform 1 0 5664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_60
timestamp 1679581782
transform 1 0 6336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_67
timestamp 1679581782
transform 1 0 7008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_74
timestamp 1679581782
transform 1 0 7680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_81
timestamp 1679581782
transform 1 0 8352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_88
timestamp 1679581782
transform 1 0 9024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_95
timestamp 1679581782
transform 1 0 9696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_102
timestamp 1679581782
transform 1 0 10368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_109
timestamp 1679581782
transform 1 0 11040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_116
timestamp 1679581782
transform 1 0 11712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_123
timestamp 1679581782
transform 1 0 12384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_130
timestamp 1679581782
transform 1 0 13056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_137
timestamp 1679581782
transform 1 0 13728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_144
timestamp 1679581782
transform 1 0 14400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_151
timestamp 1679581782
transform 1 0 15072 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_158
timestamp 1679581782
transform 1 0 15744 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_165
timestamp 1679581782
transform 1 0 16416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_172
timestamp 1679581782
transform 1 0 17088 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_179
timestamp 1679581782
transform 1 0 17760 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_186
timestamp 1679581782
transform 1 0 18432 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_193
timestamp 1679581782
transform 1 0 19104 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_200
timestamp 1679581782
transform 1 0 19776 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_207
timestamp 1679581782
transform 1 0 20448 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_214
timestamp 1679581782
transform 1 0 21120 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_221
timestamp 1679581782
transform 1 0 21792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_228
timestamp 1679581782
transform 1 0 22464 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_235
timestamp 1679581782
transform 1 0 23136 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_242
timestamp 1679581782
transform 1 0 23808 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_249
timestamp 1679581782
transform 1 0 24480 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_256
timestamp 1679581782
transform 1 0 25152 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_263
timestamp 1679581782
transform 1 0 25824 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_270
timestamp 1679581782
transform 1 0 26496 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_277
timestamp 1679581782
transform 1 0 27168 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_284
timestamp 1679581782
transform 1 0 27840 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_291
timestamp 1679581782
transform 1 0 28512 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_298
timestamp 1679581782
transform 1 0 29184 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_305
timestamp 1679581782
transform 1 0 29856 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_312
timestamp 1679581782
transform 1 0 30528 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_319
timestamp 1679581782
transform 1 0 31200 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_326
timestamp 1679581782
transform 1 0 31872 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_333
timestamp 1679581782
transform 1 0 32544 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_340
timestamp 1679581782
transform 1 0 33216 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_347
timestamp 1679581782
transform 1 0 33888 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_354
timestamp 1679581782
transform 1 0 34560 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_361
timestamp 1679581782
transform 1 0 35232 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_368
timestamp 1679581782
transform 1 0 35904 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_375
timestamp 1679581782
transform 1 0 36576 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_382
timestamp 1679581782
transform 1 0 37248 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_389
timestamp 1679581782
transform 1 0 37920 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_396
timestamp 1679581782
transform 1 0 38592 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_403
timestamp 1679581782
transform 1 0 39264 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_410
timestamp 1679581782
transform 1 0 39936 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_417
timestamp 1679581782
transform 1 0 40608 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_424
timestamp 1679581782
transform 1 0 41280 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_431
timestamp 1679581782
transform 1 0 41952 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_438
timestamp 1679581782
transform 1 0 42624 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_445
timestamp 1679581782
transform 1 0 43296 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_452
timestamp 1679581782
transform 1 0 43968 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_459
timestamp 1679581782
transform 1 0 44640 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_466
timestamp 1679581782
transform 1 0 45312 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_473
timestamp 1679581782
transform 1 0 45984 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_480
timestamp 1679581782
transform 1 0 46656 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_487
timestamp 1679581782
transform 1 0 47328 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_494
timestamp 1679581782
transform 1 0 48000 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_501
timestamp 1679581782
transform 1 0 48672 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_508
timestamp 1679581782
transform 1 0 49344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_515
timestamp 1679581782
transform 1 0 50016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_522
timestamp 1679581782
transform 1 0 50688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_529
timestamp 1679581782
transform 1 0 51360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_536
timestamp 1679581782
transform 1 0 52032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_543
timestamp 1679581782
transform 1 0 52704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_550
timestamp 1679581782
transform 1 0 53376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_557
timestamp 1679581782
transform 1 0 54048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_564
timestamp 1679581782
transform 1 0 54720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_571
timestamp 1679581782
transform 1 0 55392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_578
timestamp 1679581782
transform 1 0 56064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_585
timestamp 1679581782
transform 1 0 56736 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_592
timestamp 1679581782
transform 1 0 57408 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_599
timestamp 1679581782
transform 1 0 58080 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_606
timestamp 1679581782
transform 1 0 58752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_613
timestamp 1679581782
transform 1 0 59424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_620
timestamp 1679581782
transform 1 0 60096 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_627
timestamp 1679581782
transform 1 0 60768 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_634
timestamp 1679581782
transform 1 0 61440 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_641
timestamp 1679581782
transform 1 0 62112 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_648
timestamp 1679581782
transform 1 0 62784 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_655
timestamp 1679581782
transform 1 0 63456 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_662
timestamp 1679581782
transform 1 0 64128 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_669
timestamp 1679581782
transform 1 0 64800 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_676
timestamp 1679581782
transform 1 0 65472 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_683
timestamp 1679581782
transform 1 0 66144 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_690
timestamp 1679581782
transform 1 0 66816 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_697
timestamp 1679581782
transform 1 0 67488 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_704
timestamp 1679581782
transform 1 0 68160 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_711
timestamp 1677580104
transform 1 0 68832 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_713
timestamp 1677579658
transform 1 0 69024 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_17_718
timestamp 1677580104
transform 1 0 69504 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_4
timestamp 1679581782
transform 1 0 960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_15
timestamp 1679581782
transform 1 0 2016 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_22
timestamp 1679581782
transform 1 0 2688 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_29
timestamp 1679581782
transform 1 0 3360 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_36
timestamp 1679581782
transform 1 0 4032 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_43
timestamp 1679581782
transform 1 0 4704 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_50
timestamp 1679581782
transform 1 0 5376 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_57
timestamp 1679581782
transform 1 0 6048 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_64
timestamp 1679581782
transform 1 0 6720 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_71
timestamp 1679581782
transform 1 0 7392 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_78
timestamp 1679581782
transform 1 0 8064 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_85
timestamp 1679581782
transform 1 0 8736 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_92
timestamp 1679581782
transform 1 0 9408 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_99
timestamp 1679581782
transform 1 0 10080 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_106
timestamp 1679581782
transform 1 0 10752 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_113
timestamp 1679581782
transform 1 0 11424 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_120
timestamp 1679581782
transform 1 0 12096 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_127
timestamp 1679581782
transform 1 0 12768 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_134
timestamp 1679581782
transform 1 0 13440 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_141
timestamp 1679581782
transform 1 0 14112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_148
timestamp 1679581782
transform 1 0 14784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_155
timestamp 1679581782
transform 1 0 15456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_162
timestamp 1679581782
transform 1 0 16128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_169
timestamp 1679581782
transform 1 0 16800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_176
timestamp 1679581782
transform 1 0 17472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_183
timestamp 1679581782
transform 1 0 18144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_190
timestamp 1679581782
transform 1 0 18816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_197
timestamp 1679581782
transform 1 0 19488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_204
timestamp 1679581782
transform 1 0 20160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_211
timestamp 1679581782
transform 1 0 20832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_218
timestamp 1679581782
transform 1 0 21504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_225
timestamp 1679581782
transform 1 0 22176 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_232
timestamp 1679581782
transform 1 0 22848 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_239
timestamp 1679581782
transform 1 0 23520 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_246
timestamp 1679581782
transform 1 0 24192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_253
timestamp 1679581782
transform 1 0 24864 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_260
timestamp 1679581782
transform 1 0 25536 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_267
timestamp 1679581782
transform 1 0 26208 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_274
timestamp 1679581782
transform 1 0 26880 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_281
timestamp 1679581782
transform 1 0 27552 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_288
timestamp 1679581782
transform 1 0 28224 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_295
timestamp 1679581782
transform 1 0 28896 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_302
timestamp 1679581782
transform 1 0 29568 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_309
timestamp 1679581782
transform 1 0 30240 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_316
timestamp 1679581782
transform 1 0 30912 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_323
timestamp 1679581782
transform 1 0 31584 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_330
timestamp 1679581782
transform 1 0 32256 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_337
timestamp 1679581782
transform 1 0 32928 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_344
timestamp 1679581782
transform 1 0 33600 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_351
timestamp 1679581782
transform 1 0 34272 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_358
timestamp 1679581782
transform 1 0 34944 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_365
timestamp 1679581782
transform 1 0 35616 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_372
timestamp 1679581782
transform 1 0 36288 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_379
timestamp 1679581782
transform 1 0 36960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_386
timestamp 1679581782
transform 1 0 37632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_393
timestamp 1679581782
transform 1 0 38304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_400
timestamp 1679581782
transform 1 0 38976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_407
timestamp 1679581782
transform 1 0 39648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_414
timestamp 1679581782
transform 1 0 40320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_421
timestamp 1679581782
transform 1 0 40992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_428
timestamp 1679581782
transform 1 0 41664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_435
timestamp 1679581782
transform 1 0 42336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_442
timestamp 1679581782
transform 1 0 43008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_449
timestamp 1679581782
transform 1 0 43680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_456
timestamp 1679581782
transform 1 0 44352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_463
timestamp 1679581782
transform 1 0 45024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_470
timestamp 1679581782
transform 1 0 45696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_477
timestamp 1679581782
transform 1 0 46368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_484
timestamp 1679581782
transform 1 0 47040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_491
timestamp 1679581782
transform 1 0 47712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_498
timestamp 1679581782
transform 1 0 48384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_505
timestamp 1679581782
transform 1 0 49056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_512
timestamp 1679581782
transform 1 0 49728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_519
timestamp 1679581782
transform 1 0 50400 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_526
timestamp 1679581782
transform 1 0 51072 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_533
timestamp 1679581782
transform 1 0 51744 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_540
timestamp 1679581782
transform 1 0 52416 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_547
timestamp 1679581782
transform 1 0 53088 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_554
timestamp 1679581782
transform 1 0 53760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_561
timestamp 1679581782
transform 1 0 54432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_568
timestamp 1679581782
transform 1 0 55104 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_575
timestamp 1679581782
transform 1 0 55776 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_582
timestamp 1679581782
transform 1 0 56448 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_589
timestamp 1679581782
transform 1 0 57120 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_596
timestamp 1679581782
transform 1 0 57792 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_603
timestamp 1679581782
transform 1 0 58464 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_610
timestamp 1679581782
transform 1 0 59136 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_617
timestamp 1679581782
transform 1 0 59808 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_624
timestamp 1679581782
transform 1 0 60480 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_631
timestamp 1679581782
transform 1 0 61152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_638
timestamp 1679581782
transform 1 0 61824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_645
timestamp 1679581782
transform 1 0 62496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_652
timestamp 1679581782
transform 1 0 63168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_659
timestamp 1679581782
transform 1 0 63840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_666
timestamp 1679581782
transform 1 0 64512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_673
timestamp 1679581782
transform 1 0 65184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_680
timestamp 1679581782
transform 1 0 65856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_687
timestamp 1679581782
transform 1 0 66528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_694
timestamp 1679581782
transform 1 0 67200 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_701
timestamp 1677579658
transform 1 0 67872 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_705
timestamp 1677580104
transform 1 0 68256 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_707
timestamp 1677579658
transform 1 0 68448 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_711
timestamp 1677579658
transform 1 0 68832 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_715
timestamp 1677579658
transform 1 0 69216 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_4
timestamp 1679581782
transform 1 0 960 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_11
timestamp 1677579658
transform 1 0 1632 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_16
timestamp 1679581782
transform 1 0 2112 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_23
timestamp 1679581782
transform 1 0 2784 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_30
timestamp 1679581782
transform 1 0 3456 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_37
timestamp 1679581782
transform 1 0 4128 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_44
timestamp 1679581782
transform 1 0 4800 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_51
timestamp 1679581782
transform 1 0 5472 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_58
timestamp 1679581782
transform 1 0 6144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_65
timestamp 1679581782
transform 1 0 6816 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_72
timestamp 1679581782
transform 1 0 7488 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_79
timestamp 1679581782
transform 1 0 8160 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_86
timestamp 1679581782
transform 1 0 8832 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_93
timestamp 1679581782
transform 1 0 9504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_100
timestamp 1679581782
transform 1 0 10176 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_107
timestamp 1679581782
transform 1 0 10848 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_114
timestamp 1679581782
transform 1 0 11520 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_121
timestamp 1679581782
transform 1 0 12192 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_128
timestamp 1679581782
transform 1 0 12864 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_135
timestamp 1679581782
transform 1 0 13536 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_142
timestamp 1679581782
transform 1 0 14208 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_149
timestamp 1679581782
transform 1 0 14880 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_156
timestamp 1679581782
transform 1 0 15552 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_163
timestamp 1679581782
transform 1 0 16224 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_170
timestamp 1679581782
transform 1 0 16896 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_177
timestamp 1679581782
transform 1 0 17568 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_184
timestamp 1679581782
transform 1 0 18240 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_191
timestamp 1679581782
transform 1 0 18912 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_198
timestamp 1679581782
transform 1 0 19584 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_205
timestamp 1679581782
transform 1 0 20256 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_212
timestamp 1679581782
transform 1 0 20928 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_219
timestamp 1679581782
transform 1 0 21600 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_226
timestamp 1679581782
transform 1 0 22272 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_233
timestamp 1679581782
transform 1 0 22944 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_240
timestamp 1679581782
transform 1 0 23616 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_247
timestamp 1679581782
transform 1 0 24288 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_254
timestamp 1679581782
transform 1 0 24960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_261
timestamp 1679581782
transform 1 0 25632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_268
timestamp 1679581782
transform 1 0 26304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_275
timestamp 1679581782
transform 1 0 26976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_282
timestamp 1679581782
transform 1 0 27648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_289
timestamp 1679581782
transform 1 0 28320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_296
timestamp 1679581782
transform 1 0 28992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_303
timestamp 1679581782
transform 1 0 29664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_310
timestamp 1679581782
transform 1 0 30336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_317
timestamp 1679581782
transform 1 0 31008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_324
timestamp 1679581782
transform 1 0 31680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_331
timestamp 1679581782
transform 1 0 32352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_338
timestamp 1679581782
transform 1 0 33024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_345
timestamp 1679581782
transform 1 0 33696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_352
timestamp 1679581782
transform 1 0 34368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_359
timestamp 1679581782
transform 1 0 35040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_366
timestamp 1679581782
transform 1 0 35712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_373
timestamp 1679581782
transform 1 0 36384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_380
timestamp 1679581782
transform 1 0 37056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_387
timestamp 1679581782
transform 1 0 37728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_394
timestamp 1679581782
transform 1 0 38400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_401
timestamp 1679581782
transform 1 0 39072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_408
timestamp 1679581782
transform 1 0 39744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_415
timestamp 1679581782
transform 1 0 40416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_422
timestamp 1679581782
transform 1 0 41088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_429
timestamp 1679581782
transform 1 0 41760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_436
timestamp 1679581782
transform 1 0 42432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_443
timestamp 1679581782
transform 1 0 43104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_450
timestamp 1679581782
transform 1 0 43776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_457
timestamp 1679581782
transform 1 0 44448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_464
timestamp 1679581782
transform 1 0 45120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_471
timestamp 1679581782
transform 1 0 45792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_478
timestamp 1679581782
transform 1 0 46464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_485
timestamp 1679581782
transform 1 0 47136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_492
timestamp 1679581782
transform 1 0 47808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_499
timestamp 1679581782
transform 1 0 48480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_506
timestamp 1679581782
transform 1 0 49152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_513
timestamp 1679581782
transform 1 0 49824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_520
timestamp 1679581782
transform 1 0 50496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_527
timestamp 1679581782
transform 1 0 51168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_534
timestamp 1679581782
transform 1 0 51840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_541
timestamp 1679581782
transform 1 0 52512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_548
timestamp 1679581782
transform 1 0 53184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_555
timestamp 1679581782
transform 1 0 53856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_562
timestamp 1679581782
transform 1 0 54528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_569
timestamp 1679581782
transform 1 0 55200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_576
timestamp 1679581782
transform 1 0 55872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_583
timestamp 1679581782
transform 1 0 56544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_590
timestamp 1679581782
transform 1 0 57216 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_597
timestamp 1679581782
transform 1 0 57888 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_604
timestamp 1679581782
transform 1 0 58560 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_611
timestamp 1679581782
transform 1 0 59232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_618
timestamp 1679581782
transform 1 0 59904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_625
timestamp 1679581782
transform 1 0 60576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_632
timestamp 1679581782
transform 1 0 61248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_639
timestamp 1679581782
transform 1 0 61920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_646
timestamp 1679581782
transform 1 0 62592 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_653
timestamp 1679581782
transform 1 0 63264 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_660
timestamp 1679581782
transform 1 0 63936 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_667
timestamp 1679581782
transform 1 0 64608 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_674
timestamp 1679581782
transform 1 0 65280 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_681
timestamp 1679581782
transform 1 0 65952 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_19_688
timestamp 1679577901
transform 1 0 66624 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_692
timestamp 1677579658
transform 1 0 67008 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_701
timestamp 1677580104
transform 1 0 67872 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_19_708
timestamp 1679581782
transform 1 0 68544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_715
timestamp 1679581782
transform 1 0 69216 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_722
timestamp 1677579658
transform 1 0 69888 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_4
timestamp 1679581782
transform 1 0 960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_11
timestamp 1679581782
transform 1 0 1632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_18
timestamp 1679581782
transform 1 0 2304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_25
timestamp 1679581782
transform 1 0 2976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_32
timestamp 1679581782
transform 1 0 3648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_39
timestamp 1679581782
transform 1 0 4320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_46
timestamp 1679581782
transform 1 0 4992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_53
timestamp 1679581782
transform 1 0 5664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_60
timestamp 1679581782
transform 1 0 6336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_67
timestamp 1679581782
transform 1 0 7008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_74
timestamp 1679581782
transform 1 0 7680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_81
timestamp 1679581782
transform 1 0 8352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_88
timestamp 1679581782
transform 1 0 9024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_95
timestamp 1679581782
transform 1 0 9696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_102
timestamp 1679581782
transform 1 0 10368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_109
timestamp 1679581782
transform 1 0 11040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_116
timestamp 1679581782
transform 1 0 11712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_123
timestamp 1679581782
transform 1 0 12384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_130
timestamp 1679581782
transform 1 0 13056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_137
timestamp 1679581782
transform 1 0 13728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_144
timestamp 1679581782
transform 1 0 14400 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_151
timestamp 1679581782
transform 1 0 15072 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_158
timestamp 1679581782
transform 1 0 15744 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_165
timestamp 1679581782
transform 1 0 16416 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_172
timestamp 1679581782
transform 1 0 17088 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_179
timestamp 1679581782
transform 1 0 17760 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_186
timestamp 1679581782
transform 1 0 18432 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_193
timestamp 1679581782
transform 1 0 19104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_200
timestamp 1679581782
transform 1 0 19776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_207
timestamp 1679581782
transform 1 0 20448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_214
timestamp 1679581782
transform 1 0 21120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_221
timestamp 1679581782
transform 1 0 21792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_228
timestamp 1679581782
transform 1 0 22464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_235
timestamp 1679581782
transform 1 0 23136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_242
timestamp 1679581782
transform 1 0 23808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_249
timestamp 1679581782
transform 1 0 24480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_256
timestamp 1679581782
transform 1 0 25152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_263
timestamp 1679581782
transform 1 0 25824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_270
timestamp 1679581782
transform 1 0 26496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_277
timestamp 1679581782
transform 1 0 27168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_284
timestamp 1679581782
transform 1 0 27840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_291
timestamp 1679581782
transform 1 0 28512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_298
timestamp 1679581782
transform 1 0 29184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_305
timestamp 1679581782
transform 1 0 29856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_312
timestamp 1679581782
transform 1 0 30528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_319
timestamp 1679581782
transform 1 0 31200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_326
timestamp 1679581782
transform 1 0 31872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_333
timestamp 1679581782
transform 1 0 32544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_340
timestamp 1679581782
transform 1 0 33216 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_347
timestamp 1679581782
transform 1 0 33888 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_354
timestamp 1679581782
transform 1 0 34560 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_361
timestamp 1679581782
transform 1 0 35232 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_368
timestamp 1679581782
transform 1 0 35904 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_375
timestamp 1679581782
transform 1 0 36576 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_382
timestamp 1679581782
transform 1 0 37248 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_389
timestamp 1679581782
transform 1 0 37920 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_396
timestamp 1679581782
transform 1 0 38592 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_403
timestamp 1679581782
transform 1 0 39264 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_410
timestamp 1679581782
transform 1 0 39936 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_417
timestamp 1679581782
transform 1 0 40608 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_424
timestamp 1679581782
transform 1 0 41280 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_431
timestamp 1679581782
transform 1 0 41952 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_438
timestamp 1679581782
transform 1 0 42624 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_445
timestamp 1679581782
transform 1 0 43296 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_452
timestamp 1679581782
transform 1 0 43968 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_459
timestamp 1679581782
transform 1 0 44640 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_466
timestamp 1679581782
transform 1 0 45312 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_473
timestamp 1679581782
transform 1 0 45984 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_480
timestamp 1679581782
transform 1 0 46656 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_487
timestamp 1679581782
transform 1 0 47328 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_494
timestamp 1679581782
transform 1 0 48000 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_501
timestamp 1679581782
transform 1 0 48672 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_508
timestamp 1679581782
transform 1 0 49344 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_515
timestamp 1679581782
transform 1 0 50016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_522
timestamp 1679581782
transform 1 0 50688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_529
timestamp 1679581782
transform 1 0 51360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_536
timestamp 1679581782
transform 1 0 52032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_543
timestamp 1679581782
transform 1 0 52704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_550
timestamp 1679581782
transform 1 0 53376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_557
timestamp 1679581782
transform 1 0 54048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_564
timestamp 1679581782
transform 1 0 54720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_571
timestamp 1679581782
transform 1 0 55392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_578
timestamp 1679581782
transform 1 0 56064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_585
timestamp 1679581782
transform 1 0 56736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_592
timestamp 1679581782
transform 1 0 57408 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_599
timestamp 1679581782
transform 1 0 58080 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_606
timestamp 1679581782
transform 1 0 58752 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_613
timestamp 1679581782
transform 1 0 59424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_620
timestamp 1679581782
transform 1 0 60096 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_627
timestamp 1679581782
transform 1 0 60768 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_634
timestamp 1679581782
transform 1 0 61440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_641
timestamp 1679581782
transform 1 0 62112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_648
timestamp 1679581782
transform 1 0 62784 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_655
timestamp 1679581782
transform 1 0 63456 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_662
timestamp 1679581782
transform 1 0 64128 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_669
timestamp 1679581782
transform 1 0 64800 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_676
timestamp 1679581782
transform 1 0 65472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_683
timestamp 1679581782
transform 1 0 66144 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_690
timestamp 1679581782
transform 1 0 66816 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_697
timestamp 1679581782
transform 1 0 67488 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_704
timestamp 1679581782
transform 1 0 68160 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_711
timestamp 1677580104
transform 1 0 68832 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_717
timestamp 1679577901
transform 1 0 69408 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_721
timestamp 1677580104
transform 1 0 69792 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679581782
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_11
timestamp 1679581782
transform 1 0 1632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_18
timestamp 1679581782
transform 1 0 2304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_25
timestamp 1679581782
transform 1 0 2976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_32
timestamp 1679581782
transform 1 0 3648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_39
timestamp 1679581782
transform 1 0 4320 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_46
timestamp 1679581782
transform 1 0 4992 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_53
timestamp 1679581782
transform 1 0 5664 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_60
timestamp 1679581782
transform 1 0 6336 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_67
timestamp 1679581782
transform 1 0 7008 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_74
timestamp 1679581782
transform 1 0 7680 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_81
timestamp 1679581782
transform 1 0 8352 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_88
timestamp 1679581782
transform 1 0 9024 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_95
timestamp 1679581782
transform 1 0 9696 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_102
timestamp 1679581782
transform 1 0 10368 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_109
timestamp 1679581782
transform 1 0 11040 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_116
timestamp 1679581782
transform 1 0 11712 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_123
timestamp 1679581782
transform 1 0 12384 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_130
timestamp 1679581782
transform 1 0 13056 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_137
timestamp 1679581782
transform 1 0 13728 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_144
timestamp 1679581782
transform 1 0 14400 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_151
timestamp 1679581782
transform 1 0 15072 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_158
timestamp 1679581782
transform 1 0 15744 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_165
timestamp 1679581782
transform 1 0 16416 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_172
timestamp 1679581782
transform 1 0 17088 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_179
timestamp 1679581782
transform 1 0 17760 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_186
timestamp 1679581782
transform 1 0 18432 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_193
timestamp 1679581782
transform 1 0 19104 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_200
timestamp 1679581782
transform 1 0 19776 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_207
timestamp 1679581782
transform 1 0 20448 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_214
timestamp 1679581782
transform 1 0 21120 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_221
timestamp 1679581782
transform 1 0 21792 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_228
timestamp 1679581782
transform 1 0 22464 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_235
timestamp 1679581782
transform 1 0 23136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_242
timestamp 1679581782
transform 1 0 23808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_249
timestamp 1679581782
transform 1 0 24480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_256
timestamp 1679581782
transform 1 0 25152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_263
timestamp 1679581782
transform 1 0 25824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_270
timestamp 1679581782
transform 1 0 26496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_277
timestamp 1679581782
transform 1 0 27168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_284
timestamp 1679581782
transform 1 0 27840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_291
timestamp 1679581782
transform 1 0 28512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_298
timestamp 1679581782
transform 1 0 29184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_305
timestamp 1679581782
transform 1 0 29856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_312
timestamp 1679581782
transform 1 0 30528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_319
timestamp 1679581782
transform 1 0 31200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_326
timestamp 1679581782
transform 1 0 31872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_333
timestamp 1679581782
transform 1 0 32544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_340
timestamp 1679581782
transform 1 0 33216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_347
timestamp 1679581782
transform 1 0 33888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_354
timestamp 1679581782
transform 1 0 34560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_361
timestamp 1679581782
transform 1 0 35232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_368
timestamp 1679581782
transform 1 0 35904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_375
timestamp 1679581782
transform 1 0 36576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_382
timestamp 1679581782
transform 1 0 37248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_389
timestamp 1679581782
transform 1 0 37920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_396
timestamp 1679581782
transform 1 0 38592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_403
timestamp 1679581782
transform 1 0 39264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_410
timestamp 1679581782
transform 1 0 39936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_417
timestamp 1679581782
transform 1 0 40608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_424
timestamp 1679581782
transform 1 0 41280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_431
timestamp 1679581782
transform 1 0 41952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_438
timestamp 1679581782
transform 1 0 42624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_445
timestamp 1679581782
transform 1 0 43296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_452
timestamp 1679581782
transform 1 0 43968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_459
timestamp 1679581782
transform 1 0 44640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_466
timestamp 1679581782
transform 1 0 45312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_473
timestamp 1679581782
transform 1 0 45984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_480
timestamp 1679581782
transform 1 0 46656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_487
timestamp 1679581782
transform 1 0 47328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_494
timestamp 1679581782
transform 1 0 48000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_501
timestamp 1679581782
transform 1 0 48672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_508
timestamp 1679581782
transform 1 0 49344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_515
timestamp 1679581782
transform 1 0 50016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_522
timestamp 1679581782
transform 1 0 50688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_529
timestamp 1679581782
transform 1 0 51360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_536
timestamp 1679581782
transform 1 0 52032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_543
timestamp 1679581782
transform 1 0 52704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_550
timestamp 1679581782
transform 1 0 53376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_557
timestamp 1679581782
transform 1 0 54048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_564
timestamp 1679581782
transform 1 0 54720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_571
timestamp 1679581782
transform 1 0 55392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_578
timestamp 1679581782
transform 1 0 56064 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_585
timestamp 1679581782
transform 1 0 56736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_592
timestamp 1679581782
transform 1 0 57408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_599
timestamp 1679581782
transform 1 0 58080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_606
timestamp 1679581782
transform 1 0 58752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_613
timestamp 1679581782
transform 1 0 59424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_620
timestamp 1679581782
transform 1 0 60096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_627
timestamp 1679581782
transform 1 0 60768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_634
timestamp 1679581782
transform 1 0 61440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_641
timestamp 1679581782
transform 1 0 62112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_648
timestamp 1679581782
transform 1 0 62784 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_655
timestamp 1679581782
transform 1 0 63456 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_662
timestamp 1679581782
transform 1 0 64128 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_669
timestamp 1679581782
transform 1 0 64800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_676
timestamp 1679581782
transform 1 0 65472 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_683
timestamp 1679581782
transform 1 0 66144 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_690
timestamp 1679581782
transform 1 0 66816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_697
timestamp 1679581782
transform 1 0 67488 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_704
timestamp 1679581782
transform 1 0 68160 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_711
timestamp 1679581782
transform 1 0 68832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_21_718
timestamp 1679577901
transform 1 0 69504 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_722
timestamp 1677579658
transform 1 0 69888 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_4
timestamp 1679581782
transform 1 0 960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_11
timestamp 1679581782
transform 1 0 1632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_18
timestamp 1679581782
transform 1 0 2304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_25
timestamp 1679581782
transform 1 0 2976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_32
timestamp 1679581782
transform 1 0 3648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_39
timestamp 1679581782
transform 1 0 4320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_46
timestamp 1679581782
transform 1 0 4992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_53
timestamp 1679581782
transform 1 0 5664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_60
timestamp 1679581782
transform 1 0 6336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_67
timestamp 1679581782
transform 1 0 7008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_74
timestamp 1679581782
transform 1 0 7680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_81
timestamp 1679581782
transform 1 0 8352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_88
timestamp 1679581782
transform 1 0 9024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_95
timestamp 1679581782
transform 1 0 9696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_102
timestamp 1679581782
transform 1 0 10368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_109
timestamp 1679581782
transform 1 0 11040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_116
timestamp 1679581782
transform 1 0 11712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_123
timestamp 1679581782
transform 1 0 12384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_130
timestamp 1679581782
transform 1 0 13056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_137
timestamp 1679581782
transform 1 0 13728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_144
timestamp 1679581782
transform 1 0 14400 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_151
timestamp 1679581782
transform 1 0 15072 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_158
timestamp 1679581782
transform 1 0 15744 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_165
timestamp 1679581782
transform 1 0 16416 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_172
timestamp 1679581782
transform 1 0 17088 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_179
timestamp 1679581782
transform 1 0 17760 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_186
timestamp 1679581782
transform 1 0 18432 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_193
timestamp 1679581782
transform 1 0 19104 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_200
timestamp 1679581782
transform 1 0 19776 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_207
timestamp 1679581782
transform 1 0 20448 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_214
timestamp 1679581782
transform 1 0 21120 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_221
timestamp 1679581782
transform 1 0 21792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_228
timestamp 1679581782
transform 1 0 22464 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_235
timestamp 1679581782
transform 1 0 23136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_242
timestamp 1679581782
transform 1 0 23808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_249
timestamp 1679581782
transform 1 0 24480 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_256
timestamp 1679581782
transform 1 0 25152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_263
timestamp 1679581782
transform 1 0 25824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_270
timestamp 1679581782
transform 1 0 26496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_277
timestamp 1679581782
transform 1 0 27168 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_284
timestamp 1679581782
transform 1 0 27840 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_291
timestamp 1679581782
transform 1 0 28512 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_298
timestamp 1679581782
transform 1 0 29184 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_305
timestamp 1679581782
transform 1 0 29856 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_312
timestamp 1679581782
transform 1 0 30528 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_319
timestamp 1679581782
transform 1 0 31200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_326
timestamp 1679581782
transform 1 0 31872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_333
timestamp 1679581782
transform 1 0 32544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_340
timestamp 1679581782
transform 1 0 33216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_347
timestamp 1679581782
transform 1 0 33888 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_354
timestamp 1679581782
transform 1 0 34560 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_361
timestamp 1679581782
transform 1 0 35232 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_368
timestamp 1679581782
transform 1 0 35904 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_375
timestamp 1679581782
transform 1 0 36576 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_382
timestamp 1679581782
transform 1 0 37248 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_389
timestamp 1679581782
transform 1 0 37920 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_396
timestamp 1679581782
transform 1 0 38592 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_403
timestamp 1679581782
transform 1 0 39264 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_410
timestamp 1679581782
transform 1 0 39936 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_417
timestamp 1679581782
transform 1 0 40608 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_424
timestamp 1679581782
transform 1 0 41280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_431
timestamp 1679581782
transform 1 0 41952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_438
timestamp 1679581782
transform 1 0 42624 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_445
timestamp 1679581782
transform 1 0 43296 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_452
timestamp 1679581782
transform 1 0 43968 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_459
timestamp 1679581782
transform 1 0 44640 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_466
timestamp 1679581782
transform 1 0 45312 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_473
timestamp 1679581782
transform 1 0 45984 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_480
timestamp 1679581782
transform 1 0 46656 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_487
timestamp 1679581782
transform 1 0 47328 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_494
timestamp 1679581782
transform 1 0 48000 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_501
timestamp 1679581782
transform 1 0 48672 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_508
timestamp 1679581782
transform 1 0 49344 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_515
timestamp 1679581782
transform 1 0 50016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_522
timestamp 1679581782
transform 1 0 50688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_529
timestamp 1679581782
transform 1 0 51360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_536
timestamp 1679581782
transform 1 0 52032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_543
timestamp 1679581782
transform 1 0 52704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_550
timestamp 1679581782
transform 1 0 53376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_557
timestamp 1679581782
transform 1 0 54048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_564
timestamp 1679581782
transform 1 0 54720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_571
timestamp 1679581782
transform 1 0 55392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_578
timestamp 1679581782
transform 1 0 56064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_585
timestamp 1679581782
transform 1 0 56736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_592
timestamp 1679581782
transform 1 0 57408 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_599
timestamp 1679581782
transform 1 0 58080 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_606
timestamp 1679581782
transform 1 0 58752 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_613
timestamp 1679581782
transform 1 0 59424 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_620
timestamp 1679581782
transform 1 0 60096 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_627
timestamp 1679581782
transform 1 0 60768 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_634
timestamp 1679581782
transform 1 0 61440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_641
timestamp 1679581782
transform 1 0 62112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_648
timestamp 1679581782
transform 1 0 62784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_655
timestamp 1679581782
transform 1 0 63456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_662
timestamp 1679581782
transform 1 0 64128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_669
timestamp 1679581782
transform 1 0 64800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_676
timestamp 1679581782
transform 1 0 65472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_683
timestamp 1679581782
transform 1 0 66144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_690
timestamp 1679581782
transform 1 0 66816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_697
timestamp 1679581782
transform 1 0 67488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_704
timestamp 1679581782
transform 1 0 68160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_711
timestamp 1679581782
transform 1 0 68832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_718
timestamp 1679581782
transform 1 0 69504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_725
timestamp 1679581782
transform 1 0 70176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_732
timestamp 1679581782
transform 1 0 70848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_739
timestamp 1679581782
transform 1 0 71520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_746
timestamp 1679581782
transform 1 0 72192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_753
timestamp 1679581782
transform 1 0 72864 0 1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_760
timestamp 1677579658
transform 1 0 73536 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_773
timestamp 1677580104
transform 1 0 74784 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_785
timestamp 1677580104
transform 1 0 75936 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_806
timestamp 1677580104
transform 1 0 77952 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_812
timestamp 1677579658
transform 1 0 78528 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_820
timestamp 1677579658
transform 1 0 79296 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_824
timestamp 1677579658
transform 1 0 79680 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_845
timestamp 1677579658
transform 1 0 81696 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_849
timestamp 1677579658
transform 1 0 82080 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_853
timestamp 1677579658
transform 1 0 82464 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_861
timestamp 1677579658
transform 1 0 83232 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_865
timestamp 1677579658
transform 1 0 83616 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_869
timestamp 1677579658
transform 1 0 84000 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_873
timestamp 1677580104
transform 1 0 84384 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_882
timestamp 1677579658
transform 1 0 85248 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_886
timestamp 1677579658
transform 1 0 85632 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_890
timestamp 1677579658
transform 1 0 86016 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_898
timestamp 1677580104
transform 1 0 86784 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_903
timestamp 1677579658
transform 1 0 87264 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_907
timestamp 1679577901
transform 1 0 87648 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_911
timestamp 1677579658
transform 1 0 88032 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_915
timestamp 1677579658
transform 1 0 88416 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_919
timestamp 1677580104
transform 1 0 88800 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_924
timestamp 1677579658
transform 1 0 89280 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_932
timestamp 1677579658
transform 1 0 90048 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_936
timestamp 1677579658
transform 1 0 90432 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_940
timestamp 1677579658
transform 1 0 90816 0 1 17388
box -48 -56 144 834
use sg13g2_fill_1  FILLER_22_944
timestamp 1677579658
transform 1 0 91200 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_948
timestamp 1677580104
transform 1 0 91584 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_953
timestamp 1677579658
transform 1 0 92064 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_957
timestamp 1677580104
transform 1 0 92448 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_959
timestamp 1677579658
transform 1 0 92640 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_966
timestamp 1677580104
transform 1 0 93312 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_978
timestamp 1677580104
transform 1 0 94464 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_990
timestamp 1677580104
transform 1 0 95616 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_999
timestamp 1677579658
transform 1 0 96480 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_1015
timestamp 1677580104
transform 1 0 98016 0 1 17388
box -48 -56 240 834
use sg13g2_decap_4  FILLER_22_1024
timestamp 1679577901
transform 1 0 98880 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_1028
timestamp 1677579658
transform 1 0 99264 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679581782
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_11
timestamp 1679581782
transform 1 0 1632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_18
timestamp 1679581782
transform 1 0 2304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_25
timestamp 1679581782
transform 1 0 2976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_32
timestamp 1679581782
transform 1 0 3648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_39
timestamp 1679581782
transform 1 0 4320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_46
timestamp 1679581782
transform 1 0 4992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_53
timestamp 1679581782
transform 1 0 5664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_60
timestamp 1679581782
transform 1 0 6336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_67
timestamp 1679581782
transform 1 0 7008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_74
timestamp 1679581782
transform 1 0 7680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_81
timestamp 1679581782
transform 1 0 8352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_88
timestamp 1679581782
transform 1 0 9024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_95
timestamp 1679581782
transform 1 0 9696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_102
timestamp 1679581782
transform 1 0 10368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_109
timestamp 1679581782
transform 1 0 11040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_116
timestamp 1679581782
transform 1 0 11712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_123
timestamp 1679581782
transform 1 0 12384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_130
timestamp 1679581782
transform 1 0 13056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_137
timestamp 1679581782
transform 1 0 13728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_144
timestamp 1679581782
transform 1 0 14400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_151
timestamp 1679581782
transform 1 0 15072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_158
timestamp 1679581782
transform 1 0 15744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_165
timestamp 1679581782
transform 1 0 16416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_172
timestamp 1679581782
transform 1 0 17088 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_179
timestamp 1679581782
transform 1 0 17760 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_186
timestamp 1679581782
transform 1 0 18432 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_193
timestamp 1679581782
transform 1 0 19104 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_200
timestamp 1679581782
transform 1 0 19776 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_207
timestamp 1679581782
transform 1 0 20448 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_214
timestamp 1679581782
transform 1 0 21120 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_221
timestamp 1679581782
transform 1 0 21792 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_228
timestamp 1679581782
transform 1 0 22464 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_235
timestamp 1679581782
transform 1 0 23136 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_242
timestamp 1679581782
transform 1 0 23808 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_249
timestamp 1679581782
transform 1 0 24480 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_256
timestamp 1679581782
transform 1 0 25152 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_263
timestamp 1679581782
transform 1 0 25824 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_270
timestamp 1679581782
transform 1 0 26496 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_277
timestamp 1679581782
transform 1 0 27168 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_284
timestamp 1679581782
transform 1 0 27840 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_291
timestamp 1679581782
transform 1 0 28512 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_298
timestamp 1679581782
transform 1 0 29184 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_305
timestamp 1679581782
transform 1 0 29856 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_312
timestamp 1679581782
transform 1 0 30528 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_319
timestamp 1679581782
transform 1 0 31200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_326
timestamp 1679581782
transform 1 0 31872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_333
timestamp 1679581782
transform 1 0 32544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_340
timestamp 1679581782
transform 1 0 33216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_347
timestamp 1679581782
transform 1 0 33888 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_354
timestamp 1679581782
transform 1 0 34560 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_361
timestamp 1679581782
transform 1 0 35232 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_368
timestamp 1679581782
transform 1 0 35904 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_375
timestamp 1679581782
transform 1 0 36576 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_382
timestamp 1679581782
transform 1 0 37248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_389
timestamp 1679581782
transform 1 0 37920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_396
timestamp 1679581782
transform 1 0 38592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_403
timestamp 1679581782
transform 1 0 39264 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_410
timestamp 1679581782
transform 1 0 39936 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_417
timestamp 1679581782
transform 1 0 40608 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_424
timestamp 1679581782
transform 1 0 41280 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_431
timestamp 1679581782
transform 1 0 41952 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_438
timestamp 1679581782
transform 1 0 42624 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_445
timestamp 1679581782
transform 1 0 43296 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_452
timestamp 1679581782
transform 1 0 43968 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_459
timestamp 1679581782
transform 1 0 44640 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_466
timestamp 1679581782
transform 1 0 45312 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_473
timestamp 1679581782
transform 1 0 45984 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_480
timestamp 1679581782
transform 1 0 46656 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_487
timestamp 1679581782
transform 1 0 47328 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_494
timestamp 1679581782
transform 1 0 48000 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_501
timestamp 1679581782
transform 1 0 48672 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_508
timestamp 1679581782
transform 1 0 49344 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_515
timestamp 1679581782
transform 1 0 50016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_522
timestamp 1679581782
transform 1 0 50688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_529
timestamp 1679581782
transform 1 0 51360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_536
timestamp 1679581782
transform 1 0 52032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_543
timestamp 1679581782
transform 1 0 52704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_550
timestamp 1679581782
transform 1 0 53376 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_557
timestamp 1679581782
transform 1 0 54048 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_564
timestamp 1679581782
transform 1 0 54720 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_571
timestamp 1679581782
transform 1 0 55392 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_578
timestamp 1679581782
transform 1 0 56064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_585
timestamp 1679581782
transform 1 0 56736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_592
timestamp 1679581782
transform 1 0 57408 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_599
timestamp 1679581782
transform 1 0 58080 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_606
timestamp 1679581782
transform 1 0 58752 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_613
timestamp 1679581782
transform 1 0 59424 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_620
timestamp 1679581782
transform 1 0 60096 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_627
timestamp 1679581782
transform 1 0 60768 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_634
timestamp 1679581782
transform 1 0 61440 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_641
timestamp 1679581782
transform 1 0 62112 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_648
timestamp 1679581782
transform 1 0 62784 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_655
timestamp 1679581782
transform 1 0 63456 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_662
timestamp 1679581782
transform 1 0 64128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_669
timestamp 1679581782
transform 1 0 64800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_676
timestamp 1679581782
transform 1 0 65472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_683
timestamp 1679581782
transform 1 0 66144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_690
timestamp 1679581782
transform 1 0 66816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_697
timestamp 1679581782
transform 1 0 67488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_704
timestamp 1679581782
transform 1 0 68160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_711
timestamp 1679581782
transform 1 0 68832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_718
timestamp 1679581782
transform 1 0 69504 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_725
timestamp 1679581782
transform 1 0 70176 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_732
timestamp 1679581782
transform 1 0 70848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_739
timestamp 1679581782
transform 1 0 71520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_746
timestamp 1679581782
transform 1 0 72192 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_756
timestamp 1679581782
transform 1 0 73152 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_763
timestamp 1677580104
transform 1 0 73824 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_765
timestamp 1677579658
transform 1 0 74016 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_769
timestamp 1677579658
transform 1 0 74400 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_778
timestamp 1679577901
transform 1 0 75264 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_782
timestamp 1677579658
transform 1 0 75648 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_787
timestamp 1677580104
transform 1 0 76128 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_789
timestamp 1677579658
transform 1 0 76320 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_793
timestamp 1679581782
transform 1 0 76704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_803
timestamp 1679577901
transform 1 0 77664 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_818
timestamp 1677580104
transform 1 0 79104 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_824
timestamp 1677579658
transform 1 0 79680 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_829
timestamp 1679581782
transform 1 0 80160 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_836
timestamp 1677579658
transform 1 0 80832 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_849
timestamp 1677579658
transform 1 0 82080 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_854
timestamp 1679577901
transform 1 0 82560 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_870
timestamp 1677579658
transform 1 0 84096 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_882
timestamp 1677580104
transform 1 0 85248 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_899
timestamp 1677579658
transform 1 0 86880 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_904
timestamp 1677580104
transform 1 0 87360 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_906
timestamp 1677579658
transform 1 0 87552 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_911
timestamp 1677579658
transform 1 0 88032 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_924
timestamp 1677579658
transform 1 0 89280 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_936
timestamp 1677579658
transform 1 0 90432 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_941
timestamp 1677580104
transform 1 0 90912 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_943
timestamp 1677579658
transform 1 0 91104 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_967
timestamp 1679577901
transform 1 0 93408 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_979
timestamp 1677579658
transform 1 0 94560 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_987
timestamp 1677579658
transform 1 0 95328 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_23_995
timestamp 1677579658
transform 1 0 96096 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_1000
timestamp 1677580104
transform 1 0 96576 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_1012
timestamp 1679581782
transform 1 0 97728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1019
timestamp 1679581782
transform 1 0 98400 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_1026
timestamp 1677580104
transform 1 0 99072 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_1028
timestamp 1677579658
transform 1 0 99264 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679581782
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_18
timestamp 1679581782
transform 1 0 2304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_25
timestamp 1679581782
transform 1 0 2976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_32
timestamp 1679581782
transform 1 0 3648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_39
timestamp 1679581782
transform 1 0 4320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_46
timestamp 1679581782
transform 1 0 4992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_53
timestamp 1679581782
transform 1 0 5664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_60
timestamp 1679581782
transform 1 0 6336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_67
timestamp 1679581782
transform 1 0 7008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_74
timestamp 1679581782
transform 1 0 7680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_81
timestamp 1679581782
transform 1 0 8352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_88
timestamp 1679581782
transform 1 0 9024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_95
timestamp 1679581782
transform 1 0 9696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_102
timestamp 1679581782
transform 1 0 10368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_109
timestamp 1679581782
transform 1 0 11040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_116
timestamp 1679581782
transform 1 0 11712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_123
timestamp 1679581782
transform 1 0 12384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_130
timestamp 1679581782
transform 1 0 13056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_137
timestamp 1679581782
transform 1 0 13728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_144
timestamp 1679581782
transform 1 0 14400 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_151
timestamp 1679581782
transform 1 0 15072 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_158
timestamp 1679581782
transform 1 0 15744 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_165
timestamp 1679581782
transform 1 0 16416 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_172
timestamp 1679581782
transform 1 0 17088 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_179
timestamp 1679581782
transform 1 0 17760 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_186
timestamp 1679581782
transform 1 0 18432 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_193
timestamp 1679581782
transform 1 0 19104 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_200
timestamp 1679581782
transform 1 0 19776 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_207
timestamp 1679581782
transform 1 0 20448 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_214
timestamp 1679581782
transform 1 0 21120 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_221
timestamp 1679581782
transform 1 0 21792 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_228
timestamp 1679581782
transform 1 0 22464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_235
timestamp 1679581782
transform 1 0 23136 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_242
timestamp 1679581782
transform 1 0 23808 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_249
timestamp 1679581782
transform 1 0 24480 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_256
timestamp 1679581782
transform 1 0 25152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_263
timestamp 1679581782
transform 1 0 25824 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_270
timestamp 1679581782
transform 1 0 26496 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_277
timestamp 1679581782
transform 1 0 27168 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_284
timestamp 1679581782
transform 1 0 27840 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_291
timestamp 1679581782
transform 1 0 28512 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_298
timestamp 1679581782
transform 1 0 29184 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_305
timestamp 1679581782
transform 1 0 29856 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_312
timestamp 1679581782
transform 1 0 30528 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_319
timestamp 1679581782
transform 1 0 31200 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_326
timestamp 1679581782
transform 1 0 31872 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_333
timestamp 1679581782
transform 1 0 32544 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_340
timestamp 1679581782
transform 1 0 33216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_347
timestamp 1679581782
transform 1 0 33888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_354
timestamp 1679581782
transform 1 0 34560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_361
timestamp 1679581782
transform 1 0 35232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_368
timestamp 1679581782
transform 1 0 35904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_375
timestamp 1679581782
transform 1 0 36576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_382
timestamp 1679581782
transform 1 0 37248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_389
timestamp 1679581782
transform 1 0 37920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_396
timestamp 1679581782
transform 1 0 38592 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_403
timestamp 1679581782
transform 1 0 39264 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_410
timestamp 1679581782
transform 1 0 39936 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_417
timestamp 1679581782
transform 1 0 40608 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_424
timestamp 1679581782
transform 1 0 41280 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_431
timestamp 1679581782
transform 1 0 41952 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_438
timestamp 1679581782
transform 1 0 42624 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_445
timestamp 1679581782
transform 1 0 43296 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_452
timestamp 1679581782
transform 1 0 43968 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_459
timestamp 1679581782
transform 1 0 44640 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_466
timestamp 1679581782
transform 1 0 45312 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_473
timestamp 1679581782
transform 1 0 45984 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_480
timestamp 1679581782
transform 1 0 46656 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_487
timestamp 1679581782
transform 1 0 47328 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_494
timestamp 1679581782
transform 1 0 48000 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_501
timestamp 1679581782
transform 1 0 48672 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_508
timestamp 1679581782
transform 1 0 49344 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_515
timestamp 1679581782
transform 1 0 50016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_522
timestamp 1679581782
transform 1 0 50688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_529
timestamp 1679581782
transform 1 0 51360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_536
timestamp 1679581782
transform 1 0 52032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_543
timestamp 1679581782
transform 1 0 52704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_550
timestamp 1679581782
transform 1 0 53376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_557
timestamp 1679581782
transform 1 0 54048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_564
timestamp 1679581782
transform 1 0 54720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_571
timestamp 1679581782
transform 1 0 55392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_578
timestamp 1679581782
transform 1 0 56064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_585
timestamp 1679581782
transform 1 0 56736 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_592
timestamp 1679581782
transform 1 0 57408 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_599
timestamp 1679581782
transform 1 0 58080 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_606
timestamp 1679581782
transform 1 0 58752 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_613
timestamp 1679581782
transform 1 0 59424 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_620
timestamp 1679581782
transform 1 0 60096 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_627
timestamp 1679581782
transform 1 0 60768 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_634
timestamp 1679581782
transform 1 0 61440 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_641
timestamp 1679581782
transform 1 0 62112 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_648
timestamp 1679581782
transform 1 0 62784 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_655
timestamp 1679581782
transform 1 0 63456 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_662
timestamp 1679581782
transform 1 0 64128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_669
timestamp 1679581782
transform 1 0 64800 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_676
timestamp 1679581782
transform 1 0 65472 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_683
timestamp 1679581782
transform 1 0 66144 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_690
timestamp 1679581782
transform 1 0 66816 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_697
timestamp 1679581782
transform 1 0 67488 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_704
timestamp 1679581782
transform 1 0 68160 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_711
timestamp 1679581782
transform 1 0 68832 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_718
timestamp 1679581782
transform 1 0 69504 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_725
timestamp 1679581782
transform 1 0 70176 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_732
timestamp 1679581782
transform 1 0 70848 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_739
timestamp 1679581782
transform 1 0 71520 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_746
timestamp 1679581782
transform 1 0 72192 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_753
timestamp 1679581782
transform 1 0 72864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_760
timestamp 1679581782
transform 1 0 73536 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_767
timestamp 1679577901
transform 1 0 74208 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_771
timestamp 1677579658
transform 1 0 74592 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_784
timestamp 1679581782
transform 1 0 75840 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_794
timestamp 1677580104
transform 1 0 76800 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_799
timestamp 1677580104
transform 1 0 77280 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_801
timestamp 1677579658
transform 1 0 77472 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_810
timestamp 1677580104
transform 1 0 78336 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_815
timestamp 1679581782
transform 1 0 78816 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_822
timestamp 1679577901
transform 1 0 79488 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_826
timestamp 1677579658
transform 1 0 79872 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_834
timestamp 1679581782
transform 1 0 80640 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_841
timestamp 1679577901
transform 1 0 81312 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_845
timestamp 1677579658
transform 1 0 81696 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_850
timestamp 1679577901
transform 1 0 82176 0 1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_857
timestamp 1679581782
transform 1 0 82848 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_864
timestamp 1677580104
transform 1 0 83520 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_866
timestamp 1677579658
transform 1 0 83712 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_871
timestamp 1679581782
transform 1 0 84192 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_878
timestamp 1679581782
transform 1 0 84864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_889
timestamp 1679577901
transform 1 0 85920 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_901
timestamp 1677580104
transform 1 0 87072 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_903
timestamp 1677579658
transform 1 0 87264 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_908
timestamp 1677580104
transform 1 0 87744 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_917
timestamp 1679581782
transform 1 0 88608 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_924
timestamp 1677580104
transform 1 0 89280 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_934
timestamp 1679581782
transform 1 0 90240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_941
timestamp 1679577901
transform 1 0 90912 0 1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_24_949
timestamp 1679581782
transform 1 0 91680 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_956
timestamp 1677579658
transform 1 0 92352 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_965
timestamp 1679581782
transform 1 0 93216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_976
timestamp 1679581782
transform 1 0 94272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_24_983
timestamp 1679577901
transform 1 0 94944 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_987
timestamp 1677580104
transform 1 0 95328 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_24_993
timestamp 1679581782
transform 1 0 95904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1000
timestamp 1679581782
transform 1 0 96576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1007
timestamp 1679581782
transform 1 0 97248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1014
timestamp 1679581782
transform 1 0 97920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1021
timestamp 1679581782
transform 1 0 98592 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_1028
timestamp 1677579658
transform 1 0 99264 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679581782
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679581782
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679581782
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_25
timestamp 1679581782
transform 1 0 2976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_32
timestamp 1679581782
transform 1 0 3648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_39
timestamp 1679581782
transform 1 0 4320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_46
timestamp 1679581782
transform 1 0 4992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_53
timestamp 1679581782
transform 1 0 5664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_60
timestamp 1679581782
transform 1 0 6336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_67
timestamp 1679581782
transform 1 0 7008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_74
timestamp 1679581782
transform 1 0 7680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_81
timestamp 1679581782
transform 1 0 8352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_88
timestamp 1679581782
transform 1 0 9024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_95
timestamp 1679581782
transform 1 0 9696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_102
timestamp 1679581782
transform 1 0 10368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_109
timestamp 1679581782
transform 1 0 11040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_116
timestamp 1679581782
transform 1 0 11712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_123
timestamp 1679581782
transform 1 0 12384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_130
timestamp 1679581782
transform 1 0 13056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_137
timestamp 1679581782
transform 1 0 13728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_144
timestamp 1679581782
transform 1 0 14400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_151
timestamp 1679581782
transform 1 0 15072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_158
timestamp 1679581782
transform 1 0 15744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_165
timestamp 1679581782
transform 1 0 16416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_172
timestamp 1679581782
transform 1 0 17088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_179
timestamp 1679581782
transform 1 0 17760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_186
timestamp 1679581782
transform 1 0 18432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_193
timestamp 1679581782
transform 1 0 19104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_200
timestamp 1679581782
transform 1 0 19776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_207
timestamp 1679581782
transform 1 0 20448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_214
timestamp 1679581782
transform 1 0 21120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_221
timestamp 1679581782
transform 1 0 21792 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_228
timestamp 1679581782
transform 1 0 22464 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_235
timestamp 1679581782
transform 1 0 23136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_242
timestamp 1679581782
transform 1 0 23808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_249
timestamp 1679581782
transform 1 0 24480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_256
timestamp 1679581782
transform 1 0 25152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_263
timestamp 1679581782
transform 1 0 25824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_270
timestamp 1679581782
transform 1 0 26496 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_277
timestamp 1679581782
transform 1 0 27168 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_284
timestamp 1679581782
transform 1 0 27840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_291
timestamp 1679581782
transform 1 0 28512 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_298
timestamp 1679581782
transform 1 0 29184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_305
timestamp 1679581782
transform 1 0 29856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_312
timestamp 1679581782
transform 1 0 30528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_319
timestamp 1679581782
transform 1 0 31200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_326
timestamp 1679581782
transform 1 0 31872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_333
timestamp 1679581782
transform 1 0 32544 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_340
timestamp 1679581782
transform 1 0 33216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_347
timestamp 1679581782
transform 1 0 33888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_354
timestamp 1679581782
transform 1 0 34560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_361
timestamp 1679581782
transform 1 0 35232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_368
timestamp 1679581782
transform 1 0 35904 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_375
timestamp 1679581782
transform 1 0 36576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_382
timestamp 1679581782
transform 1 0 37248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_389
timestamp 1679581782
transform 1 0 37920 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_396
timestamp 1679581782
transform 1 0 38592 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_403
timestamp 1679581782
transform 1 0 39264 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_410
timestamp 1679581782
transform 1 0 39936 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_417
timestamp 1679581782
transform 1 0 40608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_424
timestamp 1679581782
transform 1 0 41280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_431
timestamp 1679581782
transform 1 0 41952 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_438
timestamp 1679581782
transform 1 0 42624 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_445
timestamp 1679581782
transform 1 0 43296 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_452
timestamp 1679581782
transform 1 0 43968 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_459
timestamp 1679581782
transform 1 0 44640 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_466
timestamp 1679581782
transform 1 0 45312 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_473
timestamp 1679581782
transform 1 0 45984 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_480
timestamp 1679581782
transform 1 0 46656 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_487
timestamp 1679581782
transform 1 0 47328 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_494
timestamp 1679581782
transform 1 0 48000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_501
timestamp 1679581782
transform 1 0 48672 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_508
timestamp 1679581782
transform 1 0 49344 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_515
timestamp 1679581782
transform 1 0 50016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_522
timestamp 1679581782
transform 1 0 50688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_529
timestamp 1679581782
transform 1 0 51360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_536
timestamp 1679581782
transform 1 0 52032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_543
timestamp 1679581782
transform 1 0 52704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_550
timestamp 1679581782
transform 1 0 53376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_557
timestamp 1679581782
transform 1 0 54048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_564
timestamp 1679581782
transform 1 0 54720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_571
timestamp 1679581782
transform 1 0 55392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_578
timestamp 1679581782
transform 1 0 56064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_585
timestamp 1679581782
transform 1 0 56736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_592
timestamp 1679581782
transform 1 0 57408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_599
timestamp 1679581782
transform 1 0 58080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_606
timestamp 1679581782
transform 1 0 58752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_613
timestamp 1679581782
transform 1 0 59424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_620
timestamp 1679581782
transform 1 0 60096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_627
timestamp 1679581782
transform 1 0 60768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_634
timestamp 1679581782
transform 1 0 61440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_641
timestamp 1679581782
transform 1 0 62112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_648
timestamp 1679581782
transform 1 0 62784 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_655
timestamp 1679581782
transform 1 0 63456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_662
timestamp 1679581782
transform 1 0 64128 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_669
timestamp 1679581782
transform 1 0 64800 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_676
timestamp 1679581782
transform 1 0 65472 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_683
timestamp 1679581782
transform 1 0 66144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_690
timestamp 1679581782
transform 1 0 66816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_697
timestamp 1679581782
transform 1 0 67488 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_704
timestamp 1679581782
transform 1 0 68160 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_711
timestamp 1679581782
transform 1 0 68832 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_718
timestamp 1679581782
transform 1 0 69504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_725
timestamp 1679581782
transform 1 0 70176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_732
timestamp 1679581782
transform 1 0 70848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_739
timestamp 1679581782
transform 1 0 71520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_746
timestamp 1679581782
transform 1 0 72192 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_753
timestamp 1679581782
transform 1 0 72864 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_760
timestamp 1679581782
transform 1 0 73536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_767
timestamp 1679581782
transform 1 0 74208 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_774
timestamp 1679577901
transform 1 0 74880 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_778
timestamp 1677580104
transform 1 0 75264 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_784
timestamp 1679581782
transform 1 0 75840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_791
timestamp 1679581782
transform 1 0 76512 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_798
timestamp 1679581782
transform 1 0 77184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_805
timestamp 1679581782
transform 1 0 77856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_812
timestamp 1679581782
transform 1 0 78528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_819
timestamp 1679581782
transform 1 0 79200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_826
timestamp 1679577901
transform 1 0 79872 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_830
timestamp 1677579658
transform 1 0 80256 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_835
timestamp 1679581782
transform 1 0 80736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_842
timestamp 1679581782
transform 1 0 81408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_849
timestamp 1679581782
transform 1 0 82080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_856
timestamp 1679581782
transform 1 0 82752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_863
timestamp 1679581782
transform 1 0 83424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_870
timestamp 1679581782
transform 1 0 84096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_877
timestamp 1679581782
transform 1 0 84768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_884
timestamp 1679581782
transform 1 0 85440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_891
timestamp 1679581782
transform 1 0 86112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_902
timestamp 1679581782
transform 1 0 87168 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_909
timestamp 1679581782
transform 1 0 87840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_916
timestamp 1679581782
transform 1 0 88512 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_923
timestamp 1679581782
transform 1 0 89184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_930
timestamp 1679581782
transform 1 0 89856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_937
timestamp 1679581782
transform 1 0 90528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_944
timestamp 1679581782
transform 1 0 91200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_951
timestamp 1679581782
transform 1 0 91872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_25_958
timestamp 1679577901
transform 1 0 92544 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_25_966
timestamp 1679581782
transform 1 0 93312 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_973
timestamp 1679581782
transform 1 0 93984 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_980
timestamp 1679581782
transform 1 0 94656 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_987
timestamp 1679581782
transform 1 0 95328 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_994
timestamp 1679581782
transform 1 0 96000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1001
timestamp 1679581782
transform 1 0 96672 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1008
timestamp 1679581782
transform 1 0 97344 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1015
timestamp 1679581782
transform 1 0 98016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1022
timestamp 1679581782
transform 1 0 98688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679581782
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_18
timestamp 1679581782
transform 1 0 2304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_25
timestamp 1679581782
transform 1 0 2976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_32
timestamp 1679581782
transform 1 0 3648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_39
timestamp 1679581782
transform 1 0 4320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_46
timestamp 1679581782
transform 1 0 4992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_53
timestamp 1679581782
transform 1 0 5664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_60
timestamp 1679581782
transform 1 0 6336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_67
timestamp 1679581782
transform 1 0 7008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_74
timestamp 1679581782
transform 1 0 7680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_81
timestamp 1679581782
transform 1 0 8352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_88
timestamp 1679581782
transform 1 0 9024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_95
timestamp 1679581782
transform 1 0 9696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_102
timestamp 1679581782
transform 1 0 10368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_109
timestamp 1679581782
transform 1 0 11040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_116
timestamp 1679581782
transform 1 0 11712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_123
timestamp 1679581782
transform 1 0 12384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_130
timestamp 1679581782
transform 1 0 13056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_137
timestamp 1679581782
transform 1 0 13728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_144
timestamp 1679581782
transform 1 0 14400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_151
timestamp 1679581782
transform 1 0 15072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_158
timestamp 1679581782
transform 1 0 15744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_165
timestamp 1679581782
transform 1 0 16416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_172
timestamp 1679581782
transform 1 0 17088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_179
timestamp 1679581782
transform 1 0 17760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_186
timestamp 1679581782
transform 1 0 18432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_193
timestamp 1679581782
transform 1 0 19104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_200
timestamp 1679581782
transform 1 0 19776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_207
timestamp 1679581782
transform 1 0 20448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_214
timestamp 1679581782
transform 1 0 21120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_221
timestamp 1679581782
transform 1 0 21792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_228
timestamp 1679581782
transform 1 0 22464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_235
timestamp 1679581782
transform 1 0 23136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_242
timestamp 1679581782
transform 1 0 23808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_249
timestamp 1679581782
transform 1 0 24480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_256
timestamp 1679581782
transform 1 0 25152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_263
timestamp 1679581782
transform 1 0 25824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_270
timestamp 1679581782
transform 1 0 26496 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_277
timestamp 1679581782
transform 1 0 27168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_284
timestamp 1679581782
transform 1 0 27840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_291
timestamp 1679581782
transform 1 0 28512 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_298
timestamp 1679581782
transform 1 0 29184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_305
timestamp 1679581782
transform 1 0 29856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_312
timestamp 1679581782
transform 1 0 30528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_319
timestamp 1679581782
transform 1 0 31200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_326
timestamp 1679581782
transform 1 0 31872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_333
timestamp 1679581782
transform 1 0 32544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_340
timestamp 1679581782
transform 1 0 33216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_347
timestamp 1679581782
transform 1 0 33888 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_354
timestamp 1679581782
transform 1 0 34560 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_361
timestamp 1679581782
transform 1 0 35232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_368
timestamp 1679581782
transform 1 0 35904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_375
timestamp 1679581782
transform 1 0 36576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_382
timestamp 1679581782
transform 1 0 37248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_389
timestamp 1679581782
transform 1 0 37920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_396
timestamp 1679581782
transform 1 0 38592 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_403
timestamp 1679581782
transform 1 0 39264 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_410
timestamp 1679581782
transform 1 0 39936 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_417
timestamp 1679581782
transform 1 0 40608 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_424
timestamp 1679581782
transform 1 0 41280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_431
timestamp 1679581782
transform 1 0 41952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_438
timestamp 1679581782
transform 1 0 42624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_445
timestamp 1679581782
transform 1 0 43296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_452
timestamp 1679581782
transform 1 0 43968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_459
timestamp 1679581782
transform 1 0 44640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_466
timestamp 1679581782
transform 1 0 45312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_473
timestamp 1679581782
transform 1 0 45984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_480
timestamp 1679581782
transform 1 0 46656 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_487
timestamp 1679581782
transform 1 0 47328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_494
timestamp 1679581782
transform 1 0 48000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_501
timestamp 1679581782
transform 1 0 48672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_508
timestamp 1679581782
transform 1 0 49344 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_515
timestamp 1679581782
transform 1 0 50016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_522
timestamp 1679581782
transform 1 0 50688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_529
timestamp 1679581782
transform 1 0 51360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_536
timestamp 1679581782
transform 1 0 52032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_543
timestamp 1679581782
transform 1 0 52704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_550
timestamp 1679581782
transform 1 0 53376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_557
timestamp 1679581782
transform 1 0 54048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_564
timestamp 1679581782
transform 1 0 54720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_571
timestamp 1679581782
transform 1 0 55392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_578
timestamp 1679581782
transform 1 0 56064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_585
timestamp 1679581782
transform 1 0 56736 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_592
timestamp 1679581782
transform 1 0 57408 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_599
timestamp 1679581782
transform 1 0 58080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_606
timestamp 1679581782
transform 1 0 58752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_613
timestamp 1679581782
transform 1 0 59424 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_620
timestamp 1679581782
transform 1 0 60096 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_627
timestamp 1679581782
transform 1 0 60768 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_634
timestamp 1679581782
transform 1 0 61440 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_641
timestamp 1679581782
transform 1 0 62112 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_648
timestamp 1679581782
transform 1 0 62784 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_655
timestamp 1679581782
transform 1 0 63456 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_662
timestamp 1679581782
transform 1 0 64128 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_669
timestamp 1679581782
transform 1 0 64800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_676
timestamp 1679581782
transform 1 0 65472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_683
timestamp 1679581782
transform 1 0 66144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_690
timestamp 1679581782
transform 1 0 66816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_697
timestamp 1679581782
transform 1 0 67488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_704
timestamp 1679581782
transform 1 0 68160 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_711
timestamp 1679581782
transform 1 0 68832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_718
timestamp 1679581782
transform 1 0 69504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_725
timestamp 1679581782
transform 1 0 70176 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_732
timestamp 1679581782
transform 1 0 70848 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_739
timestamp 1679581782
transform 1 0 71520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_746
timestamp 1679581782
transform 1 0 72192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_753
timestamp 1679581782
transform 1 0 72864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_760
timestamp 1679581782
transform 1 0 73536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_767
timestamp 1679581782
transform 1 0 74208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_774
timestamp 1679581782
transform 1 0 74880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_781
timestamp 1679581782
transform 1 0 75552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_788
timestamp 1679581782
transform 1 0 76224 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_795
timestamp 1679581782
transform 1 0 76896 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_802
timestamp 1679581782
transform 1 0 77568 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_809
timestamp 1679581782
transform 1 0 78240 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_816
timestamp 1679581782
transform 1 0 78912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_823
timestamp 1679581782
transform 1 0 79584 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_830
timestamp 1679581782
transform 1 0 80256 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_837
timestamp 1679581782
transform 1 0 80928 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_844
timestamp 1679581782
transform 1 0 81600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_851
timestamp 1679581782
transform 1 0 82272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_858
timestamp 1679581782
transform 1 0 82944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_865
timestamp 1679581782
transform 1 0 83616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_872
timestamp 1679581782
transform 1 0 84288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_879
timestamp 1679581782
transform 1 0 84960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_886
timestamp 1679581782
transform 1 0 85632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_893
timestamp 1679581782
transform 1 0 86304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_900
timestamp 1679581782
transform 1 0 86976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_907
timestamp 1679581782
transform 1 0 87648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_914
timestamp 1679581782
transform 1 0 88320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_921
timestamp 1679581782
transform 1 0 88992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_928
timestamp 1679581782
transform 1 0 89664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_935
timestamp 1679581782
transform 1 0 90336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_942
timestamp 1679581782
transform 1 0 91008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_949
timestamp 1679581782
transform 1 0 91680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_956
timestamp 1679581782
transform 1 0 92352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_963
timestamp 1679581782
transform 1 0 93024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_970
timestamp 1679581782
transform 1 0 93696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_977
timestamp 1679581782
transform 1 0 94368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_984
timestamp 1679581782
transform 1 0 95040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_991
timestamp 1679581782
transform 1 0 95712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_998
timestamp 1679581782
transform 1 0 96384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1005
timestamp 1679581782
transform 1 0 97056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1012
timestamp 1679581782
transform 1 0 97728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1019
timestamp 1679581782
transform 1 0 98400 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_1026
timestamp 1677580104
transform 1 0 99072 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_1028
timestamp 1677579658
transform 1 0 99264 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679581782
transform 1 0 2592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_28
timestamp 1679581782
transform 1 0 3264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_35
timestamp 1679581782
transform 1 0 3936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_42
timestamp 1679581782
transform 1 0 4608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_49
timestamp 1679581782
transform 1 0 5280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_56
timestamp 1679581782
transform 1 0 5952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_63
timestamp 1679581782
transform 1 0 6624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_70
timestamp 1679581782
transform 1 0 7296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_77
timestamp 1679581782
transform 1 0 7968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_84
timestamp 1679581782
transform 1 0 8640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_91
timestamp 1679581782
transform 1 0 9312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_98
timestamp 1679581782
transform 1 0 9984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_105
timestamp 1679581782
transform 1 0 10656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_112
timestamp 1679581782
transform 1 0 11328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_119
timestamp 1679581782
transform 1 0 12000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_126
timestamp 1679581782
transform 1 0 12672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_133
timestamp 1679581782
transform 1 0 13344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_140
timestamp 1679581782
transform 1 0 14016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_147
timestamp 1679581782
transform 1 0 14688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_154
timestamp 1679581782
transform 1 0 15360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_161
timestamp 1679581782
transform 1 0 16032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_168
timestamp 1679581782
transform 1 0 16704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_175
timestamp 1679581782
transform 1 0 17376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_182
timestamp 1679581782
transform 1 0 18048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_189
timestamp 1679581782
transform 1 0 18720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_196
timestamp 1679581782
transform 1 0 19392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_203
timestamp 1679581782
transform 1 0 20064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_210
timestamp 1679581782
transform 1 0 20736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_217
timestamp 1679581782
transform 1 0 21408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_224
timestamp 1679581782
transform 1 0 22080 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_231
timestamp 1679581782
transform 1 0 22752 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_238
timestamp 1679581782
transform 1 0 23424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_245
timestamp 1679581782
transform 1 0 24096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_252
timestamp 1679581782
transform 1 0 24768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_259
timestamp 1679581782
transform 1 0 25440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_266
timestamp 1679581782
transform 1 0 26112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_273
timestamp 1679581782
transform 1 0 26784 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_280
timestamp 1679581782
transform 1 0 27456 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_287
timestamp 1679581782
transform 1 0 28128 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_294
timestamp 1679581782
transform 1 0 28800 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_301
timestamp 1679581782
transform 1 0 29472 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_308
timestamp 1679581782
transform 1 0 30144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_315
timestamp 1679581782
transform 1 0 30816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_322
timestamp 1679581782
transform 1 0 31488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_329
timestamp 1679581782
transform 1 0 32160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_336
timestamp 1679581782
transform 1 0 32832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_343
timestamp 1679581782
transform 1 0 33504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_350
timestamp 1679581782
transform 1 0 34176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_357
timestamp 1679581782
transform 1 0 34848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_364
timestamp 1679581782
transform 1 0 35520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_371
timestamp 1679581782
transform 1 0 36192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_378
timestamp 1679581782
transform 1 0 36864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_385
timestamp 1679581782
transform 1 0 37536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_392
timestamp 1679581782
transform 1 0 38208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_399
timestamp 1679581782
transform 1 0 38880 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_406
timestamp 1679581782
transform 1 0 39552 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_413
timestamp 1679581782
transform 1 0 40224 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_420
timestamp 1679581782
transform 1 0 40896 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_427
timestamp 1679581782
transform 1 0 41568 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_434
timestamp 1679581782
transform 1 0 42240 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_441
timestamp 1679581782
transform 1 0 42912 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_448
timestamp 1679581782
transform 1 0 43584 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_455
timestamp 1679581782
transform 1 0 44256 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_462
timestamp 1679581782
transform 1 0 44928 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_469
timestamp 1679581782
transform 1 0 45600 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_476
timestamp 1679581782
transform 1 0 46272 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_483
timestamp 1679581782
transform 1 0 46944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_490
timestamp 1679581782
transform 1 0 47616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_497
timestamp 1679581782
transform 1 0 48288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_504
timestamp 1679581782
transform 1 0 48960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_511
timestamp 1679581782
transform 1 0 49632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_518
timestamp 1679581782
transform 1 0 50304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_525
timestamp 1679581782
transform 1 0 50976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_532
timestamp 1679581782
transform 1 0 51648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_539
timestamp 1679581782
transform 1 0 52320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_546
timestamp 1679581782
transform 1 0 52992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_553
timestamp 1679581782
transform 1 0 53664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_560
timestamp 1679581782
transform 1 0 54336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_567
timestamp 1679581782
transform 1 0 55008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_574
timestamp 1679581782
transform 1 0 55680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_581
timestamp 1679581782
transform 1 0 56352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_588
timestamp 1679581782
transform 1 0 57024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_595
timestamp 1679581782
transform 1 0 57696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_602
timestamp 1679581782
transform 1 0 58368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_609
timestamp 1679581782
transform 1 0 59040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_616
timestamp 1679581782
transform 1 0 59712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_623
timestamp 1679581782
transform 1 0 60384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_630
timestamp 1679581782
transform 1 0 61056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_637
timestamp 1679581782
transform 1 0 61728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_644
timestamp 1679581782
transform 1 0 62400 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_651
timestamp 1679581782
transform 1 0 63072 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_658
timestamp 1679581782
transform 1 0 63744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_665
timestamp 1679581782
transform 1 0 64416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_672
timestamp 1679581782
transform 1 0 65088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_679
timestamp 1679581782
transform 1 0 65760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_686
timestamp 1679581782
transform 1 0 66432 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_693
timestamp 1679581782
transform 1 0 67104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_700
timestamp 1679581782
transform 1 0 67776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_707
timestamp 1679581782
transform 1 0 68448 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_714
timestamp 1679581782
transform 1 0 69120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_721
timestamp 1679581782
transform 1 0 69792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_728
timestamp 1679581782
transform 1 0 70464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_735
timestamp 1679581782
transform 1 0 71136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_742
timestamp 1679581782
transform 1 0 71808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_749
timestamp 1679581782
transform 1 0 72480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_756
timestamp 1679581782
transform 1 0 73152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_763
timestamp 1679581782
transform 1 0 73824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_770
timestamp 1679581782
transform 1 0 74496 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_777
timestamp 1679577901
transform 1 0 75168 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_781
timestamp 1677579658
transform 1 0 75552 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_785
timestamp 1679577901
transform 1 0 75936 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_789
timestamp 1677580104
transform 1 0 76320 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_27_795
timestamp 1679577901
transform 1 0 76896 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_799
timestamp 1677580104
transform 1 0 77280 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_804
timestamp 1679581782
transform 1 0 77760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_811
timestamp 1679577901
transform 1 0 78432 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_27_823
timestamp 1679581782
transform 1 0 79584 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_830
timestamp 1679577901
transform 1 0 80256 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_834
timestamp 1677579658
transform 1 0 80640 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_839
timestamp 1679581782
transform 1 0 81120 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_846
timestamp 1677580104
transform 1 0 81792 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_848
timestamp 1677579658
transform 1 0 81984 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_856
timestamp 1679577901
transform 1 0 82752 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_860
timestamp 1677580104
transform 1 0 83136 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_27_866
timestamp 1679577901
transform 1 0 83712 0 -1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_27_874
timestamp 1679581782
transform 1 0 84480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_881
timestamp 1679581782
transform 1 0 85152 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_891
timestamp 1677580104
transform 1 0 86112 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_896
timestamp 1677579658
transform 1 0 86592 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_900
timestamp 1679581782
transform 1 0 86976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_907
timestamp 1679581782
transform 1 0 87648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_914
timestamp 1679581782
transform 1 0 88320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_928
timestamp 1679581782
transform 1 0 89664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_935
timestamp 1679581782
transform 1 0 90336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_945
timestamp 1679581782
transform 1 0 91296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_952
timestamp 1679581782
transform 1 0 91968 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_962
timestamp 1677580104
transform 1 0 92928 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_964
timestamp 1677579658
transform 1 0 93120 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_968
timestamp 1679581782
transform 1 0 93504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_975
timestamp 1679581782
transform 1 0 94176 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_982
timestamp 1677580104
transform 1 0 94848 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_984
timestamp 1677579658
transform 1 0 95040 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_988
timestamp 1679581782
transform 1 0 95424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_995
timestamp 1679581782
transform 1 0 96096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1002
timestamp 1679581782
transform 1 0 96768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1009
timestamp 1679581782
transform 1 0 97440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1016
timestamp 1679581782
transform 1 0 98112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_1023
timestamp 1679577901
transform 1 0 98784 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_1027
timestamp 1677580104
transform 1 0 99168 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679581782
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679581782
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679581782
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_25
timestamp 1679581782
transform 1 0 2976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_32
timestamp 1679581782
transform 1 0 3648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_39
timestamp 1679581782
transform 1 0 4320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_46
timestamp 1679581782
transform 1 0 4992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_53
timestamp 1679581782
transform 1 0 5664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_60
timestamp 1679581782
transform 1 0 6336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_67
timestamp 1679581782
transform 1 0 7008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_74
timestamp 1679581782
transform 1 0 7680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_81
timestamp 1679581782
transform 1 0 8352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_88
timestamp 1679581782
transform 1 0 9024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_95
timestamp 1679581782
transform 1 0 9696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_102
timestamp 1679581782
transform 1 0 10368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_109
timestamp 1679581782
transform 1 0 11040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_116
timestamp 1679581782
transform 1 0 11712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_123
timestamp 1679581782
transform 1 0 12384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_130
timestamp 1679581782
transform 1 0 13056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_137
timestamp 1679581782
transform 1 0 13728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_144
timestamp 1679581782
transform 1 0 14400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_151
timestamp 1679581782
transform 1 0 15072 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_158
timestamp 1679581782
transform 1 0 15744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_165
timestamp 1679581782
transform 1 0 16416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_172
timestamp 1679581782
transform 1 0 17088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_179
timestamp 1679581782
transform 1 0 17760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_186
timestamp 1679581782
transform 1 0 18432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_193
timestamp 1679581782
transform 1 0 19104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_200
timestamp 1679581782
transform 1 0 19776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_207
timestamp 1679581782
transform 1 0 20448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_214
timestamp 1679581782
transform 1 0 21120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_221
timestamp 1679581782
transform 1 0 21792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_228
timestamp 1679581782
transform 1 0 22464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_235
timestamp 1679581782
transform 1 0 23136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_242
timestamp 1679581782
transform 1 0 23808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_249
timestamp 1679581782
transform 1 0 24480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_256
timestamp 1679581782
transform 1 0 25152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_263
timestamp 1679581782
transform 1 0 25824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_270
timestamp 1679581782
transform 1 0 26496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_277
timestamp 1679581782
transform 1 0 27168 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_284
timestamp 1679581782
transform 1 0 27840 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_291
timestamp 1679581782
transform 1 0 28512 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_298
timestamp 1679581782
transform 1 0 29184 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_305
timestamp 1679581782
transform 1 0 29856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_312
timestamp 1679581782
transform 1 0 30528 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_319
timestamp 1679581782
transform 1 0 31200 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_326
timestamp 1679581782
transform 1 0 31872 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_333
timestamp 1679581782
transform 1 0 32544 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_340
timestamp 1679581782
transform 1 0 33216 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_347
timestamp 1679581782
transform 1 0 33888 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_354
timestamp 1679581782
transform 1 0 34560 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_361
timestamp 1679581782
transform 1 0 35232 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_368
timestamp 1679581782
transform 1 0 35904 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_375
timestamp 1679581782
transform 1 0 36576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_382
timestamp 1679581782
transform 1 0 37248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_389
timestamp 1679581782
transform 1 0 37920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_396
timestamp 1679581782
transform 1 0 38592 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_403
timestamp 1679581782
transform 1 0 39264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_410
timestamp 1679581782
transform 1 0 39936 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_417
timestamp 1679581782
transform 1 0 40608 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_424
timestamp 1679581782
transform 1 0 41280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_431
timestamp 1679581782
transform 1 0 41952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_438
timestamp 1679581782
transform 1 0 42624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_445
timestamp 1679581782
transform 1 0 43296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_452
timestamp 1679581782
transform 1 0 43968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_459
timestamp 1679581782
transform 1 0 44640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_466
timestamp 1679581782
transform 1 0 45312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_473
timestamp 1679581782
transform 1 0 45984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_480
timestamp 1679581782
transform 1 0 46656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_487
timestamp 1679581782
transform 1 0 47328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_494
timestamp 1679581782
transform 1 0 48000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_501
timestamp 1679581782
transform 1 0 48672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_508
timestamp 1679581782
transform 1 0 49344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_515
timestamp 1679581782
transform 1 0 50016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_522
timestamp 1679581782
transform 1 0 50688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_529
timestamp 1679581782
transform 1 0 51360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_536
timestamp 1679581782
transform 1 0 52032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_543
timestamp 1679581782
transform 1 0 52704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_550
timestamp 1679581782
transform 1 0 53376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_557
timestamp 1679581782
transform 1 0 54048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_564
timestamp 1679581782
transform 1 0 54720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_571
timestamp 1679581782
transform 1 0 55392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_578
timestamp 1679581782
transform 1 0 56064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_585
timestamp 1679581782
transform 1 0 56736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_592
timestamp 1679581782
transform 1 0 57408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_599
timestamp 1679581782
transform 1 0 58080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_606
timestamp 1679581782
transform 1 0 58752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_613
timestamp 1679581782
transform 1 0 59424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_620
timestamp 1679581782
transform 1 0 60096 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_627
timestamp 1679581782
transform 1 0 60768 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_634
timestamp 1679581782
transform 1 0 61440 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_641
timestamp 1679581782
transform 1 0 62112 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_648
timestamp 1679581782
transform 1 0 62784 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_655
timestamp 1679581782
transform 1 0 63456 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_662
timestamp 1679581782
transform 1 0 64128 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_669
timestamp 1679581782
transform 1 0 64800 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_676
timestamp 1679581782
transform 1 0 65472 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_683
timestamp 1679581782
transform 1 0 66144 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_690
timestamp 1679581782
transform 1 0 66816 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_697
timestamp 1679581782
transform 1 0 67488 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_704
timestamp 1679581782
transform 1 0 68160 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_711
timestamp 1679581782
transform 1 0 68832 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_718
timestamp 1679581782
transform 1 0 69504 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_725
timestamp 1679581782
transform 1 0 70176 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_732
timestamp 1679581782
transform 1 0 70848 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_739
timestamp 1679581782
transform 1 0 71520 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_746
timestamp 1679581782
transform 1 0 72192 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_753
timestamp 1679581782
transform 1 0 72864 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_760
timestamp 1677580104
transform 1 0 73536 0 1 21924
box -48 -56 240 834
use sg13g2_decap_4  FILLER_28_765
timestamp 1679577901
transform 1 0 74016 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_769
timestamp 1677579658
transform 1 0 74400 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_774
timestamp 1677579658
transform 1 0 74880 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_790
timestamp 1677579658
transform 1 0 76416 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_794
timestamp 1677580104
transform 1 0 76800 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_796
timestamp 1677579658
transform 1 0 76992 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_800
timestamp 1677580104
transform 1 0 77376 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_802
timestamp 1677579658
transform 1 0 77568 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_811
timestamp 1677580104
transform 1 0 78432 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_813
timestamp 1677579658
transform 1 0 78624 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_817
timestamp 1679577901
transform 1 0 79008 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_821
timestamp 1677579658
transform 1 0 79392 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_830
timestamp 1677579658
transform 1 0 80256 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_838
timestamp 1677580104
transform 1 0 81024 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_848
timestamp 1679581782
transform 1 0 81984 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_855
timestamp 1677580104
transform 1 0 82656 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_857
timestamp 1677579658
transform 1 0 82848 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_862
timestamp 1677579658
transform 1 0 83328 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_873
timestamp 1677579658
transform 1 0 84384 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_882
timestamp 1677579658
transform 1 0 85248 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_918
timestamp 1677579658
transform 1 0 88704 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_923
timestamp 1679577901
transform 1 0 89184 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_927
timestamp 1677579658
transform 1 0 89568 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_932
timestamp 1677579658
transform 1 0 90048 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_964
timestamp 1677580104
transform 1 0 93120 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_966
timestamp 1677579658
transform 1 0 93312 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_981
timestamp 1677579658
transform 1 0 94752 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_998
timestamp 1677579658
transform 1 0 96384 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_1003
timestamp 1677579658
transform 1 0 96864 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_1008
timestamp 1677580104
transform 1 0 97344 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_1018
timestamp 1679581782
transform 1 0 98304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_28_1025
timestamp 1679577901
transform 1 0 98976 0 1 21924
box -48 -56 432 834
use sg13g2_decap_8  FILLER_29_5
timestamp 1679581782
transform 1 0 1056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_12
timestamp 1679581782
transform 1 0 1728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_19
timestamp 1679581782
transform 1 0 2400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_26
timestamp 1679581782
transform 1 0 3072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_33
timestamp 1679581782
transform 1 0 3744 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_40
timestamp 1679581782
transform 1 0 4416 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_47
timestamp 1679581782
transform 1 0 5088 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_54
timestamp 1679581782
transform 1 0 5760 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_61
timestamp 1679581782
transform 1 0 6432 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_68
timestamp 1679581782
transform 1 0 7104 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_75
timestamp 1679581782
transform 1 0 7776 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_82
timestamp 1679581782
transform 1 0 8448 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_89
timestamp 1679581782
transform 1 0 9120 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_96
timestamp 1679581782
transform 1 0 9792 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_103
timestamp 1679581782
transform 1 0 10464 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_110
timestamp 1679581782
transform 1 0 11136 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_117
timestamp 1679581782
transform 1 0 11808 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_124
timestamp 1679581782
transform 1 0 12480 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_131
timestamp 1679581782
transform 1 0 13152 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_138
timestamp 1679581782
transform 1 0 13824 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_145
timestamp 1679581782
transform 1 0 14496 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_152
timestamp 1679581782
transform 1 0 15168 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_159
timestamp 1679581782
transform 1 0 15840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_166
timestamp 1679581782
transform 1 0 16512 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_173
timestamp 1679581782
transform 1 0 17184 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_180
timestamp 1679581782
transform 1 0 17856 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_187
timestamp 1679581782
transform 1 0 18528 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_194
timestamp 1679581782
transform 1 0 19200 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_201
timestamp 1679581782
transform 1 0 19872 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_208
timestamp 1679581782
transform 1 0 20544 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_215
timestamp 1679581782
transform 1 0 21216 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_222
timestamp 1679581782
transform 1 0 21888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_229
timestamp 1679581782
transform 1 0 22560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_236
timestamp 1679581782
transform 1 0 23232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_243
timestamp 1679581782
transform 1 0 23904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_250
timestamp 1679581782
transform 1 0 24576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_257
timestamp 1679581782
transform 1 0 25248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_264
timestamp 1679581782
transform 1 0 25920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_271
timestamp 1679581782
transform 1 0 26592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_278
timestamp 1679581782
transform 1 0 27264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_285
timestamp 1679581782
transform 1 0 27936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_292
timestamp 1679581782
transform 1 0 28608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_299
timestamp 1679581782
transform 1 0 29280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_306
timestamp 1679581782
transform 1 0 29952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_313
timestamp 1679581782
transform 1 0 30624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_320
timestamp 1679581782
transform 1 0 31296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_327
timestamp 1679581782
transform 1 0 31968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_334
timestamp 1679581782
transform 1 0 32640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_341
timestamp 1679581782
transform 1 0 33312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_348
timestamp 1679581782
transform 1 0 33984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_355
timestamp 1679581782
transform 1 0 34656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_362
timestamp 1679581782
transform 1 0 35328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_369
timestamp 1679581782
transform 1 0 36000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_376
timestamp 1679581782
transform 1 0 36672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_383
timestamp 1679581782
transform 1 0 37344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_390
timestamp 1679581782
transform 1 0 38016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_397
timestamp 1679581782
transform 1 0 38688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_404
timestamp 1679581782
transform 1 0 39360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_411
timestamp 1679581782
transform 1 0 40032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_418
timestamp 1679581782
transform 1 0 40704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_425
timestamp 1679581782
transform 1 0 41376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_432
timestamp 1679581782
transform 1 0 42048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_439
timestamp 1679581782
transform 1 0 42720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_446
timestamp 1679581782
transform 1 0 43392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_453
timestamp 1679581782
transform 1 0 44064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_460
timestamp 1679581782
transform 1 0 44736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_467
timestamp 1679581782
transform 1 0 45408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_474
timestamp 1679581782
transform 1 0 46080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_481
timestamp 1679581782
transform 1 0 46752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_488
timestamp 1679581782
transform 1 0 47424 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_495
timestamp 1679581782
transform 1 0 48096 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_502
timestamp 1679581782
transform 1 0 48768 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_509
timestamp 1679581782
transform 1 0 49440 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_516
timestamp 1679581782
transform 1 0 50112 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_523
timestamp 1679581782
transform 1 0 50784 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_530
timestamp 1679581782
transform 1 0 51456 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_537
timestamp 1679581782
transform 1 0 52128 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_544
timestamp 1679581782
transform 1 0 52800 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_551
timestamp 1679581782
transform 1 0 53472 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_558
timestamp 1679581782
transform 1 0 54144 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_565
timestamp 1679581782
transform 1 0 54816 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_572
timestamp 1679581782
transform 1 0 55488 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_579
timestamp 1679581782
transform 1 0 56160 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_586
timestamp 1679581782
transform 1 0 56832 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_593
timestamp 1679581782
transform 1 0 57504 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_600
timestamp 1679581782
transform 1 0 58176 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_607
timestamp 1679581782
transform 1 0 58848 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_614
timestamp 1679581782
transform 1 0 59520 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_621
timestamp 1679581782
transform 1 0 60192 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_628
timestamp 1679581782
transform 1 0 60864 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_635
timestamp 1679581782
transform 1 0 61536 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_642
timestamp 1679581782
transform 1 0 62208 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_649
timestamp 1679581782
transform 1 0 62880 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_656
timestamp 1679581782
transform 1 0 63552 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_663
timestamp 1679581782
transform 1 0 64224 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_670
timestamp 1679581782
transform 1 0 64896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_677
timestamp 1679581782
transform 1 0 65568 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_684
timestamp 1679581782
transform 1 0 66240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_691
timestamp 1679581782
transform 1 0 66912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_698
timestamp 1679581782
transform 1 0 67584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_705
timestamp 1679581782
transform 1 0 68256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_712
timestamp 1679581782
transform 1 0 68928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_719
timestamp 1679581782
transform 1 0 69600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_726
timestamp 1679581782
transform 1 0 70272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_733
timestamp 1679581782
transform 1 0 70944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_740
timestamp 1679581782
transform 1 0 71616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_747
timestamp 1679581782
transform 1 0 72288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_29_760
timestamp 1679577901
transform 1 0 73536 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_764
timestamp 1677579658
transform 1 0 73920 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_792
timestamp 1677580104
transform 1 0 76608 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_809
timestamp 1677579658
transform 1 0 78240 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_851
timestamp 1677579658
transform 1 0 82272 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_871
timestamp 1677579658
transform 1 0 84192 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_875
timestamp 1677579658
transform 1 0 84576 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_879
timestamp 1677579658
transform 1 0 84960 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_913
timestamp 1677579658
transform 1 0 88224 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_917
timestamp 1677579658
transform 1 0 88608 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_921
timestamp 1677580104
transform 1 0 88992 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_923
timestamp 1677579658
transform 1 0 89184 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_960
timestamp 1677579658
transform 1 0 92736 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_975
timestamp 1677580104
transform 1 0 94176 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_984
timestamp 1677580104
transform 1 0 95040 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_1010
timestamp 1677579658
transform 1 0 97536 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_1014
timestamp 1677579658
transform 1 0 97920 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_1018
timestamp 1677579658
transform 1 0 98304 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_1026
timestamp 1677580104
transform 1 0 99072 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_1028
timestamp 1677579658
transform 1 0 99264 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_5
timestamp 1679581782
transform 1 0 1056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_12
timestamp 1679581782
transform 1 0 1728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_19
timestamp 1679581782
transform 1 0 2400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_26
timestamp 1679581782
transform 1 0 3072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_33
timestamp 1679581782
transform 1 0 3744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_40
timestamp 1679581782
transform 1 0 4416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_47
timestamp 1679581782
transform 1 0 5088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_54
timestamp 1679581782
transform 1 0 5760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_61
timestamp 1679581782
transform 1 0 6432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_68
timestamp 1679581782
transform 1 0 7104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_75
timestamp 1679581782
transform 1 0 7776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_82
timestamp 1679581782
transform 1 0 8448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_89
timestamp 1679581782
transform 1 0 9120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_96
timestamp 1679581782
transform 1 0 9792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_103
timestamp 1679581782
transform 1 0 10464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_110
timestamp 1679581782
transform 1 0 11136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_117
timestamp 1679581782
transform 1 0 11808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_124
timestamp 1679581782
transform 1 0 12480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_131
timestamp 1679581782
transform 1 0 13152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_138
timestamp 1679581782
transform 1 0 13824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_145
timestamp 1679581782
transform 1 0 14496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_152
timestamp 1679581782
transform 1 0 15168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_159
timestamp 1679581782
transform 1 0 15840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_166
timestamp 1679581782
transform 1 0 16512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_173
timestamp 1679581782
transform 1 0 17184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_180
timestamp 1679581782
transform 1 0 17856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_187
timestamp 1679581782
transform 1 0 18528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_194
timestamp 1679581782
transform 1 0 19200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_201
timestamp 1679581782
transform 1 0 19872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_208
timestamp 1679581782
transform 1 0 20544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_215
timestamp 1679581782
transform 1 0 21216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_222
timestamp 1679581782
transform 1 0 21888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_229
timestamp 1679581782
transform 1 0 22560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_236
timestamp 1679581782
transform 1 0 23232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_243
timestamp 1679581782
transform 1 0 23904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_250
timestamp 1679581782
transform 1 0 24576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_257
timestamp 1679581782
transform 1 0 25248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_264
timestamp 1679581782
transform 1 0 25920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_271
timestamp 1679581782
transform 1 0 26592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_278
timestamp 1679581782
transform 1 0 27264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_285
timestamp 1679581782
transform 1 0 27936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_292
timestamp 1679581782
transform 1 0 28608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_299
timestamp 1679581782
transform 1 0 29280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_306
timestamp 1679581782
transform 1 0 29952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_313
timestamp 1679581782
transform 1 0 30624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_320
timestamp 1679581782
transform 1 0 31296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_327
timestamp 1679581782
transform 1 0 31968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_334
timestamp 1679581782
transform 1 0 32640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_341
timestamp 1679581782
transform 1 0 33312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_348
timestamp 1679581782
transform 1 0 33984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_355
timestamp 1679581782
transform 1 0 34656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_362
timestamp 1679581782
transform 1 0 35328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_369
timestamp 1679581782
transform 1 0 36000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_376
timestamp 1679581782
transform 1 0 36672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_383
timestamp 1679581782
transform 1 0 37344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_390
timestamp 1679581782
transform 1 0 38016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_397
timestamp 1679581782
transform 1 0 38688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_404
timestamp 1679581782
transform 1 0 39360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_411
timestamp 1679581782
transform 1 0 40032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_418
timestamp 1679581782
transform 1 0 40704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_425
timestamp 1679581782
transform 1 0 41376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_432
timestamp 1679581782
transform 1 0 42048 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_439
timestamp 1679581782
transform 1 0 42720 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_446
timestamp 1679581782
transform 1 0 43392 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_453
timestamp 1679581782
transform 1 0 44064 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_460
timestamp 1679581782
transform 1 0 44736 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_467
timestamp 1679581782
transform 1 0 45408 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_474
timestamp 1679581782
transform 1 0 46080 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_481
timestamp 1679581782
transform 1 0 46752 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_488
timestamp 1679581782
transform 1 0 47424 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_495
timestamp 1679581782
transform 1 0 48096 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_502
timestamp 1679581782
transform 1 0 48768 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_509
timestamp 1679581782
transform 1 0 49440 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_516
timestamp 1679581782
transform 1 0 50112 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_523
timestamp 1679581782
transform 1 0 50784 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_530
timestamp 1679581782
transform 1 0 51456 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_537
timestamp 1679581782
transform 1 0 52128 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_544
timestamp 1679581782
transform 1 0 52800 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_551
timestamp 1679581782
transform 1 0 53472 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_558
timestamp 1679581782
transform 1 0 54144 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_565
timestamp 1679581782
transform 1 0 54816 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_572
timestamp 1679581782
transform 1 0 55488 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_579
timestamp 1679581782
transform 1 0 56160 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_586
timestamp 1679581782
transform 1 0 56832 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_593
timestamp 1679581782
transform 1 0 57504 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_600
timestamp 1679581782
transform 1 0 58176 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_607
timestamp 1679581782
transform 1 0 58848 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_614
timestamp 1679581782
transform 1 0 59520 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_621
timestamp 1679581782
transform 1 0 60192 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_628
timestamp 1679581782
transform 1 0 60864 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_635
timestamp 1679581782
transform 1 0 61536 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_642
timestamp 1679581782
transform 1 0 62208 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_649
timestamp 1679581782
transform 1 0 62880 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_656
timestamp 1679581782
transform 1 0 63552 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_663
timestamp 1679581782
transform 1 0 64224 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_670
timestamp 1679581782
transform 1 0 64896 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_677
timestamp 1679581782
transform 1 0 65568 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_684
timestamp 1679581782
transform 1 0 66240 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_691
timestamp 1679581782
transform 1 0 66912 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_698
timestamp 1679581782
transform 1 0 67584 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_705
timestamp 1679581782
transform 1 0 68256 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_712
timestamp 1679581782
transform 1 0 68928 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_719
timestamp 1679577901
transform 1 0 69600 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_31_5
timestamp 1679581782
transform 1 0 1056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_12
timestamp 1679581782
transform 1 0 1728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_19
timestamp 1679581782
transform 1 0 2400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_26
timestamp 1679581782
transform 1 0 3072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_33
timestamp 1679581782
transform 1 0 3744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_40
timestamp 1679581782
transform 1 0 4416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_47
timestamp 1679581782
transform 1 0 5088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_54
timestamp 1679581782
transform 1 0 5760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_61
timestamp 1679581782
transform 1 0 6432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_68
timestamp 1679581782
transform 1 0 7104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_75
timestamp 1679581782
transform 1 0 7776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_82
timestamp 1679581782
transform 1 0 8448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_89
timestamp 1679581782
transform 1 0 9120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_96
timestamp 1679581782
transform 1 0 9792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_103
timestamp 1679581782
transform 1 0 10464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_110
timestamp 1679581782
transform 1 0 11136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_117
timestamp 1679581782
transform 1 0 11808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_124
timestamp 1679581782
transform 1 0 12480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_131
timestamp 1679581782
transform 1 0 13152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_138
timestamp 1679581782
transform 1 0 13824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_145
timestamp 1679581782
transform 1 0 14496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_152
timestamp 1679581782
transform 1 0 15168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_159
timestamp 1679581782
transform 1 0 15840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_166
timestamp 1679581782
transform 1 0 16512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_173
timestamp 1679581782
transform 1 0 17184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_180
timestamp 1679581782
transform 1 0 17856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_187
timestamp 1679581782
transform 1 0 18528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_194
timestamp 1679581782
transform 1 0 19200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_201
timestamp 1679581782
transform 1 0 19872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_208
timestamp 1679581782
transform 1 0 20544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_215
timestamp 1679581782
transform 1 0 21216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_222
timestamp 1679581782
transform 1 0 21888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_229
timestamp 1679581782
transform 1 0 22560 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_236
timestamp 1679581782
transform 1 0 23232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_243
timestamp 1679581782
transform 1 0 23904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_250
timestamp 1679581782
transform 1 0 24576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_257
timestamp 1679581782
transform 1 0 25248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_264
timestamp 1679581782
transform 1 0 25920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_271
timestamp 1679581782
transform 1 0 26592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_278
timestamp 1679581782
transform 1 0 27264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_285
timestamp 1679581782
transform 1 0 27936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_292
timestamp 1679581782
transform 1 0 28608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_299
timestamp 1679581782
transform 1 0 29280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_306
timestamp 1679581782
transform 1 0 29952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_313
timestamp 1679581782
transform 1 0 30624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_320
timestamp 1679581782
transform 1 0 31296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_327
timestamp 1679581782
transform 1 0 31968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_334
timestamp 1679581782
transform 1 0 32640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_341
timestamp 1679581782
transform 1 0 33312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_348
timestamp 1679581782
transform 1 0 33984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_355
timestamp 1679581782
transform 1 0 34656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_362
timestamp 1679581782
transform 1 0 35328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_369
timestamp 1679581782
transform 1 0 36000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_376
timestamp 1679581782
transform 1 0 36672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_383
timestamp 1679581782
transform 1 0 37344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_390
timestamp 1679581782
transform 1 0 38016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_397
timestamp 1679581782
transform 1 0 38688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_404
timestamp 1679581782
transform 1 0 39360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_411
timestamp 1679581782
transform 1 0 40032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_418
timestamp 1679581782
transform 1 0 40704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_425
timestamp 1679581782
transform 1 0 41376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_432
timestamp 1679581782
transform 1 0 42048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_439
timestamp 1679581782
transform 1 0 42720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_446
timestamp 1679581782
transform 1 0 43392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_453
timestamp 1679581782
transform 1 0 44064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_460
timestamp 1679581782
transform 1 0 44736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_467
timestamp 1679581782
transform 1 0 45408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_474
timestamp 1679581782
transform 1 0 46080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_481
timestamp 1679581782
transform 1 0 46752 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_488
timestamp 1679581782
transform 1 0 47424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_495
timestamp 1679581782
transform 1 0 48096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_502
timestamp 1679581782
transform 1 0 48768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_509
timestamp 1679581782
transform 1 0 49440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_516
timestamp 1679581782
transform 1 0 50112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_523
timestamp 1679581782
transform 1 0 50784 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_530
timestamp 1679581782
transform 1 0 51456 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_537
timestamp 1679581782
transform 1 0 52128 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_544
timestamp 1679581782
transform 1 0 52800 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_551
timestamp 1679581782
transform 1 0 53472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_558
timestamp 1679581782
transform 1 0 54144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_565
timestamp 1679581782
transform 1 0 54816 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_572
timestamp 1679581782
transform 1 0 55488 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_579
timestamp 1679581782
transform 1 0 56160 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_586
timestamp 1679581782
transform 1 0 56832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_593
timestamp 1679581782
transform 1 0 57504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_600
timestamp 1679581782
transform 1 0 58176 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_607
timestamp 1679581782
transform 1 0 58848 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_614
timestamp 1679581782
transform 1 0 59520 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_621
timestamp 1679581782
transform 1 0 60192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_628
timestamp 1679581782
transform 1 0 60864 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_635
timestamp 1679581782
transform 1 0 61536 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_642
timestamp 1679581782
transform 1 0 62208 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_649
timestamp 1679581782
transform 1 0 62880 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_656
timestamp 1679581782
transform 1 0 63552 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_663
timestamp 1679581782
transform 1 0 64224 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_670
timestamp 1679581782
transform 1 0 64896 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_677
timestamp 1679581782
transform 1 0 65568 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_684
timestamp 1679581782
transform 1 0 66240 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_691
timestamp 1679581782
transform 1 0 66912 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_698
timestamp 1679581782
transform 1 0 67584 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_705
timestamp 1679581782
transform 1 0 68256 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_712
timestamp 1679581782
transform 1 0 68928 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_4  FILLER_31_719
timestamp 1679577901
transform 1 0 69600 0 -1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_32_5
timestamp 1679581782
transform 1 0 1056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_12
timestamp 1679581782
transform 1 0 1728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_19
timestamp 1679581782
transform 1 0 2400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_26
timestamp 1679581782
transform 1 0 3072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_33
timestamp 1679581782
transform 1 0 3744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_40
timestamp 1679581782
transform 1 0 4416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_47
timestamp 1679581782
transform 1 0 5088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_54
timestamp 1679581782
transform 1 0 5760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_61
timestamp 1679581782
transform 1 0 6432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_68
timestamp 1679581782
transform 1 0 7104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_75
timestamp 1679581782
transform 1 0 7776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_82
timestamp 1679581782
transform 1 0 8448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_89
timestamp 1679581782
transform 1 0 9120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_96
timestamp 1679581782
transform 1 0 9792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_103
timestamp 1679581782
transform 1 0 10464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_110
timestamp 1679581782
transform 1 0 11136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_117
timestamp 1679581782
transform 1 0 11808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_124
timestamp 1679581782
transform 1 0 12480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_131
timestamp 1679581782
transform 1 0 13152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_138
timestamp 1679581782
transform 1 0 13824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_145
timestamp 1679581782
transform 1 0 14496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_152
timestamp 1679581782
transform 1 0 15168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_159
timestamp 1679581782
transform 1 0 15840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_166
timestamp 1679581782
transform 1 0 16512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_173
timestamp 1679581782
transform 1 0 17184 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_180
timestamp 1679581782
transform 1 0 17856 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_187
timestamp 1679581782
transform 1 0 18528 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_194
timestamp 1679581782
transform 1 0 19200 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_201
timestamp 1679581782
transform 1 0 19872 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_208
timestamp 1679581782
transform 1 0 20544 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_215
timestamp 1679581782
transform 1 0 21216 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_222
timestamp 1679581782
transform 1 0 21888 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_229
timestamp 1679581782
transform 1 0 22560 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_236
timestamp 1679581782
transform 1 0 23232 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_243
timestamp 1679581782
transform 1 0 23904 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_250
timestamp 1679581782
transform 1 0 24576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_257
timestamp 1679581782
transform 1 0 25248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_264
timestamp 1679581782
transform 1 0 25920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_271
timestamp 1679581782
transform 1 0 26592 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_278
timestamp 1679581782
transform 1 0 27264 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_285
timestamp 1679581782
transform 1 0 27936 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_292
timestamp 1679581782
transform 1 0 28608 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_299
timestamp 1679581782
transform 1 0 29280 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_306
timestamp 1679581782
transform 1 0 29952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_313
timestamp 1679581782
transform 1 0 30624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_320
timestamp 1679581782
transform 1 0 31296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_327
timestamp 1679581782
transform 1 0 31968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_334
timestamp 1679581782
transform 1 0 32640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_341
timestamp 1679581782
transform 1 0 33312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_348
timestamp 1679581782
transform 1 0 33984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_355
timestamp 1679581782
transform 1 0 34656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_362
timestamp 1679581782
transform 1 0 35328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_369
timestamp 1679581782
transform 1 0 36000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_376
timestamp 1679581782
transform 1 0 36672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_383
timestamp 1679581782
transform 1 0 37344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_390
timestamp 1679581782
transform 1 0 38016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_397
timestamp 1679581782
transform 1 0 38688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_404
timestamp 1679581782
transform 1 0 39360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_411
timestamp 1679581782
transform 1 0 40032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_418
timestamp 1679581782
transform 1 0 40704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_425
timestamp 1679581782
transform 1 0 41376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_432
timestamp 1679581782
transform 1 0 42048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_439
timestamp 1679581782
transform 1 0 42720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_446
timestamp 1679581782
transform 1 0 43392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_453
timestamp 1679581782
transform 1 0 44064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_460
timestamp 1679581782
transform 1 0 44736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_467
timestamp 1679581782
transform 1 0 45408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_474
timestamp 1679581782
transform 1 0 46080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_481
timestamp 1679581782
transform 1 0 46752 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_488
timestamp 1679581782
transform 1 0 47424 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_495
timestamp 1679581782
transform 1 0 48096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_502
timestamp 1679581782
transform 1 0 48768 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_509
timestamp 1679581782
transform 1 0 49440 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_516
timestamp 1679581782
transform 1 0 50112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_523
timestamp 1679581782
transform 1 0 50784 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_530
timestamp 1679581782
transform 1 0 51456 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_537
timestamp 1679581782
transform 1 0 52128 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_544
timestamp 1679581782
transform 1 0 52800 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_551
timestamp 1679581782
transform 1 0 53472 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_558
timestamp 1679581782
transform 1 0 54144 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_565
timestamp 1679581782
transform 1 0 54816 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_572
timestamp 1679581782
transform 1 0 55488 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_579
timestamp 1679581782
transform 1 0 56160 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_586
timestamp 1679581782
transform 1 0 56832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_593
timestamp 1679581782
transform 1 0 57504 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_600
timestamp 1679581782
transform 1 0 58176 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_607
timestamp 1679581782
transform 1 0 58848 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_614
timestamp 1679581782
transform 1 0 59520 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_621
timestamp 1679581782
transform 1 0 60192 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_628
timestamp 1679581782
transform 1 0 60864 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_635
timestamp 1679581782
transform 1 0 61536 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_642
timestamp 1679581782
transform 1 0 62208 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_649
timestamp 1679581782
transform 1 0 62880 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_656
timestamp 1679581782
transform 1 0 63552 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_663
timestamp 1679581782
transform 1 0 64224 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_670
timestamp 1679581782
transform 1 0 64896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_677
timestamp 1679581782
transform 1 0 65568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_684
timestamp 1679581782
transform 1 0 66240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_691
timestamp 1679581782
transform 1 0 66912 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_698
timestamp 1679581782
transform 1 0 67584 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_705
timestamp 1677580104
transform 1 0 68256 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_707
timestamp 1677579658
transform 1 0 68448 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_712
timestamp 1677580104
transform 1 0 68928 0 1 24948
box -48 -56 240 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679581782
transform 1 0 576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1679581782
transform 1 0 1248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1679581782
transform 1 0 1920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_21
timestamp 1679581782
transform 1 0 2592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_28
timestamp 1679581782
transform 1 0 3264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_35
timestamp 1679581782
transform 1 0 3936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_42
timestamp 1679581782
transform 1 0 4608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_49
timestamp 1679581782
transform 1 0 5280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_56
timestamp 1679581782
transform 1 0 5952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_63
timestamp 1679581782
transform 1 0 6624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_70
timestamp 1679581782
transform 1 0 7296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_77
timestamp 1679581782
transform 1 0 7968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_84
timestamp 1679581782
transform 1 0 8640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_91
timestamp 1679581782
transform 1 0 9312 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_98
timestamp 1679581782
transform 1 0 9984 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_105
timestamp 1679581782
transform 1 0 10656 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_112
timestamp 1679581782
transform 1 0 11328 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_119
timestamp 1679581782
transform 1 0 12000 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_126
timestamp 1679581782
transform 1 0 12672 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_133
timestamp 1679581782
transform 1 0 13344 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_140
timestamp 1679581782
transform 1 0 14016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_147
timestamp 1679581782
transform 1 0 14688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_154
timestamp 1679581782
transform 1 0 15360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_161
timestamp 1679581782
transform 1 0 16032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_168
timestamp 1679581782
transform 1 0 16704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_175
timestamp 1679581782
transform 1 0 17376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_182
timestamp 1679581782
transform 1 0 18048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_189
timestamp 1679581782
transform 1 0 18720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_196
timestamp 1679581782
transform 1 0 19392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_203
timestamp 1679581782
transform 1 0 20064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_210
timestamp 1679581782
transform 1 0 20736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_217
timestamp 1679581782
transform 1 0 21408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_224
timestamp 1679581782
transform 1 0 22080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_231
timestamp 1679581782
transform 1 0 22752 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_238
timestamp 1679581782
transform 1 0 23424 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_245
timestamp 1679581782
transform 1 0 24096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_252
timestamp 1679581782
transform 1 0 24768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_259
timestamp 1679581782
transform 1 0 25440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_266
timestamp 1679581782
transform 1 0 26112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_273
timestamp 1679581782
transform 1 0 26784 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_280
timestamp 1679581782
transform 1 0 27456 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_287
timestamp 1679581782
transform 1 0 28128 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_294
timestamp 1679581782
transform 1 0 28800 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_301
timestamp 1679581782
transform 1 0 29472 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_308
timestamp 1679581782
transform 1 0 30144 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_315
timestamp 1679581782
transform 1 0 30816 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_322
timestamp 1679581782
transform 1 0 31488 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_329
timestamp 1679581782
transform 1 0 32160 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_336
timestamp 1679581782
transform 1 0 32832 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_343
timestamp 1679581782
transform 1 0 33504 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_350
timestamp 1679581782
transform 1 0 34176 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_357
timestamp 1679581782
transform 1 0 34848 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_364
timestamp 1679581782
transform 1 0 35520 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_371
timestamp 1679581782
transform 1 0 36192 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_378
timestamp 1679581782
transform 1 0 36864 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_385
timestamp 1679581782
transform 1 0 37536 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_392
timestamp 1679581782
transform 1 0 38208 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_399
timestamp 1679581782
transform 1 0 38880 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_406
timestamp 1679581782
transform 1 0 39552 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_413
timestamp 1679581782
transform 1 0 40224 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_420
timestamp 1679581782
transform 1 0 40896 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_427
timestamp 1679581782
transform 1 0 41568 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_434
timestamp 1679581782
transform 1 0 42240 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_441
timestamp 1679581782
transform 1 0 42912 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_448
timestamp 1679581782
transform 1 0 43584 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_455
timestamp 1679581782
transform 1 0 44256 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_462
timestamp 1679581782
transform 1 0 44928 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_469
timestamp 1679581782
transform 1 0 45600 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_476
timestamp 1679581782
transform 1 0 46272 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_483
timestamp 1679581782
transform 1 0 46944 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_490
timestamp 1679581782
transform 1 0 47616 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_497
timestamp 1679581782
transform 1 0 48288 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_504
timestamp 1679581782
transform 1 0 48960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_511
timestamp 1679581782
transform 1 0 49632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_518
timestamp 1679581782
transform 1 0 50304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_525
timestamp 1679581782
transform 1 0 50976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_532
timestamp 1679581782
transform 1 0 51648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_539
timestamp 1679581782
transform 1 0 52320 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_546
timestamp 1679581782
transform 1 0 52992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_553
timestamp 1679581782
transform 1 0 53664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_560
timestamp 1679581782
transform 1 0 54336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_567
timestamp 1679581782
transform 1 0 55008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_574
timestamp 1679581782
transform 1 0 55680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_581
timestamp 1679581782
transform 1 0 56352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_588
timestamp 1679581782
transform 1 0 57024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_595
timestamp 1679581782
transform 1 0 57696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_602
timestamp 1679581782
transform 1 0 58368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_609
timestamp 1679581782
transform 1 0 59040 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_616
timestamp 1679581782
transform 1 0 59712 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_623
timestamp 1679581782
transform 1 0 60384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_630
timestamp 1679581782
transform 1 0 61056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_637
timestamp 1679581782
transform 1 0 61728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_644
timestamp 1679581782
transform 1 0 62400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_651
timestamp 1679581782
transform 1 0 63072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_658
timestamp 1679581782
transform 1 0 63744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_665
timestamp 1679581782
transform 1 0 64416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_672
timestamp 1679581782
transform 1 0 65088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_679
timestamp 1679581782
transform 1 0 65760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_686
timestamp 1679581782
transform 1 0 66432 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_693
timestamp 1677580104
transform 1 0 67104 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_695
timestamp 1677579658
transform 1 0 67296 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_33_703
timestamp 1679577901
transform 1 0 68064 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679581782
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679581782
transform 1 0 1920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679581782
transform 1 0 2592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679581782
transform 1 0 3264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_35
timestamp 1679581782
transform 1 0 3936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_42
timestamp 1679581782
transform 1 0 4608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679581782
transform 1 0 5280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_56
timestamp 1679581782
transform 1 0 5952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_63
timestamp 1679581782
transform 1 0 6624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_70
timestamp 1679581782
transform 1 0 7296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_77
timestamp 1679581782
transform 1 0 7968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_84
timestamp 1679581782
transform 1 0 8640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_91
timestamp 1679581782
transform 1 0 9312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_98
timestamp 1679581782
transform 1 0 9984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_105
timestamp 1679581782
transform 1 0 10656 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_112
timestamp 1679581782
transform 1 0 11328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_119
timestamp 1679581782
transform 1 0 12000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_126
timestamp 1679581782
transform 1 0 12672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_133
timestamp 1679581782
transform 1 0 13344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_140
timestamp 1679581782
transform 1 0 14016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_147
timestamp 1679581782
transform 1 0 14688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_154
timestamp 1679581782
transform 1 0 15360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_161
timestamp 1679581782
transform 1 0 16032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_168
timestamp 1679581782
transform 1 0 16704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_175
timestamp 1679581782
transform 1 0 17376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_182
timestamp 1679581782
transform 1 0 18048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_189
timestamp 1679581782
transform 1 0 18720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_196
timestamp 1679581782
transform 1 0 19392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_203
timestamp 1679581782
transform 1 0 20064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_210
timestamp 1679581782
transform 1 0 20736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_217
timestamp 1679581782
transform 1 0 21408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_224
timestamp 1679581782
transform 1 0 22080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_231
timestamp 1679581782
transform 1 0 22752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_238
timestamp 1679581782
transform 1 0 23424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_245
timestamp 1679581782
transform 1 0 24096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_252
timestamp 1679581782
transform 1 0 24768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_259
timestamp 1679581782
transform 1 0 25440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_266
timestamp 1679581782
transform 1 0 26112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_273
timestamp 1679581782
transform 1 0 26784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_280
timestamp 1679581782
transform 1 0 27456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_287
timestamp 1679581782
transform 1 0 28128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_294
timestamp 1679581782
transform 1 0 28800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_301
timestamp 1679581782
transform 1 0 29472 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_308
timestamp 1679581782
transform 1 0 30144 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_315
timestamp 1679581782
transform 1 0 30816 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_322
timestamp 1679581782
transform 1 0 31488 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_329
timestamp 1679581782
transform 1 0 32160 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_336
timestamp 1679581782
transform 1 0 32832 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_343
timestamp 1679581782
transform 1 0 33504 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_350
timestamp 1679581782
transform 1 0 34176 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_357
timestamp 1679581782
transform 1 0 34848 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_364
timestamp 1679581782
transform 1 0 35520 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_371
timestamp 1679581782
transform 1 0 36192 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_378
timestamp 1679581782
transform 1 0 36864 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_385
timestamp 1679581782
transform 1 0 37536 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_392
timestamp 1679581782
transform 1 0 38208 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_399
timestamp 1679581782
transform 1 0 38880 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_406
timestamp 1679581782
transform 1 0 39552 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_413
timestamp 1679581782
transform 1 0 40224 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_420
timestamp 1679581782
transform 1 0 40896 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_427
timestamp 1679581782
transform 1 0 41568 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_434
timestamp 1679581782
transform 1 0 42240 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_441
timestamp 1679581782
transform 1 0 42912 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_448
timestamp 1679581782
transform 1 0 43584 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_455
timestamp 1679581782
transform 1 0 44256 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_462
timestamp 1679581782
transform 1 0 44928 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_469
timestamp 1679581782
transform 1 0 45600 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_476
timestamp 1679581782
transform 1 0 46272 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_483
timestamp 1679581782
transform 1 0 46944 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_490
timestamp 1679581782
transform 1 0 47616 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_497
timestamp 1679581782
transform 1 0 48288 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_504
timestamp 1679581782
transform 1 0 48960 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_511
timestamp 1679581782
transform 1 0 49632 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_518
timestamp 1679581782
transform 1 0 50304 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_525
timestamp 1679581782
transform 1 0 50976 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_532
timestamp 1679581782
transform 1 0 51648 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_539
timestamp 1679581782
transform 1 0 52320 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_546
timestamp 1679581782
transform 1 0 52992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_553
timestamp 1679581782
transform 1 0 53664 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_560
timestamp 1679581782
transform 1 0 54336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_567
timestamp 1679581782
transform 1 0 55008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_574
timestamp 1679581782
transform 1 0 55680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_581
timestamp 1679581782
transform 1 0 56352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_588
timestamp 1679581782
transform 1 0 57024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_595
timestamp 1679581782
transform 1 0 57696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_602
timestamp 1679581782
transform 1 0 58368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_609
timestamp 1679581782
transform 1 0 59040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_616
timestamp 1679581782
transform 1 0 59712 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_623
timestamp 1679581782
transform 1 0 60384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_630
timestamp 1679581782
transform 1 0 61056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_637
timestamp 1679581782
transform 1 0 61728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_644
timestamp 1679581782
transform 1 0 62400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_651
timestamp 1679581782
transform 1 0 63072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_658
timestamp 1679581782
transform 1 0 63744 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_665
timestamp 1679581782
transform 1 0 64416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_672
timestamp 1679581782
transform 1 0 65088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_679
timestamp 1679581782
transform 1 0 65760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_686
timestamp 1679581782
transform 1 0 66432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_693
timestamp 1679577901
transform 1 0 67104 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_697
timestamp 1677580104
transform 1 0 67488 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_34_707
timestamp 1679581782
transform 1 0 68448 0 1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_34_714
timestamp 1677580104
transform 1 0 69120 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_716
timestamp 1677579658
transform 1 0 69312 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_721
timestamp 1677580104
transform 1 0 69792 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679581782
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679581782
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679581782
transform 1 0 2592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_28
timestamp 1679581782
transform 1 0 3264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_35
timestamp 1679581782
transform 1 0 3936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_42
timestamp 1679581782
transform 1 0 4608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_49
timestamp 1679581782
transform 1 0 5280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_56
timestamp 1679581782
transform 1 0 5952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_63
timestamp 1679581782
transform 1 0 6624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_70
timestamp 1679581782
transform 1 0 7296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_77
timestamp 1679581782
transform 1 0 7968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_84
timestamp 1679581782
transform 1 0 8640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_91
timestamp 1679581782
transform 1 0 9312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_98
timestamp 1679581782
transform 1 0 9984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_105
timestamp 1679581782
transform 1 0 10656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_112
timestamp 1679581782
transform 1 0 11328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_119
timestamp 1679581782
transform 1 0 12000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_126
timestamp 1679581782
transform 1 0 12672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_133
timestamp 1679581782
transform 1 0 13344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_140
timestamp 1679581782
transform 1 0 14016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_147
timestamp 1679581782
transform 1 0 14688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_154
timestamp 1679581782
transform 1 0 15360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_161
timestamp 1679581782
transform 1 0 16032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_168
timestamp 1679581782
transform 1 0 16704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_175
timestamp 1679581782
transform 1 0 17376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_182
timestamp 1679581782
transform 1 0 18048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_189
timestamp 1679581782
transform 1 0 18720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_196
timestamp 1679581782
transform 1 0 19392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_203
timestamp 1679581782
transform 1 0 20064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_210
timestamp 1679581782
transform 1 0 20736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_217
timestamp 1679581782
transform 1 0 21408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_224
timestamp 1679581782
transform 1 0 22080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_231
timestamp 1679581782
transform 1 0 22752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_238
timestamp 1679581782
transform 1 0 23424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_245
timestamp 1679581782
transform 1 0 24096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_252
timestamp 1679581782
transform 1 0 24768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_259
timestamp 1679581782
transform 1 0 25440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_266
timestamp 1679581782
transform 1 0 26112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_273
timestamp 1679581782
transform 1 0 26784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_280
timestamp 1679581782
transform 1 0 27456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_287
timestamp 1679581782
transform 1 0 28128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_294
timestamp 1679581782
transform 1 0 28800 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_301
timestamp 1679581782
transform 1 0 29472 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_308
timestamp 1679581782
transform 1 0 30144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_315
timestamp 1679581782
transform 1 0 30816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_322
timestamp 1679581782
transform 1 0 31488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_329
timestamp 1679581782
transform 1 0 32160 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_336
timestamp 1679581782
transform 1 0 32832 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_343
timestamp 1679581782
transform 1 0 33504 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_350
timestamp 1679581782
transform 1 0 34176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_357
timestamp 1679581782
transform 1 0 34848 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_364
timestamp 1679581782
transform 1 0 35520 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_371
timestamp 1679581782
transform 1 0 36192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_378
timestamp 1679581782
transform 1 0 36864 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_385
timestamp 1679581782
transform 1 0 37536 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_392
timestamp 1679581782
transform 1 0 38208 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_399
timestamp 1679581782
transform 1 0 38880 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_406
timestamp 1679581782
transform 1 0 39552 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_413
timestamp 1679581782
transform 1 0 40224 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_420
timestamp 1679581782
transform 1 0 40896 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_427
timestamp 1679581782
transform 1 0 41568 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_434
timestamp 1679581782
transform 1 0 42240 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_441
timestamp 1679581782
transform 1 0 42912 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_448
timestamp 1679581782
transform 1 0 43584 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_455
timestamp 1679581782
transform 1 0 44256 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_462
timestamp 1679581782
transform 1 0 44928 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_469
timestamp 1679581782
transform 1 0 45600 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_476
timestamp 1679581782
transform 1 0 46272 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_483
timestamp 1679581782
transform 1 0 46944 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_490
timestamp 1679581782
transform 1 0 47616 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_497
timestamp 1679581782
transform 1 0 48288 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_504
timestamp 1679581782
transform 1 0 48960 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_511
timestamp 1679581782
transform 1 0 49632 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_518
timestamp 1679581782
transform 1 0 50304 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_525
timestamp 1679581782
transform 1 0 50976 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_532
timestamp 1679581782
transform 1 0 51648 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_539
timestamp 1679581782
transform 1 0 52320 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_546
timestamp 1679581782
transform 1 0 52992 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_553
timestamp 1679581782
transform 1 0 53664 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_560
timestamp 1679581782
transform 1 0 54336 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_567
timestamp 1679581782
transform 1 0 55008 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_574
timestamp 1679581782
transform 1 0 55680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_581
timestamp 1679581782
transform 1 0 56352 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_588
timestamp 1679581782
transform 1 0 57024 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_595
timestamp 1679581782
transform 1 0 57696 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_602
timestamp 1679581782
transform 1 0 58368 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_609
timestamp 1679581782
transform 1 0 59040 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_616
timestamp 1679581782
transform 1 0 59712 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_623
timestamp 1679581782
transform 1 0 60384 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_630
timestamp 1679581782
transform 1 0 61056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_637
timestamp 1679581782
transform 1 0 61728 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_644
timestamp 1679581782
transform 1 0 62400 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_651
timestamp 1679581782
transform 1 0 63072 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_658
timestamp 1679581782
transform 1 0 63744 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_665
timestamp 1679581782
transform 1 0 64416 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_672
timestamp 1679581782
transform 1 0 65088 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_679
timestamp 1679581782
transform 1 0 65760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_686
timestamp 1679581782
transform 1 0 66432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_693
timestamp 1679581782
transform 1 0 67104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_700
timestamp 1679581782
transform 1 0 67776 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_707
timestamp 1677580104
transform 1 0 68448 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_709
timestamp 1677579658
transform 1 0 68640 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_714
timestamp 1679581782
transform 1 0 69120 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_721
timestamp 1677580104
transform 1 0 69792 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679581782
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679581782
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679581782
transform 1 0 2592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679581782
transform 1 0 3264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679581782
transform 1 0 3936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679581782
transform 1 0 4608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679581782
transform 1 0 5280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_56
timestamp 1679581782
transform 1 0 5952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_63
timestamp 1679581782
transform 1 0 6624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_70
timestamp 1679581782
transform 1 0 7296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_77
timestamp 1679581782
transform 1 0 7968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_84
timestamp 1679581782
transform 1 0 8640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_91
timestamp 1679581782
transform 1 0 9312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_98
timestamp 1679581782
transform 1 0 9984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_105
timestamp 1679581782
transform 1 0 10656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_112
timestamp 1679581782
transform 1 0 11328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_119
timestamp 1679581782
transform 1 0 12000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679581782
transform 1 0 12672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_133
timestamp 1679581782
transform 1 0 13344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_140
timestamp 1679581782
transform 1 0 14016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_147
timestamp 1679581782
transform 1 0 14688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_154
timestamp 1679581782
transform 1 0 15360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_161
timestamp 1679581782
transform 1 0 16032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_168
timestamp 1679581782
transform 1 0 16704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_175
timestamp 1679581782
transform 1 0 17376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_182
timestamp 1679581782
transform 1 0 18048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_189
timestamp 1679581782
transform 1 0 18720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_196
timestamp 1679581782
transform 1 0 19392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_203
timestamp 1679581782
transform 1 0 20064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_210
timestamp 1679581782
transform 1 0 20736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_217
timestamp 1679581782
transform 1 0 21408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_224
timestamp 1679581782
transform 1 0 22080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_231
timestamp 1679581782
transform 1 0 22752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_238
timestamp 1679581782
transform 1 0 23424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_245
timestamp 1679581782
transform 1 0 24096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_252
timestamp 1679581782
transform 1 0 24768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_259
timestamp 1679581782
transform 1 0 25440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_266
timestamp 1679581782
transform 1 0 26112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_273
timestamp 1679581782
transform 1 0 26784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_280
timestamp 1679581782
transform 1 0 27456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_287
timestamp 1679581782
transform 1 0 28128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_294
timestamp 1679581782
transform 1 0 28800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_301
timestamp 1679581782
transform 1 0 29472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_308
timestamp 1679581782
transform 1 0 30144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_315
timestamp 1679581782
transform 1 0 30816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_322
timestamp 1679581782
transform 1 0 31488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_329
timestamp 1679581782
transform 1 0 32160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_336
timestamp 1679581782
transform 1 0 32832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_343
timestamp 1679581782
transform 1 0 33504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_350
timestamp 1679581782
transform 1 0 34176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_357
timestamp 1679581782
transform 1 0 34848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_364
timestamp 1679581782
transform 1 0 35520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_371
timestamp 1679581782
transform 1 0 36192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_378
timestamp 1679581782
transform 1 0 36864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_385
timestamp 1679581782
transform 1 0 37536 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_392
timestamp 1679581782
transform 1 0 38208 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_399
timestamp 1679581782
transform 1 0 38880 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_406
timestamp 1679581782
transform 1 0 39552 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_413
timestamp 1679581782
transform 1 0 40224 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_420
timestamp 1679581782
transform 1 0 40896 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_427
timestamp 1679581782
transform 1 0 41568 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_434
timestamp 1679581782
transform 1 0 42240 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_441
timestamp 1679581782
transform 1 0 42912 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_448
timestamp 1679581782
transform 1 0 43584 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_455
timestamp 1679581782
transform 1 0 44256 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_462
timestamp 1679581782
transform 1 0 44928 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_469
timestamp 1679581782
transform 1 0 45600 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_476
timestamp 1679581782
transform 1 0 46272 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_483
timestamp 1679581782
transform 1 0 46944 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_490
timestamp 1679581782
transform 1 0 47616 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_497
timestamp 1679581782
transform 1 0 48288 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_504
timestamp 1679581782
transform 1 0 48960 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_511
timestamp 1679581782
transform 1 0 49632 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_518
timestamp 1679581782
transform 1 0 50304 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_525
timestamp 1679581782
transform 1 0 50976 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_532
timestamp 1679581782
transform 1 0 51648 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_539
timestamp 1679581782
transform 1 0 52320 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_546
timestamp 1679581782
transform 1 0 52992 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_553
timestamp 1679581782
transform 1 0 53664 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_560
timestamp 1679581782
transform 1 0 54336 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_567
timestamp 1679581782
transform 1 0 55008 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_574
timestamp 1679581782
transform 1 0 55680 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_581
timestamp 1679581782
transform 1 0 56352 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_588
timestamp 1679581782
transform 1 0 57024 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_595
timestamp 1679581782
transform 1 0 57696 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_602
timestamp 1679581782
transform 1 0 58368 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_609
timestamp 1679581782
transform 1 0 59040 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_616
timestamp 1679581782
transform 1 0 59712 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_623
timestamp 1679581782
transform 1 0 60384 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_630
timestamp 1679581782
transform 1 0 61056 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_637
timestamp 1679581782
transform 1 0 61728 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_644
timestamp 1679581782
transform 1 0 62400 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_651
timestamp 1679581782
transform 1 0 63072 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_658
timestamp 1679581782
transform 1 0 63744 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_665
timestamp 1679581782
transform 1 0 64416 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_672
timestamp 1679581782
transform 1 0 65088 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_679
timestamp 1679581782
transform 1 0 65760 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_686
timestamp 1679581782
transform 1 0 66432 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_693
timestamp 1679581782
transform 1 0 67104 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_700
timestamp 1679581782
transform 1 0 67776 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_707
timestamp 1679581782
transform 1 0 68448 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_714
timestamp 1679581782
transform 1 0 69120 0 1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_36_721
timestamp 1677580104
transform 1 0 69792 0 1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679581782
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679581782
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679581782
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679581782
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679581782
transform 1 0 3936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679581782
transform 1 0 4608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679581782
transform 1 0 5280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679581782
transform 1 0 5952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679581782
transform 1 0 6624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_70
timestamp 1679581782
transform 1 0 7296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_77
timestamp 1679581782
transform 1 0 7968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_84
timestamp 1679581782
transform 1 0 8640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_91
timestamp 1679581782
transform 1 0 9312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679581782
transform 1 0 9984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679581782
transform 1 0 10656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679581782
transform 1 0 11328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679581782
transform 1 0 12000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679581782
transform 1 0 12672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679581782
transform 1 0 13344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679581782
transform 1 0 14016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_147
timestamp 1679581782
transform 1 0 14688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_154
timestamp 1679581782
transform 1 0 15360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_161
timestamp 1679581782
transform 1 0 16032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_168
timestamp 1679581782
transform 1 0 16704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_175
timestamp 1679581782
transform 1 0 17376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_182
timestamp 1679581782
transform 1 0 18048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_189
timestamp 1679581782
transform 1 0 18720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_196
timestamp 1679581782
transform 1 0 19392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_203
timestamp 1679581782
transform 1 0 20064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_210
timestamp 1679581782
transform 1 0 20736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_217
timestamp 1679581782
transform 1 0 21408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_224
timestamp 1679581782
transform 1 0 22080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_231
timestamp 1679581782
transform 1 0 22752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_238
timestamp 1679581782
transform 1 0 23424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_245
timestamp 1679581782
transform 1 0 24096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_252
timestamp 1679581782
transform 1 0 24768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_259
timestamp 1679581782
transform 1 0 25440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_266
timestamp 1679581782
transform 1 0 26112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_273
timestamp 1679581782
transform 1 0 26784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_280
timestamp 1679581782
transform 1 0 27456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_287
timestamp 1679581782
transform 1 0 28128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_294
timestamp 1679581782
transform 1 0 28800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_301
timestamp 1679581782
transform 1 0 29472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_308
timestamp 1679581782
transform 1 0 30144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_315
timestamp 1679581782
transform 1 0 30816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_322
timestamp 1679581782
transform 1 0 31488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_329
timestamp 1679581782
transform 1 0 32160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_336
timestamp 1679581782
transform 1 0 32832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_343
timestamp 1679581782
transform 1 0 33504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_350
timestamp 1679581782
transform 1 0 34176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_357
timestamp 1679581782
transform 1 0 34848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_364
timestamp 1679581782
transform 1 0 35520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_371
timestamp 1679581782
transform 1 0 36192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_378
timestamp 1679581782
transform 1 0 36864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_385
timestamp 1679581782
transform 1 0 37536 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_392
timestamp 1679581782
transform 1 0 38208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_399
timestamp 1679581782
transform 1 0 38880 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_406
timestamp 1679581782
transform 1 0 39552 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_413
timestamp 1679581782
transform 1 0 40224 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_420
timestamp 1679581782
transform 1 0 40896 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_427
timestamp 1679581782
transform 1 0 41568 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_434
timestamp 1679581782
transform 1 0 42240 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_441
timestamp 1679581782
transform 1 0 42912 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_448
timestamp 1679581782
transform 1 0 43584 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_455
timestamp 1679581782
transform 1 0 44256 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_462
timestamp 1679581782
transform 1 0 44928 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_469
timestamp 1679581782
transform 1 0 45600 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_476
timestamp 1679581782
transform 1 0 46272 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_483
timestamp 1679581782
transform 1 0 46944 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_490
timestamp 1679581782
transform 1 0 47616 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_497
timestamp 1679581782
transform 1 0 48288 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_504
timestamp 1679581782
transform 1 0 48960 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_511
timestamp 1679581782
transform 1 0 49632 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_518
timestamp 1679581782
transform 1 0 50304 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_525
timestamp 1679581782
transform 1 0 50976 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_532
timestamp 1679581782
transform 1 0 51648 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_539
timestamp 1679581782
transform 1 0 52320 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_546
timestamp 1679581782
transform 1 0 52992 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_553
timestamp 1679581782
transform 1 0 53664 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_560
timestamp 1679581782
transform 1 0 54336 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_567
timestamp 1679581782
transform 1 0 55008 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_574
timestamp 1679581782
transform 1 0 55680 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_581
timestamp 1679581782
transform 1 0 56352 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_588
timestamp 1679581782
transform 1 0 57024 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_595
timestamp 1679581782
transform 1 0 57696 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_602
timestamp 1679581782
transform 1 0 58368 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_609
timestamp 1679581782
transform 1 0 59040 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_616
timestamp 1679581782
transform 1 0 59712 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_623
timestamp 1679581782
transform 1 0 60384 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_630
timestamp 1679581782
transform 1 0 61056 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_637
timestamp 1679581782
transform 1 0 61728 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_644
timestamp 1679581782
transform 1 0 62400 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_651
timestamp 1679581782
transform 1 0 63072 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_658
timestamp 1679581782
transform 1 0 63744 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_665
timestamp 1679581782
transform 1 0 64416 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_672
timestamp 1679581782
transform 1 0 65088 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_679
timestamp 1679581782
transform 1 0 65760 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_686
timestamp 1679581782
transform 1 0 66432 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_693
timestamp 1679581782
transform 1 0 67104 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_700
timestamp 1679581782
transform 1 0 67776 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_707
timestamp 1679581782
transform 1 0 68448 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_714
timestamp 1679581782
transform 1 0 69120 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_721
timestamp 1677580104
transform 1 0 69792 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679581782
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679581782
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679581782
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679581782
transform 1 0 3264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679581782
transform 1 0 3936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679581782
transform 1 0 4608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679581782
transform 1 0 5280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_56
timestamp 1679581782
transform 1 0 5952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_63
timestamp 1679581782
transform 1 0 6624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_70
timestamp 1679581782
transform 1 0 7296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_77
timestamp 1679581782
transform 1 0 7968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_84
timestamp 1679581782
transform 1 0 8640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_91
timestamp 1679581782
transform 1 0 9312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_98
timestamp 1679581782
transform 1 0 9984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_105
timestamp 1679581782
transform 1 0 10656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_112
timestamp 1679581782
transform 1 0 11328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_119
timestamp 1679581782
transform 1 0 12000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_126
timestamp 1679581782
transform 1 0 12672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_133
timestamp 1679581782
transform 1 0 13344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_140
timestamp 1679581782
transform 1 0 14016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_147
timestamp 1679581782
transform 1 0 14688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_154
timestamp 1679581782
transform 1 0 15360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_161
timestamp 1679581782
transform 1 0 16032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_168
timestamp 1679581782
transform 1 0 16704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_175
timestamp 1679581782
transform 1 0 17376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_182
timestamp 1679581782
transform 1 0 18048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_189
timestamp 1679581782
transform 1 0 18720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_196
timestamp 1679581782
transform 1 0 19392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_203
timestamp 1679581782
transform 1 0 20064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_210
timestamp 1679581782
transform 1 0 20736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_217
timestamp 1679581782
transform 1 0 21408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_224
timestamp 1679581782
transform 1 0 22080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_231
timestamp 1679581782
transform 1 0 22752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_238
timestamp 1679581782
transform 1 0 23424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_245
timestamp 1679581782
transform 1 0 24096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_252
timestamp 1679581782
transform 1 0 24768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_259
timestamp 1679581782
transform 1 0 25440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_266
timestamp 1679581782
transform 1 0 26112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_273
timestamp 1679581782
transform 1 0 26784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_280
timestamp 1679581782
transform 1 0 27456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_287
timestamp 1679581782
transform 1 0 28128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_294
timestamp 1679581782
transform 1 0 28800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_301
timestamp 1679581782
transform 1 0 29472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_308
timestamp 1679581782
transform 1 0 30144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_315
timestamp 1679581782
transform 1 0 30816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_322
timestamp 1679581782
transform 1 0 31488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_329
timestamp 1679581782
transform 1 0 32160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_336
timestamp 1679581782
transform 1 0 32832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_343
timestamp 1679581782
transform 1 0 33504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_350
timestamp 1679581782
transform 1 0 34176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_357
timestamp 1679581782
transform 1 0 34848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_364
timestamp 1679581782
transform 1 0 35520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_371
timestamp 1679581782
transform 1 0 36192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_378
timestamp 1679581782
transform 1 0 36864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_385
timestamp 1679581782
transform 1 0 37536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_392
timestamp 1679581782
transform 1 0 38208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_399
timestamp 1679581782
transform 1 0 38880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_406
timestamp 1679581782
transform 1 0 39552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_413
timestamp 1679581782
transform 1 0 40224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_420
timestamp 1679581782
transform 1 0 40896 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_427
timestamp 1679581782
transform 1 0 41568 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_434
timestamp 1679581782
transform 1 0 42240 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_441
timestamp 1679581782
transform 1 0 42912 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_448
timestamp 1679581782
transform 1 0 43584 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_455
timestamp 1679581782
transform 1 0 44256 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_462
timestamp 1679581782
transform 1 0 44928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_469
timestamp 1679581782
transform 1 0 45600 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_476
timestamp 1679581782
transform 1 0 46272 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_483
timestamp 1679581782
transform 1 0 46944 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_490
timestamp 1679581782
transform 1 0 47616 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_497
timestamp 1679581782
transform 1 0 48288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_504
timestamp 1679581782
transform 1 0 48960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_511
timestamp 1679581782
transform 1 0 49632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_518
timestamp 1679581782
transform 1 0 50304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_525
timestamp 1679581782
transform 1 0 50976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_532
timestamp 1679581782
transform 1 0 51648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_539
timestamp 1679581782
transform 1 0 52320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_546
timestamp 1679581782
transform 1 0 52992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_553
timestamp 1679581782
transform 1 0 53664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_560
timestamp 1679581782
transform 1 0 54336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_567
timestamp 1679581782
transform 1 0 55008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_574
timestamp 1679581782
transform 1 0 55680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_581
timestamp 1679581782
transform 1 0 56352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_588
timestamp 1679581782
transform 1 0 57024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_595
timestamp 1679581782
transform 1 0 57696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_602
timestamp 1679581782
transform 1 0 58368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_609
timestamp 1679581782
transform 1 0 59040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_616
timestamp 1679581782
transform 1 0 59712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_623
timestamp 1679581782
transform 1 0 60384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_630
timestamp 1679581782
transform 1 0 61056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_637
timestamp 1679581782
transform 1 0 61728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_644
timestamp 1679581782
transform 1 0 62400 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_651
timestamp 1679581782
transform 1 0 63072 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_658
timestamp 1679581782
transform 1 0 63744 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_665
timestamp 1679581782
transform 1 0 64416 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_672
timestamp 1679581782
transform 1 0 65088 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_679
timestamp 1679581782
transform 1 0 65760 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_686
timestamp 1679581782
transform 1 0 66432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_693
timestamp 1679581782
transform 1 0 67104 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_700
timestamp 1679581782
transform 1 0 67776 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_707
timestamp 1679581782
transform 1 0 68448 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_714
timestamp 1679581782
transform 1 0 69120 0 1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_38_721
timestamp 1677580104
transform 1 0 69792 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679581782
transform 1 0 1248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679581782
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679581782
transform 1 0 2592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_28
timestamp 1679581782
transform 1 0 3264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_35
timestamp 1679581782
transform 1 0 3936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_42
timestamp 1679581782
transform 1 0 4608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_49
timestamp 1679581782
transform 1 0 5280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_56
timestamp 1679581782
transform 1 0 5952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_63
timestamp 1679581782
transform 1 0 6624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_70
timestamp 1679581782
transform 1 0 7296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_77
timestamp 1679581782
transform 1 0 7968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_84
timestamp 1679581782
transform 1 0 8640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_91
timestamp 1679581782
transform 1 0 9312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_98
timestamp 1679581782
transform 1 0 9984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_105
timestamp 1679581782
transform 1 0 10656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_112
timestamp 1679581782
transform 1 0 11328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_119
timestamp 1679581782
transform 1 0 12000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_126
timestamp 1679581782
transform 1 0 12672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_133
timestamp 1679581782
transform 1 0 13344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_140
timestamp 1679581782
transform 1 0 14016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_147
timestamp 1679581782
transform 1 0 14688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_154
timestamp 1679581782
transform 1 0 15360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_161
timestamp 1679581782
transform 1 0 16032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_168
timestamp 1679581782
transform 1 0 16704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_175
timestamp 1679581782
transform 1 0 17376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_182
timestamp 1679581782
transform 1 0 18048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_189
timestamp 1679581782
transform 1 0 18720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_196
timestamp 1679581782
transform 1 0 19392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_203
timestamp 1679581782
transform 1 0 20064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_210
timestamp 1679581782
transform 1 0 20736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_217
timestamp 1679581782
transform 1 0 21408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_224
timestamp 1679581782
transform 1 0 22080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_231
timestamp 1679581782
transform 1 0 22752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_238
timestamp 1679581782
transform 1 0 23424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_245
timestamp 1679581782
transform 1 0 24096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_252
timestamp 1679581782
transform 1 0 24768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_259
timestamp 1679581782
transform 1 0 25440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_266
timestamp 1679581782
transform 1 0 26112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_273
timestamp 1679581782
transform 1 0 26784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_280
timestamp 1679581782
transform 1 0 27456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_287
timestamp 1679581782
transform 1 0 28128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_294
timestamp 1679581782
transform 1 0 28800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_301
timestamp 1679581782
transform 1 0 29472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_308
timestamp 1679581782
transform 1 0 30144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_315
timestamp 1679581782
transform 1 0 30816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_322
timestamp 1679581782
transform 1 0 31488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_329
timestamp 1679581782
transform 1 0 32160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_336
timestamp 1679581782
transform 1 0 32832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_343
timestamp 1679581782
transform 1 0 33504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_350
timestamp 1679581782
transform 1 0 34176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_357
timestamp 1679581782
transform 1 0 34848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_364
timestamp 1679581782
transform 1 0 35520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_371
timestamp 1679581782
transform 1 0 36192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_378
timestamp 1679581782
transform 1 0 36864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_385
timestamp 1679581782
transform 1 0 37536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_392
timestamp 1679581782
transform 1 0 38208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_399
timestamp 1679581782
transform 1 0 38880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_406
timestamp 1679581782
transform 1 0 39552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_413
timestamp 1679581782
transform 1 0 40224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_420
timestamp 1679581782
transform 1 0 40896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_427
timestamp 1679581782
transform 1 0 41568 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_434
timestamp 1679581782
transform 1 0 42240 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_441
timestamp 1679581782
transform 1 0 42912 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_448
timestamp 1679581782
transform 1 0 43584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_455
timestamp 1679581782
transform 1 0 44256 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_462
timestamp 1679581782
transform 1 0 44928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_469
timestamp 1679581782
transform 1 0 45600 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_476
timestamp 1679581782
transform 1 0 46272 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_483
timestamp 1679581782
transform 1 0 46944 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_490
timestamp 1679581782
transform 1 0 47616 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_497
timestamp 1679581782
transform 1 0 48288 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_504
timestamp 1679581782
transform 1 0 48960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_511
timestamp 1679581782
transform 1 0 49632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_518
timestamp 1679581782
transform 1 0 50304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_525
timestamp 1679581782
transform 1 0 50976 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_532
timestamp 1679581782
transform 1 0 51648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_539
timestamp 1679581782
transform 1 0 52320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_546
timestamp 1679581782
transform 1 0 52992 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_553
timestamp 1679581782
transform 1 0 53664 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_560
timestamp 1679581782
transform 1 0 54336 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_567
timestamp 1679581782
transform 1 0 55008 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_574
timestamp 1679581782
transform 1 0 55680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_581
timestamp 1679581782
transform 1 0 56352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_588
timestamp 1679581782
transform 1 0 57024 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_595
timestamp 1679581782
transform 1 0 57696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_602
timestamp 1679581782
transform 1 0 58368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_609
timestamp 1679581782
transform 1 0 59040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_616
timestamp 1679581782
transform 1 0 59712 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_623
timestamp 1679581782
transform 1 0 60384 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_630
timestamp 1679581782
transform 1 0 61056 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_637
timestamp 1679581782
transform 1 0 61728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_644
timestamp 1679581782
transform 1 0 62400 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_651
timestamp 1679581782
transform 1 0 63072 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_658
timestamp 1679581782
transform 1 0 63744 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_665
timestamp 1679581782
transform 1 0 64416 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_672
timestamp 1679581782
transform 1 0 65088 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_679
timestamp 1679581782
transform 1 0 65760 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_686
timestamp 1679581782
transform 1 0 66432 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_693
timestamp 1677580104
transform 1 0 67104 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_39_699
timestamp 1679581782
transform 1 0 67680 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_706
timestamp 1677579658
transform 1 0 68352 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_710
timestamp 1677580104
transform 1 0 68736 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_721
timestamp 1677580104
transform 1 0 69792 0 -1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679581782
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679581782
transform 1 0 1920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679581782
transform 1 0 2592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_28
timestamp 1679581782
transform 1 0 3264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_35
timestamp 1679581782
transform 1 0 3936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_42
timestamp 1679581782
transform 1 0 4608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_49
timestamp 1679581782
transform 1 0 5280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_56
timestamp 1679581782
transform 1 0 5952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_63
timestamp 1679581782
transform 1 0 6624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_70
timestamp 1679581782
transform 1 0 7296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_77
timestamp 1679581782
transform 1 0 7968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_84
timestamp 1679581782
transform 1 0 8640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_91
timestamp 1679581782
transform 1 0 9312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_98
timestamp 1679581782
transform 1 0 9984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_105
timestamp 1679581782
transform 1 0 10656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_112
timestamp 1679581782
transform 1 0 11328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_119
timestamp 1679581782
transform 1 0 12000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_126
timestamp 1679581782
transform 1 0 12672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_133
timestamp 1679581782
transform 1 0 13344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_140
timestamp 1679581782
transform 1 0 14016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_147
timestamp 1679581782
transform 1 0 14688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_154
timestamp 1679581782
transform 1 0 15360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_161
timestamp 1679581782
transform 1 0 16032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_168
timestamp 1679581782
transform 1 0 16704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_175
timestamp 1679581782
transform 1 0 17376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_182
timestamp 1679581782
transform 1 0 18048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_189
timestamp 1679581782
transform 1 0 18720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_196
timestamp 1679581782
transform 1 0 19392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_203
timestamp 1679581782
transform 1 0 20064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_210
timestamp 1679581782
transform 1 0 20736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_217
timestamp 1679581782
transform 1 0 21408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_224
timestamp 1679581782
transform 1 0 22080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_231
timestamp 1679581782
transform 1 0 22752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_238
timestamp 1679581782
transform 1 0 23424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_245
timestamp 1679581782
transform 1 0 24096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_252
timestamp 1679581782
transform 1 0 24768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_259
timestamp 1679581782
transform 1 0 25440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_266
timestamp 1679581782
transform 1 0 26112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_273
timestamp 1679581782
transform 1 0 26784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_280
timestamp 1679581782
transform 1 0 27456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_287
timestamp 1679581782
transform 1 0 28128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_294
timestamp 1679581782
transform 1 0 28800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_301
timestamp 1679581782
transform 1 0 29472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_308
timestamp 1679581782
transform 1 0 30144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_315
timestamp 1679581782
transform 1 0 30816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_322
timestamp 1679581782
transform 1 0 31488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_329
timestamp 1679581782
transform 1 0 32160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_336
timestamp 1679581782
transform 1 0 32832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_343
timestamp 1679581782
transform 1 0 33504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_350
timestamp 1679581782
transform 1 0 34176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_357
timestamp 1679581782
transform 1 0 34848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_364
timestamp 1679581782
transform 1 0 35520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_371
timestamp 1679581782
transform 1 0 36192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_378
timestamp 1679581782
transform 1 0 36864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_385
timestamp 1679581782
transform 1 0 37536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_392
timestamp 1679581782
transform 1 0 38208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_399
timestamp 1679581782
transform 1 0 38880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_406
timestamp 1679581782
transform 1 0 39552 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_413
timestamp 1679581782
transform 1 0 40224 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_420
timestamp 1679581782
transform 1 0 40896 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_427
timestamp 1679581782
transform 1 0 41568 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_434
timestamp 1679581782
transform 1 0 42240 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_441
timestamp 1679581782
transform 1 0 42912 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_448
timestamp 1679581782
transform 1 0 43584 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_455
timestamp 1679581782
transform 1 0 44256 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_462
timestamp 1679581782
transform 1 0 44928 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_469
timestamp 1679581782
transform 1 0 45600 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_476
timestamp 1679581782
transform 1 0 46272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_483
timestamp 1679581782
transform 1 0 46944 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_490
timestamp 1679581782
transform 1 0 47616 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_497
timestamp 1679581782
transform 1 0 48288 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_504
timestamp 1679581782
transform 1 0 48960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_511
timestamp 1679581782
transform 1 0 49632 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_518
timestamp 1679581782
transform 1 0 50304 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_525
timestamp 1679581782
transform 1 0 50976 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_532
timestamp 1679581782
transform 1 0 51648 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_539
timestamp 1679581782
transform 1 0 52320 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_546
timestamp 1679581782
transform 1 0 52992 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_553
timestamp 1679581782
transform 1 0 53664 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_560
timestamp 1679581782
transform 1 0 54336 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_567
timestamp 1679581782
transform 1 0 55008 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_574
timestamp 1679581782
transform 1 0 55680 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_581
timestamp 1679581782
transform 1 0 56352 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_588
timestamp 1679581782
transform 1 0 57024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_595
timestamp 1679581782
transform 1 0 57696 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_602
timestamp 1679581782
transform 1 0 58368 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_609
timestamp 1679581782
transform 1 0 59040 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_616
timestamp 1679581782
transform 1 0 59712 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_623
timestamp 1679581782
transform 1 0 60384 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_630
timestamp 1679581782
transform 1 0 61056 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_637
timestamp 1679581782
transform 1 0 61728 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_644
timestamp 1679581782
transform 1 0 62400 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_651
timestamp 1679581782
transform 1 0 63072 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_658
timestamp 1679581782
transform 1 0 63744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_665
timestamp 1679581782
transform 1 0 64416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_672
timestamp 1679581782
transform 1 0 65088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_679
timestamp 1679581782
transform 1 0 65760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_686
timestamp 1679581782
transform 1 0 66432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_701
timestamp 1679581782
transform 1 0 67872 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679581782
transform 1 0 1248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679581782
transform 1 0 1920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679581782
transform 1 0 2592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679581782
transform 1 0 3264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679581782
transform 1 0 3936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679581782
transform 1 0 4608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679581782
transform 1 0 5280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679581782
transform 1 0 5952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_63
timestamp 1679581782
transform 1 0 6624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_70
timestamp 1679581782
transform 1 0 7296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_77
timestamp 1679581782
transform 1 0 7968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_84
timestamp 1679581782
transform 1 0 8640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_91
timestamp 1679581782
transform 1 0 9312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_98
timestamp 1679581782
transform 1 0 9984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_105
timestamp 1679581782
transform 1 0 10656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_112
timestamp 1679581782
transform 1 0 11328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_119
timestamp 1679581782
transform 1 0 12000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_126
timestamp 1679581782
transform 1 0 12672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_133
timestamp 1679581782
transform 1 0 13344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_140
timestamp 1679581782
transform 1 0 14016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_147
timestamp 1679581782
transform 1 0 14688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_154
timestamp 1679581782
transform 1 0 15360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679581782
transform 1 0 16032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_168
timestamp 1679581782
transform 1 0 16704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_175
timestamp 1679581782
transform 1 0 17376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_182
timestamp 1679581782
transform 1 0 18048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_189
timestamp 1679581782
transform 1 0 18720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_196
timestamp 1679581782
transform 1 0 19392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_203
timestamp 1679581782
transform 1 0 20064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_210
timestamp 1679581782
transform 1 0 20736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_217
timestamp 1679581782
transform 1 0 21408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_224
timestamp 1679581782
transform 1 0 22080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_231
timestamp 1679581782
transform 1 0 22752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_238
timestamp 1679581782
transform 1 0 23424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_245
timestamp 1679581782
transform 1 0 24096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_252
timestamp 1679581782
transform 1 0 24768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_259
timestamp 1679581782
transform 1 0 25440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_266
timestamp 1679581782
transform 1 0 26112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_273
timestamp 1679581782
transform 1 0 26784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_280
timestamp 1679581782
transform 1 0 27456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_287
timestamp 1679581782
transform 1 0 28128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_294
timestamp 1679581782
transform 1 0 28800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_301
timestamp 1679581782
transform 1 0 29472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_308
timestamp 1679581782
transform 1 0 30144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_315
timestamp 1679581782
transform 1 0 30816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_322
timestamp 1679581782
transform 1 0 31488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_329
timestamp 1679581782
transform 1 0 32160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_336
timestamp 1679581782
transform 1 0 32832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_343
timestamp 1679581782
transform 1 0 33504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_350
timestamp 1679581782
transform 1 0 34176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_357
timestamp 1679581782
transform 1 0 34848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_364
timestamp 1679581782
transform 1 0 35520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_371
timestamp 1679581782
transform 1 0 36192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_378
timestamp 1679581782
transform 1 0 36864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_385
timestamp 1679581782
transform 1 0 37536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_392
timestamp 1679581782
transform 1 0 38208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_399
timestamp 1679581782
transform 1 0 38880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_406
timestamp 1679581782
transform 1 0 39552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_413
timestamp 1679581782
transform 1 0 40224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_420
timestamp 1679581782
transform 1 0 40896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_427
timestamp 1679581782
transform 1 0 41568 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_434
timestamp 1679581782
transform 1 0 42240 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_441
timestamp 1679581782
transform 1 0 42912 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_448
timestamp 1679581782
transform 1 0 43584 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_455
timestamp 1679581782
transform 1 0 44256 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_462
timestamp 1679581782
transform 1 0 44928 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_469
timestamp 1679581782
transform 1 0 45600 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_476
timestamp 1679581782
transform 1 0 46272 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_483
timestamp 1679581782
transform 1 0 46944 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_490
timestamp 1679581782
transform 1 0 47616 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_497
timestamp 1679581782
transform 1 0 48288 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_504
timestamp 1679581782
transform 1 0 48960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_511
timestamp 1679581782
transform 1 0 49632 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_518
timestamp 1679581782
transform 1 0 50304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_525
timestamp 1679581782
transform 1 0 50976 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_532
timestamp 1679581782
transform 1 0 51648 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_539
timestamp 1679581782
transform 1 0 52320 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_546
timestamp 1679581782
transform 1 0 52992 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_553
timestamp 1679581782
transform 1 0 53664 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_560
timestamp 1679581782
transform 1 0 54336 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_567
timestamp 1679581782
transform 1 0 55008 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_574
timestamp 1679581782
transform 1 0 55680 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_581
timestamp 1679581782
transform 1 0 56352 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_588
timestamp 1679581782
transform 1 0 57024 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_595
timestamp 1679581782
transform 1 0 57696 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_602
timestamp 1679581782
transform 1 0 58368 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_609
timestamp 1679581782
transform 1 0 59040 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_616
timestamp 1679581782
transform 1 0 59712 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_623
timestamp 1679581782
transform 1 0 60384 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_630
timestamp 1679581782
transform 1 0 61056 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_637
timestamp 1679581782
transform 1 0 61728 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_644
timestamp 1679581782
transform 1 0 62400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_651
timestamp 1679581782
transform 1 0 63072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_658
timestamp 1679581782
transform 1 0 63744 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_665
timestamp 1679581782
transform 1 0 64416 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_672
timestamp 1679581782
transform 1 0 65088 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_679
timestamp 1679581782
transform 1 0 65760 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_686
timestamp 1679581782
transform 1 0 66432 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_693
timestamp 1679581782
transform 1 0 67104 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_700
timestamp 1679581782
transform 1 0 67776 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_707
timestamp 1679581782
transform 1 0 68448 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_41_714
timestamp 1679577901
transform 1 0 69120 0 -1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_41_718
timestamp 1677580104
transform 1 0 69504 0 -1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679581782
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679581782
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679581782
transform 1 0 3264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679581782
transform 1 0 3936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679581782
transform 1 0 4608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_49
timestamp 1679581782
transform 1 0 5280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_56
timestamp 1679581782
transform 1 0 5952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_63
timestamp 1679581782
transform 1 0 6624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_70
timestamp 1679581782
transform 1 0 7296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_77
timestamp 1679581782
transform 1 0 7968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_84
timestamp 1679581782
transform 1 0 8640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_91
timestamp 1679581782
transform 1 0 9312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_98
timestamp 1679581782
transform 1 0 9984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_105
timestamp 1679581782
transform 1 0 10656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_112
timestamp 1679581782
transform 1 0 11328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_119
timestamp 1679581782
transform 1 0 12000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_126
timestamp 1679581782
transform 1 0 12672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_133
timestamp 1679581782
transform 1 0 13344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_140
timestamp 1679581782
transform 1 0 14016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_147
timestamp 1679581782
transform 1 0 14688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_154
timestamp 1679581782
transform 1 0 15360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_161
timestamp 1679581782
transform 1 0 16032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_168
timestamp 1679581782
transform 1 0 16704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_175
timestamp 1679581782
transform 1 0 17376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_182
timestamp 1679581782
transform 1 0 18048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_189
timestamp 1679581782
transform 1 0 18720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_196
timestamp 1679581782
transform 1 0 19392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_203
timestamp 1679581782
transform 1 0 20064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_210
timestamp 1679581782
transform 1 0 20736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_217
timestamp 1679581782
transform 1 0 21408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_224
timestamp 1679581782
transform 1 0 22080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_231
timestamp 1679581782
transform 1 0 22752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_238
timestamp 1679581782
transform 1 0 23424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_245
timestamp 1679581782
transform 1 0 24096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_252
timestamp 1679581782
transform 1 0 24768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_259
timestamp 1679581782
transform 1 0 25440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_266
timestamp 1679581782
transform 1 0 26112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_273
timestamp 1679581782
transform 1 0 26784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_280
timestamp 1679581782
transform 1 0 27456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_287
timestamp 1679581782
transform 1 0 28128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_294
timestamp 1679581782
transform 1 0 28800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_301
timestamp 1679581782
transform 1 0 29472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_308
timestamp 1679581782
transform 1 0 30144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_315
timestamp 1679581782
transform 1 0 30816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_322
timestamp 1679581782
transform 1 0 31488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_329
timestamp 1679581782
transform 1 0 32160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_336
timestamp 1679581782
transform 1 0 32832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_343
timestamp 1679581782
transform 1 0 33504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_350
timestamp 1679581782
transform 1 0 34176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_357
timestamp 1679581782
transform 1 0 34848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_364
timestamp 1679581782
transform 1 0 35520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_371
timestamp 1679581782
transform 1 0 36192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_378
timestamp 1679581782
transform 1 0 36864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_385
timestamp 1679581782
transform 1 0 37536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_392
timestamp 1679581782
transform 1 0 38208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_399
timestamp 1679581782
transform 1 0 38880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_406
timestamp 1679581782
transform 1 0 39552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_413
timestamp 1679581782
transform 1 0 40224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_420
timestamp 1679581782
transform 1 0 40896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_427
timestamp 1679581782
transform 1 0 41568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_434
timestamp 1679581782
transform 1 0 42240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_441
timestamp 1679581782
transform 1 0 42912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_448
timestamp 1679581782
transform 1 0 43584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_455
timestamp 1679581782
transform 1 0 44256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_462
timestamp 1679581782
transform 1 0 44928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_469
timestamp 1679581782
transform 1 0 45600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_476
timestamp 1679581782
transform 1 0 46272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_483
timestamp 1679581782
transform 1 0 46944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_490
timestamp 1679581782
transform 1 0 47616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_497
timestamp 1679581782
transform 1 0 48288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_504
timestamp 1679581782
transform 1 0 48960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_511
timestamp 1679581782
transform 1 0 49632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_518
timestamp 1679581782
transform 1 0 50304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_525
timestamp 1679581782
transform 1 0 50976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_532
timestamp 1679581782
transform 1 0 51648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_539
timestamp 1679581782
transform 1 0 52320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_546
timestamp 1679581782
transform 1 0 52992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_553
timestamp 1679581782
transform 1 0 53664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_560
timestamp 1679581782
transform 1 0 54336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_567
timestamp 1679581782
transform 1 0 55008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_574
timestamp 1679581782
transform 1 0 55680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_581
timestamp 1679581782
transform 1 0 56352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_588
timestamp 1679581782
transform 1 0 57024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_595
timestamp 1679581782
transform 1 0 57696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_602
timestamp 1679581782
transform 1 0 58368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_609
timestamp 1679581782
transform 1 0 59040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_616
timestamp 1679581782
transform 1 0 59712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_623
timestamp 1679581782
transform 1 0 60384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_630
timestamp 1679581782
transform 1 0 61056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_637
timestamp 1679581782
transform 1 0 61728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_644
timestamp 1679581782
transform 1 0 62400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_651
timestamp 1679581782
transform 1 0 63072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_658
timestamp 1679581782
transform 1 0 63744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_665
timestamp 1679581782
transform 1 0 64416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_672
timestamp 1679581782
transform 1 0 65088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_679
timestamp 1679581782
transform 1 0 65760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_686
timestamp 1679581782
transform 1 0 66432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_693
timestamp 1679581782
transform 1 0 67104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_700
timestamp 1679581782
transform 1 0 67776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_707
timestamp 1679581782
transform 1 0 68448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_714
timestamp 1679581782
transform 1 0 69120 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_721
timestamp 1677580104
transform 1 0 69792 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679581782
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679581782
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679581782
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679581782
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679581782
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679581782
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679581782
transform 1 0 5952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679581782
transform 1 0 6624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679581782
transform 1 0 7296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679581782
transform 1 0 7968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679581782
transform 1 0 8640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679581782
transform 1 0 9312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679581782
transform 1 0 9984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679581782
transform 1 0 10656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_112
timestamp 1679581782
transform 1 0 11328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_119
timestamp 1679581782
transform 1 0 12000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_126
timestamp 1679581782
transform 1 0 12672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_133
timestamp 1679581782
transform 1 0 13344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_140
timestamp 1679581782
transform 1 0 14016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_147
timestamp 1679581782
transform 1 0 14688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_154
timestamp 1679581782
transform 1 0 15360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_161
timestamp 1679581782
transform 1 0 16032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_168
timestamp 1679581782
transform 1 0 16704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_175
timestamp 1679581782
transform 1 0 17376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_182
timestamp 1679581782
transform 1 0 18048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_189
timestamp 1679581782
transform 1 0 18720 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_196
timestamp 1679581782
transform 1 0 19392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_203
timestamp 1679581782
transform 1 0 20064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_210
timestamp 1679581782
transform 1 0 20736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_217
timestamp 1679581782
transform 1 0 21408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_224
timestamp 1679581782
transform 1 0 22080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_231
timestamp 1679581782
transform 1 0 22752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_238
timestamp 1679581782
transform 1 0 23424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_245
timestamp 1679581782
transform 1 0 24096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_252
timestamp 1679581782
transform 1 0 24768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_259
timestamp 1679581782
transform 1 0 25440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_266
timestamp 1679581782
transform 1 0 26112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_273
timestamp 1679581782
transform 1 0 26784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_280
timestamp 1679581782
transform 1 0 27456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_287
timestamp 1679581782
transform 1 0 28128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_294
timestamp 1679581782
transform 1 0 28800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_301
timestamp 1679581782
transform 1 0 29472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_308
timestamp 1679581782
transform 1 0 30144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_315
timestamp 1679581782
transform 1 0 30816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_322
timestamp 1679581782
transform 1 0 31488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_329
timestamp 1679581782
transform 1 0 32160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_336
timestamp 1679581782
transform 1 0 32832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_343
timestamp 1679581782
transform 1 0 33504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_350
timestamp 1679581782
transform 1 0 34176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_357
timestamp 1679581782
transform 1 0 34848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_364
timestamp 1679581782
transform 1 0 35520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_371
timestamp 1679581782
transform 1 0 36192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_378
timestamp 1679581782
transform 1 0 36864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_385
timestamp 1679581782
transform 1 0 37536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_392
timestamp 1679581782
transform 1 0 38208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_399
timestamp 1679581782
transform 1 0 38880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_406
timestamp 1679581782
transform 1 0 39552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_413
timestamp 1679581782
transform 1 0 40224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_420
timestamp 1679581782
transform 1 0 40896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_427
timestamp 1679581782
transform 1 0 41568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_434
timestamp 1679581782
transform 1 0 42240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_441
timestamp 1679581782
transform 1 0 42912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_448
timestamp 1679581782
transform 1 0 43584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_455
timestamp 1679581782
transform 1 0 44256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_462
timestamp 1679581782
transform 1 0 44928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_469
timestamp 1679581782
transform 1 0 45600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_476
timestamp 1679581782
transform 1 0 46272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_483
timestamp 1679581782
transform 1 0 46944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_490
timestamp 1679581782
transform 1 0 47616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_497
timestamp 1679581782
transform 1 0 48288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_504
timestamp 1679581782
transform 1 0 48960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_511
timestamp 1679581782
transform 1 0 49632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_518
timestamp 1679581782
transform 1 0 50304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_525
timestamp 1679581782
transform 1 0 50976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_532
timestamp 1679581782
transform 1 0 51648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_539
timestamp 1679581782
transform 1 0 52320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_546
timestamp 1679581782
transform 1 0 52992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_553
timestamp 1679581782
transform 1 0 53664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_560
timestamp 1679581782
transform 1 0 54336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_567
timestamp 1679581782
transform 1 0 55008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_574
timestamp 1679581782
transform 1 0 55680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_581
timestamp 1679581782
transform 1 0 56352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_588
timestamp 1679581782
transform 1 0 57024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_595
timestamp 1679581782
transform 1 0 57696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_602
timestamp 1679581782
transform 1 0 58368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_609
timestamp 1679581782
transform 1 0 59040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_616
timestamp 1679581782
transform 1 0 59712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_623
timestamp 1679581782
transform 1 0 60384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_630
timestamp 1679581782
transform 1 0 61056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_637
timestamp 1679581782
transform 1 0 61728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_644
timestamp 1679581782
transform 1 0 62400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_651
timestamp 1679581782
transform 1 0 63072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_658
timestamp 1679581782
transform 1 0 63744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_665
timestamp 1679581782
transform 1 0 64416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_672
timestamp 1679581782
transform 1 0 65088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_679
timestamp 1679581782
transform 1 0 65760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_686
timestamp 1679581782
transform 1 0 66432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_693
timestamp 1679581782
transform 1 0 67104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_700
timestamp 1679581782
transform 1 0 67776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_707
timestamp 1679581782
transform 1 0 68448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_714
timestamp 1679581782
transform 1 0 69120 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_721
timestamp 1677580104
transform 1 0 69792 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679581782
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679581782
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679581782
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679581782
transform 1 0 3264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679581782
transform 1 0 3936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679581782
transform 1 0 4608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679581782
transform 1 0 5280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679581782
transform 1 0 5952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_63
timestamp 1679581782
transform 1 0 6624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_70
timestamp 1679581782
transform 1 0 7296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_77
timestamp 1679581782
transform 1 0 7968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_84
timestamp 1679581782
transform 1 0 8640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_91
timestamp 1679581782
transform 1 0 9312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_98
timestamp 1679581782
transform 1 0 9984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_105
timestamp 1679581782
transform 1 0 10656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_112
timestamp 1679581782
transform 1 0 11328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_119
timestamp 1679581782
transform 1 0 12000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_126
timestamp 1679581782
transform 1 0 12672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_133
timestamp 1679581782
transform 1 0 13344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_140
timestamp 1679581782
transform 1 0 14016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_147
timestamp 1679581782
transform 1 0 14688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_154
timestamp 1679581782
transform 1 0 15360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_161
timestamp 1679581782
transform 1 0 16032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_168
timestamp 1679581782
transform 1 0 16704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_175
timestamp 1679581782
transform 1 0 17376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_182
timestamp 1679581782
transform 1 0 18048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_189
timestamp 1679581782
transform 1 0 18720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_196
timestamp 1679581782
transform 1 0 19392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_203
timestamp 1679581782
transform 1 0 20064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_210
timestamp 1679581782
transform 1 0 20736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_217
timestamp 1679581782
transform 1 0 21408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_224
timestamp 1679581782
transform 1 0 22080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_231
timestamp 1679581782
transform 1 0 22752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_238
timestamp 1679581782
transform 1 0 23424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_245
timestamp 1679581782
transform 1 0 24096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_252
timestamp 1679581782
transform 1 0 24768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_259
timestamp 1679581782
transform 1 0 25440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_266
timestamp 1679581782
transform 1 0 26112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_273
timestamp 1679581782
transform 1 0 26784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_280
timestamp 1679581782
transform 1 0 27456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_287
timestamp 1679581782
transform 1 0 28128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_294
timestamp 1679581782
transform 1 0 28800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_301
timestamp 1679581782
transform 1 0 29472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_308
timestamp 1679581782
transform 1 0 30144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_315
timestamp 1679581782
transform 1 0 30816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_322
timestamp 1679581782
transform 1 0 31488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_329
timestamp 1679581782
transform 1 0 32160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_336
timestamp 1679581782
transform 1 0 32832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_343
timestamp 1679581782
transform 1 0 33504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_350
timestamp 1679581782
transform 1 0 34176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_357
timestamp 1679581782
transform 1 0 34848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_364
timestamp 1679581782
transform 1 0 35520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_371
timestamp 1679581782
transform 1 0 36192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_378
timestamp 1679581782
transform 1 0 36864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_385
timestamp 1679581782
transform 1 0 37536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_392
timestamp 1679581782
transform 1 0 38208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_399
timestamp 1679581782
transform 1 0 38880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_406
timestamp 1679581782
transform 1 0 39552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_413
timestamp 1679581782
transform 1 0 40224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_420
timestamp 1679581782
transform 1 0 40896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_427
timestamp 1679581782
transform 1 0 41568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_434
timestamp 1679581782
transform 1 0 42240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_441
timestamp 1679581782
transform 1 0 42912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_448
timestamp 1679581782
transform 1 0 43584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_455
timestamp 1679581782
transform 1 0 44256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_462
timestamp 1679581782
transform 1 0 44928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_469
timestamp 1679581782
transform 1 0 45600 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_476
timestamp 1679581782
transform 1 0 46272 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_483
timestamp 1679581782
transform 1 0 46944 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_490
timestamp 1679581782
transform 1 0 47616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_497
timestamp 1679581782
transform 1 0 48288 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_504
timestamp 1679581782
transform 1 0 48960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_511
timestamp 1679581782
transform 1 0 49632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_518
timestamp 1679581782
transform 1 0 50304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_525
timestamp 1679581782
transform 1 0 50976 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_532
timestamp 1679581782
transform 1 0 51648 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_539
timestamp 1679581782
transform 1 0 52320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_546
timestamp 1679581782
transform 1 0 52992 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_553
timestamp 1679581782
transform 1 0 53664 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_560
timestamp 1679581782
transform 1 0 54336 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_567
timestamp 1679581782
transform 1 0 55008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_574
timestamp 1679581782
transform 1 0 55680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_581
timestamp 1679581782
transform 1 0 56352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_588
timestamp 1679581782
transform 1 0 57024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_595
timestamp 1679581782
transform 1 0 57696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_602
timestamp 1679581782
transform 1 0 58368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_609
timestamp 1679581782
transform 1 0 59040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_616
timestamp 1679581782
transform 1 0 59712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_623
timestamp 1679581782
transform 1 0 60384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_630
timestamp 1679581782
transform 1 0 61056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_637
timestamp 1679581782
transform 1 0 61728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_644
timestamp 1679581782
transform 1 0 62400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_651
timestamp 1679581782
transform 1 0 63072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_658
timestamp 1679581782
transform 1 0 63744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_665
timestamp 1679581782
transform 1 0 64416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_672
timestamp 1679581782
transform 1 0 65088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_679
timestamp 1679581782
transform 1 0 65760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_686
timestamp 1679581782
transform 1 0 66432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_693
timestamp 1679581782
transform 1 0 67104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_700
timestamp 1679581782
transform 1 0 67776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_707
timestamp 1679581782
transform 1 0 68448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_714
timestamp 1679581782
transform 1 0 69120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_721
timestamp 1679581782
transform 1 0 69792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_728
timestamp 1679581782
transform 1 0 70464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_735
timestamp 1679581782
transform 1 0 71136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_742
timestamp 1679581782
transform 1 0 71808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_749
timestamp 1679581782
transform 1 0 72480 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_756
timestamp 1677580104
transform 1 0 73152 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_762
timestamp 1677579658
transform 1 0 73728 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_767
timestamp 1677580104
transform 1 0 74208 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_783
timestamp 1677579658
transform 1 0 75744 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_791
timestamp 1677579658
transform 1 0 76512 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_799
timestamp 1677580104
transform 1 0 77280 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_818
timestamp 1677580104
transform 1 0 79104 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_823
timestamp 1677579658
transform 1 0 79584 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_857
timestamp 1677580104
transform 1 0 82848 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_886
timestamp 1677579658
transform 1 0 85632 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_891
timestamp 1677580104
transform 1 0 86112 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_906
timestamp 1677580104
transform 1 0 87552 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_912
timestamp 1677579658
transform 1 0 88128 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_920
timestamp 1677580104
transform 1 0 88896 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_932
timestamp 1677579658
transform 1 0 90048 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_940
timestamp 1677579658
transform 1 0 90816 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_970
timestamp 1677579658
transform 1 0 93696 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_978
timestamp 1677579658
transform 1 0 94464 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_987
timestamp 1677579658
transform 1 0 95328 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_991
timestamp 1677579658
transform 1 0 95712 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_1000
timestamp 1677579658
transform 1 0 96576 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_1008
timestamp 1677579658
transform 1 0 97344 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679581782
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679581782
transform 1 0 5280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679581782
transform 1 0 5952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679581782
transform 1 0 6624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679581782
transform 1 0 7296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679581782
transform 1 0 7968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679581782
transform 1 0 8640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679581782
transform 1 0 9312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679581782
transform 1 0 9984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679581782
transform 1 0 10656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679581782
transform 1 0 11328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_119
timestamp 1679581782
transform 1 0 12000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_126
timestamp 1679581782
transform 1 0 12672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_133
timestamp 1679581782
transform 1 0 13344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_140
timestamp 1679581782
transform 1 0 14016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_147
timestamp 1679581782
transform 1 0 14688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_154
timestamp 1679581782
transform 1 0 15360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_161
timestamp 1679581782
transform 1 0 16032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_168
timestamp 1679581782
transform 1 0 16704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_175
timestamp 1679581782
transform 1 0 17376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_182
timestamp 1679581782
transform 1 0 18048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_189
timestamp 1679581782
transform 1 0 18720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_196
timestamp 1679581782
transform 1 0 19392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_203
timestamp 1679581782
transform 1 0 20064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_210
timestamp 1679581782
transform 1 0 20736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_217
timestamp 1679581782
transform 1 0 21408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_224
timestamp 1679581782
transform 1 0 22080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_231
timestamp 1679581782
transform 1 0 22752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_238
timestamp 1679581782
transform 1 0 23424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_245
timestamp 1679581782
transform 1 0 24096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_252
timestamp 1679581782
transform 1 0 24768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_259
timestamp 1679581782
transform 1 0 25440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_266
timestamp 1679581782
transform 1 0 26112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_273
timestamp 1679581782
transform 1 0 26784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_280
timestamp 1679581782
transform 1 0 27456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_287
timestamp 1679581782
transform 1 0 28128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_294
timestamp 1679581782
transform 1 0 28800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_301
timestamp 1679581782
transform 1 0 29472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_308
timestamp 1679581782
transform 1 0 30144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_315
timestamp 1679581782
transform 1 0 30816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_322
timestamp 1679581782
transform 1 0 31488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_329
timestamp 1679581782
transform 1 0 32160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_336
timestamp 1679581782
transform 1 0 32832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_343
timestamp 1679581782
transform 1 0 33504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_350
timestamp 1679581782
transform 1 0 34176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_357
timestamp 1679581782
transform 1 0 34848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_364
timestamp 1679581782
transform 1 0 35520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_371
timestamp 1679581782
transform 1 0 36192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_378
timestamp 1679581782
transform 1 0 36864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_385
timestamp 1679581782
transform 1 0 37536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_392
timestamp 1679581782
transform 1 0 38208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_399
timestamp 1679581782
transform 1 0 38880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_406
timestamp 1679581782
transform 1 0 39552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_413
timestamp 1679581782
transform 1 0 40224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_420
timestamp 1679581782
transform 1 0 40896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_427
timestamp 1679581782
transform 1 0 41568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_434
timestamp 1679581782
transform 1 0 42240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_441
timestamp 1679581782
transform 1 0 42912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_448
timestamp 1679581782
transform 1 0 43584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_455
timestamp 1679581782
transform 1 0 44256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_462
timestamp 1679581782
transform 1 0 44928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_469
timestamp 1679581782
transform 1 0 45600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_476
timestamp 1679581782
transform 1 0 46272 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_483
timestamp 1679581782
transform 1 0 46944 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_490
timestamp 1679581782
transform 1 0 47616 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_497
timestamp 1679581782
transform 1 0 48288 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_504
timestamp 1679581782
transform 1 0 48960 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_511
timestamp 1679581782
transform 1 0 49632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_518
timestamp 1679581782
transform 1 0 50304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_525
timestamp 1679581782
transform 1 0 50976 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_532
timestamp 1679581782
transform 1 0 51648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_539
timestamp 1679581782
transform 1 0 52320 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_546
timestamp 1679581782
transform 1 0 52992 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_553
timestamp 1679581782
transform 1 0 53664 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_560
timestamp 1679581782
transform 1 0 54336 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_567
timestamp 1679581782
transform 1 0 55008 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_574
timestamp 1679581782
transform 1 0 55680 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_581
timestamp 1679581782
transform 1 0 56352 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_588
timestamp 1679581782
transform 1 0 57024 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_595
timestamp 1679581782
transform 1 0 57696 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_602
timestamp 1679581782
transform 1 0 58368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_609
timestamp 1679581782
transform 1 0 59040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_616
timestamp 1679581782
transform 1 0 59712 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_623
timestamp 1679581782
transform 1 0 60384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_630
timestamp 1679581782
transform 1 0 61056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_637
timestamp 1679581782
transform 1 0 61728 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_644
timestamp 1679581782
transform 1 0 62400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_651
timestamp 1679581782
transform 1 0 63072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_658
timestamp 1679581782
transform 1 0 63744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_665
timestamp 1679581782
transform 1 0 64416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_672
timestamp 1679581782
transform 1 0 65088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_679
timestamp 1679581782
transform 1 0 65760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_686
timestamp 1679581782
transform 1 0 66432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_693
timestamp 1679581782
transform 1 0 67104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_700
timestamp 1679581782
transform 1 0 67776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_707
timestamp 1679581782
transform 1 0 68448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_714
timestamp 1679581782
transform 1 0 69120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_721
timestamp 1679581782
transform 1 0 69792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_728
timestamp 1679581782
transform 1 0 70464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_735
timestamp 1679581782
transform 1 0 71136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_742
timestamp 1679581782
transform 1 0 71808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_749
timestamp 1679581782
transform 1 0 72480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_756
timestamp 1679577901
transform 1 0 73152 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_760
timestamp 1677579658
transform 1 0 73536 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_773
timestamp 1679581782
transform 1 0 74784 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_780
timestamp 1677579658
transform 1 0 75456 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_45_788
timestamp 1679577901
transform 1 0 76224 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_795
timestamp 1677579658
transform 1 0 76896 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_803
timestamp 1679581782
transform 1 0 77664 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_810
timestamp 1677579658
transform 1 0 78336 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_814
timestamp 1677580104
transform 1 0 78720 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_827
timestamp 1677579658
transform 1 0 79968 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_832
timestamp 1677579658
transform 1 0 80448 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_840
timestamp 1677580104
transform 1 0 81216 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_45_849
timestamp 1677580104
transform 1 0 82080 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_858
timestamp 1677579658
transform 1 0 82944 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_878
timestamp 1677579658
transform 1 0 84864 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_45_882
timestamp 1679577901
transform 1 0 85248 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_45_886
timestamp 1677579658
transform 1 0 85632 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_937
timestamp 1677579658
transform 1 0 90528 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_953
timestamp 1677579658
transform 1 0 92064 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_957
timestamp 1677579658
transform 1 0 92448 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_962
timestamp 1677579658
transform 1 0 92928 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_970
timestamp 1677580104
transform 1 0 93696 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_983
timestamp 1677579658
transform 1 0 94944 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_45_1006
timestamp 1679577901
transform 1 0 97152 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_1010
timestamp 1677580104
transform 1 0 97536 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_1016
timestamp 1679581782
transform 1 0 98112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_45_1023
timestamp 1679577901
transform 1 0 98784 0 -1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_45_1027
timestamp 1677580104
transform 1 0 99168 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679581782
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679581782
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679581782
transform 1 0 13344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679581782
transform 1 0 14016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679581782
transform 1 0 14688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679581782
transform 1 0 15360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679581782
transform 1 0 16032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679581782
transform 1 0 16704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679581782
transform 1 0 17376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_182
timestamp 1679581782
transform 1 0 18048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_189
timestamp 1679581782
transform 1 0 18720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_196
timestamp 1679581782
transform 1 0 19392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679581782
transform 1 0 20064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_210
timestamp 1679581782
transform 1 0 20736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_217
timestamp 1679581782
transform 1 0 21408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679581782
transform 1 0 22080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679581782
transform 1 0 22752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679581782
transform 1 0 23424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679581782
transform 1 0 24096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679581782
transform 1 0 24768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679581782
transform 1 0 25440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_266
timestamp 1679581782
transform 1 0 26112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_273
timestamp 1679581782
transform 1 0 26784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_280
timestamp 1679581782
transform 1 0 27456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679581782
transform 1 0 28128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679581782
transform 1 0 28800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679581782
transform 1 0 29472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679581782
transform 1 0 30144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_315
timestamp 1679581782
transform 1 0 30816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_322
timestamp 1679581782
transform 1 0 31488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_329
timestamp 1679581782
transform 1 0 32160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_336
timestamp 1679581782
transform 1 0 32832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_343
timestamp 1679581782
transform 1 0 33504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_350
timestamp 1679581782
transform 1 0 34176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_357
timestamp 1679581782
transform 1 0 34848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_364
timestamp 1679581782
transform 1 0 35520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_371
timestamp 1679581782
transform 1 0 36192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_378
timestamp 1679581782
transform 1 0 36864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_385
timestamp 1679581782
transform 1 0 37536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_392
timestamp 1679581782
transform 1 0 38208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_399
timestamp 1679581782
transform 1 0 38880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_406
timestamp 1679581782
transform 1 0 39552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_413
timestamp 1679581782
transform 1 0 40224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_420
timestamp 1679581782
transform 1 0 40896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679581782
transform 1 0 41568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679581782
transform 1 0 42240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679581782
transform 1 0 42912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679581782
transform 1 0 43584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679581782
transform 1 0 44256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679581782
transform 1 0 44928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679581782
transform 1 0 45600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679581782
transform 1 0 46272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679581782
transform 1 0 46944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679581782
transform 1 0 47616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_497
timestamp 1679581782
transform 1 0 48288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_504
timestamp 1679581782
transform 1 0 48960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_511
timestamp 1679581782
transform 1 0 49632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_518
timestamp 1679581782
transform 1 0 50304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_525
timestamp 1679581782
transform 1 0 50976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_532
timestamp 1679581782
transform 1 0 51648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_539
timestamp 1679581782
transform 1 0 52320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_546
timestamp 1679581782
transform 1 0 52992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_553
timestamp 1679581782
transform 1 0 53664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_560
timestamp 1679581782
transform 1 0 54336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_567
timestamp 1679581782
transform 1 0 55008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_574
timestamp 1679581782
transform 1 0 55680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_581
timestamp 1679581782
transform 1 0 56352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_588
timestamp 1679581782
transform 1 0 57024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_595
timestamp 1679581782
transform 1 0 57696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_602
timestamp 1679581782
transform 1 0 58368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_609
timestamp 1679581782
transform 1 0 59040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_616
timestamp 1679581782
transform 1 0 59712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_623
timestamp 1679581782
transform 1 0 60384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_630
timestamp 1679581782
transform 1 0 61056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_637
timestamp 1679581782
transform 1 0 61728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_644
timestamp 1679581782
transform 1 0 62400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_651
timestamp 1679581782
transform 1 0 63072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_658
timestamp 1679581782
transform 1 0 63744 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_665
timestamp 1679581782
transform 1 0 64416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_672
timestamp 1679581782
transform 1 0 65088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_679
timestamp 1679581782
transform 1 0 65760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_686
timestamp 1679581782
transform 1 0 66432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_693
timestamp 1679581782
transform 1 0 67104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_700
timestamp 1679581782
transform 1 0 67776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_707
timestamp 1679581782
transform 1 0 68448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_714
timestamp 1679581782
transform 1 0 69120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_721
timestamp 1679581782
transform 1 0 69792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_728
timestamp 1679581782
transform 1 0 70464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_735
timestamp 1679581782
transform 1 0 71136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_742
timestamp 1679581782
transform 1 0 71808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_749
timestamp 1679581782
transform 1 0 72480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_756
timestamp 1679581782
transform 1 0 73152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_763
timestamp 1679581782
transform 1 0 73824 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_770
timestamp 1677580104
transform 1 0 74496 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_772
timestamp 1677579658
transform 1 0 74688 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_777
timestamp 1679581782
transform 1 0 75168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_784
timestamp 1679581782
transform 1 0 75840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_795
timestamp 1679577901
transform 1 0 76896 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_799
timestamp 1677579658
transform 1 0 77280 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_804
timestamp 1679581782
transform 1 0 77760 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_811
timestamp 1677579658
transform 1 0 78432 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_816
timestamp 1677580104
transform 1 0 78912 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_822
timestamp 1679581782
transform 1 0 79488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_832
timestamp 1679581782
transform 1 0 80448 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_839
timestamp 1677580104
transform 1 0 81120 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_845
timestamp 1679581782
transform 1 0 81696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_852
timestamp 1679581782
transform 1 0 82368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_859
timestamp 1679581782
transform 1 0 83040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_866
timestamp 1679581782
transform 1 0 83712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_873
timestamp 1679577901
transform 1 0 84384 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_877
timestamp 1677580104
transform 1 0 84768 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_887
timestamp 1679581782
transform 1 0 85728 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_894
timestamp 1677579658
transform 1 0 86400 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_898
timestamp 1679581782
transform 1 0 86784 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_905
timestamp 1677580104
transform 1 0 87456 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_907
timestamp 1677579658
transform 1 0 87648 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_911
timestamp 1679581782
transform 1 0 88032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_918
timestamp 1679581782
transform 1 0 88704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_925
timestamp 1679577901
transform 1 0 89376 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_932
timestamp 1677579658
transform 1 0 90048 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_936
timestamp 1679581782
transform 1 0 90432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_943
timestamp 1679581782
transform 1 0 91104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_950
timestamp 1679577901
transform 1 0 91776 0 1 35532
box -48 -56 432 834
use sg13g2_decap_8  FILLER_46_958
timestamp 1679581782
transform 1 0 92544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_965
timestamp 1679577901
transform 1 0 93216 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_969
timestamp 1677580104
transform 1 0 93600 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_974
timestamp 1679581782
transform 1 0 94080 0 1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_981
timestamp 1677579658
transform 1 0 94752 0 1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_985
timestamp 1679581782
transform 1 0 95136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_992
timestamp 1679581782
transform 1 0 95808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_999
timestamp 1679581782
transform 1 0 96480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1006
timestamp 1679581782
transform 1 0 97152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1013
timestamp 1679581782
transform 1 0 97824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1020
timestamp 1679581782
transform 1 0 98496 0 1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_46_1027
timestamp 1677580104
transform 1 0 99168 0 1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679581782
transform 1 0 18048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679581782
transform 1 0 18720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679581782
transform 1 0 19392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679581782
transform 1 0 20064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679581782
transform 1 0 20736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679581782
transform 1 0 21408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679581782
transform 1 0 22080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679581782
transform 1 0 22752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679581782
transform 1 0 23424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679581782
transform 1 0 24096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679581782
transform 1 0 24768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679581782
transform 1 0 25440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679581782
transform 1 0 26112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679581782
transform 1 0 26784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679581782
transform 1 0 27456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679581782
transform 1 0 28128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679581782
transform 1 0 28800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679581782
transform 1 0 29472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679581782
transform 1 0 30144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679581782
transform 1 0 30816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679581782
transform 1 0 31488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679581782
transform 1 0 32160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679581782
transform 1 0 32832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679581782
transform 1 0 33504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679581782
transform 1 0 34176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679581782
transform 1 0 34848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679581782
transform 1 0 35520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679581782
transform 1 0 36192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679581782
transform 1 0 36864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679581782
transform 1 0 37536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679581782
transform 1 0 38208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679581782
transform 1 0 38880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679581782
transform 1 0 39552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679581782
transform 1 0 40224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679581782
transform 1 0 40896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679581782
transform 1 0 41568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679581782
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679581782
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679581782
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679581782
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679581782
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679581782
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679581782
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679581782
transform 1 0 54336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679581782
transform 1 0 55008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679581782
transform 1 0 55680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679581782
transform 1 0 56352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679581782
transform 1 0 57024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679581782
transform 1 0 57696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679581782
transform 1 0 58368 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679581782
transform 1 0 59040 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679581782
transform 1 0 59712 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679581782
transform 1 0 60384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679581782
transform 1 0 61056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679581782
transform 1 0 61728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679581782
transform 1 0 62400 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679581782
transform 1 0 63072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679581782
transform 1 0 63744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679581782
transform 1 0 64416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679581782
transform 1 0 65088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679581782
transform 1 0 65760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679581782
transform 1 0 66432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679581782
transform 1 0 67104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679581782
transform 1 0 67776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679581782
transform 1 0 68448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679581782
transform 1 0 69120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679581782
transform 1 0 69792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679581782
transform 1 0 70464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679581782
transform 1 0 71136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679581782
transform 1 0 71808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679581782
transform 1 0 72480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_756
timestamp 1679581782
transform 1 0 73152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_763
timestamp 1679581782
transform 1 0 73824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_770
timestamp 1679581782
transform 1 0 74496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_777
timestamp 1679581782
transform 1 0 75168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_784
timestamp 1679581782
transform 1 0 75840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_791
timestamp 1679581782
transform 1 0 76512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_798
timestamp 1679581782
transform 1 0 77184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_805
timestamp 1679581782
transform 1 0 77856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_812
timestamp 1679581782
transform 1 0 78528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_819
timestamp 1679581782
transform 1 0 79200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_826
timestamp 1679581782
transform 1 0 79872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_833
timestamp 1679581782
transform 1 0 80544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_840
timestamp 1679581782
transform 1 0 81216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_847
timestamp 1679581782
transform 1 0 81888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_854
timestamp 1679581782
transform 1 0 82560 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_861
timestamp 1679581782
transform 1 0 83232 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_868
timestamp 1679581782
transform 1 0 83904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_875
timestamp 1679581782
transform 1 0 84576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_882
timestamp 1679581782
transform 1 0 85248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_889
timestamp 1679581782
transform 1 0 85920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_896
timestamp 1679581782
transform 1 0 86592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_903
timestamp 1679581782
transform 1 0 87264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_910
timestamp 1679581782
transform 1 0 87936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_917
timestamp 1679581782
transform 1 0 88608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_924
timestamp 1679581782
transform 1 0 89280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_931
timestamp 1679581782
transform 1 0 89952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_938
timestamp 1679581782
transform 1 0 90624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_945
timestamp 1679581782
transform 1 0 91296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_952
timestamp 1679581782
transform 1 0 91968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_959
timestamp 1679581782
transform 1 0 92640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_966
timestamp 1679581782
transform 1 0 93312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_973
timestamp 1679581782
transform 1 0 93984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_980
timestamp 1679581782
transform 1 0 94656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_987
timestamp 1679581782
transform 1 0 95328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_994
timestamp 1679581782
transform 1 0 96000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1001
timestamp 1679581782
transform 1 0 96672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1008
timestamp 1679581782
transform 1 0 97344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1015
timestamp 1679581782
transform 1 0 98016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1022
timestamp 1679581782
transform 1 0 98688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679581782
transform 1 0 27456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679581782
transform 1 0 30816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679581782
transform 1 0 31488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679581782
transform 1 0 32160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679581782
transform 1 0 32832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679581782
transform 1 0 33504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679581782
transform 1 0 34176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679581782
transform 1 0 34848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679581782
transform 1 0 35520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679581782
transform 1 0 36192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679581782
transform 1 0 36864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679581782
transform 1 0 37536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679581782
transform 1 0 38208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679581782
transform 1 0 38880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679581782
transform 1 0 39552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679581782
transform 1 0 40224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679581782
transform 1 0 40896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679581782
transform 1 0 41568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679581782
transform 1 0 42240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679581782
transform 1 0 42912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679581782
transform 1 0 43584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679581782
transform 1 0 44256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679581782
transform 1 0 44928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679581782
transform 1 0 45600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679581782
transform 1 0 46272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679581782
transform 1 0 46944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679581782
transform 1 0 47616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679581782
transform 1 0 48288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679581782
transform 1 0 48960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679581782
transform 1 0 49632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679581782
transform 1 0 50304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679581782
transform 1 0 50976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679581782
transform 1 0 51648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679581782
transform 1 0 52320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679581782
transform 1 0 52992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679581782
transform 1 0 53664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679581782
transform 1 0 54336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_567
timestamp 1679581782
transform 1 0 55008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_574
timestamp 1679581782
transform 1 0 55680 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_581
timestamp 1679581782
transform 1 0 56352 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_588
timestamp 1679581782
transform 1 0 57024 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_595
timestamp 1679581782
transform 1 0 57696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_602
timestamp 1679581782
transform 1 0 58368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_609
timestamp 1679581782
transform 1 0 59040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_616
timestamp 1679581782
transform 1 0 59712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_623
timestamp 1679581782
transform 1 0 60384 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_630
timestamp 1679581782
transform 1 0 61056 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_637
timestamp 1679581782
transform 1 0 61728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_644
timestamp 1679581782
transform 1 0 62400 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_651
timestamp 1679581782
transform 1 0 63072 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_658
timestamp 1679581782
transform 1 0 63744 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_665
timestamp 1679581782
transform 1 0 64416 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_672
timestamp 1679581782
transform 1 0 65088 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_679
timestamp 1679581782
transform 1 0 65760 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_686
timestamp 1679581782
transform 1 0 66432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_693
timestamp 1679581782
transform 1 0 67104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_700
timestamp 1679581782
transform 1 0 67776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_707
timestamp 1679581782
transform 1 0 68448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_714
timestamp 1679581782
transform 1 0 69120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_721
timestamp 1679581782
transform 1 0 69792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_728
timestamp 1679581782
transform 1 0 70464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_735
timestamp 1679581782
transform 1 0 71136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_742
timestamp 1679581782
transform 1 0 71808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_749
timestamp 1679581782
transform 1 0 72480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_756
timestamp 1679581782
transform 1 0 73152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_763
timestamp 1679581782
transform 1 0 73824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_770
timestamp 1679581782
transform 1 0 74496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_777
timestamp 1679581782
transform 1 0 75168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_784
timestamp 1679581782
transform 1 0 75840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_791
timestamp 1679581782
transform 1 0 76512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_798
timestamp 1679581782
transform 1 0 77184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_805
timestamp 1679581782
transform 1 0 77856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_812
timestamp 1679581782
transform 1 0 78528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_819
timestamp 1679581782
transform 1 0 79200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_826
timestamp 1679581782
transform 1 0 79872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_833
timestamp 1679581782
transform 1 0 80544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_840
timestamp 1679581782
transform 1 0 81216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_847
timestamp 1679581782
transform 1 0 81888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_854
timestamp 1679581782
transform 1 0 82560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_861
timestamp 1679581782
transform 1 0 83232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_868
timestamp 1679581782
transform 1 0 83904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_875
timestamp 1679581782
transform 1 0 84576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_882
timestamp 1679581782
transform 1 0 85248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_889
timestamp 1679581782
transform 1 0 85920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_896
timestamp 1679581782
transform 1 0 86592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_903
timestamp 1679581782
transform 1 0 87264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_910
timestamp 1679581782
transform 1 0 87936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_917
timestamp 1679581782
transform 1 0 88608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_924
timestamp 1679581782
transform 1 0 89280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_931
timestamp 1679581782
transform 1 0 89952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_938
timestamp 1679581782
transform 1 0 90624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_945
timestamp 1679581782
transform 1 0 91296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_952
timestamp 1679581782
transform 1 0 91968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_959
timestamp 1679581782
transform 1 0 92640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_966
timestamp 1679581782
transform 1 0 93312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_973
timestamp 1679581782
transform 1 0 93984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_980
timestamp 1679581782
transform 1 0 94656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_987
timestamp 1679581782
transform 1 0 95328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_994
timestamp 1679581782
transform 1 0 96000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1001
timestamp 1679581782
transform 1 0 96672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1008
timestamp 1679581782
transform 1 0 97344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1015
timestamp 1679581782
transform 1 0 98016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1022
timestamp 1679581782
transform 1 0 98688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_0
timestamp 1679581782
transform 1 0 576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_7
timestamp 1679581782
transform 1 0 1248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_14
timestamp 1679581782
transform 1 0 1920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679581782
transform 1 0 2592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_28
timestamp 1679581782
transform 1 0 3264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_35
timestamp 1679581782
transform 1 0 3936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_42
timestamp 1679581782
transform 1 0 4608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_49
timestamp 1679581782
transform 1 0 5280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_56
timestamp 1679581782
transform 1 0 5952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_63
timestamp 1679581782
transform 1 0 6624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_70
timestamp 1679581782
transform 1 0 7296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_77
timestamp 1679581782
transform 1 0 7968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_84
timestamp 1679581782
transform 1 0 8640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_91
timestamp 1679581782
transform 1 0 9312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_98
timestamp 1679581782
transform 1 0 9984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_105
timestamp 1679581782
transform 1 0 10656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_112
timestamp 1679581782
transform 1 0 11328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_119
timestamp 1679581782
transform 1 0 12000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_126
timestamp 1679581782
transform 1 0 12672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_133
timestamp 1679581782
transform 1 0 13344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_140
timestamp 1679581782
transform 1 0 14016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_147
timestamp 1679581782
transform 1 0 14688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_154
timestamp 1679581782
transform 1 0 15360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_161
timestamp 1679581782
transform 1 0 16032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_168
timestamp 1679581782
transform 1 0 16704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_175
timestamp 1679581782
transform 1 0 17376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_182
timestamp 1679581782
transform 1 0 18048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_189
timestamp 1679581782
transform 1 0 18720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_196
timestamp 1679581782
transform 1 0 19392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_203
timestamp 1679581782
transform 1 0 20064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_210
timestamp 1679581782
transform 1 0 20736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_217
timestamp 1679581782
transform 1 0 21408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_224
timestamp 1679581782
transform 1 0 22080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_231
timestamp 1679581782
transform 1 0 22752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_238
timestamp 1679581782
transform 1 0 23424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_245
timestamp 1679581782
transform 1 0 24096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_252
timestamp 1679581782
transform 1 0 24768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_259
timestamp 1679581782
transform 1 0 25440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_266
timestamp 1679581782
transform 1 0 26112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_273
timestamp 1679581782
transform 1 0 26784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_280
timestamp 1679581782
transform 1 0 27456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_287
timestamp 1679581782
transform 1 0 28128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_294
timestamp 1679581782
transform 1 0 28800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_301
timestamp 1679581782
transform 1 0 29472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_308
timestamp 1679581782
transform 1 0 30144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_315
timestamp 1679581782
transform 1 0 30816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_322
timestamp 1679581782
transform 1 0 31488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_329
timestamp 1679581782
transform 1 0 32160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_336
timestamp 1679581782
transform 1 0 32832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_343
timestamp 1679581782
transform 1 0 33504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_350
timestamp 1679581782
transform 1 0 34176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_357
timestamp 1679581782
transform 1 0 34848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_364
timestamp 1679581782
transform 1 0 35520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_371
timestamp 1679581782
transform 1 0 36192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_378
timestamp 1679581782
transform 1 0 36864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_385
timestamp 1679581782
transform 1 0 37536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_392
timestamp 1679581782
transform 1 0 38208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_399
timestamp 1679581782
transform 1 0 38880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_406
timestamp 1679581782
transform 1 0 39552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_413
timestamp 1679581782
transform 1 0 40224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_420
timestamp 1679581782
transform 1 0 40896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_427
timestamp 1679581782
transform 1 0 41568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_434
timestamp 1679581782
transform 1 0 42240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_441
timestamp 1679581782
transform 1 0 42912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_448
timestamp 1679581782
transform 1 0 43584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_455
timestamp 1679581782
transform 1 0 44256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_462
timestamp 1679581782
transform 1 0 44928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_469
timestamp 1679581782
transform 1 0 45600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_476
timestamp 1679581782
transform 1 0 46272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_483
timestamp 1679581782
transform 1 0 46944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_490
timestamp 1679581782
transform 1 0 47616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_497
timestamp 1679581782
transform 1 0 48288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_504
timestamp 1679581782
transform 1 0 48960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_511
timestamp 1679581782
transform 1 0 49632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_518
timestamp 1679581782
transform 1 0 50304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_525
timestamp 1679581782
transform 1 0 50976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_532
timestamp 1679581782
transform 1 0 51648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_539
timestamp 1679581782
transform 1 0 52320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_546
timestamp 1679581782
transform 1 0 52992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_553
timestamp 1679581782
transform 1 0 53664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_560
timestamp 1679581782
transform 1 0 54336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_567
timestamp 1679581782
transform 1 0 55008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_574
timestamp 1679581782
transform 1 0 55680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_581
timestamp 1679581782
transform 1 0 56352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_588
timestamp 1679581782
transform 1 0 57024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_595
timestamp 1679581782
transform 1 0 57696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_602
timestamp 1679581782
transform 1 0 58368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_609
timestamp 1679581782
transform 1 0 59040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_616
timestamp 1679581782
transform 1 0 59712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_623
timestamp 1679581782
transform 1 0 60384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_630
timestamp 1679581782
transform 1 0 61056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_637
timestamp 1679581782
transform 1 0 61728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_644
timestamp 1679581782
transform 1 0 62400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_651
timestamp 1679581782
transform 1 0 63072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_658
timestamp 1679581782
transform 1 0 63744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_665
timestamp 1679581782
transform 1 0 64416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_672
timestamp 1679581782
transform 1 0 65088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_679
timestamp 1679581782
transform 1 0 65760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_686
timestamp 1679581782
transform 1 0 66432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_693
timestamp 1679581782
transform 1 0 67104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_700
timestamp 1679581782
transform 1 0 67776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_707
timestamp 1679581782
transform 1 0 68448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_714
timestamp 1679581782
transform 1 0 69120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_721
timestamp 1679581782
transform 1 0 69792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_728
timestamp 1679581782
transform 1 0 70464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_735
timestamp 1679581782
transform 1 0 71136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_742
timestamp 1679581782
transform 1 0 71808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_749
timestamp 1679581782
transform 1 0 72480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_756
timestamp 1679581782
transform 1 0 73152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_763
timestamp 1679581782
transform 1 0 73824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_770
timestamp 1679581782
transform 1 0 74496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_777
timestamp 1679581782
transform 1 0 75168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_784
timestamp 1679581782
transform 1 0 75840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_791
timestamp 1679581782
transform 1 0 76512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_798
timestamp 1679581782
transform 1 0 77184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_805
timestamp 1679581782
transform 1 0 77856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_812
timestamp 1679581782
transform 1 0 78528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_819
timestamp 1679581782
transform 1 0 79200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_826
timestamp 1679581782
transform 1 0 79872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_833
timestamp 1679581782
transform 1 0 80544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_840
timestamp 1679581782
transform 1 0 81216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_847
timestamp 1679581782
transform 1 0 81888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_854
timestamp 1679581782
transform 1 0 82560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_861
timestamp 1679581782
transform 1 0 83232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_868
timestamp 1679581782
transform 1 0 83904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_875
timestamp 1679581782
transform 1 0 84576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_882
timestamp 1679581782
transform 1 0 85248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_889
timestamp 1679581782
transform 1 0 85920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_896
timestamp 1679581782
transform 1 0 86592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_903
timestamp 1679581782
transform 1 0 87264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_910
timestamp 1679581782
transform 1 0 87936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_917
timestamp 1679581782
transform 1 0 88608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_924
timestamp 1679581782
transform 1 0 89280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_931
timestamp 1679581782
transform 1 0 89952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_938
timestamp 1679581782
transform 1 0 90624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_945
timestamp 1679581782
transform 1 0 91296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_952
timestamp 1679581782
transform 1 0 91968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_959
timestamp 1679581782
transform 1 0 92640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_966
timestamp 1679581782
transform 1 0 93312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_973
timestamp 1679581782
transform 1 0 93984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_980
timestamp 1679581782
transform 1 0 94656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_987
timestamp 1679581782
transform 1 0 95328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_994
timestamp 1679581782
transform 1 0 96000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1001
timestamp 1679581782
transform 1 0 96672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1008
timestamp 1679581782
transform 1 0 97344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1015
timestamp 1679581782
transform 1 0 98016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1022
timestamp 1679581782
transform 1 0 98688 0 -1 38556
box -48 -56 720 834
use sg13g2_tiehi  heichips25_pudding_118
timestamp 1680000651
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_119
timestamp 1680000651
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_120
timestamp 1680000651
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_121
timestamp 1680000651
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_122
timestamp 1680000651
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_123
timestamp 1680000651
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_124
timestamp 1680000651
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_125
timestamp 1680000651
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_buf_2  input1
timestamp 1676381867
transform -1 0 1056 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_2  input2
timestamp 1676381867
transform -1 0 1056 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  input3
timestamp 1676381867
transform -1 0 1056 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_2  input4
timestamp 1676381867
transform -1 0 1056 0 1 24948
box -48 -56 528 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform -1 0 960 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform -1 0 960 0 1 8316
box -48 -56 432 834
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 8316 630 8756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 12316 630 12756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 16316 630 16756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 20316 630 20756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 24316 630 24756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 28316 630 28756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 32316 630 32756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 36316 630 36756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 40316 630 40756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 44316 630 44756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 48316 630 48756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 52316 630 52756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 56316 630 56756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 60316 630 60756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64316 630 64756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 68316 630 68756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 72316 630 72756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 76316 630 76756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 80316 630 80756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 84316 630 84756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 88316 630 88756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 92316 630 92756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 96316 630 96756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 4496 99404 4936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 8496 99404 8936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 12496 99404 12936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 16496 99404 16936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 20496 99404 20936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 24496 99404 24936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 28496 99404 28936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 32496 99404 32936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 36496 99404 36936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 7076 712 7516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 11076 712 11516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 15076 712 15516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 19076 712 19516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 23076 712 23516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 27076 712 27516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 31076 712 31516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 35076 712 35516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 39076 712 39516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 43076 712 43516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 47076 712 47516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 51076 712 51516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 55076 712 55516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 59076 712 59516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63076 712 63516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 67076 712 67516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 71076 712 71516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 75076 712 75516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 79076 712 79516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 83076 712 83516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 87076 712 87516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 91076 712 91516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 95076 712 95516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 99076 712 99516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 3256 99516 3696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 7256 99516 7696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 11256 99516 11696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 15256 99516 15696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 19256 99516 19696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 23256 99516 23696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 27256 99516 27696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 31256 99516 31696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 35256 99516 35696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel via6 96536 12716 96536 12716 0 VGND
rlabel via6 95296 15476 95296 15476 0 VPWR
rlabel metal2 68544 25746 68544 25746 0 digitalH.g\[0\].u.OUTN
rlabel metal2 72725 25904 72725 25904 0 digitalH.g\[0\].u.OUTP
rlabel metal2 83525 31426 83525 31426 0 digitalH.g\[100\].u.OUTN
rlabel metal2 83635 31300 83635 31300 0 digitalH.g\[100\].u.OUTP
rlabel metal2 83125 31468 83125 31468 0 digitalH.g\[101\].u.OUTN
rlabel metal2 83235 31468 83235 31468 0 digitalH.g\[101\].u.OUTP
rlabel metal2 82725 31426 82725 31426 0 digitalH.g\[102\].u.OUTN
rlabel metal2 82835 31468 82835 31468 0 digitalH.g\[102\].u.OUTP
rlabel metal2 82325 31426 82325 31426 0 digitalH.g\[103\].u.OUTN
rlabel metal2 82435 31468 82435 31468 0 digitalH.g\[103\].u.OUTP
rlabel metal2 81984 32172 81984 32172 0 digitalH.g\[104\].u.OUTN
rlabel metal2 82035 31426 82035 31426 0 digitalH.g\[104\].u.OUTP
rlabel metal2 81525 31468 81525 31468 0 digitalH.g\[105\].u.OUTN
rlabel metal2 81635 31426 81635 31426 0 digitalH.g\[105\].u.OUTP
rlabel metal2 81125 31426 81125 31426 0 digitalH.g\[106\].u.OUTN
rlabel metal2 81235 31468 81235 31468 0 digitalH.g\[106\].u.OUTP
rlabel metal2 80725 31468 80725 31468 0 digitalH.g\[107\].u.OUTN
rlabel metal2 80835 31468 80835 31468 0 digitalH.g\[107\].u.OUTP
rlabel metal2 80325 31468 80325 31468 0 digitalH.g\[108\].u.OUTN
rlabel metal2 80435 31468 80435 31468 0 digitalH.g\[108\].u.OUTP
rlabel metal2 79925 31300 79925 31300 0 digitalH.g\[109\].u.OUTN
rlabel metal2 80035 31300 80035 31300 0 digitalH.g\[109\].u.OUTP
rlabel metal2 76704 22890 76704 22890 0 digitalH.g\[10\].u.OUTN
rlabel metal2 76800 23688 76800 23688 0 digitalH.g\[10\].u.OUTP
rlabel metal2 79525 31468 79525 31468 0 digitalH.g\[110\].u.OUTN
rlabel metal2 79635 31468 79635 31468 0 digitalH.g\[110\].u.OUTP
rlabel metal2 79125 31468 79125 31468 0 digitalH.g\[111\].u.OUTN
rlabel metal2 79235 31510 79235 31510 0 digitalH.g\[111\].u.OUTP
rlabel metal2 78725 31468 78725 31468 0 digitalH.g\[112\].u.OUTN
rlabel metal2 78835 31468 78835 31468 0 digitalH.g\[112\].u.OUTP
rlabel metal2 78325 31468 78325 31468 0 digitalH.g\[113\].u.OUTN
rlabel metal2 78435 31468 78435 31468 0 digitalH.g\[113\].u.OUTP
rlabel metal2 77925 31468 77925 31468 0 digitalH.g\[114\].u.OUTN
rlabel metal2 78035 31468 78035 31468 0 digitalH.g\[114\].u.OUTP
rlabel metal2 77525 31426 77525 31426 0 digitalH.g\[115\].u.OUTN
rlabel metal2 77635 31468 77635 31468 0 digitalH.g\[115\].u.OUTP
rlabel metal2 77125 31300 77125 31300 0 digitalH.g\[116\].u.OUTN
rlabel metal2 77235 31300 77235 31300 0 digitalH.g\[116\].u.OUTP
rlabel metal2 76725 31468 76725 31468 0 digitalH.g\[117\].u.OUTN
rlabel metal2 76835 31384 76835 31384 0 digitalH.g\[117\].u.OUTP
rlabel metal2 76325 31426 76325 31426 0 digitalH.g\[118\].u.OUTN
rlabel metal2 76435 31468 76435 31468 0 digitalH.g\[118\].u.OUTP
rlabel metal2 75925 31468 75925 31468 0 digitalH.g\[119\].u.OUTN
rlabel metal2 76035 31300 76035 31300 0 digitalH.g\[119\].u.OUTP
rlabel metal2 77232 22512 77232 22512 0 digitalH.g\[11\].u.OUTN
rlabel metal2 77088 24444 77088 24444 0 digitalH.g\[11\].u.OUTP
rlabel metal2 75525 31468 75525 31468 0 digitalH.g\[120\].u.OUTN
rlabel metal2 75635 31468 75635 31468 0 digitalH.g\[120\].u.OUTP
rlabel metal2 75125 31468 75125 31468 0 digitalH.g\[121\].u.OUTN
rlabel metal2 75235 31510 75235 31510 0 digitalH.g\[121\].u.OUTP
rlabel metal2 74688 31668 74688 31668 0 digitalH.g\[122\].u.OUTN
rlabel metal2 74835 31384 74835 31384 0 digitalH.g\[122\].u.OUTP
rlabel metal2 68784 30828 68784 30828 0 digitalH.g\[123\].u.OUTN
rlabel metal2 74435 31468 74435 31468 0 digitalH.g\[123\].u.OUTP
rlabel metal2 67200 31542 67200 31542 0 digitalH.g\[124\].u.OUTN
rlabel metal2 74035 31468 74035 31468 0 digitalH.g\[124\].u.OUTP
rlabel metal3 71484 31584 71484 31584 0 digitalH.g\[125\].u.OUTN
rlabel metal3 68736 31752 68736 31752 0 digitalH.g\[125\].u.OUTP
rlabel metal2 69456 30828 69456 30828 0 digitalH.g\[126\].u.OUTN
rlabel metal3 68832 31626 68832 31626 0 digitalH.g\[126\].u.OUTP
rlabel metal3 70512 30828 70512 30828 0 digitalH.g\[127\].u.OUTN
rlabel metal2 72835 31342 72835 31342 0 digitalH.g\[127\].u.OUTP
rlabel metal2 77616 21756 77616 21756 0 digitalH.g\[12\].u.OUTN
rlabel metal2 77472 24444 77472 24444 0 digitalH.g\[12\].u.OUTP
rlabel metal2 78048 24444 78048 24444 0 digitalH.g\[13\].u.OUTN
rlabel metal2 77952 24066 77952 24066 0 digitalH.g\[13\].u.OUTP
rlabel metal3 78816 23268 78816 23268 0 digitalH.g\[14\].u.OUTN
rlabel metal2 78336 24066 78336 24066 0 digitalH.g\[14\].u.OUTP
rlabel metal2 78816 22092 78816 22092 0 digitalH.g\[15\].u.OUTN
rlabel metal2 78624 24528 78624 24528 0 digitalH.g\[15\].u.OUTP
rlabel metal2 79488 23856 79488 23856 0 digitalH.g\[16\].u.OUTN
rlabel metal2 79104 22050 79104 22050 0 digitalH.g\[16\].u.OUTP
rlabel metal2 79872 24486 79872 24486 0 digitalH.g\[17\].u.OUTN
rlabel metal2 79584 21756 79584 21756 0 digitalH.g\[17\].u.OUTP
rlabel metal2 80928 23856 80928 23856 0 digitalH.g\[18\].u.OUTN
rlabel metal2 79872 22512 79872 22512 0 digitalH.g\[18\].u.OUTP
rlabel metal2 81216 23814 81216 23814 0 digitalH.g\[19\].u.OUTN
rlabel metal2 80160 24066 80160 24066 0 digitalH.g\[19\].u.OUTP
rlabel metal2 68928 25494 68928 25494 0 digitalH.g\[1\].u.OUTN
rlabel metal2 73248 25620 73248 25620 0 digitalH.g\[1\].u.OUTP
rlabel metal2 80832 24066 80832 24066 0 digitalH.g\[20\].u.OUTN
rlabel metal2 80640 22890 80640 22890 0 digitalH.g\[20\].u.OUTP
rlabel metal2 81408 23268 81408 23268 0 digitalH.g\[21\].u.OUTN
rlabel metal2 81072 21756 81072 21756 0 digitalH.g\[21\].u.OUTP
rlabel metal2 81792 24444 81792 24444 0 digitalH.g\[22\].u.OUTN
rlabel metal2 81600 22512 81600 22512 0 digitalH.g\[22\].u.OUTP
rlabel metal2 82080 24444 82080 24444 0 digitalH.g\[23\].u.OUTN
rlabel metal2 81984 24024 81984 24024 0 digitalH.g\[23\].u.OUTP
rlabel metal2 82560 23730 82560 23730 0 digitalH.g\[24\].u.OUTN
rlabel metal2 82368 23688 82368 23688 0 digitalH.g\[24\].u.OUTP
rlabel metal2 82944 24444 82944 24444 0 digitalH.g\[25\].u.OUTN
rlabel metal2 82656 24444 82656 24444 0 digitalH.g\[25\].u.OUTP
rlabel metal3 83664 22848 83664 22848 0 digitalH.g\[26\].u.OUTN
rlabel metal2 83040 24066 83040 24066 0 digitalH.g\[26\].u.OUTP
rlabel metal2 83664 22512 83664 22512 0 digitalH.g\[27\].u.OUTN
rlabel metal2 83616 22050 83616 22050 0 digitalH.g\[27\].u.OUTP
rlabel metal2 84288 22092 84288 22092 0 digitalH.g\[28\].u.OUTN
rlabel metal2 83952 22512 83952 22512 0 digitalH.g\[28\].u.OUTP
rlabel metal2 84384 23268 84384 23268 0 digitalH.g\[29\].u.OUTN
rlabel metal3 84336 21756 84336 21756 0 digitalH.g\[29\].u.OUTP
rlabel metal2 73536 23268 73536 23268 0 digitalH.g\[2\].u.OUTN
rlabel metal2 69792 25368 69792 25368 0 digitalH.g\[2\].u.OUTP
rlabel metal2 84864 24444 84864 24444 0 digitalH.g\[30\].u.OUTN
rlabel metal2 84864 22512 84864 22512 0 digitalH.g\[30\].u.OUTP
rlabel metal2 85248 24444 85248 24444 0 digitalH.g\[31\].u.OUTN
rlabel metal2 85104 22512 85104 22512 0 digitalH.g\[31\].u.OUTP
rlabel metal2 85536 24444 85536 24444 0 digitalH.g\[32\].u.OUTN
rlabel metal4 85440 23226 85440 23226 0 digitalH.g\[32\].u.OUTP
rlabel metal2 86016 22050 86016 22050 0 digitalH.g\[33\].u.OUTN
rlabel metal2 86016 24066 86016 24066 0 digitalH.g\[33\].u.OUTP
rlabel metal2 86448 21756 86448 21756 0 digitalH.g\[34\].u.OUTN
rlabel metal2 86304 24486 86304 24486 0 digitalH.g\[34\].u.OUTP
rlabel metal2 86880 23688 86880 23688 0 digitalH.g\[35\].u.OUTN
rlabel metal2 86784 24024 86784 24024 0 digitalH.g\[35\].u.OUTP
rlabel metal2 87744 24486 87744 24486 0 digitalH.g\[36\].u.OUTN
rlabel metal2 87168 24444 87168 24444 0 digitalH.g\[36\].u.OUTP
rlabel metal3 87360 22512 87360 22512 0 digitalH.g\[37\].u.OUTN
rlabel metal2 87504 22512 87504 22512 0 digitalH.g\[37\].u.OUTP
rlabel metal2 88032 24444 88032 24444 0 digitalH.g\[38\].u.OUTN
rlabel metal2 87888 22512 87888 22512 0 digitalH.g\[38\].u.OUTP
rlabel metal3 88320 23268 88320 23268 0 digitalH.g\[39\].u.OUTN
rlabel metal2 88224 24150 88224 24150 0 digitalH.g\[39\].u.OUTP
rlabel metal2 69936 25872 69936 25872 0 digitalH.g\[3\].u.OUTN
rlabel metal3 68448 25494 68448 25494 0 digitalH.g\[3\].u.OUTP
rlabel metal2 88896 24444 88896 24444 0 digitalH.g\[40\].u.OUTN
rlabel metal2 88608 22890 88608 22890 0 digitalH.g\[40\].u.OUTP
rlabel metal2 89136 21756 89136 21756 0 digitalH.g\[41\].u.OUTN
rlabel metal2 89088 24066 89088 24066 0 digitalH.g\[41\].u.OUTP
rlabel metal3 89520 23268 89520 23268 0 digitalH.g\[42\].u.OUTN
rlabel metal2 89568 23688 89568 23688 0 digitalH.g\[42\].u.OUTP
rlabel metal2 90528 24486 90528 24486 0 digitalH.g\[43\].u.OUTN
rlabel metal2 89952 24066 89952 24066 0 digitalH.g\[43\].u.OUTP
rlabel metal2 90816 23562 90816 23562 0 digitalH.g\[44\].u.OUTN
rlabel metal2 90240 24066 90240 24066 0 digitalH.g\[44\].u.OUTP
rlabel metal2 91104 23604 91104 23604 0 digitalH.g\[45\].u.OUTN
rlabel metal2 90725 25820 90725 25820 0 digitalH.g\[45\].u.OUTP
rlabel metal2 91200 22134 91200 22134 0 digitalH.g\[46\].u.OUTN
rlabel metal2 91728 22512 91728 22512 0 digitalH.g\[46\].u.OUTP
rlabel metal3 91536 22260 91536 22260 0 digitalH.g\[47\].u.OUTN
rlabel metal2 91536 22512 91536 22512 0 digitalH.g\[47\].u.OUTP
rlabel metal2 91440 23268 91440 23268 0 digitalH.g\[48\].u.OUTN
rlabel metal2 92112 22512 92112 22512 0 digitalH.g\[48\].u.OUTP
rlabel metal2 93648 23100 93648 23100 0 digitalH.g\[49\].u.OUTN
rlabel metal2 92400 22512 92400 22512 0 digitalH.g\[49\].u.OUTP
rlabel metal2 73920 24108 73920 24108 0 digitalH.g\[4\].u.OUTN
rlabel metal2 68832 25746 68832 25746 0 digitalH.g\[4\].u.OUTP
rlabel metal2 92880 21756 92880 21756 0 digitalH.g\[50\].u.OUTN
rlabel metal2 92778 25620 92778 25620 0 digitalH.g\[50\].u.OUTP
rlabel metal2 93360 21756 93360 21756 0 digitalH.g\[51\].u.OUTN
rlabel metal2 93122 25620 93122 25620 0 digitalH.g\[51\].u.OUTP
rlabel metal3 93840 23268 93840 23268 0 digitalH.g\[52\].u.OUTN
rlabel metal2 93514 25620 93514 25620 0 digitalH.g\[52\].u.OUTP
rlabel metal2 93792 22176 93792 22176 0 digitalH.g\[53\].u.OUTN
rlabel metal2 93936 22512 93936 22512 0 digitalH.g\[53\].u.OUTP
rlabel metal2 94435 25862 94435 25862 0 digitalH.g\[54\].u.OUTN
rlabel metal2 94346 25620 94346 25620 0 digitalH.g\[54\].u.OUTP
rlabel metal2 94841 25620 94841 25620 0 digitalH.g\[55\].u.OUTN
rlabel metal2 94690 25620 94690 25620 0 digitalH.g\[55\].u.OUTP
rlabel metal3 95136 21756 95136 21756 0 digitalH.g\[56\].u.OUTN
rlabel metal3 95040 22428 95040 22428 0 digitalH.g\[56\].u.OUTP
rlabel metal3 95568 24696 95568 24696 0 digitalH.g\[57\].u.OUTN
rlabel metal2 95568 22512 95568 22512 0 digitalH.g\[57\].u.OUTP
rlabel metal3 96288 23268 96288 23268 0 digitalH.g\[58\].u.OUTN
rlabel metal2 95952 22512 95952 22512 0 digitalH.g\[58\].u.OUTP
rlabel metal2 96816 23268 96816 23268 0 digitalH.g\[59\].u.OUTN
rlabel metal2 96240 22512 96240 22512 0 digitalH.g\[59\].u.OUTP
rlabel metal2 73152 23688 73152 23688 0 digitalH.g\[5\].u.OUTN
rlabel metal2 74640 22512 74640 22512 0 digitalH.g\[5\].u.OUTP
rlabel metal2 97008 24948 97008 24948 0 digitalH.g\[60\].u.OUTN
rlabel metal2 96864 22512 96864 22512 0 digitalH.g\[60\].u.OUTP
rlabel metal2 97289 25620 97289 25620 0 digitalH.g\[61\].u.OUTN
rlabel metal2 97152 22512 97152 22512 0 digitalH.g\[61\].u.OUTP
rlabel metal2 97681 25620 97681 25620 0 digitalH.g\[62\].u.OUTN
rlabel metal2 97584 22512 97584 22512 0 digitalH.g\[62\].u.OUTP
rlabel metal2 98073 25620 98073 25620 0 digitalH.g\[63\].u.OUTN
rlabel metal2 97968 22512 97968 22512 0 digitalH.g\[63\].u.OUTP
rlabel metal3 98448 34188 98448 34188 0 digitalH.g\[64\].u.OUTN
rlabel metal2 98064 34944 98064 34944 0 digitalH.g\[64\].u.OUTP
rlabel metal2 97525 31426 97525 31426 0 digitalH.g\[65\].u.OUTN
rlabel metal2 97635 31426 97635 31426 0 digitalH.g\[65\].u.OUTP
rlabel metal3 97008 34524 97008 34524 0 digitalH.g\[66\].u.OUTN
rlabel metal2 97235 31468 97235 31468 0 digitalH.g\[66\].u.OUTP
rlabel metal3 97440 34020 97440 34020 0 digitalH.g\[67\].u.OUTN
rlabel metal3 96816 34104 96816 34104 0 digitalH.g\[67\].u.OUTP
rlabel metal3 96576 34944 96576 34944 0 digitalH.g\[68\].u.OUTN
rlabel metal2 96336 34188 96336 34188 0 digitalH.g\[68\].u.OUTP
rlabel metal3 95472 34944 95472 34944 0 digitalH.g\[69\].u.OUTN
rlabel metal2 96017 31668 96017 31668 0 digitalH.g\[69\].u.OUTP
rlabel metal2 67584 25368 67584 25368 0 digitalH.g\[6\].u.OUTN
rlabel metal2 74976 24444 74976 24444 0 digitalH.g\[6\].u.OUTP
rlabel metal2 95522 31668 95522 31668 0 digitalH.g\[70\].u.OUTN
rlabel metal2 95664 34944 95664 34944 0 digitalH.g\[70\].u.OUTP
rlabel metal2 95088 34608 95088 34608 0 digitalH.g\[71\].u.OUTN
rlabel metal2 95233 31668 95233 31668 0 digitalH.g\[71\].u.OUTP
rlabel metal2 94725 31468 94725 31468 0 digitalH.g\[72\].u.OUTN
rlabel metal2 94835 31468 94835 31468 0 digitalH.g\[72\].u.OUTP
rlabel metal2 94325 31468 94325 31468 0 digitalH.g\[73\].u.OUTN
rlabel metal2 94416 34944 94416 34944 0 digitalH.g\[73\].u.OUTP
rlabel metal2 93936 34608 93936 34608 0 digitalH.g\[74\].u.OUTN
rlabel metal2 94035 31468 94035 31468 0 digitalH.g\[74\].u.OUTP
rlabel metal2 93312 34944 93312 34944 0 digitalH.g\[75\].u.OUTN
rlabel metal2 93648 34944 93648 34944 0 digitalH.g\[75\].u.OUTP
rlabel metal3 93312 34188 93312 34188 0 digitalH.g\[76\].u.OUTN
rlabel metal2 93264 34188 93264 34188 0 digitalH.g\[76\].u.OUTP
rlabel metal3 92400 34188 92400 34188 0 digitalH.g\[77\].u.OUTN
rlabel metal2 92880 34944 92880 34944 0 digitalH.g\[77\].u.OUTP
rlabel metal2 92304 34188 92304 34188 0 digitalH.g\[78\].u.OUTN
rlabel metal3 92352 35700 92352 35700 0 digitalH.g\[78\].u.OUTP
rlabel metal2 91728 34944 91728 34944 0 digitalH.g\[79\].u.OUTN
rlabel metal2 92064 34944 92064 34944 0 digitalH.g\[79\].u.OUTP
rlabel metal2 74112 24234 74112 24234 0 digitalH.g\[7\].u.OUTN
rlabel metal2 75552 24444 75552 24444 0 digitalH.g\[7\].u.OUTP
rlabel metal2 91680 33474 91680 33474 0 digitalH.g\[80\].u.OUTN
rlabel metal2 90912 33852 90912 33852 0 digitalH.g\[80\].u.OUTP
rlabel metal2 91125 31384 91125 31384 0 digitalH.g\[81\].u.OUTN
rlabel metal2 91056 34608 91056 34608 0 digitalH.g\[81\].u.OUTP
rlabel metal2 90725 31468 90725 31468 0 digitalH.g\[82\].u.OUTN
rlabel metal2 90825 31668 90825 31668 0 digitalH.g\[82\].u.OUTP
rlabel metal2 90325 31468 90325 31468 0 digitalH.g\[83\].u.OUTN
rlabel metal2 90435 31468 90435 31468 0 digitalH.g\[83\].u.OUTP
rlabel metal2 89952 35490 89952 35490 0 digitalH.g\[84\].u.OUTN
rlabel metal2 90035 31468 90035 31468 0 digitalH.g\[84\].u.OUTP
rlabel metal2 89525 31342 89525 31342 0 digitalH.g\[85\].u.OUTN
rlabel metal2 89635 31468 89635 31468 0 digitalH.g\[85\].u.OUTP
rlabel metal2 89125 31468 89125 31468 0 digitalH.g\[86\].u.OUTN
rlabel metal2 89235 31300 89235 31300 0 digitalH.g\[86\].u.OUTP
rlabel metal2 88725 31300 88725 31300 0 digitalH.g\[87\].u.OUTN
rlabel metal2 88835 31300 88835 31300 0 digitalH.g\[87\].u.OUTP
rlabel metal2 88325 31426 88325 31426 0 digitalH.g\[88\].u.OUTN
rlabel metal2 88435 31426 88435 31426 0 digitalH.g\[88\].u.OUTP
rlabel metal2 87925 31468 87925 31468 0 digitalH.g\[89\].u.OUTN
rlabel metal2 88035 31468 88035 31468 0 digitalH.g\[89\].u.OUTP
rlabel metal2 75936 21756 75936 21756 0 digitalH.g\[8\].u.OUTN
rlabel metal2 75936 24444 75936 24444 0 digitalH.g\[8\].u.OUTP
rlabel metal2 87525 31300 87525 31300 0 digitalH.g\[90\].u.OUTN
rlabel metal2 87635 31468 87635 31468 0 digitalH.g\[90\].u.OUTP
rlabel metal2 87125 31384 87125 31384 0 digitalH.g\[91\].u.OUTN
rlabel metal2 87235 31426 87235 31426 0 digitalH.g\[91\].u.OUTP
rlabel metal2 86725 31468 86725 31468 0 digitalH.g\[92\].u.OUTN
rlabel metal2 86835 31384 86835 31384 0 digitalH.g\[92\].u.OUTP
rlabel metal2 86325 31426 86325 31426 0 digitalH.g\[93\].u.OUTN
rlabel metal2 86435 31468 86435 31468 0 digitalH.g\[93\].u.OUTP
rlabel metal2 85925 31468 85925 31468 0 digitalH.g\[94\].u.OUTN
rlabel metal2 86035 31468 86035 31468 0 digitalH.g\[94\].u.OUTP
rlabel metal2 85525 31468 85525 31468 0 digitalH.g\[95\].u.OUTN
rlabel metal2 85635 31468 85635 31468 0 digitalH.g\[95\].u.OUTP
rlabel metal2 85125 31468 85125 31468 0 digitalH.g\[96\].u.OUTN
rlabel metal2 85235 31384 85235 31384 0 digitalH.g\[96\].u.OUTP
rlabel metal2 84725 31426 84725 31426 0 digitalH.g\[97\].u.OUTN
rlabel metal2 84835 31468 84835 31468 0 digitalH.g\[97\].u.OUTP
rlabel metal2 84325 31468 84325 31468 0 digitalH.g\[98\].u.OUTN
rlabel metal2 84435 31468 84435 31468 0 digitalH.g\[98\].u.OUTP
rlabel metal2 83925 31426 83925 31426 0 digitalH.g\[99\].u.OUTN
rlabel metal2 84035 31468 84035 31468 0 digitalH.g\[99\].u.OUTP
rlabel metal2 75888 22512 75888 22512 0 digitalH.g\[9\].u.OUTN
rlabel metal2 76272 22512 76272 22512 0 digitalH.g\[9\].u.OUTP
rlabel metal2 68256 9828 68256 9828 0 digitalL.g\[0\].u.OUTN
rlabel metal3 70944 9324 70944 9324 0 digitalL.g\[0\].u.OUTP
rlabel metal2 83525 15424 83525 15424 0 digitalL.g\[100\].u.OUTN
rlabel metal2 83635 15424 83635 15424 0 digitalL.g\[100\].u.OUTP
rlabel metal2 83125 15424 83125 15424 0 digitalL.g\[101\].u.OUTN
rlabel metal2 83235 15424 83235 15424 0 digitalL.g\[101\].u.OUTP
rlabel metal2 82725 15424 82725 15424 0 digitalL.g\[102\].u.OUTN
rlabel metal2 82835 15340 82835 15340 0 digitalL.g\[102\].u.OUTP
rlabel metal2 82325 15424 82325 15424 0 digitalL.g\[103\].u.OUTN
rlabel metal2 82435 15424 82435 15424 0 digitalL.g\[103\].u.OUTP
rlabel metal2 81984 16590 81984 16590 0 digitalL.g\[104\].u.OUTN
rlabel metal2 82035 15382 82035 15382 0 digitalL.g\[104\].u.OUTP
rlabel metal2 81525 15424 81525 15424 0 digitalL.g\[105\].u.OUTN
rlabel metal2 81635 15424 81635 15424 0 digitalL.g\[105\].u.OUTP
rlabel metal2 81125 15424 81125 15424 0 digitalL.g\[106\].u.OUTN
rlabel metal2 81235 15382 81235 15382 0 digitalL.g\[106\].u.OUTP
rlabel metal2 80725 15424 80725 15424 0 digitalL.g\[107\].u.OUTN
rlabel metal2 80835 15298 80835 15298 0 digitalL.g\[107\].u.OUTP
rlabel metal2 80325 15340 80325 15340 0 digitalL.g\[108\].u.OUTN
rlabel metal2 80435 15382 80435 15382 0 digitalL.g\[108\].u.OUTP
rlabel metal2 79925 15424 79925 15424 0 digitalL.g\[109\].u.OUTN
rlabel metal2 80035 15424 80035 15424 0 digitalL.g\[109\].u.OUTP
rlabel metal2 76800 8148 76800 8148 0 digitalL.g\[10\].u.OUTN
rlabel metal2 76666 9744 76666 9744 0 digitalL.g\[10\].u.OUTP
rlabel metal2 79525 15424 79525 15424 0 digitalL.g\[110\].u.OUTN
rlabel metal2 79635 15424 79635 15424 0 digitalL.g\[110\].u.OUTP
rlabel metal2 79125 15424 79125 15424 0 digitalL.g\[111\].u.OUTN
rlabel metal2 79235 15382 79235 15382 0 digitalL.g\[111\].u.OUTP
rlabel metal2 78725 15424 78725 15424 0 digitalL.g\[112\].u.OUTN
rlabel metal2 78835 15298 78835 15298 0 digitalL.g\[112\].u.OUTP
rlabel metal2 78325 15424 78325 15424 0 digitalL.g\[113\].u.OUTN
rlabel metal2 78435 15340 78435 15340 0 digitalL.g\[113\].u.OUTP
rlabel metal2 77925 15298 77925 15298 0 digitalL.g\[114\].u.OUTN
rlabel metal2 77904 19068 77904 19068 0 digitalL.g\[114\].u.OUTP
rlabel metal2 77525 15424 77525 15424 0 digitalL.g\[115\].u.OUTN
rlabel metal2 77635 15424 77635 15424 0 digitalL.g\[115\].u.OUTP
rlabel metal2 77125 15424 77125 15424 0 digitalL.g\[116\].u.OUTN
rlabel metal2 77235 15424 77235 15424 0 digitalL.g\[116\].u.OUTP
rlabel metal2 76725 15298 76725 15298 0 digitalL.g\[117\].u.OUTN
rlabel metal2 76835 15340 76835 15340 0 digitalL.g\[117\].u.OUTP
rlabel metal2 76325 15340 76325 15340 0 digitalL.g\[118\].u.OUTN
rlabel metal2 76435 15382 76435 15382 0 digitalL.g\[118\].u.OUTP
rlabel metal2 75925 15424 75925 15424 0 digitalL.g\[119\].u.OUTN
rlabel metal2 76035 15424 76035 15424 0 digitalL.g\[119\].u.OUTP
rlabel metal3 76608 7182 76608 7182 0 digitalL.g\[11\].u.OUTN
rlabel metal2 77184 8148 77184 8148 0 digitalL.g\[11\].u.OUTP
rlabel metal2 75525 15424 75525 15424 0 digitalL.g\[120\].u.OUTN
rlabel metal2 75635 15424 75635 15424 0 digitalL.g\[120\].u.OUTP
rlabel metal2 75125 15298 75125 15298 0 digitalL.g\[121\].u.OUTN
rlabel metal2 74832 18312 74832 18312 0 digitalL.g\[121\].u.OUTP
rlabel metal2 74725 15382 74725 15382 0 digitalL.g\[122\].u.OUTN
rlabel metal2 74835 15424 74835 15424 0 digitalL.g\[122\].u.OUTP
rlabel metal2 69936 14196 69936 14196 0 digitalL.g\[123\].u.OUTN
rlabel metal2 74435 15424 74435 15424 0 digitalL.g\[123\].u.OUTP
rlabel metal2 68784 14952 68784 14952 0 digitalL.g\[124\].u.OUTN
rlabel metal2 74035 15424 74035 15424 0 digitalL.g\[124\].u.OUTP
rlabel metal2 73056 16926 73056 16926 0 digitalL.g\[125\].u.OUTN
rlabel metal2 69888 15330 69888 15330 0 digitalL.g\[125\].u.OUTP
rlabel metal2 69504 15288 69504 15288 0 digitalL.g\[126\].u.OUTN
rlabel metal2 67392 15834 67392 15834 0 digitalL.g\[126\].u.OUTP
rlabel metal3 71856 15204 71856 15204 0 digitalL.g\[127\].u.OUTN
rlabel metal3 72321 15540 72321 15540 0 digitalL.g\[127\].u.OUTP
rlabel metal3 77856 7392 77856 7392 0 digitalL.g\[12\].u.OUTN
rlabel metal3 77280 7392 77280 7392 0 digitalL.g\[12\].u.OUTP
rlabel metal2 78336 7476 78336 7476 0 digitalL.g\[13\].u.OUTN
rlabel metal2 77952 8148 77952 8148 0 digitalL.g\[13\].u.OUTP
rlabel metal2 78336 6090 78336 6090 0 digitalL.g\[14\].u.OUTN
rlabel metal2 78288 6636 78288 6636 0 digitalL.g\[14\].u.OUTP
rlabel metal2 78816 8568 78816 8568 0 digitalL.g\[15\].u.OUTN
rlabel metal2 78768 7224 78768 7224 0 digitalL.g\[15\].u.OUTP
rlabel metal2 79104 7392 79104 7392 0 digitalL.g\[16\].u.OUTN
rlabel metal2 79104 6804 79104 6804 0 digitalL.g\[16\].u.OUTP
rlabel metal2 79536 7392 79536 7392 0 digitalL.g\[17\].u.OUTN
rlabel metal2 79392 6426 79392 6426 0 digitalL.g\[17\].u.OUTP
rlabel metal2 80016 6636 80016 6636 0 digitalL.g\[18\].u.OUTN
rlabel metal2 79872 8526 79872 8526 0 digitalL.g\[18\].u.OUTP
rlabel metal2 80304 5880 80304 5880 0 digitalL.g\[19\].u.OUTN
rlabel metal3 80242 9744 80242 9744 0 digitalL.g\[19\].u.OUTP
rlabel metal2 69792 9996 69792 9996 0 digitalL.g\[1\].u.OUTN
rlabel metal2 69216 9912 69216 9912 0 digitalL.g\[1\].u.OUTP
rlabel metal3 81312 7392 81312 7392 0 digitalL.g\[20\].u.OUTN
rlabel metal2 80736 6636 80736 6636 0 digitalL.g\[20\].u.OUTP
rlabel metal2 81225 9660 81225 9660 0 digitalL.g\[21\].u.OUTN
rlabel metal2 81072 6636 81072 6636 0 digitalL.g\[21\].u.OUTP
rlabel metal2 81696 8610 81696 8610 0 digitalL.g\[22\].u.OUTN
rlabel metal2 81504 8526 81504 8526 0 digitalL.g\[22\].u.OUTP
rlabel metal2 81552 6636 81552 6636 0 digitalL.g\[23\].u.OUTN
rlabel metal2 81888 6972 81888 6972 0 digitalL.g\[23\].u.OUTP
rlabel metal2 82368 8526 82368 8526 0 digitalL.g\[24\].u.OUTN
rlabel metal2 82320 6636 82320 6636 0 digitalL.g\[24\].u.OUTP
rlabel metal2 82992 7224 82992 7224 0 digitalL.g\[25\].u.OUTN
rlabel metal2 82656 6342 82656 6342 0 digitalL.g\[25\].u.OUTP
rlabel metal2 83232 7392 83232 7392 0 digitalL.g\[26\].u.OUTN
rlabel metal2 82944 6846 82944 6846 0 digitalL.g\[26\].u.OUTP
rlabel metal4 83616 7812 83616 7812 0 digitalL.g\[27\].u.OUTN
rlabel metal2 83520 6636 83520 6636 0 digitalL.g\[27\].u.OUTP
rlabel metal3 84000 7392 84000 7392 0 digitalL.g\[28\].u.OUTN
rlabel metal2 83952 6636 83952 6636 0 digitalL.g\[28\].u.OUTP
rlabel metal2 85728 7476 85728 7476 0 digitalL.g\[29\].u.OUTN
rlabel metal2 84336 6636 84336 6636 0 digitalL.g\[29\].u.OUTP
rlabel metal2 69504 9744 69504 9744 0 digitalL.g\[2\].u.OUTN
rlabel metal2 70752 9870 70752 9870 0 digitalL.g\[2\].u.OUTP
rlabel metal3 84768 7392 84768 7392 0 digitalL.g\[30\].u.OUTN
rlabel metal2 84816 6636 84816 6636 0 digitalL.g\[30\].u.OUTP
rlabel metal2 85056 6636 85056 6636 0 digitalL.g\[31\].u.OUTN
rlabel metal2 85056 8526 85056 8526 0 digitalL.g\[31\].u.OUTP
rlabel metal2 85633 9660 85633 9660 0 digitalL.g\[32\].u.OUTN
rlabel metal2 85488 6636 85488 6636 0 digitalL.g\[32\].u.OUTP
rlabel metal3 86496 6972 86496 6972 0 digitalL.g\[33\].u.OUTN
rlabel metal2 85824 8148 85824 8148 0 digitalL.g\[33\].u.OUTP
rlabel metal3 87072 7392 87072 7392 0 digitalL.g\[34\].u.OUTN
rlabel metal2 86352 6636 86352 6636 0 digitalL.g\[34\].u.OUTP
rlabel metal3 87216 7140 87216 7140 0 digitalL.g\[35\].u.OUTN
rlabel metal2 86784 7770 86784 7770 0 digitalL.g\[35\].u.OUTP
rlabel metal2 87744 8568 87744 8568 0 digitalL.g\[36\].u.OUTN
rlabel metal2 87072 7014 87072 7014 0 digitalL.g\[36\].u.OUTP
rlabel metal2 87648 7770 87648 7770 0 digitalL.g\[37\].u.OUTN
rlabel metal2 87456 6636 87456 6636 0 digitalL.g\[37\].u.OUTP
rlabel metal2 88992 7476 88992 7476 0 digitalL.g\[38\].u.OUTN
rlabel metal2 87936 8148 87936 8148 0 digitalL.g\[38\].u.OUTP
rlabel metal2 88425 9660 88425 9660 0 digitalL.g\[39\].u.OUTN
rlabel metal2 88272 6636 88272 6636 0 digitalL.g\[39\].u.OUTP
rlabel metal2 73584 7392 73584 7392 0 digitalL.g\[3\].u.OUTN
rlabel metal2 73925 9986 73925 9986 0 digitalL.g\[3\].u.OUTP
rlabel metal2 88800 6552 88800 6552 0 digitalL.g\[40\].u.OUTN
rlabel metal2 88800 8526 88800 8526 0 digitalL.g\[40\].u.OUTP
rlabel metal2 89280 8148 89280 8148 0 digitalL.g\[41\].u.OUTN
rlabel metal4 89088 7812 89088 7812 0 digitalL.g\[41\].u.OUTP
rlabel metal2 89712 5880 89712 5880 0 digitalL.g\[42\].u.OUTN
rlabel metal2 89520 6300 89520 6300 0 digitalL.g\[42\].u.OUTP
rlabel metal3 90336 7392 90336 7392 0 digitalL.g\[43\].u.OUTN
rlabel metal3 89760 7392 89760 7392 0 digitalL.g\[43\].u.OUTP
rlabel metal2 90432 8526 90432 8526 0 digitalL.g\[44\].u.OUTN
rlabel metal2 90240 7770 90240 7770 0 digitalL.g\[44\].u.OUTP
rlabel metal3 91392 7392 91392 7392 0 digitalL.g\[45\].u.OUTN
rlabel metal2 90576 6636 90576 6636 0 digitalL.g\[45\].u.OUTP
rlabel metal2 91296 7014 91296 7014 0 digitalL.g\[46\].u.OUTN
rlabel metal2 91104 7014 91104 7014 0 digitalL.g\[46\].u.OUTP
rlabel metal2 91632 5880 91632 5880 0 digitalL.g\[47\].u.OUTN
rlabel metal3 91488 7308 91488 7308 0 digitalL.g\[47\].u.OUTP
rlabel metal2 92544 6636 92544 6636 0 digitalL.g\[48\].u.OUTN
rlabel metal2 91920 6636 91920 6636 0 digitalL.g\[48\].u.OUTP
rlabel metal2 93312 7476 93312 7476 0 digitalL.g\[49\].u.OUTN
rlabel metal2 92304 6636 92304 6636 0 digitalL.g\[49\].u.OUTP
rlabel metal2 74435 9818 74435 9818 0 digitalL.g\[4\].u.OUTN
rlabel metal2 73824 8526 73824 8526 0 digitalL.g\[4\].u.OUTP
rlabel metal2 92832 7770 92832 7770 0 digitalL.g\[50\].u.OUTN
rlabel metal2 92928 8568 92928 8568 0 digitalL.g\[50\].u.OUTP
rlabel metal2 93168 5880 93168 5880 0 digitalL.g\[51\].u.OUTN
rlabel metal2 93216 8148 93216 8148 0 digitalL.g\[51\].u.OUTP
rlabel metal2 93552 5880 93552 5880 0 digitalL.g\[52\].u.OUTN
rlabel metal2 93600 8148 93600 8148 0 digitalL.g\[52\].u.OUTP
rlabel metal2 93984 6342 93984 6342 0 digitalL.g\[53\].u.OUTN
rlabel metal2 94128 6636 94128 6636 0 digitalL.g\[53\].u.OUTP
rlabel metal3 94128 6972 94128 6972 0 digitalL.g\[54\].u.OUTN
rlabel metal2 94272 8148 94272 8148 0 digitalL.g\[54\].u.OUTP
rlabel metal2 94848 8148 94848 8148 0 digitalL.g\[55\].u.OUTN
rlabel metal2 94752 8526 94752 8526 0 digitalL.g\[55\].u.OUTP
rlabel metal3 96096 6216 96096 6216 0 digitalL.g\[56\].u.OUTN
rlabel metal2 95088 7392 95088 7392 0 digitalL.g\[56\].u.OUTP
rlabel metal2 95616 8148 95616 8148 0 digitalL.g\[57\].u.OUTN
rlabel metal2 95474 9660 95474 9660 0 digitalL.g\[57\].u.OUTP
rlabel metal2 96048 5880 96048 5880 0 digitalL.g\[58\].u.OUTN
rlabel metal2 95760 5880 95760 5880 0 digitalL.g\[58\].u.OUTP
rlabel metal3 96672 7392 96672 7392 0 digitalL.g\[59\].u.OUTN
rlabel metal2 95904 8568 95904 8568 0 digitalL.g\[59\].u.OUTP
rlabel metal2 74208 7098 74208 7098 0 digitalL.g\[5\].u.OUTN
rlabel metal3 74976 7392 74976 7392 0 digitalL.g\[5\].u.OUTP
rlabel metal2 97152 7476 97152 7476 0 digitalL.g\[60\].u.OUTN
rlabel metal2 96672 6636 96672 6636 0 digitalL.g\[60\].u.OUTP
rlabel metal2 97392 6636 97392 6636 0 digitalL.g\[61\].u.OUTN
rlabel metal2 97104 6636 97104 6636 0 digitalL.g\[61\].u.OUTP
rlabel metal2 97728 8148 97728 8148 0 digitalL.g\[62\].u.OUTN
rlabel metal2 97440 8526 97440 8526 0 digitalL.g\[62\].u.OUTP
rlabel metal2 98112 8190 98112 8190 0 digitalL.g\[63\].u.OUTN
rlabel metal2 98016 8526 98016 8526 0 digitalL.g\[63\].u.OUTP
rlabel metal2 97925 15424 97925 15424 0 digitalL.g\[64\].u.OUTN
rlabel metal2 98035 15424 98035 15424 0 digitalL.g\[64\].u.OUTP
rlabel metal2 97525 15424 97525 15424 0 digitalL.g\[65\].u.OUTN
rlabel metal2 97635 15424 97635 15424 0 digitalL.g\[65\].u.OUTP
rlabel metal2 97125 15424 97125 15424 0 digitalL.g\[66\].u.OUTN
rlabel metal2 97235 15340 97235 15340 0 digitalL.g\[66\].u.OUTP
rlabel metal2 96725 15424 96725 15424 0 digitalL.g\[67\].u.OUTN
rlabel metal2 96835 15340 96835 15340 0 digitalL.g\[67\].u.OUTP
rlabel metal2 96325 15424 96325 15424 0 digitalL.g\[68\].u.OUTN
rlabel metal2 96435 15382 96435 15382 0 digitalL.g\[68\].u.OUTP
rlabel metal2 95952 18312 95952 18312 0 digitalL.g\[69\].u.OUTN
rlabel metal2 96035 15298 96035 15298 0 digitalL.g\[69\].u.OUTP
rlabel metal2 75120 6636 75120 6636 0 digitalL.g\[6\].u.OUTN
rlabel metal2 74928 6300 74928 6300 0 digitalL.g\[6\].u.OUTP
rlabel metal2 95525 15424 95525 15424 0 digitalL.g\[70\].u.OUTN
rlabel metal2 95635 15298 95635 15298 0 digitalL.g\[70\].u.OUTP
rlabel metal2 95125 15424 95125 15424 0 digitalL.g\[71\].u.OUTN
rlabel metal2 95235 15340 95235 15340 0 digitalL.g\[71\].u.OUTP
rlabel metal2 94725 15382 94725 15382 0 digitalL.g\[72\].u.OUTN
rlabel metal2 94835 15424 94835 15424 0 digitalL.g\[72\].u.OUTP
rlabel metal2 94325 15424 94325 15424 0 digitalL.g\[73\].u.OUTN
rlabel metal2 94435 15424 94435 15424 0 digitalL.g\[73\].u.OUTP
rlabel metal2 93925 15424 93925 15424 0 digitalL.g\[74\].u.OUTN
rlabel metal2 94035 15424 94035 15424 0 digitalL.g\[74\].u.OUTP
rlabel metal2 93525 15298 93525 15298 0 digitalL.g\[75\].u.OUTN
rlabel metal2 93635 15340 93635 15340 0 digitalL.g\[75\].u.OUTP
rlabel metal2 93125 15424 93125 15424 0 digitalL.g\[76\].u.OUTN
rlabel metal2 93235 15298 93235 15298 0 digitalL.g\[76\].u.OUTP
rlabel metal2 92725 15424 92725 15424 0 digitalL.g\[77\].u.OUTN
rlabel metal2 92835 15382 92835 15382 0 digitalL.g\[77\].u.OUTP
rlabel metal2 92325 15382 92325 15382 0 digitalL.g\[78\].u.OUTN
rlabel metal2 92435 15382 92435 15382 0 digitalL.g\[78\].u.OUTP
rlabel metal2 91925 15424 91925 15424 0 digitalL.g\[79\].u.OUTN
rlabel metal2 92035 15424 92035 15424 0 digitalL.g\[79\].u.OUTP
rlabel metal2 75552 7392 75552 7392 0 digitalL.g\[7\].u.OUTN
rlabel metal2 75168 5880 75168 5880 0 digitalL.g\[7\].u.OUTP
rlabel metal2 91525 15424 91525 15424 0 digitalL.g\[80\].u.OUTN
rlabel metal2 91635 15466 91635 15466 0 digitalL.g\[80\].u.OUTP
rlabel metal2 91125 15424 91125 15424 0 digitalL.g\[81\].u.OUTN
rlabel metal2 91235 15466 91235 15466 0 digitalL.g\[81\].u.OUTP
rlabel metal2 90624 16380 90624 16380 0 digitalL.g\[82\].u.OUTN
rlabel metal2 90835 15424 90835 15424 0 digitalL.g\[82\].u.OUTP
rlabel metal2 90325 15424 90325 15424 0 digitalL.g\[83\].u.OUTN
rlabel metal2 90435 15424 90435 15424 0 digitalL.g\[83\].u.OUTP
rlabel metal2 89925 15382 89925 15382 0 digitalL.g\[84\].u.OUTN
rlabel metal2 90035 15424 90035 15424 0 digitalL.g\[84\].u.OUTP
rlabel metal2 89525 15340 89525 15340 0 digitalL.g\[85\].u.OUTN
rlabel metal2 89635 15340 89635 15340 0 digitalL.g\[85\].u.OUTP
rlabel metal2 89125 15424 89125 15424 0 digitalL.g\[86\].u.OUTN
rlabel metal2 89235 15424 89235 15424 0 digitalL.g\[86\].u.OUTP
rlabel metal2 88725 15424 88725 15424 0 digitalL.g\[87\].u.OUTN
rlabel metal2 88835 15382 88835 15382 0 digitalL.g\[87\].u.OUTP
rlabel metal2 88325 15424 88325 15424 0 digitalL.g\[88\].u.OUTN
rlabel metal3 88320 17556 88320 17556 0 digitalL.g\[88\].u.OUTP
rlabel metal2 87925 15424 87925 15424 0 digitalL.g\[89\].u.OUTN
rlabel metal2 88035 15424 88035 15424 0 digitalL.g\[89\].u.OUTP
rlabel metal2 75936 6636 75936 6636 0 digitalL.g\[8\].u.OUTN
rlabel metal2 75936 8526 75936 8526 0 digitalL.g\[8\].u.OUTP
rlabel metal2 87525 15424 87525 15424 0 digitalL.g\[90\].u.OUTN
rlabel metal2 87635 15424 87635 15424 0 digitalL.g\[90\].u.OUTP
rlabel metal2 87125 15382 87125 15382 0 digitalL.g\[91\].u.OUTN
rlabel metal2 87235 15424 87235 15424 0 digitalL.g\[91\].u.OUTP
rlabel metal2 86725 15424 86725 15424 0 digitalL.g\[92\].u.OUTN
rlabel metal2 86835 15424 86835 15424 0 digitalL.g\[92\].u.OUTP
rlabel metal2 86325 15298 86325 15298 0 digitalL.g\[93\].u.OUTN
rlabel metal2 86435 15340 86435 15340 0 digitalL.g\[93\].u.OUTP
rlabel metal2 85925 15424 85925 15424 0 digitalL.g\[94\].u.OUTN
rlabel metal2 86035 15424 86035 15424 0 digitalL.g\[94\].u.OUTP
rlabel metal2 85525 15424 85525 15424 0 digitalL.g\[95\].u.OUTN
rlabel metal2 85635 15424 85635 15424 0 digitalL.g\[95\].u.OUTP
rlabel metal2 85125 15298 85125 15298 0 digitalL.g\[96\].u.OUTN
rlabel metal2 85152 16590 85152 16590 0 digitalL.g\[96\].u.OUTP
rlabel metal2 84725 15382 84725 15382 0 digitalL.g\[97\].u.OUTN
rlabel metal2 84835 15424 84835 15424 0 digitalL.g\[97\].u.OUTP
rlabel metal2 84325 15424 84325 15424 0 digitalL.g\[98\].u.OUTN
rlabel metal2 84435 15382 84435 15382 0 digitalL.g\[98\].u.OUTP
rlabel metal2 83925 15424 83925 15424 0 digitalL.g\[99\].u.OUTN
rlabel metal2 84035 15466 84035 15466 0 digitalL.g\[99\].u.OUTP
rlabel metal2 76320 6636 76320 6636 0 digitalL.g\[9\].u.OUTN
rlabel metal2 76320 8526 76320 8526 0 digitalL.g\[9\].u.OUTP
rlabel metal2 69216 25830 69216 25830 0 digitalenH.g\[0\].u.OUTN
rlabel metal3 70962 25872 70962 25872 0 digitalenH.g\[0\].u.OUTP
rlabel metal2 98657 25704 98657 25704 0 digitalenH.g\[1\].u.OUTN
rlabel metal2 98410 25620 98410 25620 0 digitalenH.g\[1\].u.OUTP
rlabel metal2 98325 31426 98325 31426 0 digitalenH.g\[2\].u.OUTN
rlabel metal2 98435 31468 98435 31468 0 digitalenH.g\[2\].u.OUTP
rlabel metal2 69696 31080 69696 31080 0 digitalenH.g\[3\].u.OUTN
rlabel metal2 72435 31384 72435 31384 0 digitalenH.g\[3\].u.OUTP
rlabel metal2 69888 9702 69888 9702 0 digitalenL.g\[0\].u.OUTN
rlabel metal2 69600 9744 69600 9744 0 digitalenL.g\[0\].u.OUTP
rlabel metal2 98784 7812 98784 7812 0 digitalenL.g\[1\].u.OUTN
rlabel metal2 98496 8526 98496 8526 0 digitalenL.g\[1\].u.OUTP
rlabel metal2 98592 5460 98592 5460 0 digitalenL.g\[2\].u.OUTN
rlabel metal2 97152 4872 97152 4872 0 digitalenL.g\[2\].u.OUTP
rlabel metal2 72114 15372 72114 15372 0 digitalenL.g\[3\].u.OUTN
rlabel metal3 72169 15372 72169 15372 0 digitalenL.g\[3\].u.OUTP
rlabel metal2 2016 19278 2016 19278 0 net1
rlabel metal2 864 13314 864 13314 0 net10
rlabel metal2 95904 5670 95904 5670 0 net100
rlabel metal2 96672 7266 96672 7266 0 net101
rlabel metal3 94224 7224 94224 7224 0 net102
rlabel metal2 95712 6552 95712 6552 0 net103
rlabel metal2 87072 18522 87072 18522 0 net104
rlabel metal2 88416 19236 88416 19236 0 net105
rlabel metal3 91632 18480 91632 18480 0 net106
rlabel metal2 91296 18522 91296 18522 0 net107
rlabel metal2 89952 19488 89952 19488 0 net108
rlabel metal2 92928 19362 92928 19362 0 net109
rlabel metal3 1104 14196 1104 14196 0 net11
rlabel metal2 93936 18480 93936 18480 0 net110
rlabel metal2 96672 17892 96672 17892 0 net111
rlabel metal3 98304 17808 98304 17808 0 net112
rlabel metal2 97152 18102 97152 18102 0 net113
rlabel metal2 89952 19278 89952 19278 0 net114
rlabel metal5 86648 19320 86648 19320 0 net115
rlabel metal3 73248 7224 73248 7224 0 net116
rlabel metal2 1536 9828 1536 9828 0 net117
rlabel metal3 366 15708 366 15708 0 net118
rlabel metal3 366 16548 366 16548 0 net119
rlabel metal3 1296 14952 1296 14952 0 net12
rlabel metal3 366 17388 366 17388 0 net120
rlabel metal3 366 18228 366 18228 0 net121
rlabel metal3 366 19068 366 19068 0 net122
rlabel metal3 366 19908 366 19908 0 net123
rlabel metal3 366 20748 366 20748 0 net124
rlabel metal3 366 21588 366 21588 0 net125
rlabel metal2 816 2688 816 2688 0 net13
rlabel metal2 912 3360 912 3360 0 net14
rlabel metal3 1248 4200 1248 4200 0 net15
rlabel metal2 864 5166 864 5166 0 net16
rlabel metal2 864 5754 864 5754 0 net17
rlabel metal3 1104 6636 1104 6636 0 net18
rlabel metal2 864 7854 864 7854 0 net19
rlabel metal3 1488 23772 1488 23772 0 net2
rlabel metal2 864 8778 864 8778 0 net20
rlabel metal2 69696 25200 69696 25200 0 net21
rlabel metal3 71280 25284 71280 25284 0 net22
rlabel metal2 69792 31752 69792 31752 0 net23
rlabel metal2 68064 28812 68064 28812 0 net24
rlabel metal2 76608 22176 76608 22176 0 net25
rlabel metal3 79104 21504 79104 21504 0 net26
rlabel metal2 79008 22974 79008 22974 0 net27
rlabel metal2 77856 22932 77856 22932 0 net28
rlabel metal3 78000 22260 78000 22260 0 net29
rlabel metal2 960 22974 960 22974 0 net3
rlabel metal2 82464 23058 82464 23058 0 net30
rlabel via2 82656 22344 82656 22344 0 net31
rlabel metal2 83520 22302 83520 22302 0 net32
rlabel metal2 83520 22932 83520 22932 0 net33
rlabel metal2 83808 23100 83808 23100 0 net34
rlabel metal2 76752 35196 76752 35196 0 net35
rlabel metal2 79776 34818 79776 34818 0 net36
rlabel metal2 79008 35952 79008 35952 0 net37
rlabel metal3 78048 35112 78048 35112 0 net38
rlabel metal2 77568 34314 77568 34314 0 net39
rlabel metal3 70608 26040 70608 26040 0 net4
rlabel metal3 82656 35070 82656 35070 0 net40
rlabel metal2 82272 34487 82272 34487 0 net41
rlabel metal2 84288 35154 84288 35154 0 net42
rlabel metal2 84672 34398 84672 34398 0 net43
rlabel metal3 84096 34440 84096 34440 0 net44
rlabel metal2 86112 22848 86112 22848 0 net45
rlabel metal2 88512 22974 88512 22974 0 net46
rlabel metal2 91872 22386 91872 22386 0 net47
rlabel metal2 91296 22428 91296 22428 0 net48
rlabel metal2 90912 22218 90912 22218 0 net49
rlabel metal2 864 9366 864 9366 0 net5
rlabel metal2 94176 22302 94176 22302 0 net50
rlabel metal2 93456 21588 93456 21588 0 net51
rlabel metal2 97440 23016 97440 23016 0 net52
rlabel metal3 98016 23100 98016 23100 0 net53
rlabel metal2 93504 22386 93504 22386 0 net54
rlabel metal3 87264 35112 87264 35112 0 net55
rlabel metal2 88128 35616 88128 35616 0 net56
rlabel metal2 90048 35868 90048 35868 0 net57
rlabel metal2 91200 34482 91200 34482 0 net58
rlabel metal2 91008 34356 91008 34356 0 net59
rlabel metal2 864 10290 864 10290 0 net6
rlabel metal2 93600 34314 93600 34314 0 net60
rlabel metal2 94032 34944 94032 34944 0 net61
rlabel metal3 98592 34356 98592 34356 0 net62
rlabel metal2 97056 34398 97056 34398 0 net63
rlabel metal2 94224 35112 94224 35112 0 net64
rlabel metal2 91680 23100 91680 23100 0 net65
rlabel metal3 71808 32802 71808 32802 0 net66
rlabel metal2 2016 5838 2016 5838 0 net67
rlabel metal2 73344 7182 73344 7182 0 net68
rlabel metal3 70608 18564 70608 18564 0 net69
rlabel metal2 864 10878 864 10878 0 net7
rlabel metal3 68784 15540 68784 15540 0 net70
rlabel metal2 74592 5964 74592 5964 0 net71
rlabel metal3 74640 6972 74640 6972 0 net72
rlabel metal2 78192 5628 78192 5628 0 net73
rlabel metal2 79680 7266 79680 7266 0 net74
rlabel metal2 79104 7182 79104 7182 0 net75
rlabel metal2 75744 6720 75744 6720 0 net76
rlabel metal2 80784 5628 80784 5628 0 net77
rlabel metal2 82752 6048 82752 6048 0 net78
rlabel metal2 84864 7182 84864 7182 0 net79
rlabel metal3 1248 11760 1248 11760 0 net8
rlabel metal2 86112 6468 86112 6468 0 net80
rlabel metal2 80736 7266 80736 7266 0 net81
rlabel metal3 74832 7308 74832 7308 0 net82
rlabel metal2 75648 19026 75648 19026 0 net83
rlabel metal2 75168 18774 75168 18774 0 net84
rlabel metal2 77760 17766 77760 17766 0 net85
rlabel metal2 78816 18438 78816 18438 0 net86
rlabel metal2 79008 18354 79008 18354 0 net87
rlabel metal2 80352 19152 80352 19152 0 net88
rlabel metal2 82272 18102 82272 18102 0 net89
rlabel metal3 1440 11928 1440 11928 0 net9
rlabel metal2 83856 18480 83856 18480 0 net90
rlabel metal2 85920 18774 85920 18774 0 net91
rlabel metal3 84864 19320 84864 19320 0 net92
rlabel metal2 87264 7224 87264 7224 0 net93
rlabel metal3 88464 7224 88464 7224 0 net94
rlabel metal2 89856 7056 89856 7056 0 net95
rlabel metal2 91584 7098 91584 7098 0 net96
rlabel metal2 90048 7140 90048 7140 0 net97
rlabel metal2 93120 7266 93120 7266 0 net98
rlabel metal3 94272 6384 94272 6384 0 net99
rlabel metal3 318 22428 318 22428 0 ui_in[0]
rlabel metal3 366 23268 366 23268 0 ui_in[1]
rlabel metal3 366 24108 366 24108 0 ui_in[2]
rlabel metal3 366 24948 366 24948 0 ui_in[3]
rlabel metal3 366 8988 366 8988 0 uio_out[0]
rlabel metal3 366 9828 366 9828 0 uio_out[1]
rlabel metal3 366 10668 366 10668 0 uio_out[2]
rlabel metal3 366 11508 366 11508 0 uio_out[3]
rlabel metal3 366 12348 366 12348 0 uio_out[4]
rlabel metal3 366 13188 366 13188 0 uio_out[5]
rlabel metal3 366 14028 366 14028 0 uio_out[6]
rlabel metal3 366 14868 366 14868 0 uio_out[7]
rlabel metal3 366 2268 366 2268 0 uo_out[0]
rlabel metal3 366 3108 366 3108 0 uo_out[1]
rlabel metal3 366 3948 366 3948 0 uo_out[2]
rlabel metal3 366 4788 366 4788 0 uo_out[3]
rlabel metal3 366 5628 366 5628 0 uo_out[4]
rlabel metal3 366 6468 366 6468 0 uo_out[5]
rlabel metal3 366 7308 366 7308 0 uo_out[6]
rlabel metal3 366 8148 366 8148 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
