module heichips25_pudding (VGND,
    VPWR,
    clk,
    ena,
    i_in,
    i_out,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 inout VGND;
 inout VPWR;
 input clk;
 input ena;
 inout i_in;
 inout i_out;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire \bias[0] ;
 wire \bias[1] ;
 wire \daisychain[0] ;
 wire \daisychain[100] ;
 wire \daisychain[101] ;
 wire \daisychain[102] ;
 wire \daisychain[103] ;
 wire \daisychain[104] ;
 wire \daisychain[105] ;
 wire \daisychain[106] ;
 wire \daisychain[107] ;
 wire \daisychain[108] ;
 wire \daisychain[109] ;
 wire \daisychain[10] ;
 wire \daisychain[110] ;
 wire \daisychain[111] ;
 wire \daisychain[112] ;
 wire \daisychain[113] ;
 wire \daisychain[114] ;
 wire \daisychain[115] ;
 wire \daisychain[116] ;
 wire \daisychain[117] ;
 wire \daisychain[118] ;
 wire \daisychain[119] ;
 wire \daisychain[11] ;
 wire \daisychain[120] ;
 wire \daisychain[121] ;
 wire \daisychain[122] ;
 wire \daisychain[123] ;
 wire \daisychain[124] ;
 wire \daisychain[125] ;
 wire \daisychain[126] ;
 wire \daisychain[127] ;
 wire \daisychain[12] ;
 wire \daisychain[13] ;
 wire \daisychain[14] ;
 wire \daisychain[15] ;
 wire \daisychain[16] ;
 wire \daisychain[17] ;
 wire \daisychain[18] ;
 wire \daisychain[19] ;
 wire \daisychain[1] ;
 wire \daisychain[20] ;
 wire \daisychain[21] ;
 wire \daisychain[22] ;
 wire \daisychain[23] ;
 wire \daisychain[24] ;
 wire \daisychain[25] ;
 wire \daisychain[26] ;
 wire \daisychain[27] ;
 wire \daisychain[28] ;
 wire \daisychain[29] ;
 wire \daisychain[2] ;
 wire \daisychain[30] ;
 wire \daisychain[31] ;
 wire \daisychain[32] ;
 wire \daisychain[33] ;
 wire \daisychain[34] ;
 wire \daisychain[35] ;
 wire \daisychain[36] ;
 wire \daisychain[37] ;
 wire \daisychain[38] ;
 wire \daisychain[39] ;
 wire \daisychain[3] ;
 wire \daisychain[40] ;
 wire \daisychain[41] ;
 wire \daisychain[42] ;
 wire \daisychain[43] ;
 wire \daisychain[44] ;
 wire \daisychain[45] ;
 wire \daisychain[46] ;
 wire \daisychain[47] ;
 wire \daisychain[48] ;
 wire \daisychain[49] ;
 wire \daisychain[4] ;
 wire \daisychain[50] ;
 wire \daisychain[51] ;
 wire \daisychain[52] ;
 wire \daisychain[53] ;
 wire \daisychain[54] ;
 wire \daisychain[55] ;
 wire \daisychain[56] ;
 wire \daisychain[57] ;
 wire \daisychain[58] ;
 wire \daisychain[59] ;
 wire \daisychain[5] ;
 wire \daisychain[60] ;
 wire \daisychain[61] ;
 wire \daisychain[62] ;
 wire \daisychain[63] ;
 wire \daisychain[64] ;
 wire \daisychain[65] ;
 wire \daisychain[66] ;
 wire \daisychain[67] ;
 wire \daisychain[68] ;
 wire \daisychain[69] ;
 wire \daisychain[6] ;
 wire \daisychain[70] ;
 wire \daisychain[71] ;
 wire \daisychain[72] ;
 wire \daisychain[73] ;
 wire \daisychain[74] ;
 wire \daisychain[75] ;
 wire \daisychain[76] ;
 wire \daisychain[77] ;
 wire \daisychain[78] ;
 wire \daisychain[79] ;
 wire \daisychain[7] ;
 wire \daisychain[80] ;
 wire \daisychain[81] ;
 wire \daisychain[82] ;
 wire \daisychain[83] ;
 wire \daisychain[84] ;
 wire \daisychain[85] ;
 wire \daisychain[86] ;
 wire \daisychain[87] ;
 wire \daisychain[88] ;
 wire \daisychain[89] ;
 wire \daisychain[8] ;
 wire \daisychain[90] ;
 wire \daisychain[91] ;
 wire \daisychain[92] ;
 wire \daisychain[93] ;
 wire \daisychain[94] ;
 wire \daisychain[95] ;
 wire \daisychain[96] ;
 wire \daisychain[97] ;
 wire \daisychain[98] ;
 wire \daisychain[99] ;
 wire \daisychain[9] ;
 wire \digitalen.g[0].u.OUTN ;
 wire \digitalen.g[0].u.OUTP ;
 wire \digitalen.g[1].u.OUTN ;
 wire \digitalen.g[1].u.OUTP ;
 wire \digitalen.g[2].u.OUTN ;
 wire \digitalen.g[2].u.OUTP ;
 wire \digitalen.g[3].u.OUTN ;
 wire \digitalen.g[3].u.OUTP ;
 wire net1;
 wire \state[0] ;
 wire \state[100] ;
 wire \state[101] ;
 wire \state[102] ;
 wire \state[103] ;
 wire \state[104] ;
 wire \state[105] ;
 wire \state[106] ;
 wire \state[107] ;
 wire \state[108] ;
 wire \state[109] ;
 wire \state[10] ;
 wire \state[110] ;
 wire \state[111] ;
 wire \state[112] ;
 wire \state[113] ;
 wire \state[114] ;
 wire \state[115] ;
 wire \state[116] ;
 wire \state[117] ;
 wire \state[118] ;
 wire \state[119] ;
 wire \state[11] ;
 wire \state[120] ;
 wire \state[121] ;
 wire \state[122] ;
 wire \state[123] ;
 wire \state[124] ;
 wire \state[125] ;
 wire \state[126] ;
 wire \state[127] ;
 wire \state[12] ;
 wire \state[13] ;
 wire \state[14] ;
 wire \state[15] ;
 wire \state[16] ;
 wire \state[17] ;
 wire \state[18] ;
 wire \state[19] ;
 wire \state[1] ;
 wire \state[20] ;
 wire \state[21] ;
 wire \state[22] ;
 wire \state[23] ;
 wire \state[24] ;
 wire \state[25] ;
 wire \state[26] ;
 wire \state[27] ;
 wire \state[28] ;
 wire \state[29] ;
 wire \state[2] ;
 wire \state[30] ;
 wire \state[31] ;
 wire \state[32] ;
 wire \state[33] ;
 wire \state[34] ;
 wire \state[35] ;
 wire \state[36] ;
 wire \state[37] ;
 wire \state[38] ;
 wire \state[39] ;
 wire \state[3] ;
 wire \state[40] ;
 wire \state[41] ;
 wire \state[42] ;
 wire \state[43] ;
 wire \state[44] ;
 wire \state[45] ;
 wire \state[46] ;
 wire \state[47] ;
 wire \state[48] ;
 wire \state[49] ;
 wire \state[4] ;
 wire \state[50] ;
 wire \state[51] ;
 wire \state[52] ;
 wire \state[53] ;
 wire \state[54] ;
 wire \state[55] ;
 wire \state[56] ;
 wire \state[57] ;
 wire \state[58] ;
 wire \state[59] ;
 wire \state[5] ;
 wire \state[60] ;
 wire \state[61] ;
 wire \state[62] ;
 wire \state[63] ;
 wire \state[64] ;
 wire \state[65] ;
 wire \state[66] ;
 wire \state[67] ;
 wire \state[68] ;
 wire \state[69] ;
 wire \state[6] ;
 wire \state[70] ;
 wire \state[71] ;
 wire \state[72] ;
 wire \state[73] ;
 wire \state[74] ;
 wire \state[75] ;
 wire \state[76] ;
 wire \state[77] ;
 wire \state[78] ;
 wire \state[79] ;
 wire \state[7] ;
 wire \state[80] ;
 wire \state[81] ;
 wire \state[82] ;
 wire \state[83] ;
 wire \state[84] ;
 wire \state[85] ;
 wire \state[86] ;
 wire \state[87] ;
 wire \state[88] ;
 wire \state[89] ;
 wire \state[8] ;
 wire \state[90] ;
 wire \state[91] ;
 wire \state[92] ;
 wire \state[93] ;
 wire \state[94] ;
 wire \state[95] ;
 wire \state[96] ;
 wire \state[97] ;
 wire \state[98] ;
 wire \state[99] ;
 wire \state[9] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire clknet_leaf_0_clk;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_inv_1 _1284_ (.VDD(VPWR),
    .Y(_0030_),
    .A(\state[127] ),
    .VSS(VGND));
 sg13g2_inv_1 _1285_ (.VDD(VPWR),
    .Y(_0846_),
    .A(net156),
    .VSS(VGND));
 sg13g2_inv_1 _1286_ (.VDD(VPWR),
    .Y(_0029_),
    .A(\state[126] ),
    .VSS(VGND));
 sg13g2_inv_1 _1287_ (.VDD(VPWR),
    .Y(_0028_),
    .A(\state[125] ),
    .VSS(VGND));
 sg13g2_inv_1 _1288_ (.VDD(VPWR),
    .Y(_0027_),
    .A(\state[124] ),
    .VSS(VGND));
 sg13g2_inv_1 _1289_ (.VDD(VPWR),
    .Y(_0026_),
    .A(\state[123] ),
    .VSS(VGND));
 sg13g2_inv_1 _1290_ (.VDD(VPWR),
    .Y(_0025_),
    .A(\state[122] ),
    .VSS(VGND));
 sg13g2_inv_1 _1291_ (.VDD(VPWR),
    .Y(_0024_),
    .A(\state[121] ),
    .VSS(VGND));
 sg13g2_inv_1 _1292_ (.VDD(VPWR),
    .Y(_0023_),
    .A(\state[120] ),
    .VSS(VGND));
 sg13g2_inv_1 _1293_ (.VDD(VPWR),
    .Y(_0021_),
    .A(\state[119] ),
    .VSS(VGND));
 sg13g2_inv_1 _1294_ (.VDD(VPWR),
    .Y(_0020_),
    .A(\state[118] ),
    .VSS(VGND));
 sg13g2_inv_1 _1295_ (.VDD(VPWR),
    .Y(_0019_),
    .A(\state[117] ),
    .VSS(VGND));
 sg13g2_inv_1 _1296_ (.VDD(VPWR),
    .Y(_0018_),
    .A(\state[116] ),
    .VSS(VGND));
 sg13g2_inv_1 _1297_ (.VDD(VPWR),
    .Y(_0017_),
    .A(\state[115] ),
    .VSS(VGND));
 sg13g2_inv_1 _1298_ (.VDD(VPWR),
    .Y(_0016_),
    .A(\state[114] ),
    .VSS(VGND));
 sg13g2_inv_1 _1299_ (.VDD(VPWR),
    .Y(_0015_),
    .A(\state[113] ),
    .VSS(VGND));
 sg13g2_inv_1 _1300_ (.VDD(VPWR),
    .Y(_0014_),
    .A(\state[112] ),
    .VSS(VGND));
 sg13g2_inv_1 _1301_ (.VDD(VPWR),
    .Y(_0013_),
    .A(\state[111] ),
    .VSS(VGND));
 sg13g2_inv_1 _1302_ (.VDD(VPWR),
    .Y(_0012_),
    .A(\state[110] ),
    .VSS(VGND));
 sg13g2_inv_1 _1303_ (.VDD(VPWR),
    .Y(_0010_),
    .A(\state[109] ),
    .VSS(VGND));
 sg13g2_inv_1 _1304_ (.VDD(VPWR),
    .Y(_0009_),
    .A(\state[108] ),
    .VSS(VGND));
 sg13g2_inv_1 _1305_ (.VDD(VPWR),
    .Y(_0008_),
    .A(\state[107] ),
    .VSS(VGND));
 sg13g2_inv_1 _1306_ (.VDD(VPWR),
    .Y(_0007_),
    .A(\state[106] ),
    .VSS(VGND));
 sg13g2_inv_1 _1307_ (.VDD(VPWR),
    .Y(_0006_),
    .A(\state[105] ),
    .VSS(VGND));
 sg13g2_inv_1 _1308_ (.VDD(VPWR),
    .Y(_0005_),
    .A(\state[104] ),
    .VSS(VGND));
 sg13g2_inv_1 _1309_ (.VDD(VPWR),
    .Y(_0004_),
    .A(\state[103] ),
    .VSS(VGND));
 sg13g2_inv_1 _1310_ (.VDD(VPWR),
    .Y(_0003_),
    .A(\state[102] ),
    .VSS(VGND));
 sg13g2_inv_1 _1311_ (.VDD(VPWR),
    .Y(_0002_),
    .A(\state[101] ),
    .VSS(VGND));
 sg13g2_inv_1 _1312_ (.VDD(VPWR),
    .Y(_0001_),
    .A(\state[100] ),
    .VSS(VGND));
 sg13g2_inv_1 _1313_ (.VDD(VPWR),
    .Y(_0126_),
    .A(\state[99] ),
    .VSS(VGND));
 sg13g2_inv_1 _1314_ (.VDD(VPWR),
    .Y(_0125_),
    .A(\state[98] ),
    .VSS(VGND));
 sg13g2_inv_1 _1315_ (.VDD(VPWR),
    .Y(_0124_),
    .A(\state[97] ),
    .VSS(VGND));
 sg13g2_inv_1 _1316_ (.VDD(VPWR),
    .Y(_0123_),
    .A(\state[96] ),
    .VSS(VGND));
 sg13g2_inv_1 _1317_ (.VDD(VPWR),
    .Y(_0122_),
    .A(\state[95] ),
    .VSS(VGND));
 sg13g2_inv_1 _1318_ (.VDD(VPWR),
    .Y(_0121_),
    .A(\state[94] ),
    .VSS(VGND));
 sg13g2_inv_1 _1319_ (.VDD(VPWR),
    .Y(_0120_),
    .A(\state[93] ),
    .VSS(VGND));
 sg13g2_inv_1 _1320_ (.VDD(VPWR),
    .Y(_0119_),
    .A(\state[92] ),
    .VSS(VGND));
 sg13g2_inv_1 _1321_ (.VDD(VPWR),
    .Y(_0118_),
    .A(\state[91] ),
    .VSS(VGND));
 sg13g2_inv_1 _1322_ (.VDD(VPWR),
    .Y(_0117_),
    .A(\state[90] ),
    .VSS(VGND));
 sg13g2_inv_1 _1323_ (.VDD(VPWR),
    .Y(_0115_),
    .A(\state[89] ),
    .VSS(VGND));
 sg13g2_inv_1 _1324_ (.VDD(VPWR),
    .Y(_0114_),
    .A(\state[88] ),
    .VSS(VGND));
 sg13g2_inv_1 _1325_ (.VDD(VPWR),
    .Y(_0113_),
    .A(\state[87] ),
    .VSS(VGND));
 sg13g2_inv_1 _1326_ (.VDD(VPWR),
    .Y(_0112_),
    .A(\state[86] ),
    .VSS(VGND));
 sg13g2_inv_1 _1327_ (.VDD(VPWR),
    .Y(_0111_),
    .A(\state[85] ),
    .VSS(VGND));
 sg13g2_inv_1 _1328_ (.VDD(VPWR),
    .Y(_0110_),
    .A(\state[84] ),
    .VSS(VGND));
 sg13g2_inv_1 _1329_ (.VDD(VPWR),
    .Y(_0109_),
    .A(\state[83] ),
    .VSS(VGND));
 sg13g2_inv_1 _1330_ (.VDD(VPWR),
    .Y(_0108_),
    .A(\state[82] ),
    .VSS(VGND));
 sg13g2_inv_1 _1331_ (.VDD(VPWR),
    .Y(_0107_),
    .A(\state[81] ),
    .VSS(VGND));
 sg13g2_inv_1 _1332_ (.VDD(VPWR),
    .Y(_0106_),
    .A(\state[80] ),
    .VSS(VGND));
 sg13g2_inv_1 _1333_ (.VDD(VPWR),
    .Y(_0104_),
    .A(\state[79] ),
    .VSS(VGND));
 sg13g2_inv_1 _1334_ (.VDD(VPWR),
    .Y(_0103_),
    .A(\state[78] ),
    .VSS(VGND));
 sg13g2_inv_1 _1335_ (.VDD(VPWR),
    .Y(_0102_),
    .A(\state[77] ),
    .VSS(VGND));
 sg13g2_inv_1 _1336_ (.VDD(VPWR),
    .Y(_0101_),
    .A(\state[76] ),
    .VSS(VGND));
 sg13g2_inv_1 _1337_ (.VDD(VPWR),
    .Y(_0100_),
    .A(\state[75] ),
    .VSS(VGND));
 sg13g2_inv_1 _1338_ (.VDD(VPWR),
    .Y(_0099_),
    .A(\state[74] ),
    .VSS(VGND));
 sg13g2_inv_1 _1339_ (.VDD(VPWR),
    .Y(_0098_),
    .A(\state[73] ),
    .VSS(VGND));
 sg13g2_inv_1 _1340_ (.VDD(VPWR),
    .Y(_0097_),
    .A(\state[72] ),
    .VSS(VGND));
 sg13g2_inv_1 _1341_ (.VDD(VPWR),
    .Y(_0096_),
    .A(\state[71] ),
    .VSS(VGND));
 sg13g2_inv_1 _1342_ (.VDD(VPWR),
    .Y(_0095_),
    .A(\state[70] ),
    .VSS(VGND));
 sg13g2_inv_1 _1343_ (.VDD(VPWR),
    .Y(_0093_),
    .A(\state[69] ),
    .VSS(VGND));
 sg13g2_inv_1 _1344_ (.VDD(VPWR),
    .Y(_0092_),
    .A(\state[68] ),
    .VSS(VGND));
 sg13g2_inv_1 _1345_ (.VDD(VPWR),
    .Y(_0091_),
    .A(\state[67] ),
    .VSS(VGND));
 sg13g2_inv_1 _1346_ (.VDD(VPWR),
    .Y(_0090_),
    .A(\state[66] ),
    .VSS(VGND));
 sg13g2_inv_1 _1347_ (.VDD(VPWR),
    .Y(_0089_),
    .A(\state[65] ),
    .VSS(VGND));
 sg13g2_inv_1 _1348_ (.VDD(VPWR),
    .Y(_0088_),
    .A(\state[64] ),
    .VSS(VGND));
 sg13g2_inv_1 _1349_ (.VDD(VPWR),
    .Y(_0087_),
    .A(\state[63] ),
    .VSS(VGND));
 sg13g2_inv_1 _1350_ (.VDD(VPWR),
    .Y(_0086_),
    .A(\state[62] ),
    .VSS(VGND));
 sg13g2_inv_1 _1351_ (.VDD(VPWR),
    .Y(_0085_),
    .A(\state[61] ),
    .VSS(VGND));
 sg13g2_inv_1 _1352_ (.VDD(VPWR),
    .Y(_0084_),
    .A(\state[60] ),
    .VSS(VGND));
 sg13g2_inv_1 _1353_ (.VDD(VPWR),
    .Y(_0082_),
    .A(\state[59] ),
    .VSS(VGND));
 sg13g2_inv_1 _1354_ (.VDD(VPWR),
    .Y(_0081_),
    .A(\state[58] ),
    .VSS(VGND));
 sg13g2_inv_1 _1355_ (.VDD(VPWR),
    .Y(_0080_),
    .A(\state[57] ),
    .VSS(VGND));
 sg13g2_inv_1 _1356_ (.VDD(VPWR),
    .Y(_0079_),
    .A(\state[56] ),
    .VSS(VGND));
 sg13g2_inv_1 _1357_ (.VDD(VPWR),
    .Y(_0078_),
    .A(\state[55] ),
    .VSS(VGND));
 sg13g2_inv_1 _1358_ (.VDD(VPWR),
    .Y(_0077_),
    .A(\state[54] ),
    .VSS(VGND));
 sg13g2_inv_1 _1359_ (.VDD(VPWR),
    .Y(_0076_),
    .A(\state[53] ),
    .VSS(VGND));
 sg13g2_inv_1 _1360_ (.VDD(VPWR),
    .Y(_0075_),
    .A(\state[52] ),
    .VSS(VGND));
 sg13g2_inv_1 _1361_ (.VDD(VPWR),
    .Y(_0074_),
    .A(\state[51] ),
    .VSS(VGND));
 sg13g2_inv_1 _1362_ (.VDD(VPWR),
    .Y(_0073_),
    .A(\state[50] ),
    .VSS(VGND));
 sg13g2_inv_1 _1363_ (.VDD(VPWR),
    .Y(_0071_),
    .A(\state[49] ),
    .VSS(VGND));
 sg13g2_inv_1 _1364_ (.VDD(VPWR),
    .Y(_0070_),
    .A(\state[48] ),
    .VSS(VGND));
 sg13g2_inv_1 _1365_ (.VDD(VPWR),
    .Y(_0069_),
    .A(\state[47] ),
    .VSS(VGND));
 sg13g2_inv_1 _1366_ (.VDD(VPWR),
    .Y(_0068_),
    .A(\state[46] ),
    .VSS(VGND));
 sg13g2_inv_1 _1367_ (.VDD(VPWR),
    .Y(_0067_),
    .A(\state[45] ),
    .VSS(VGND));
 sg13g2_inv_1 _1368_ (.VDD(VPWR),
    .Y(_0066_),
    .A(\state[44] ),
    .VSS(VGND));
 sg13g2_inv_1 _1369_ (.VDD(VPWR),
    .Y(_0065_),
    .A(\state[43] ),
    .VSS(VGND));
 sg13g2_inv_1 _1370_ (.VDD(VPWR),
    .Y(_0064_),
    .A(\state[42] ),
    .VSS(VGND));
 sg13g2_inv_1 _1371_ (.VDD(VPWR),
    .Y(_0063_),
    .A(\state[41] ),
    .VSS(VGND));
 sg13g2_inv_1 _1372_ (.VDD(VPWR),
    .Y(_0062_),
    .A(\state[40] ),
    .VSS(VGND));
 sg13g2_inv_1 _1373_ (.VDD(VPWR),
    .Y(_0060_),
    .A(\state[39] ),
    .VSS(VGND));
 sg13g2_inv_1 _1374_ (.VDD(VPWR),
    .Y(_0059_),
    .A(\state[38] ),
    .VSS(VGND));
 sg13g2_inv_1 _1375_ (.VDD(VPWR),
    .Y(_0058_),
    .A(\state[37] ),
    .VSS(VGND));
 sg13g2_inv_1 _1376_ (.VDD(VPWR),
    .Y(_0057_),
    .A(\state[36] ),
    .VSS(VGND));
 sg13g2_inv_1 _1377_ (.VDD(VPWR),
    .Y(_0056_),
    .A(\state[35] ),
    .VSS(VGND));
 sg13g2_inv_1 _1378_ (.VDD(VPWR),
    .Y(_0055_),
    .A(\state[34] ),
    .VSS(VGND));
 sg13g2_inv_1 _1379_ (.VDD(VPWR),
    .Y(_0054_),
    .A(\state[33] ),
    .VSS(VGND));
 sg13g2_inv_1 _1380_ (.VDD(VPWR),
    .Y(_0053_),
    .A(\state[32] ),
    .VSS(VGND));
 sg13g2_inv_1 _1381_ (.VDD(VPWR),
    .Y(_0052_),
    .A(\state[31] ),
    .VSS(VGND));
 sg13g2_inv_1 _1382_ (.VDD(VPWR),
    .Y(_0051_),
    .A(\state[30] ),
    .VSS(VGND));
 sg13g2_inv_1 _1383_ (.VDD(VPWR),
    .Y(_0049_),
    .A(\state[29] ),
    .VSS(VGND));
 sg13g2_inv_1 _1384_ (.VDD(VPWR),
    .Y(_0048_),
    .A(\state[28] ),
    .VSS(VGND));
 sg13g2_inv_1 _1385_ (.VDD(VPWR),
    .Y(_0047_),
    .A(\state[27] ),
    .VSS(VGND));
 sg13g2_inv_1 _1386_ (.VDD(VPWR),
    .Y(_0046_),
    .A(\state[26] ),
    .VSS(VGND));
 sg13g2_inv_1 _1387_ (.VDD(VPWR),
    .Y(_0045_),
    .A(\state[25] ),
    .VSS(VGND));
 sg13g2_inv_1 _1388_ (.VDD(VPWR),
    .Y(_0044_),
    .A(\state[24] ),
    .VSS(VGND));
 sg13g2_inv_1 _1389_ (.VDD(VPWR),
    .Y(_0043_),
    .A(\state[23] ),
    .VSS(VGND));
 sg13g2_inv_1 _1390_ (.VDD(VPWR),
    .Y(_0042_),
    .A(\state[22] ),
    .VSS(VGND));
 sg13g2_inv_1 _1391_ (.VDD(VPWR),
    .Y(_0041_),
    .A(\state[21] ),
    .VSS(VGND));
 sg13g2_inv_1 _1392_ (.VDD(VPWR),
    .Y(_0040_),
    .A(\state[20] ),
    .VSS(VGND));
 sg13g2_inv_1 _1393_ (.VDD(VPWR),
    .Y(_0038_),
    .A(\state[19] ),
    .VSS(VGND));
 sg13g2_inv_1 _1394_ (.VDD(VPWR),
    .Y(_0037_),
    .A(\state[18] ),
    .VSS(VGND));
 sg13g2_inv_1 _1395_ (.VDD(VPWR),
    .Y(_0036_),
    .A(\state[17] ),
    .VSS(VGND));
 sg13g2_inv_1 _1396_ (.VDD(VPWR),
    .Y(_0035_),
    .A(\state[16] ),
    .VSS(VGND));
 sg13g2_inv_1 _1397_ (.VDD(VPWR),
    .Y(_0034_),
    .A(\state[15] ),
    .VSS(VGND));
 sg13g2_inv_1 _1398_ (.VDD(VPWR),
    .Y(_0033_),
    .A(\state[14] ),
    .VSS(VGND));
 sg13g2_inv_1 _1399_ (.VDD(VPWR),
    .Y(_0032_),
    .A(\state[13] ),
    .VSS(VGND));
 sg13g2_inv_1 _1400_ (.VDD(VPWR),
    .Y(_0031_),
    .A(\state[12] ),
    .VSS(VGND));
 sg13g2_inv_1 _1401_ (.VDD(VPWR),
    .Y(_0022_),
    .A(\state[11] ),
    .VSS(VGND));
 sg13g2_inv_1 _1402_ (.VDD(VPWR),
    .Y(_0011_),
    .A(\state[10] ),
    .VSS(VGND));
 sg13g2_inv_1 _1403_ (.VDD(VPWR),
    .Y(_0127_),
    .A(\state[9] ),
    .VSS(VGND));
 sg13g2_inv_1 _1404_ (.VDD(VPWR),
    .Y(_0116_),
    .A(\state[8] ),
    .VSS(VGND));
 sg13g2_inv_1 _1405_ (.VDD(VPWR),
    .Y(_0105_),
    .A(\state[7] ),
    .VSS(VGND));
 sg13g2_inv_1 _1406_ (.VDD(VPWR),
    .Y(_0094_),
    .A(\state[6] ),
    .VSS(VGND));
 sg13g2_inv_1 _1407_ (.VDD(VPWR),
    .Y(_0083_),
    .A(\state[5] ),
    .VSS(VGND));
 sg13g2_inv_1 _1408_ (.VDD(VPWR),
    .Y(_0072_),
    .A(\state[4] ),
    .VSS(VGND));
 sg13g2_inv_1 _1409_ (.VDD(VPWR),
    .Y(_0061_),
    .A(\state[3] ),
    .VSS(VGND));
 sg13g2_inv_1 _1410_ (.VDD(VPWR),
    .Y(_0050_),
    .A(\state[2] ),
    .VSS(VGND));
 sg13g2_inv_1 _1411_ (.VDD(VPWR),
    .Y(_0039_),
    .A(\state[1] ),
    .VSS(VGND));
 sg13g2_inv_1 _1412_ (.VDD(VPWR),
    .Y(_0000_),
    .A(\state[0] ),
    .VSS(VGND));
 sg13g2_inv_1 _1413_ (.VDD(VPWR),
    .Y(_0847_),
    .A(net178),
    .VSS(VGND));
 sg13g2_mux2_1 _1414_ (.A0(\state[0] ),
    .A1(\daisychain[0] ),
    .S(net134),
    .X(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1415_ (.Y(_0849_),
    .A(net157),
    .B(_0848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _1416_ (.A(net157),
    .B(net3),
    .Y(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _1417_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0851_),
    .B(net3),
    .A(net157));
 sg13g2_a21oi_1 _1418_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net92),
    .A2(net2),
    .Y(_0852_),
    .B1(net46));
 sg13g2_o21ai_1 _1419_ (.B1(net179),
    .VDD(VPWR),
    .Y(_0853_),
    .VSS(VGND),
    .A1(\daisychain[0] ),
    .A2(net24));
 sg13g2_a21oi_1 _1420_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0849_),
    .A2(_0852_),
    .Y(_0128_),
    .B1(_0853_));
 sg13g2_mux2_1 _1421_ (.A0(\state[1] ),
    .A1(\daisychain[1] ),
    .S(net134),
    .X(_0854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1422_ (.Y(_0855_),
    .A(net157),
    .B(_0854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1423_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net92),
    .A2(\daisychain[0] ),
    .Y(_0856_),
    .B1(net67));
 sg13g2_o21ai_1 _1424_ (.B1(net179),
    .VDD(VPWR),
    .Y(_0857_),
    .VSS(VGND),
    .A1(\daisychain[1] ),
    .A2(net24));
 sg13g2_a21oi_1 _1425_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0855_),
    .A2(_0856_),
    .Y(_0129_),
    .B1(_0857_));
 sg13g2_mux2_1 _1426_ (.A0(\state[2] ),
    .A1(\daisychain[2] ),
    .S(net134),
    .X(_0858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1427_ (.Y(_0859_),
    .A(net157),
    .B(_0858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1428_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net92),
    .A2(\daisychain[1] ),
    .Y(_0860_),
    .B1(net67));
 sg13g2_o21ai_1 _1429_ (.B1(net179),
    .VDD(VPWR),
    .Y(_0861_),
    .VSS(VGND),
    .A1(\daisychain[2] ),
    .A2(net24));
 sg13g2_a21oi_1 _1430_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0859_),
    .A2(_0860_),
    .Y(_0130_),
    .B1(_0861_));
 sg13g2_mux2_1 _1431_ (.A0(\state[3] ),
    .A1(\daisychain[3] ),
    .S(net135),
    .X(_0862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1432_ (.Y(_0863_),
    .A(net158),
    .B(_0862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1433_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net94),
    .A2(\daisychain[2] ),
    .Y(_0864_),
    .B1(net47));
 sg13g2_o21ai_1 _1434_ (.B1(net180),
    .VDD(VPWR),
    .Y(_0865_),
    .VSS(VGND),
    .A1(\daisychain[3] ),
    .A2(net25));
 sg13g2_a21oi_1 _1435_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0863_),
    .A2(_0864_),
    .Y(_0131_),
    .B1(_0865_));
 sg13g2_mux2_1 _1436_ (.A0(\state[4] ),
    .A1(\daisychain[4] ),
    .S(net135),
    .X(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1437_ (.Y(_0867_),
    .A(net158),
    .B(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1438_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net94),
    .A2(\daisychain[3] ),
    .Y(_0868_),
    .B1(net47));
 sg13g2_o21ai_1 _1439_ (.B1(net180),
    .VDD(VPWR),
    .Y(_0869_),
    .VSS(VGND),
    .A1(\daisychain[4] ),
    .A2(net25));
 sg13g2_a21oi_1 _1440_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0867_),
    .A2(_0868_),
    .Y(_0132_),
    .B1(_0869_));
 sg13g2_mux2_1 _1441_ (.A0(\state[5] ),
    .A1(\daisychain[5] ),
    .S(net135),
    .X(_0870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1442_ (.Y(_0871_),
    .A(net158),
    .B(_0870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1443_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net102),
    .A2(\daisychain[4] ),
    .Y(_0872_),
    .B1(net51));
 sg13g2_o21ai_1 _1444_ (.B1(net184),
    .VDD(VPWR),
    .Y(_0873_),
    .VSS(VGND),
    .A1(\daisychain[5] ),
    .A2(net29));
 sg13g2_a21oi_1 _1445_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0871_),
    .A2(_0872_),
    .Y(_0133_),
    .B1(_0873_));
 sg13g2_mux2_1 _1446_ (.A0(\state[6] ),
    .A1(\daisychain[6] ),
    .S(net137),
    .X(_0874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1447_ (.Y(_0875_),
    .A(net160),
    .B(_0874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1448_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net104),
    .A2(\daisychain[5] ),
    .Y(_0876_),
    .B1(net52));
 sg13g2_o21ai_1 _1449_ (.B1(net182),
    .VDD(VPWR),
    .Y(_0877_),
    .VSS(VGND),
    .A1(\daisychain[6] ),
    .A2(net27));
 sg13g2_a21oi_1 _1450_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0875_),
    .A2(_0876_),
    .Y(_0134_),
    .B1(_0877_));
 sg13g2_mux2_1 _1451_ (.A0(\state[7] ),
    .A1(\daisychain[7] ),
    .S(net137),
    .X(_0878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1452_ (.Y(_0879_),
    .A(net160),
    .B(_0878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1453_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net99),
    .A2(\daisychain[6] ),
    .Y(_0880_),
    .B1(net49));
 sg13g2_o21ai_1 _1454_ (.B1(net182),
    .VDD(VPWR),
    .Y(_0881_),
    .VSS(VGND),
    .A1(\daisychain[7] ),
    .A2(net27));
 sg13g2_a21oi_1 _1455_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0879_),
    .A2(_0880_),
    .Y(_0135_),
    .B1(_0881_));
 sg13g2_mux2_1 _1456_ (.A0(\state[8] ),
    .A1(\daisychain[8] ),
    .S(net137),
    .X(_0882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1457_ (.Y(_0883_),
    .A(net160),
    .B(_0882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1458_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net99),
    .A2(\daisychain[7] ),
    .Y(_0884_),
    .B1(net49));
 sg13g2_o21ai_1 _1459_ (.B1(net182),
    .VDD(VPWR),
    .Y(_0885_),
    .VSS(VGND),
    .A1(\daisychain[8] ),
    .A2(net27));
 sg13g2_a21oi_1 _1460_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0883_),
    .A2(_0884_),
    .Y(_0136_),
    .B1(_0885_));
 sg13g2_mux2_1 _1461_ (.A0(\state[9] ),
    .A1(\daisychain[9] ),
    .S(net135),
    .X(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1462_ (.Y(_0887_),
    .A(net158),
    .B(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1463_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net95),
    .A2(\daisychain[8] ),
    .Y(_0888_),
    .B1(net47));
 sg13g2_o21ai_1 _1464_ (.B1(net180),
    .VDD(VPWR),
    .Y(_0889_),
    .VSS(VGND),
    .A1(\daisychain[9] ),
    .A2(net25));
 sg13g2_a21oi_1 _1465_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0887_),
    .A2(_0888_),
    .Y(_0137_),
    .B1(_0889_));
 sg13g2_mux2_1 _1466_ (.A0(\state[10] ),
    .A1(\daisychain[10] ),
    .S(net135),
    .X(_0890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1467_ (.Y(_0891_),
    .A(net158),
    .B(_0890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1468_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net95),
    .A2(\daisychain[9] ),
    .Y(_0892_),
    .B1(net47));
 sg13g2_o21ai_1 _1469_ (.B1(net180),
    .VDD(VPWR),
    .Y(_0893_),
    .VSS(VGND),
    .A1(\daisychain[10] ),
    .A2(net25));
 sg13g2_a21oi_1 _1470_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0891_),
    .A2(_0892_),
    .Y(_0138_),
    .B1(_0893_));
 sg13g2_mux2_1 _1471_ (.A0(\state[11] ),
    .A1(\daisychain[11] ),
    .S(net135),
    .X(_0894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1472_ (.Y(_0895_),
    .A(net158),
    .B(_0894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1473_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net94),
    .A2(\daisychain[10] ),
    .Y(_0896_),
    .B1(net47));
 sg13g2_o21ai_1 _1474_ (.B1(net180),
    .VDD(VPWR),
    .Y(_0897_),
    .VSS(VGND),
    .A1(\daisychain[11] ),
    .A2(net25));
 sg13g2_a21oi_1 _1475_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0895_),
    .A2(_0896_),
    .Y(_0139_),
    .B1(_0897_));
 sg13g2_mux2_1 _1476_ (.A0(\state[12] ),
    .A1(\daisychain[12] ),
    .S(net134),
    .X(_0898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1477_ (.Y(_0899_),
    .A(net158),
    .B(_0898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1478_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net94),
    .A2(\daisychain[11] ),
    .Y(_0900_),
    .B1(net47));
 sg13g2_o21ai_1 _1479_ (.B1(net180),
    .VDD(VPWR),
    .Y(_0901_),
    .VSS(VGND),
    .A1(\daisychain[12] ),
    .A2(net25));
 sg13g2_a21oi_1 _1480_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0899_),
    .A2(_0900_),
    .Y(_0140_),
    .B1(_0901_));
 sg13g2_mux2_1 _1481_ (.A0(\state[13] ),
    .A1(\daisychain[13] ),
    .S(net135),
    .X(_0902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1482_ (.Y(_0903_),
    .A(net158),
    .B(_0902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1483_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net94),
    .A2(\daisychain[12] ),
    .Y(_0904_),
    .B1(net47));
 sg13g2_o21ai_1 _1484_ (.B1(net180),
    .VDD(VPWR),
    .Y(_0905_),
    .VSS(VGND),
    .A1(\daisychain[13] ),
    .A2(net25));
 sg13g2_a21oi_1 _1485_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0903_),
    .A2(_0904_),
    .Y(_0141_),
    .B1(_0905_));
 sg13g2_mux2_1 _1486_ (.A0(\state[14] ),
    .A1(\daisychain[14] ),
    .S(net138),
    .X(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1487_ (.Y(_0907_),
    .A(net161),
    .B(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1488_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net94),
    .A2(\daisychain[13] ),
    .Y(_0908_),
    .B1(net47));
 sg13g2_o21ai_1 _1489_ (.B1(net183),
    .VDD(VPWR),
    .Y(_0909_),
    .VSS(VGND),
    .A1(\daisychain[14] ),
    .A2(net28));
 sg13g2_a21oi_1 _1490_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0907_),
    .A2(_0908_),
    .Y(_0142_),
    .B1(_0909_));
 sg13g2_mux2_1 _1491_ (.A0(\state[15] ),
    .A1(\daisychain[15] ),
    .S(net135),
    .X(_0910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1492_ (.Y(_0911_),
    .A(net161),
    .B(_0910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1493_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net95),
    .A2(\daisychain[14] ),
    .Y(_0912_),
    .B1(net50));
 sg13g2_o21ai_1 _1494_ (.B1(net180),
    .VDD(VPWR),
    .Y(_0913_),
    .VSS(VGND),
    .A1(\daisychain[15] ),
    .A2(net25));
 sg13g2_a21oi_1 _1495_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0911_),
    .A2(_0912_),
    .Y(_0143_),
    .B1(_0913_));
 sg13g2_mux2_1 _1496_ (.A0(\state[16] ),
    .A1(\daisychain[16] ),
    .S(net136),
    .X(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1497_ (.Y(_0915_),
    .A(net159),
    .B(_0914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1498_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net109),
    .A2(\daisychain[15] ),
    .Y(_0916_),
    .B1(net50));
 sg13g2_o21ai_1 _1499_ (.B1(net181),
    .VDD(VPWR),
    .Y(_0917_),
    .VSS(VGND),
    .A1(\daisychain[16] ),
    .A2(net26));
 sg13g2_a21oi_1 _1500_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0915_),
    .A2(_0916_),
    .Y(_0144_),
    .B1(_0917_));
 sg13g2_mux2_1 _1501_ (.A0(\state[17] ),
    .A1(\daisychain[17] ),
    .S(net136),
    .X(_0918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1502_ (.Y(_0919_),
    .A(net159),
    .B(_0918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1503_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net98),
    .A2(\daisychain[16] ),
    .Y(_0920_),
    .B1(net48));
 sg13g2_o21ai_1 _1504_ (.B1(net181),
    .VDD(VPWR),
    .Y(_0921_),
    .VSS(VGND),
    .A1(\daisychain[17] ),
    .A2(net26));
 sg13g2_a21oi_1 _1505_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0919_),
    .A2(_0920_),
    .Y(_0145_),
    .B1(_0921_));
 sg13g2_mux2_1 _1506_ (.A0(\state[18] ),
    .A1(\daisychain[18] ),
    .S(net136),
    .X(_0922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1507_ (.Y(_0923_),
    .A(net159),
    .B(_0922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1508_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net98),
    .A2(\daisychain[17] ),
    .Y(_0924_),
    .B1(net48));
 sg13g2_o21ai_1 _1509_ (.B1(net181),
    .VDD(VPWR),
    .Y(_0925_),
    .VSS(VGND),
    .A1(\daisychain[18] ),
    .A2(net26));
 sg13g2_a21oi_1 _1510_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0923_),
    .A2(_0924_),
    .Y(_0146_),
    .B1(_0925_));
 sg13g2_mux2_1 _1511_ (.A0(\state[19] ),
    .A1(\daisychain[19] ),
    .S(net136),
    .X(_0926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1512_ (.Y(_0927_),
    .A(net159),
    .B(_0926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1513_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net98),
    .A2(\daisychain[18] ),
    .Y(_0928_),
    .B1(net48));
 sg13g2_o21ai_1 _1514_ (.B1(net181),
    .VDD(VPWR),
    .Y(_0929_),
    .VSS(VGND),
    .A1(\daisychain[19] ),
    .A2(net26));
 sg13g2_a21oi_1 _1515_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0927_),
    .A2(_0928_),
    .Y(_0147_),
    .B1(_0929_));
 sg13g2_mux2_1 _1516_ (.A0(\state[20] ),
    .A1(\daisychain[20] ),
    .S(net136),
    .X(_0930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1517_ (.Y(_0931_),
    .A(net159),
    .B(_0930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1518_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net98),
    .A2(\daisychain[19] ),
    .Y(_0932_),
    .B1(net48));
 sg13g2_o21ai_1 _1519_ (.B1(net181),
    .VDD(VPWR),
    .Y(_0933_),
    .VSS(VGND),
    .A1(\daisychain[20] ),
    .A2(net26));
 sg13g2_a21oi_1 _1520_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0931_),
    .A2(_0932_),
    .Y(_0148_),
    .B1(_0933_));
 sg13g2_mux2_1 _1521_ (.A0(\state[21] ),
    .A1(\daisychain[21] ),
    .S(net136),
    .X(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1522_ (.Y(_0935_),
    .A(net159),
    .B(_0934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1523_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net97),
    .A2(\daisychain[20] ),
    .Y(_0936_),
    .B1(net48));
 sg13g2_o21ai_1 _1524_ (.B1(net181),
    .VDD(VPWR),
    .Y(_0937_),
    .VSS(VGND),
    .A1(\daisychain[21] ),
    .A2(net26));
 sg13g2_a21oi_1 _1525_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0935_),
    .A2(_0936_),
    .Y(_0149_),
    .B1(_0937_));
 sg13g2_mux2_1 _1526_ (.A0(\state[22] ),
    .A1(\daisychain[22] ),
    .S(net136),
    .X(_0938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1527_ (.Y(_0939_),
    .A(net159),
    .B(_0938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1528_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net97),
    .A2(\daisychain[21] ),
    .Y(_0940_),
    .B1(net48));
 sg13g2_o21ai_1 _1529_ (.B1(net181),
    .VDD(VPWR),
    .Y(_0941_),
    .VSS(VGND),
    .A1(\daisychain[22] ),
    .A2(net26));
 sg13g2_a21oi_1 _1530_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0939_),
    .A2(_0940_),
    .Y(_0150_),
    .B1(_0941_));
 sg13g2_mux2_1 _1531_ (.A0(\state[23] ),
    .A1(\daisychain[23] ),
    .S(net136),
    .X(_0942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1532_ (.Y(_0943_),
    .A(net159),
    .B(_0942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1533_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net97),
    .A2(\daisychain[22] ),
    .Y(_0944_),
    .B1(net48));
 sg13g2_o21ai_1 _1534_ (.B1(net181),
    .VDD(VPWR),
    .Y(_0945_),
    .VSS(VGND),
    .A1(\daisychain[23] ),
    .A2(net26));
 sg13g2_a21oi_1 _1535_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0943_),
    .A2(_0944_),
    .Y(_0151_),
    .B1(_0945_));
 sg13g2_mux2_1 _1536_ (.A0(\state[24] ),
    .A1(\daisychain[24] ),
    .S(net137),
    .X(_0946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1537_ (.Y(_0947_),
    .A(net160),
    .B(_0946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1538_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net97),
    .A2(\daisychain[23] ),
    .Y(_0948_),
    .B1(net48));
 sg13g2_o21ai_1 _1539_ (.B1(net182),
    .VDD(VPWR),
    .Y(_0949_),
    .VSS(VGND),
    .A1(\daisychain[24] ),
    .A2(net27));
 sg13g2_a21oi_1 _1540_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0947_),
    .A2(_0948_),
    .Y(_0152_),
    .B1(_0949_));
 sg13g2_mux2_1 _1541_ (.A0(\state[25] ),
    .A1(\daisychain[25] ),
    .S(net137),
    .X(_0950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1542_ (.Y(_0951_),
    .A(net160),
    .B(_0950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1543_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net97),
    .A2(\daisychain[24] ),
    .Y(_0952_),
    .B1(net49));
 sg13g2_o21ai_1 _1544_ (.B1(net182),
    .VDD(VPWR),
    .Y(_0953_),
    .VSS(VGND),
    .A1(\daisychain[25] ),
    .A2(net27));
 sg13g2_a21oi_1 _1545_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0951_),
    .A2(_0952_),
    .Y(_0153_),
    .B1(_0953_));
 sg13g2_mux2_1 _1546_ (.A0(\state[26] ),
    .A1(\daisychain[26] ),
    .S(net137),
    .X(_0954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1547_ (.Y(_0955_),
    .A(net160),
    .B(_0954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1548_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net100),
    .A2(\daisychain[25] ),
    .Y(_0956_),
    .B1(net49));
 sg13g2_o21ai_1 _1549_ (.B1(net182),
    .VDD(VPWR),
    .Y(_0957_),
    .VSS(VGND),
    .A1(\daisychain[26] ),
    .A2(net27));
 sg13g2_a21oi_1 _1550_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0955_),
    .A2(_0956_),
    .Y(_0154_),
    .B1(_0957_));
 sg13g2_mux2_1 _1551_ (.A0(\state[27] ),
    .A1(\daisychain[27] ),
    .S(net137),
    .X(_0958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1552_ (.Y(_0959_),
    .A(net160),
    .B(_0958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1553_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net99),
    .A2(\daisychain[26] ),
    .Y(_0960_),
    .B1(net49));
 sg13g2_o21ai_1 _1554_ (.B1(net182),
    .VDD(VPWR),
    .Y(_0961_),
    .VSS(VGND),
    .A1(\daisychain[27] ),
    .A2(net27));
 sg13g2_a21oi_1 _1555_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0959_),
    .A2(_0960_),
    .Y(_0155_),
    .B1(_0961_));
 sg13g2_mux2_1 _1556_ (.A0(\state[28] ),
    .A1(\daisychain[28] ),
    .S(net138),
    .X(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1557_ (.Y(_0963_),
    .A(net161),
    .B(_0962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1558_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net99),
    .A2(\daisychain[27] ),
    .Y(_0964_),
    .B1(net49));
 sg13g2_o21ai_1 _1559_ (.B1(net183),
    .VDD(VPWR),
    .Y(_0965_),
    .VSS(VGND),
    .A1(\daisychain[28] ),
    .A2(net28));
 sg13g2_a21oi_1 _1560_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0963_),
    .A2(_0964_),
    .Y(_0156_),
    .B1(_0965_));
 sg13g2_mux2_1 _1561_ (.A0(\state[29] ),
    .A1(\daisychain[29] ),
    .S(net138),
    .X(_0966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1562_ (.Y(_0967_),
    .A(net161),
    .B(_0966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1563_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net100),
    .A2(\daisychain[28] ),
    .Y(_0968_),
    .B1(net49));
 sg13g2_o21ai_1 _1564_ (.B1(net183),
    .VDD(VPWR),
    .Y(_0969_),
    .VSS(VGND),
    .A1(\daisychain[29] ),
    .A2(net28));
 sg13g2_a21oi_1 _1565_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0967_),
    .A2(_0968_),
    .Y(_0157_),
    .B1(_0969_));
 sg13g2_mux2_1 _1566_ (.A0(\state[30] ),
    .A1(\daisychain[30] ),
    .S(net144),
    .X(_0970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1567_ (.Y(_0971_),
    .A(net166),
    .B(_0970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1568_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net100),
    .A2(\daisychain[29] ),
    .Y(_0972_),
    .B1(net50));
 sg13g2_o21ai_1 _1569_ (.B1(net189),
    .VDD(VPWR),
    .Y(_0973_),
    .VSS(VGND),
    .A1(\daisychain[30] ),
    .A2(net34));
 sg13g2_a21oi_1 _1570_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0971_),
    .A2(_0972_),
    .Y(_0158_),
    .B1(_0973_));
 sg13g2_mux2_1 _1571_ (.A0(\state[31] ),
    .A1(\daisychain[31] ),
    .S(net144),
    .X(_0974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1572_ (.Y(_0975_),
    .A(net166),
    .B(_0974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1573_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net113),
    .A2(\daisychain[30] ),
    .Y(_0976_),
    .B1(net57));
 sg13g2_o21ai_1 _1574_ (.B1(net189),
    .VDD(VPWR),
    .Y(_0977_),
    .VSS(VGND),
    .A1(\daisychain[31] ),
    .A2(net34));
 sg13g2_a21oi_1 _1575_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0975_),
    .A2(_0976_),
    .Y(_0159_),
    .B1(_0977_));
 sg13g2_mux2_1 _1576_ (.A0(\state[32] ),
    .A1(\daisychain[32] ),
    .S(net143),
    .X(_0978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1577_ (.Y(_0979_),
    .A(net165),
    .B(_0978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1578_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net113),
    .A2(\daisychain[31] ),
    .Y(_0980_),
    .B1(net57));
 sg13g2_o21ai_1 _1579_ (.B1(net188),
    .VDD(VPWR),
    .Y(_0981_),
    .VSS(VGND),
    .A1(\daisychain[32] ),
    .A2(net33));
 sg13g2_a21oi_1 _1580_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0979_),
    .A2(_0980_),
    .Y(_0160_),
    .B1(_0981_));
 sg13g2_mux2_1 _1581_ (.A0(\state[33] ),
    .A1(\daisychain[33] ),
    .S(net143),
    .X(_0982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1582_ (.Y(_0983_),
    .A(net165),
    .B(_0982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1583_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net110),
    .A2(\daisychain[32] ),
    .Y(_0984_),
    .B1(net55));
 sg13g2_o21ai_1 _1584_ (.B1(net188),
    .VDD(VPWR),
    .Y(_0985_),
    .VSS(VGND),
    .A1(\daisychain[33] ),
    .A2(net33));
 sg13g2_a21oi_1 _1585_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0983_),
    .A2(_0984_),
    .Y(_0161_),
    .B1(_0985_));
 sg13g2_mux2_1 _1586_ (.A0(\state[34] ),
    .A1(\daisychain[34] ),
    .S(net143),
    .X(_0986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1587_ (.Y(_0987_),
    .A(net165),
    .B(_0986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1588_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net112),
    .A2(\daisychain[33] ),
    .Y(_0988_),
    .B1(net55));
 sg13g2_o21ai_1 _1589_ (.B1(net188),
    .VDD(VPWR),
    .Y(_0989_),
    .VSS(VGND),
    .A1(\daisychain[34] ),
    .A2(net33));
 sg13g2_a21oi_1 _1590_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0987_),
    .A2(_0988_),
    .Y(_0162_),
    .B1(_0989_));
 sg13g2_mux2_1 _1591_ (.A0(\state[35] ),
    .A1(\daisychain[35] ),
    .S(net143),
    .X(_0990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1592_ (.Y(_0991_),
    .A(net165),
    .B(_0990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1593_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net110),
    .A2(\daisychain[34] ),
    .Y(_0992_),
    .B1(net55));
 sg13g2_o21ai_1 _1594_ (.B1(net188),
    .VDD(VPWR),
    .Y(_0993_),
    .VSS(VGND),
    .A1(\daisychain[35] ),
    .A2(net33));
 sg13g2_a21oi_1 _1595_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0991_),
    .A2(_0992_),
    .Y(_0163_),
    .B1(_0993_));
 sg13g2_mux2_1 _1596_ (.A0(\state[36] ),
    .A1(\daisychain[36] ),
    .S(net143),
    .X(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1597_ (.Y(_0995_),
    .A(net165),
    .B(_0994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1598_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net110),
    .A2(\daisychain[35] ),
    .Y(_0996_),
    .B1(net55));
 sg13g2_o21ai_1 _1599_ (.B1(net188),
    .VDD(VPWR),
    .Y(_0997_),
    .VSS(VGND),
    .A1(\daisychain[36] ),
    .A2(net33));
 sg13g2_a21oi_1 _1600_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0995_),
    .A2(_0996_),
    .Y(_0164_),
    .B1(_0997_));
 sg13g2_mux2_1 _1601_ (.A0(\state[37] ),
    .A1(\daisychain[37] ),
    .S(net143),
    .X(_0998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1602_ (.Y(_0999_),
    .A(net165),
    .B(_0998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1603_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net110),
    .A2(\daisychain[36] ),
    .Y(_1000_),
    .B1(net55));
 sg13g2_o21ai_1 _1604_ (.B1(net188),
    .VDD(VPWR),
    .Y(_1001_),
    .VSS(VGND),
    .A1(\daisychain[37] ),
    .A2(net33));
 sg13g2_a21oi_1 _1605_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0999_),
    .A2(_1000_),
    .Y(_0165_),
    .B1(_1001_));
 sg13g2_mux2_1 _1606_ (.A0(\state[38] ),
    .A1(\daisychain[38] ),
    .S(net143),
    .X(_1002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1607_ (.Y(_1003_),
    .A(net165),
    .B(_1002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1608_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net110),
    .A2(\daisychain[37] ),
    .Y(_1004_),
    .B1(net55));
 sg13g2_o21ai_1 _1609_ (.B1(net188),
    .VDD(VPWR),
    .Y(_1005_),
    .VSS(VGND),
    .A1(\daisychain[38] ),
    .A2(net33));
 sg13g2_a21oi_1 _1610_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1003_),
    .A2(_1004_),
    .Y(_0166_),
    .B1(_1005_));
 sg13g2_mux2_1 _1611_ (.A0(\state[39] ),
    .A1(\daisychain[39] ),
    .S(net143),
    .X(_1006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1612_ (.Y(_1007_),
    .A(net165),
    .B(_1006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1613_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net111),
    .A2(\daisychain[38] ),
    .Y(_1008_),
    .B1(net55));
 sg13g2_o21ai_1 _1614_ (.B1(net188),
    .VDD(VPWR),
    .Y(_1009_),
    .VSS(VGND),
    .A1(\daisychain[39] ),
    .A2(net33));
 sg13g2_a21oi_1 _1615_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1007_),
    .A2(_1008_),
    .Y(_0167_),
    .B1(_1009_));
 sg13g2_mux2_1 _1616_ (.A0(\state[40] ),
    .A1(\daisychain[40] ),
    .S(net144),
    .X(_1010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1617_ (.Y(_1011_),
    .A(net166),
    .B(_1010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1618_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net111),
    .A2(\daisychain[39] ),
    .Y(_1012_),
    .B1(net55));
 sg13g2_o21ai_1 _1619_ (.B1(net190),
    .VDD(VPWR),
    .Y(_1013_),
    .VSS(VGND),
    .A1(\daisychain[40] ),
    .A2(net35));
 sg13g2_a21oi_1 _1620_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1011_),
    .A2(_1012_),
    .Y(_0168_),
    .B1(_1013_));
 sg13g2_mux2_1 _1621_ (.A0(\state[41] ),
    .A1(\daisychain[41] ),
    .S(net145),
    .X(_1014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1622_ (.Y(_1015_),
    .A(net167),
    .B(_1014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1623_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net111),
    .A2(\daisychain[40] ),
    .Y(_1016_),
    .B1(net56));
 sg13g2_o21ai_1 _1624_ (.B1(net190),
    .VDD(VPWR),
    .Y(_1017_),
    .VSS(VGND),
    .A1(\daisychain[41] ),
    .A2(net35));
 sg13g2_a21oi_1 _1625_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1015_),
    .A2(_1016_),
    .Y(_0169_),
    .B1(_1017_));
 sg13g2_mux2_1 _1626_ (.A0(\state[42] ),
    .A1(\daisychain[42] ),
    .S(net144),
    .X(_1018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1627_ (.Y(_1019_),
    .A(net167),
    .B(_1018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1628_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net111),
    .A2(\daisychain[41] ),
    .Y(_1020_),
    .B1(net56));
 sg13g2_o21ai_1 _1629_ (.B1(net189),
    .VDD(VPWR),
    .Y(_1021_),
    .VSS(VGND),
    .A1(\daisychain[42] ),
    .A2(net34));
 sg13g2_a21oi_1 _1630_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1019_),
    .A2(_1020_),
    .Y(_0170_),
    .B1(_1021_));
 sg13g2_mux2_1 _1631_ (.A0(\state[43] ),
    .A1(\daisychain[43] ),
    .S(net144),
    .X(_1022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1632_ (.Y(_1023_),
    .A(net166),
    .B(_1022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1633_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net111),
    .A2(\daisychain[42] ),
    .Y(_1024_),
    .B1(net56));
 sg13g2_o21ai_1 _1634_ (.B1(net189),
    .VDD(VPWR),
    .Y(_1025_),
    .VSS(VGND),
    .A1(\daisychain[43] ),
    .A2(net34));
 sg13g2_a21oi_1 _1635_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1023_),
    .A2(_1024_),
    .Y(_0171_),
    .B1(_1025_));
 sg13g2_mux2_1 _1636_ (.A0(\state[44] ),
    .A1(\daisychain[44] ),
    .S(net144),
    .X(_1026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1637_ (.Y(_1027_),
    .A(net166),
    .B(_1026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1638_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net112),
    .A2(\daisychain[43] ),
    .Y(_0384_),
    .B1(net56));
 sg13g2_o21ai_1 _1639_ (.B1(net189),
    .VDD(VPWR),
    .Y(_0385_),
    .VSS(VGND),
    .A1(\daisychain[44] ),
    .A2(net34));
 sg13g2_a21oi_1 _1640_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1027_),
    .A2(_0384_),
    .Y(_0172_),
    .B1(_0385_));
 sg13g2_mux2_1 _1641_ (.A0(\state[45] ),
    .A1(\daisychain[45] ),
    .S(net144),
    .X(_0386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1642_ (.Y(_0387_),
    .A(net166),
    .B(_0386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1643_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net113),
    .A2(\daisychain[44] ),
    .Y(_0388_),
    .B1(net57));
 sg13g2_o21ai_1 _1644_ (.B1(net189),
    .VDD(VPWR),
    .Y(_0389_),
    .VSS(VGND),
    .A1(\daisychain[45] ),
    .A2(net34));
 sg13g2_a21oi_1 _1645_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0387_),
    .A2(_0388_),
    .Y(_0173_),
    .B1(_0389_));
 sg13g2_mux2_1 _1646_ (.A0(\state[46] ),
    .A1(\daisychain[46] ),
    .S(net154),
    .X(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1647_ (.Y(_0391_),
    .A(net166),
    .B(_0390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1648_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net113),
    .A2(\daisychain[45] ),
    .Y(_0392_),
    .B1(net57));
 sg13g2_o21ai_1 _1649_ (.B1(net189),
    .VDD(VPWR),
    .Y(_0393_),
    .VSS(VGND),
    .A1(\daisychain[46] ),
    .A2(net34));
 sg13g2_a21oi_1 _1650_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0391_),
    .A2(_0392_),
    .Y(_0174_),
    .B1(_0393_));
 sg13g2_mux2_1 _1651_ (.A0(\state[47] ),
    .A1(\daisychain[47] ),
    .S(net147),
    .X(_0394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1652_ (.Y(_0395_),
    .A(net169),
    .B(_0394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1653_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net119),
    .A2(\daisychain[46] ),
    .Y(_0396_),
    .B1(net60));
 sg13g2_o21ai_1 _1654_ (.B1(net192),
    .VDD(VPWR),
    .Y(_0397_),
    .VSS(VGND),
    .A1(\daisychain[47] ),
    .A2(net37));
 sg13g2_a21oi_1 _1655_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0395_),
    .A2(_0396_),
    .Y(_0175_),
    .B1(_0397_));
 sg13g2_mux2_1 _1656_ (.A0(\state[48] ),
    .A1(\daisychain[48] ),
    .S(net147),
    .X(_0398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1657_ (.Y(_0399_),
    .A(net169),
    .B(_0398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1658_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net119),
    .A2(\daisychain[47] ),
    .Y(_0400_),
    .B1(net60));
 sg13g2_o21ai_1 _1659_ (.B1(net192),
    .VDD(VPWR),
    .Y(_0401_),
    .VSS(VGND),
    .A1(\daisychain[48] ),
    .A2(net37));
 sg13g2_a21oi_1 _1660_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0399_),
    .A2(_0400_),
    .Y(_0176_),
    .B1(_0401_));
 sg13g2_mux2_1 _1661_ (.A0(\state[49] ),
    .A1(\daisychain[49] ),
    .S(net147),
    .X(_0402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1662_ (.Y(_0403_),
    .A(net169),
    .B(_0402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1663_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net119),
    .A2(\daisychain[48] ),
    .Y(_0404_),
    .B1(net60));
 sg13g2_o21ai_1 _1664_ (.B1(net192),
    .VDD(VPWR),
    .Y(_0405_),
    .VSS(VGND),
    .A1(\daisychain[49] ),
    .A2(net37));
 sg13g2_a21oi_1 _1665_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0403_),
    .A2(_0404_),
    .Y(_0177_),
    .B1(_0405_));
 sg13g2_mux2_1 _1666_ (.A0(\state[50] ),
    .A1(\daisychain[50] ),
    .S(net145),
    .X(_0406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1667_ (.Y(_0407_),
    .A(net167),
    .B(_0406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1668_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net115),
    .A2(\daisychain[49] ),
    .Y(_0408_),
    .B1(net58));
 sg13g2_o21ai_1 _1669_ (.B1(net190),
    .VDD(VPWR),
    .Y(_0409_),
    .VSS(VGND),
    .A1(\daisychain[50] ),
    .A2(net35));
 sg13g2_a21oi_1 _1670_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0407_),
    .A2(_0408_),
    .Y(_0178_),
    .B1(_0409_));
 sg13g2_mux2_1 _1671_ (.A0(\state[51] ),
    .A1(\daisychain[51] ),
    .S(net145),
    .X(_0410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1672_ (.Y(_0411_),
    .A(net167),
    .B(_0410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1673_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net115),
    .A2(\daisychain[50] ),
    .Y(_0412_),
    .B1(net58));
 sg13g2_o21ai_1 _1674_ (.B1(net190),
    .VDD(VPWR),
    .Y(_0413_),
    .VSS(VGND),
    .A1(\daisychain[51] ),
    .A2(net35));
 sg13g2_a21oi_1 _1675_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0411_),
    .A2(_0412_),
    .Y(_0179_),
    .B1(_0413_));
 sg13g2_mux2_1 _1676_ (.A0(\state[52] ),
    .A1(\daisychain[52] ),
    .S(net145),
    .X(_0414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1677_ (.Y(_0415_),
    .A(net167),
    .B(_0414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1678_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net115),
    .A2(\daisychain[51] ),
    .Y(_0416_),
    .B1(net58));
 sg13g2_o21ai_1 _1679_ (.B1(net190),
    .VDD(VPWR),
    .Y(_0417_),
    .VSS(VGND),
    .A1(\daisychain[52] ),
    .A2(net35));
 sg13g2_a21oi_1 _1680_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0415_),
    .A2(_0416_),
    .Y(_0180_),
    .B1(_0417_));
 sg13g2_mux2_1 _1681_ (.A0(\state[53] ),
    .A1(\daisychain[53] ),
    .S(net145),
    .X(_0418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1682_ (.Y(_0419_),
    .A(net167),
    .B(_0418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1683_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net115),
    .A2(\daisychain[52] ),
    .Y(_0420_),
    .B1(net58));
 sg13g2_o21ai_1 _1684_ (.B1(net190),
    .VDD(VPWR),
    .Y(_0421_),
    .VSS(VGND),
    .A1(\daisychain[53] ),
    .A2(net35));
 sg13g2_a21oi_1 _1685_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0419_),
    .A2(_0420_),
    .Y(_0181_),
    .B1(_0421_));
 sg13g2_mux2_1 _1686_ (.A0(\state[54] ),
    .A1(\daisychain[54] ),
    .S(net145),
    .X(_0422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1687_ (.Y(_0423_),
    .A(net167),
    .B(_0422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1688_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net115),
    .A2(\daisychain[53] ),
    .Y(_0424_),
    .B1(net58));
 sg13g2_o21ai_1 _1689_ (.B1(net190),
    .VDD(VPWR),
    .Y(_0425_),
    .VSS(VGND),
    .A1(\daisychain[54] ),
    .A2(net35));
 sg13g2_a21oi_1 _1690_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0423_),
    .A2(_0424_),
    .Y(_0182_),
    .B1(_0425_));
 sg13g2_mux2_1 _1691_ (.A0(\state[55] ),
    .A1(\daisychain[55] ),
    .S(net145),
    .X(_0426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1692_ (.Y(_0427_),
    .A(net167),
    .B(_0426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1693_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net116),
    .A2(\daisychain[54] ),
    .Y(_0428_),
    .B1(net58));
 sg13g2_o21ai_1 _1694_ (.B1(net190),
    .VDD(VPWR),
    .Y(_0429_),
    .VSS(VGND),
    .A1(\daisychain[55] ),
    .A2(net35));
 sg13g2_a21oi_1 _1695_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0427_),
    .A2(_0428_),
    .Y(_0183_),
    .B1(_0429_));
 sg13g2_mux2_1 _1696_ (.A0(\state[56] ),
    .A1(\daisychain[56] ),
    .S(net145),
    .X(_0430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1697_ (.Y(_0431_),
    .A(net168),
    .B(_0430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1698_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net116),
    .A2(\daisychain[55] ),
    .Y(_0432_),
    .B1(net58));
 sg13g2_o21ai_1 _1699_ (.B1(net191),
    .VDD(VPWR),
    .Y(_0433_),
    .VSS(VGND),
    .A1(\daisychain[56] ),
    .A2(net36));
 sg13g2_a21oi_1 _1700_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0431_),
    .A2(_0432_),
    .Y(_0184_),
    .B1(_0433_));
 sg13g2_mux2_1 _1701_ (.A0(\state[57] ),
    .A1(\daisychain[57] ),
    .S(net146),
    .X(_0434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1702_ (.Y(_0435_),
    .A(net168),
    .B(_0434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1703_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net116),
    .A2(\daisychain[56] ),
    .Y(_0436_),
    .B1(net58));
 sg13g2_o21ai_1 _1704_ (.B1(net191),
    .VDD(VPWR),
    .Y(_0437_),
    .VSS(VGND),
    .A1(\daisychain[57] ),
    .A2(net36));
 sg13g2_a21oi_1 _1705_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0435_),
    .A2(_0436_),
    .Y(_0185_),
    .B1(_0437_));
 sg13g2_mux2_1 _1706_ (.A0(\state[58] ),
    .A1(\daisychain[58] ),
    .S(net146),
    .X(_0438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1707_ (.Y(_0439_),
    .A(net168),
    .B(_0438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1708_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net116),
    .A2(\daisychain[57] ),
    .Y(_0440_),
    .B1(net59));
 sg13g2_o21ai_1 _1709_ (.B1(net191),
    .VDD(VPWR),
    .Y(_0441_),
    .VSS(VGND),
    .A1(\daisychain[58] ),
    .A2(net36));
 sg13g2_a21oi_1 _1710_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0439_),
    .A2(_0440_),
    .Y(_0186_),
    .B1(_0441_));
 sg13g2_mux2_1 _1711_ (.A0(\state[59] ),
    .A1(\daisychain[59] ),
    .S(net146),
    .X(_0442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1712_ (.Y(_0443_),
    .A(net168),
    .B(_0442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1713_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net117),
    .A2(\daisychain[58] ),
    .Y(_0444_),
    .B1(net59));
 sg13g2_o21ai_1 _1714_ (.B1(net191),
    .VDD(VPWR),
    .Y(_0445_),
    .VSS(VGND),
    .A1(\daisychain[59] ),
    .A2(net36));
 sg13g2_a21oi_1 _1715_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0443_),
    .A2(_0444_),
    .Y(_0187_),
    .B1(_0445_));
 sg13g2_mux2_1 _1716_ (.A0(\state[60] ),
    .A1(\daisychain[60] ),
    .S(net146),
    .X(_0446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1717_ (.Y(_0447_),
    .A(net168),
    .B(_0446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1718_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net117),
    .A2(\daisychain[59] ),
    .Y(_0448_),
    .B1(net59));
 sg13g2_o21ai_1 _1719_ (.B1(net191),
    .VDD(VPWR),
    .Y(_0449_),
    .VSS(VGND),
    .A1(\daisychain[60] ),
    .A2(net36));
 sg13g2_a21oi_1 _1720_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0447_),
    .A2(_0448_),
    .Y(_0188_),
    .B1(_0449_));
 sg13g2_mux2_1 _1721_ (.A0(\state[61] ),
    .A1(\daisychain[61] ),
    .S(net147),
    .X(_0450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1722_ (.Y(_0451_),
    .A(net169),
    .B(_0450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1723_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net117),
    .A2(\daisychain[60] ),
    .Y(_0452_),
    .B1(net59));
 sg13g2_o21ai_1 _1724_ (.B1(net192),
    .VDD(VPWR),
    .Y(_0453_),
    .VSS(VGND),
    .A1(\daisychain[61] ),
    .A2(net37));
 sg13g2_a21oi_1 _1725_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0451_),
    .A2(_0452_),
    .Y(_0189_),
    .B1(_0453_));
 sg13g2_mux2_1 _1726_ (.A0(\state[62] ),
    .A1(\daisychain[62] ),
    .S(net147),
    .X(_0454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1727_ (.Y(_0455_),
    .A(net169),
    .B(_0454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1728_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net119),
    .A2(\daisychain[61] ),
    .Y(_0456_),
    .B1(net60));
 sg13g2_o21ai_1 _1729_ (.B1(net192),
    .VDD(VPWR),
    .Y(_0457_),
    .VSS(VGND),
    .A1(\daisychain[62] ),
    .A2(net37));
 sg13g2_a21oi_1 _1730_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0455_),
    .A2(_0456_),
    .Y(_0190_),
    .B1(_0457_));
 sg13g2_mux2_1 _1731_ (.A0(\state[63] ),
    .A1(\daisychain[63] ),
    .S(net147),
    .X(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1732_ (.Y(_0459_),
    .A(net169),
    .B(_0458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1733_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net119),
    .A2(\daisychain[62] ),
    .Y(_0460_),
    .B1(net60));
 sg13g2_o21ai_1 _1734_ (.B1(net192),
    .VDD(VPWR),
    .Y(_0461_),
    .VSS(VGND),
    .A1(\daisychain[63] ),
    .A2(net37));
 sg13g2_a21oi_1 _1735_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0459_),
    .A2(_0460_),
    .Y(_0191_),
    .B1(_0461_));
 sg13g2_mux2_1 _1736_ (.A0(\state[64] ),
    .A1(\daisychain[64] ),
    .S(net153),
    .X(_0462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1737_ (.Y(_0463_),
    .A(net175),
    .B(_0462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1738_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net119),
    .A2(\daisychain[63] ),
    .Y(_0464_),
    .B1(net60));
 sg13g2_o21ai_1 _1739_ (.B1(net198),
    .VDD(VPWR),
    .Y(_0465_),
    .VSS(VGND),
    .A1(\daisychain[64] ),
    .A2(net43));
 sg13g2_a21oi_1 _1740_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0463_),
    .A2(_0464_),
    .Y(_0192_),
    .B1(_0465_));
 sg13g2_mux2_1 _1741_ (.A0(\state[65] ),
    .A1(\daisychain[65] ),
    .S(net153),
    .X(_0466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1742_ (.Y(_0467_),
    .A(net175),
    .B(_0466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1743_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net126),
    .A2(\daisychain[64] ),
    .Y(_0468_),
    .B1(net65));
 sg13g2_o21ai_1 _1744_ (.B1(net198),
    .VDD(VPWR),
    .Y(_0469_),
    .VSS(VGND),
    .A1(\daisychain[65] ),
    .A2(net43));
 sg13g2_a21oi_1 _1745_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0467_),
    .A2(_0468_),
    .Y(_0193_),
    .B1(_0469_));
 sg13g2_mux2_1 _1746_ (.A0(\state[66] ),
    .A1(\daisychain[66] ),
    .S(net153),
    .X(_0470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1747_ (.Y(_0471_),
    .A(net175),
    .B(_0470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1748_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net126),
    .A2(\daisychain[65] ),
    .Y(_0472_),
    .B1(net65));
 sg13g2_o21ai_1 _1749_ (.B1(net196),
    .VDD(VPWR),
    .Y(_0473_),
    .VSS(VGND),
    .A1(\daisychain[66] ),
    .A2(net41));
 sg13g2_a21oi_1 _1750_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0471_),
    .A2(_0472_),
    .Y(_0194_),
    .B1(_0473_));
 sg13g2_mux2_1 _1751_ (.A0(\state[67] ),
    .A1(\daisychain[67] ),
    .S(net151),
    .X(_0474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1752_ (.Y(_0475_),
    .A(net173),
    .B(_0474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1753_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net129),
    .A2(\daisychain[66] ),
    .Y(_0476_),
    .B1(net63));
 sg13g2_o21ai_1 _1754_ (.B1(net196),
    .VDD(VPWR),
    .Y(_0477_),
    .VSS(VGND),
    .A1(\daisychain[67] ),
    .A2(net41));
 sg13g2_a21oi_1 _1755_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0475_),
    .A2(_0476_),
    .Y(_0195_),
    .B1(_0477_));
 sg13g2_mux2_1 _1756_ (.A0(\state[68] ),
    .A1(\daisychain[68] ),
    .S(net151),
    .X(_0478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1757_ (.Y(_0479_),
    .A(net173),
    .B(_0478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1758_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net129),
    .A2(\daisychain[67] ),
    .Y(_0480_),
    .B1(net63));
 sg13g2_o21ai_1 _1759_ (.B1(net196),
    .VDD(VPWR),
    .Y(_0481_),
    .VSS(VGND),
    .A1(\daisychain[68] ),
    .A2(net41));
 sg13g2_a21oi_1 _1760_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0479_),
    .A2(_0480_),
    .Y(_0196_),
    .B1(_0481_));
 sg13g2_mux2_1 _1761_ (.A0(\state[69] ),
    .A1(\daisychain[69] ),
    .S(net151),
    .X(_0482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1762_ (.Y(_0483_),
    .A(net173),
    .B(_0482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1763_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net128),
    .A2(\daisychain[68] ),
    .Y(_0484_),
    .B1(net63));
 sg13g2_o21ai_1 _1764_ (.B1(net197),
    .VDD(VPWR),
    .Y(_0485_),
    .VSS(VGND),
    .A1(\daisychain[69] ),
    .A2(net42));
 sg13g2_a21oi_1 _1765_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0483_),
    .A2(_0484_),
    .Y(_0197_),
    .B1(_0485_));
 sg13g2_mux2_1 _1766_ (.A0(\state[70] ),
    .A1(\daisychain[70] ),
    .S(net151),
    .X(_0486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1767_ (.Y(_0487_),
    .A(net173),
    .B(_0486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1768_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net128),
    .A2(\daisychain[69] ),
    .Y(_0488_),
    .B1(net64));
 sg13g2_o21ai_1 _1769_ (.B1(net197),
    .VDD(VPWR),
    .Y(_0489_),
    .VSS(VGND),
    .A1(\daisychain[70] ),
    .A2(net42));
 sg13g2_a21oi_1 _1770_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0487_),
    .A2(_0488_),
    .Y(_0198_),
    .B1(_0489_));
 sg13g2_mux2_1 _1771_ (.A0(\state[71] ),
    .A1(\daisychain[71] ),
    .S(net152),
    .X(_0490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1772_ (.Y(_0491_),
    .A(net174),
    .B(_0490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1773_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net128),
    .A2(\daisychain[70] ),
    .Y(_0492_),
    .B1(net64));
 sg13g2_o21ai_1 _1774_ (.B1(net197),
    .VDD(VPWR),
    .Y(_0493_),
    .VSS(VGND),
    .A1(\daisychain[71] ),
    .A2(net42));
 sg13g2_a21oi_1 _1775_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0491_),
    .A2(_0492_),
    .Y(_0199_),
    .B1(_0493_));
 sg13g2_mux2_1 _1776_ (.A0(\state[72] ),
    .A1(\daisychain[72] ),
    .S(net152),
    .X(_0494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1777_ (.Y(_0495_),
    .A(net174),
    .B(_0494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1778_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net128),
    .A2(\daisychain[71] ),
    .Y(_0496_),
    .B1(net64));
 sg13g2_o21ai_1 _1779_ (.B1(net197),
    .VDD(VPWR),
    .Y(_0497_),
    .VSS(VGND),
    .A1(\daisychain[72] ),
    .A2(net42));
 sg13g2_a21oi_1 _1780_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0495_),
    .A2(_0496_),
    .Y(_0200_),
    .B1(_0497_));
 sg13g2_mux2_1 _1781_ (.A0(\state[73] ),
    .A1(\daisychain[73] ),
    .S(net152),
    .X(_0498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1782_ (.Y(_0499_),
    .A(net174),
    .B(_0498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1783_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net128),
    .A2(\daisychain[72] ),
    .Y(_0500_),
    .B1(net64));
 sg13g2_o21ai_1 _1784_ (.B1(net197),
    .VDD(VPWR),
    .Y(_0501_),
    .VSS(VGND),
    .A1(\daisychain[73] ),
    .A2(net42));
 sg13g2_a21oi_1 _1785_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0499_),
    .A2(_0500_),
    .Y(_0201_),
    .B1(_0501_));
 sg13g2_mux2_1 _1786_ (.A0(\state[74] ),
    .A1(\daisychain[74] ),
    .S(net151),
    .X(_0502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1787_ (.Y(_0503_),
    .A(net173),
    .B(_0502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1788_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net127),
    .A2(\daisychain[73] ),
    .Y(_0504_),
    .B1(net63));
 sg13g2_o21ai_1 _1789_ (.B1(net196),
    .VDD(VPWR),
    .Y(_0505_),
    .VSS(VGND),
    .A1(\daisychain[74] ),
    .A2(net41));
 sg13g2_a21oi_1 _1790_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0503_),
    .A2(_0504_),
    .Y(_0202_),
    .B1(_0505_));
 sg13g2_mux2_1 _1791_ (.A0(\state[75] ),
    .A1(\daisychain[75] ),
    .S(net151),
    .X(_0506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1792_ (.Y(_0507_),
    .A(net173),
    .B(_0506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1793_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net127),
    .A2(\daisychain[74] ),
    .Y(_0508_),
    .B1(net63));
 sg13g2_o21ai_1 _1794_ (.B1(net196),
    .VDD(VPWR),
    .Y(_0509_),
    .VSS(VGND),
    .A1(\daisychain[75] ),
    .A2(net41));
 sg13g2_a21oi_1 _1795_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0507_),
    .A2(_0508_),
    .Y(_0203_),
    .B1(_0509_));
 sg13g2_mux2_1 _1796_ (.A0(\state[76] ),
    .A1(\daisychain[76] ),
    .S(net151),
    .X(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1797_ (.Y(_0511_),
    .A(net173),
    .B(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1798_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net127),
    .A2(\daisychain[75] ),
    .Y(_0512_),
    .B1(net63));
 sg13g2_o21ai_1 _1799_ (.B1(net196),
    .VDD(VPWR),
    .Y(_0513_),
    .VSS(VGND),
    .A1(\daisychain[76] ),
    .A2(net41));
 sg13g2_a21oi_1 _1800_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0511_),
    .A2(_0512_),
    .Y(_0204_),
    .B1(_0513_));
 sg13g2_mux2_1 _1801_ (.A0(\state[77] ),
    .A1(\daisychain[77] ),
    .S(net151),
    .X(_0514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1802_ (.Y(_0515_),
    .A(net173),
    .B(_0514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1803_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net127),
    .A2(\daisychain[76] ),
    .Y(_0516_),
    .B1(net63));
 sg13g2_o21ai_1 _1804_ (.B1(net196),
    .VDD(VPWR),
    .Y(_0517_),
    .VSS(VGND),
    .A1(\daisychain[77] ),
    .A2(net41));
 sg13g2_a21oi_1 _1805_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0515_),
    .A2(_0516_),
    .Y(_0205_),
    .B1(_0517_));
 sg13g2_mux2_1 _1806_ (.A0(\state[78] ),
    .A1(\daisychain[78] ),
    .S(net152),
    .X(_0518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1807_ (.Y(_0519_),
    .A(net174),
    .B(_0518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1808_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net127),
    .A2(\daisychain[77] ),
    .Y(_0520_),
    .B1(net63));
 sg13g2_o21ai_1 _1809_ (.B1(net196),
    .VDD(VPWR),
    .Y(_0521_),
    .VSS(VGND),
    .A1(\daisychain[78] ),
    .A2(net41));
 sg13g2_a21oi_1 _1810_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0519_),
    .A2(_0520_),
    .Y(_0206_),
    .B1(_0521_));
 sg13g2_mux2_1 _1811_ (.A0(\state[79] ),
    .A1(\daisychain[79] ),
    .S(net153),
    .X(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1812_ (.Y(_0523_),
    .A(net175),
    .B(_0522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1813_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net126),
    .A2(\daisychain[78] ),
    .Y(_0524_),
    .B1(net65));
 sg13g2_o21ai_1 _1814_ (.B1(net198),
    .VDD(VPWR),
    .Y(_0525_),
    .VSS(VGND),
    .A1(\daisychain[79] ),
    .A2(net43));
 sg13g2_a21oi_1 _1815_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0523_),
    .A2(_0524_),
    .Y(_0207_),
    .B1(_0525_));
 sg13g2_mux2_1 _1816_ (.A0(\state[80] ),
    .A1(\daisychain[80] ),
    .S(net153),
    .X(_0526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1817_ (.Y(_0527_),
    .A(net175),
    .B(_0526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1818_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net126),
    .A2(\daisychain[79] ),
    .Y(_0528_),
    .B1(net65));
 sg13g2_o21ai_1 _1819_ (.B1(net198),
    .VDD(VPWR),
    .Y(_0529_),
    .VSS(VGND),
    .A1(\daisychain[80] ),
    .A2(net43));
 sg13g2_a21oi_1 _1820_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0527_),
    .A2(_0528_),
    .Y(_0208_),
    .B1(_0529_));
 sg13g2_mux2_1 _1821_ (.A0(\state[81] ),
    .A1(\daisychain[81] ),
    .S(net153),
    .X(_0530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1822_ (.Y(_0531_),
    .A(net175),
    .B(_0530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1823_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net126),
    .A2(\daisychain[80] ),
    .Y(_0532_),
    .B1(net65));
 sg13g2_o21ai_1 _1824_ (.B1(net198),
    .VDD(VPWR),
    .Y(_0533_),
    .VSS(VGND),
    .A1(\daisychain[81] ),
    .A2(net43));
 sg13g2_a21oi_1 _1825_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0531_),
    .A2(_0532_),
    .Y(_0209_),
    .B1(_0533_));
 sg13g2_mux2_1 _1826_ (.A0(\state[82] ),
    .A1(\daisychain[82] ),
    .S(net150),
    .X(_0534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1827_ (.Y(_0535_),
    .A(net172),
    .B(_0534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1828_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net122),
    .A2(\daisychain[81] ),
    .Y(_0536_),
    .B1(net62));
 sg13g2_o21ai_1 _1829_ (.B1(net195),
    .VDD(VPWR),
    .Y(_0537_),
    .VSS(VGND),
    .A1(\daisychain[82] ),
    .A2(net40));
 sg13g2_a21oi_1 _1830_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0535_),
    .A2(_0536_),
    .Y(_0210_),
    .B1(_0537_));
 sg13g2_mux2_1 _1831_ (.A0(\state[83] ),
    .A1(\daisychain[83] ),
    .S(net150),
    .X(_0538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1832_ (.Y(_0539_),
    .A(net172),
    .B(_0538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1833_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net122),
    .A2(\daisychain[82] ),
    .Y(_0540_),
    .B1(net62));
 sg13g2_o21ai_1 _1834_ (.B1(net195),
    .VDD(VPWR),
    .Y(_0541_),
    .VSS(VGND),
    .A1(\daisychain[83] ),
    .A2(net40));
 sg13g2_a21oi_1 _1835_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0539_),
    .A2(_0540_),
    .Y(_0211_),
    .B1(_0541_));
 sg13g2_mux2_1 _1836_ (.A0(\state[84] ),
    .A1(\daisychain[84] ),
    .S(net150),
    .X(_0542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1837_ (.Y(_0543_),
    .A(net172),
    .B(_0542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1838_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net122),
    .A2(\daisychain[83] ),
    .Y(_0544_),
    .B1(net62));
 sg13g2_o21ai_1 _1839_ (.B1(net195),
    .VDD(VPWR),
    .Y(_0545_),
    .VSS(VGND),
    .A1(\daisychain[84] ),
    .A2(net40));
 sg13g2_a21oi_1 _1840_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0543_),
    .A2(_0544_),
    .Y(_0212_),
    .B1(_0545_));
 sg13g2_mux2_1 _1841_ (.A0(\state[85] ),
    .A1(\daisychain[85] ),
    .S(net148),
    .X(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1842_ (.Y(_0547_),
    .A(net170),
    .B(_0546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1843_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net122),
    .A2(\daisychain[84] ),
    .Y(_0548_),
    .B1(net62));
 sg13g2_o21ai_1 _1844_ (.B1(net193),
    .VDD(VPWR),
    .Y(_0549_),
    .VSS(VGND),
    .A1(\daisychain[85] ),
    .A2(net38));
 sg13g2_a21oi_1 _1845_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0547_),
    .A2(_0548_),
    .Y(_0213_),
    .B1(_0549_));
 sg13g2_mux2_1 _1846_ (.A0(\state[86] ),
    .A1(\daisychain[86] ),
    .S(net148),
    .X(_0550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1847_ (.Y(_0551_),
    .A(net170),
    .B(_0550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1848_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net123),
    .A2(\daisychain[85] ),
    .Y(_0552_),
    .B1(net61));
 sg13g2_o21ai_1 _1849_ (.B1(net193),
    .VDD(VPWR),
    .Y(_0553_),
    .VSS(VGND),
    .A1(\daisychain[86] ),
    .A2(net38));
 sg13g2_a21oi_1 _1850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0551_),
    .A2(_0552_),
    .Y(_0214_),
    .B1(_0553_));
 sg13g2_mux2_1 _1851_ (.A0(\state[87] ),
    .A1(\daisychain[87] ),
    .S(net148),
    .X(_0554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1852_ (.Y(_0555_),
    .A(net170),
    .B(_0554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1853_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net124),
    .A2(\daisychain[86] ),
    .Y(_0556_),
    .B1(net61));
 sg13g2_o21ai_1 _1854_ (.B1(net193),
    .VDD(VPWR),
    .Y(_0557_),
    .VSS(VGND),
    .A1(\daisychain[87] ),
    .A2(net38));
 sg13g2_a21oi_1 _1855_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0555_),
    .A2(_0556_),
    .Y(_0215_),
    .B1(_0557_));
 sg13g2_mux2_1 _1856_ (.A0(\state[88] ),
    .A1(\daisychain[88] ),
    .S(net149),
    .X(_0558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1857_ (.Y(_0559_),
    .A(net170),
    .B(_0558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1858_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net124),
    .A2(\daisychain[87] ),
    .Y(_0560_),
    .B1(net61));
 sg13g2_o21ai_1 _1859_ (.B1(net193),
    .VDD(VPWR),
    .Y(_0561_),
    .VSS(VGND),
    .A1(\daisychain[88] ),
    .A2(net38));
 sg13g2_a21oi_1 _1860_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0559_),
    .A2(_0560_),
    .Y(_0216_),
    .B1(_0561_));
 sg13g2_mux2_1 _1861_ (.A0(\state[89] ),
    .A1(\daisychain[89] ),
    .S(net149),
    .X(_0562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1862_ (.Y(_0563_),
    .A(net171),
    .B(_0562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1863_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net124),
    .A2(\daisychain[88] ),
    .Y(_0564_),
    .B1(net61));
 sg13g2_o21ai_1 _1864_ (.B1(net194),
    .VDD(VPWR),
    .Y(_0565_),
    .VSS(VGND),
    .A1(\daisychain[89] ),
    .A2(net39));
 sg13g2_a21oi_1 _1865_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0563_),
    .A2(_0564_),
    .Y(_0217_),
    .B1(_0565_));
 sg13g2_mux2_1 _1866_ (.A0(\state[90] ),
    .A1(\daisychain[90] ),
    .S(net149),
    .X(_0566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1867_ (.Y(_0567_),
    .A(net171),
    .B(_0566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1868_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net124),
    .A2(\daisychain[89] ),
    .Y(_0568_),
    .B1(net62));
 sg13g2_o21ai_1 _1869_ (.B1(net194),
    .VDD(VPWR),
    .Y(_0569_),
    .VSS(VGND),
    .A1(\daisychain[90] ),
    .A2(net39));
 sg13g2_a21oi_1 _1870_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0567_),
    .A2(_0568_),
    .Y(_0218_),
    .B1(_0569_));
 sg13g2_mux2_1 _1871_ (.A0(\state[91] ),
    .A1(\daisychain[91] ),
    .S(net149),
    .X(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1872_ (.Y(_0571_),
    .A(net171),
    .B(_0570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1873_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net124),
    .A2(\daisychain[90] ),
    .Y(_0572_),
    .B1(net62));
 sg13g2_o21ai_1 _1874_ (.B1(net194),
    .VDD(VPWR),
    .Y(_0573_),
    .VSS(VGND),
    .A1(\daisychain[91] ),
    .A2(net39));
 sg13g2_a21oi_1 _1875_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0571_),
    .A2(_0572_),
    .Y(_0219_),
    .B1(_0573_));
 sg13g2_mux2_1 _1876_ (.A0(\state[92] ),
    .A1(\daisychain[92] ),
    .S(net148),
    .X(_0574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1877_ (.Y(_0575_),
    .A(net171),
    .B(_0574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1878_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net125),
    .A2(\daisychain[91] ),
    .Y(_0576_),
    .B1(net62));
 sg13g2_o21ai_1 _1879_ (.B1(net194),
    .VDD(VPWR),
    .Y(_0577_),
    .VSS(VGND),
    .A1(\daisychain[92] ),
    .A2(net39));
 sg13g2_a21oi_1 _1880_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0575_),
    .A2(_0576_),
    .Y(_0220_),
    .B1(_0577_));
 sg13g2_mux2_1 _1881_ (.A0(\state[93] ),
    .A1(\daisychain[93] ),
    .S(net148),
    .X(_0578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1882_ (.Y(_0579_),
    .A(net170),
    .B(_0578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1883_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net123),
    .A2(\daisychain[92] ),
    .Y(_0580_),
    .B1(net61));
 sg13g2_o21ai_1 _1884_ (.B1(net193),
    .VDD(VPWR),
    .Y(_0581_),
    .VSS(VGND),
    .A1(\daisychain[93] ),
    .A2(net38));
 sg13g2_a21oi_1 _1885_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0579_),
    .A2(_0580_),
    .Y(_0221_),
    .B1(_0581_));
 sg13g2_mux2_1 _1886_ (.A0(\state[94] ),
    .A1(\daisychain[94] ),
    .S(net148),
    .X(_0582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1887_ (.Y(_0583_),
    .A(net170),
    .B(_0582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1888_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net123),
    .A2(\daisychain[93] ),
    .Y(_0584_),
    .B1(net61));
 sg13g2_o21ai_1 _1889_ (.B1(net193),
    .VDD(VPWR),
    .Y(_0585_),
    .VSS(VGND),
    .A1(\daisychain[94] ),
    .A2(net38));
 sg13g2_a21oi_1 _1890_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0583_),
    .A2(_0584_),
    .Y(_0222_),
    .B1(_0585_));
 sg13g2_mux2_1 _1891_ (.A0(\state[95] ),
    .A1(\daisychain[95] ),
    .S(net139),
    .X(_0586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1892_ (.Y(_0587_),
    .A(net163),
    .B(_0586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1893_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net106),
    .A2(\daisychain[94] ),
    .Y(_0588_),
    .B1(net53));
 sg13g2_o21ai_1 _1894_ (.B1(net185),
    .VDD(VPWR),
    .Y(_0589_),
    .VSS(VGND),
    .A1(\daisychain[95] ),
    .A2(net30));
 sg13g2_a21oi_1 _1895_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0587_),
    .A2(_0588_),
    .Y(_0223_),
    .B1(_0589_));
 sg13g2_mux2_1 _1896_ (.A0(\state[96] ),
    .A1(\daisychain[96] ),
    .S(net140),
    .X(_0590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1897_ (.Y(_0591_),
    .A(net163),
    .B(_0590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1898_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net106),
    .A2(\daisychain[95] ),
    .Y(_0592_),
    .B1(net53));
 sg13g2_o21ai_1 _1899_ (.B1(net186),
    .VDD(VPWR),
    .Y(_0593_),
    .VSS(VGND),
    .A1(\daisychain[96] ),
    .A2(net31));
 sg13g2_a21oi_1 _1900_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0591_),
    .A2(_0592_),
    .Y(_0224_),
    .B1(_0593_));
 sg13g2_mux2_1 _1901_ (.A0(\state[97] ),
    .A1(\daisychain[97] ),
    .S(net140),
    .X(_0594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1902_ (.Y(_0595_),
    .A(net163),
    .B(_0594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1903_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net106),
    .A2(\daisychain[96] ),
    .Y(_0596_),
    .B1(net53));
 sg13g2_o21ai_1 _1904_ (.B1(net186),
    .VDD(VPWR),
    .Y(_0597_),
    .VSS(VGND),
    .A1(\daisychain[97] ),
    .A2(net31));
 sg13g2_a21oi_1 _1905_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0595_),
    .A2(_0596_),
    .Y(_0225_),
    .B1(_0597_));
 sg13g2_mux2_1 _1906_ (.A0(\state[98] ),
    .A1(\daisychain[98] ),
    .S(net148),
    .X(_0598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1907_ (.Y(_0599_),
    .A(net170),
    .B(_0598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1908_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net123),
    .A2(\daisychain[97] ),
    .Y(_0600_),
    .B1(net61));
 sg13g2_o21ai_1 _1909_ (.B1(net193),
    .VDD(VPWR),
    .Y(_0601_),
    .VSS(VGND),
    .A1(\daisychain[98] ),
    .A2(net38));
 sg13g2_a21oi_1 _1910_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0599_),
    .A2(_0600_),
    .Y(_0226_),
    .B1(_0601_));
 sg13g2_mux2_1 _1911_ (.A0(\state[99] ),
    .A1(\daisychain[99] ),
    .S(net148),
    .X(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1912_ (.Y(_0603_),
    .A(net170),
    .B(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1913_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net123),
    .A2(\daisychain[98] ),
    .Y(_0604_),
    .B1(net61));
 sg13g2_o21ai_1 _1914_ (.B1(net193),
    .VDD(VPWR),
    .Y(_0605_),
    .VSS(VGND),
    .A1(\daisychain[99] ),
    .A2(net38));
 sg13g2_a21oi_1 _1915_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0603_),
    .A2(_0604_),
    .Y(_0227_),
    .B1(_0605_));
 sg13g2_mux2_1 _1916_ (.A0(\state[100] ),
    .A1(\daisychain[100] ),
    .S(net139),
    .X(_0606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1917_ (.Y(_0607_),
    .A(net162),
    .B(_0606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1918_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net106),
    .A2(\daisychain[99] ),
    .Y(_0608_),
    .B1(net53));
 sg13g2_o21ai_1 _1919_ (.B1(net185),
    .VDD(VPWR),
    .Y(_0609_),
    .VSS(VGND),
    .A1(\daisychain[100] ),
    .A2(net30));
 sg13g2_a21oi_1 _1920_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0607_),
    .A2(_0608_),
    .Y(_0228_),
    .B1(_0609_));
 sg13g2_mux2_1 _1921_ (.A0(\state[101] ),
    .A1(\daisychain[101] ),
    .S(net139),
    .X(_0610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1922_ (.Y(_0611_),
    .A(net162),
    .B(_0610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1923_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net105),
    .A2(\daisychain[100] ),
    .Y(_0612_),
    .B1(net52));
 sg13g2_o21ai_1 _1924_ (.B1(net185),
    .VDD(VPWR),
    .Y(_0613_),
    .VSS(VGND),
    .A1(\daisychain[101] ),
    .A2(net30));
 sg13g2_a21oi_1 _1925_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0611_),
    .A2(_0612_),
    .Y(_0229_),
    .B1(_0613_));
 sg13g2_mux2_1 _1926_ (.A0(\state[102] ),
    .A1(\daisychain[102] ),
    .S(net139),
    .X(_0614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1927_ (.Y(_0615_),
    .A(net162),
    .B(_0614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1928_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net105),
    .A2(\daisychain[101] ),
    .Y(_0616_),
    .B1(net52));
 sg13g2_o21ai_1 _1929_ (.B1(net185),
    .VDD(VPWR),
    .Y(_0617_),
    .VSS(VGND),
    .A1(\daisychain[102] ),
    .A2(net30));
 sg13g2_a21oi_1 _1930_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0615_),
    .A2(_0616_),
    .Y(_0230_),
    .B1(_0617_));
 sg13g2_mux2_1 _1931_ (.A0(\state[103] ),
    .A1(\daisychain[103] ),
    .S(net139),
    .X(_0618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1932_ (.Y(_0619_),
    .A(net163),
    .B(_0618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1933_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net105),
    .A2(\daisychain[102] ),
    .Y(_0620_),
    .B1(net52));
 sg13g2_o21ai_1 _1934_ (.B1(net185),
    .VDD(VPWR),
    .Y(_0621_),
    .VSS(VGND),
    .A1(\daisychain[103] ),
    .A2(net30));
 sg13g2_a21oi_1 _1935_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0619_),
    .A2(_0620_),
    .Y(_0231_),
    .B1(_0621_));
 sg13g2_mux2_1 _1936_ (.A0(\state[104] ),
    .A1(\daisychain[104] ),
    .S(net139),
    .X(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1937_ (.Y(_0623_),
    .A(net162),
    .B(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1938_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net104),
    .A2(\daisychain[103] ),
    .Y(_0624_),
    .B1(net52));
 sg13g2_o21ai_1 _1939_ (.B1(net185),
    .VDD(VPWR),
    .Y(_0625_),
    .VSS(VGND),
    .A1(\daisychain[104] ),
    .A2(net30));
 sg13g2_a21oi_1 _1940_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0623_),
    .A2(_0624_),
    .Y(_0232_),
    .B1(_0625_));
 sg13g2_mux2_1 _1941_ (.A0(\state[105] ),
    .A1(\daisychain[105] ),
    .S(net139),
    .X(_0626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1942_ (.Y(_0627_),
    .A(net162),
    .B(_0626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1943_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net104),
    .A2(\daisychain[104] ),
    .Y(_0628_),
    .B1(net52));
 sg13g2_o21ai_1 _1944_ (.B1(net185),
    .VDD(VPWR),
    .Y(_0629_),
    .VSS(VGND),
    .A1(\daisychain[105] ),
    .A2(net30));
 sg13g2_a21oi_1 _1945_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0627_),
    .A2(_0628_),
    .Y(_0233_),
    .B1(_0629_));
 sg13g2_mux2_1 _1946_ (.A0(\state[106] ),
    .A1(\daisychain[106] ),
    .S(net139),
    .X(_0630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1947_ (.Y(_0631_),
    .A(net162),
    .B(_0630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1948_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net104),
    .A2(\daisychain[105] ),
    .Y(_0632_),
    .B1(net52));
 sg13g2_o21ai_1 _1949_ (.B1(net185),
    .VDD(VPWR),
    .Y(_0633_),
    .VSS(VGND),
    .A1(\daisychain[106] ),
    .A2(net30));
 sg13g2_a21oi_1 _1950_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0631_),
    .A2(_0632_),
    .Y(_0234_),
    .B1(_0633_));
 sg13g2_mux2_1 _1951_ (.A0(\state[107] ),
    .A1(\daisychain[107] ),
    .S(net140),
    .X(_0634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1952_ (.Y(_0635_),
    .A(net163),
    .B(_0634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1953_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net104),
    .A2(\daisychain[106] ),
    .Y(_0636_),
    .B1(net52));
 sg13g2_o21ai_1 _1954_ (.B1(net186),
    .VDD(VPWR),
    .Y(_0637_),
    .VSS(VGND),
    .A1(\daisychain[107] ),
    .A2(net31));
 sg13g2_a21oi_1 _1955_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0635_),
    .A2(_0636_),
    .Y(_0235_),
    .B1(_0637_));
 sg13g2_mux2_1 _1956_ (.A0(\state[108] ),
    .A1(\daisychain[108] ),
    .S(net140),
    .X(_0638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1957_ (.Y(_0639_),
    .A(net163),
    .B(_0638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1958_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net107),
    .A2(\daisychain[107] ),
    .Y(_0640_),
    .B1(net53));
 sg13g2_o21ai_1 _1959_ (.B1(net186),
    .VDD(VPWR),
    .Y(_0641_),
    .VSS(VGND),
    .A1(\daisychain[108] ),
    .A2(net31));
 sg13g2_a21oi_1 _1960_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0639_),
    .A2(_0640_),
    .Y(_0236_),
    .B1(_0641_));
 sg13g2_mux2_1 _1961_ (.A0(\state[109] ),
    .A1(\daisychain[109] ),
    .S(net140),
    .X(_0642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1962_ (.Y(_0643_),
    .A(net163),
    .B(_0642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1963_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net107),
    .A2(\daisychain[108] ),
    .Y(_0644_),
    .B1(net53));
 sg13g2_o21ai_1 _1964_ (.B1(net186),
    .VDD(VPWR),
    .Y(_0645_),
    .VSS(VGND),
    .A1(\daisychain[109] ),
    .A2(net31));
 sg13g2_a21oi_1 _1965_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0643_),
    .A2(_0644_),
    .Y(_0237_),
    .B1(_0645_));
 sg13g2_mux2_1 _1966_ (.A0(\state[110] ),
    .A1(\daisychain[110] ),
    .S(net140),
    .X(_0646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1967_ (.Y(_0647_),
    .A(net164),
    .B(_0646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1968_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net107),
    .A2(\daisychain[109] ),
    .Y(_0648_),
    .B1(net53));
 sg13g2_o21ai_1 _1969_ (.B1(net186),
    .VDD(VPWR),
    .Y(_0649_),
    .VSS(VGND),
    .A1(\daisychain[110] ),
    .A2(net31));
 sg13g2_a21oi_1 _1970_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0647_),
    .A2(_0648_),
    .Y(_0238_),
    .B1(_0649_));
 sg13g2_mux2_1 _1971_ (.A0(\state[111] ),
    .A1(\daisychain[111] ),
    .S(net141),
    .X(_0650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1972_ (.Y(_0651_),
    .A(net162),
    .B(_0650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1973_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net108),
    .A2(\daisychain[110] ),
    .Y(_0652_),
    .B1(net54));
 sg13g2_o21ai_1 _1974_ (.B1(net184),
    .VDD(VPWR),
    .Y(_0653_),
    .VSS(VGND),
    .A1(\daisychain[111] ),
    .A2(net29));
 sg13g2_a21oi_1 _1975_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0651_),
    .A2(_0652_),
    .Y(_0239_),
    .B1(_0653_));
 sg13g2_mux2_1 _1976_ (.A0(\state[112] ),
    .A1(\daisychain[112] ),
    .S(net141),
    .X(_0654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1977_ (.Y(_0655_),
    .A(net164),
    .B(_0654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1978_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net102),
    .A2(\daisychain[111] ),
    .Y(_0656_),
    .B1(net51));
 sg13g2_o21ai_1 _1979_ (.B1(net184),
    .VDD(VPWR),
    .Y(_0657_),
    .VSS(VGND),
    .A1(\daisychain[112] ),
    .A2(net29));
 sg13g2_a21oi_1 _1980_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0655_),
    .A2(_0656_),
    .Y(_0240_),
    .B1(_0657_));
 sg13g2_mux2_1 _1981_ (.A0(\state[113] ),
    .A1(\daisychain[113] ),
    .S(net141),
    .X(_0658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1982_ (.Y(_0659_),
    .A(net164),
    .B(_0658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1983_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net102),
    .A2(\daisychain[112] ),
    .Y(_0660_),
    .B1(net51));
 sg13g2_o21ai_1 _1984_ (.B1(net184),
    .VDD(VPWR),
    .Y(_0661_),
    .VSS(VGND),
    .A1(\daisychain[113] ),
    .A2(net29));
 sg13g2_a21oi_1 _1985_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0659_),
    .A2(_0660_),
    .Y(_0241_),
    .B1(_0661_));
 sg13g2_mux2_1 _1986_ (.A0(\state[114] ),
    .A1(\daisychain[114] ),
    .S(net141),
    .X(_0662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1987_ (.Y(_0663_),
    .A(net162),
    .B(_0662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1988_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net102),
    .A2(\daisychain[113] ),
    .Y(_0664_),
    .B1(net51));
 sg13g2_o21ai_1 _1989_ (.B1(net184),
    .VDD(VPWR),
    .Y(_0665_),
    .VSS(VGND),
    .A1(\daisychain[114] ),
    .A2(net29));
 sg13g2_a21oi_1 _1990_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0663_),
    .A2(_0664_),
    .Y(_0242_),
    .B1(_0665_));
 sg13g2_mux2_1 _1991_ (.A0(\state[115] ),
    .A1(\daisychain[115] ),
    .S(net141),
    .X(_0666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1992_ (.Y(_0667_),
    .A(net164),
    .B(_0666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1993_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net102),
    .A2(\daisychain[114] ),
    .Y(_0668_),
    .B1(net51));
 sg13g2_o21ai_1 _1994_ (.B1(net187),
    .VDD(VPWR),
    .Y(_0669_),
    .VSS(VGND),
    .A1(\daisychain[115] ),
    .A2(net32));
 sg13g2_a21oi_1 _1995_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0667_),
    .A2(_0668_),
    .Y(_0243_),
    .B1(_0669_));
 sg13g2_mux2_1 _1996_ (.A0(\state[116] ),
    .A1(\daisychain[116] ),
    .S(net141),
    .X(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _1997_ (.Y(_0671_),
    .A(net164),
    .B(_0670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _1998_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net102),
    .A2(\daisychain[115] ),
    .Y(_0672_),
    .B1(net54));
 sg13g2_o21ai_1 _1999_ (.B1(net184),
    .VDD(VPWR),
    .Y(_0673_),
    .VSS(VGND),
    .A1(\daisychain[116] ),
    .A2(net29));
 sg13g2_a21oi_1 _2000_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0671_),
    .A2(_0672_),
    .Y(_0244_),
    .B1(_0673_));
 sg13g2_mux2_1 _2001_ (.A0(\state[117] ),
    .A1(\daisychain[117] ),
    .S(net141),
    .X(_0674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2002_ (.Y(_0675_),
    .A(net164),
    .B(_0674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2003_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net103),
    .A2(\daisychain[116] ),
    .Y(_0676_),
    .B1(net51));
 sg13g2_o21ai_1 _2004_ (.B1(net184),
    .VDD(VPWR),
    .Y(_0677_),
    .VSS(VGND),
    .A1(\daisychain[117] ),
    .A2(net29));
 sg13g2_a21oi_1 _2005_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0675_),
    .A2(_0676_),
    .Y(_0245_),
    .B1(_0677_));
 sg13g2_mux2_1 _2006_ (.A0(\state[118] ),
    .A1(\daisychain[118] ),
    .S(net141),
    .X(_0678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2007_ (.Y(_0679_),
    .A(net164),
    .B(_0678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2008_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net103),
    .A2(\daisychain[117] ),
    .Y(_0680_),
    .B1(net51));
 sg13g2_o21ai_1 _2009_ (.B1(net184),
    .VDD(VPWR),
    .Y(_0681_),
    .VSS(VGND),
    .A1(\daisychain[118] ),
    .A2(net29));
 sg13g2_a21oi_1 _2010_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0679_),
    .A2(_0680_),
    .Y(_0246_),
    .B1(_0681_));
 sg13g2_mux2_1 _2011_ (.A0(\state[119] ),
    .A1(\daisychain[119] ),
    .S(net134),
    .X(_0682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2012_ (.Y(_0683_),
    .A(net157),
    .B(_0682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2013_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net92),
    .A2(\daisychain[118] ),
    .Y(_0684_),
    .B1(net51));
 sg13g2_o21ai_1 _2014_ (.B1(net179),
    .VDD(VPWR),
    .Y(_0685_),
    .VSS(VGND),
    .A1(\daisychain[119] ),
    .A2(net24));
 sg13g2_a21oi_1 _2015_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0683_),
    .A2(_0684_),
    .Y(_0247_),
    .B1(_0685_));
 sg13g2_mux2_1 _2016_ (.A0(\state[120] ),
    .A1(\daisychain[120] ),
    .S(net133),
    .X(_0686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2017_ (.Y(_0687_),
    .A(net157),
    .B(_0686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2018_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net92),
    .A2(\daisychain[119] ),
    .Y(_0688_),
    .B1(net67));
 sg13g2_o21ai_1 _2019_ (.B1(net179),
    .VDD(VPWR),
    .Y(_0689_),
    .VSS(VGND),
    .A1(\daisychain[120] ),
    .A2(net23));
 sg13g2_a21oi_1 _2020_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0687_),
    .A2(_0688_),
    .Y(_0248_),
    .B1(_0689_));
 sg13g2_mux2_1 _2021_ (.A0(\state[121] ),
    .A1(\daisychain[121] ),
    .S(net133),
    .X(_0690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2022_ (.Y(_0691_),
    .A(net156),
    .B(_0690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2023_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net90),
    .A2(\daisychain[120] ),
    .Y(_0692_),
    .B1(net46));
 sg13g2_o21ai_1 _2024_ (.B1(net178),
    .VDD(VPWR),
    .Y(_0693_),
    .VSS(VGND),
    .A1(\daisychain[121] ),
    .A2(net23));
 sg13g2_a21oi_1 _2025_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0691_),
    .A2(_0692_),
    .Y(_0249_),
    .B1(_0693_));
 sg13g2_mux2_1 _2026_ (.A0(\state[122] ),
    .A1(\daisychain[122] ),
    .S(net133),
    .X(_0694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2027_ (.Y(_0695_),
    .A(net156),
    .B(_0694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2028_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net90),
    .A2(\daisychain[121] ),
    .Y(_0696_),
    .B1(net46));
 sg13g2_o21ai_1 _2029_ (.B1(net178),
    .VDD(VPWR),
    .Y(_0697_),
    .VSS(VGND),
    .A1(\daisychain[122] ),
    .A2(net23));
 sg13g2_a21oi_1 _2030_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0695_),
    .A2(_0696_),
    .Y(_0250_),
    .B1(_0697_));
 sg13g2_mux2_1 _2031_ (.A0(\state[123] ),
    .A1(\daisychain[123] ),
    .S(net133),
    .X(_0698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2032_ (.Y(_0699_),
    .A(net156),
    .B(_0698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2033_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net90),
    .A2(\daisychain[122] ),
    .Y(_0700_),
    .B1(net46));
 sg13g2_o21ai_1 _2034_ (.B1(net178),
    .VDD(VPWR),
    .Y(_0701_),
    .VSS(VGND),
    .A1(\daisychain[123] ),
    .A2(net23));
 sg13g2_a21oi_1 _2035_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0699_),
    .A2(_0700_),
    .Y(_0251_),
    .B1(_0701_));
 sg13g2_mux2_1 _2036_ (.A0(\state[124] ),
    .A1(\daisychain[124] ),
    .S(net133),
    .X(_0702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2037_ (.Y(_0703_),
    .A(net156),
    .B(_0702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2038_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net90),
    .A2(\daisychain[123] ),
    .Y(_0704_),
    .B1(net46));
 sg13g2_o21ai_1 _2039_ (.B1(net178),
    .VDD(VPWR),
    .Y(_0705_),
    .VSS(VGND),
    .A1(\daisychain[124] ),
    .A2(net23));
 sg13g2_a21oi_1 _2040_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0703_),
    .A2(_0704_),
    .Y(_0252_),
    .B1(_0705_));
 sg13g2_mux2_1 _2041_ (.A0(\state[125] ),
    .A1(\daisychain[125] ),
    .S(net133),
    .X(_0706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2042_ (.Y(_0707_),
    .A(net156),
    .B(_0706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2043_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net90),
    .A2(\daisychain[124] ),
    .Y(_0708_),
    .B1(net46));
 sg13g2_o21ai_1 _2044_ (.B1(net178),
    .VDD(VPWR),
    .Y(_0709_),
    .VSS(VGND),
    .A1(\daisychain[125] ),
    .A2(net23));
 sg13g2_a21oi_1 _2045_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0707_),
    .A2(_0708_),
    .Y(_0253_),
    .B1(_0709_));
 sg13g2_mux2_1 _2046_ (.A0(\state[126] ),
    .A1(\daisychain[126] ),
    .S(net133),
    .X(_0710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2047_ (.Y(_0711_),
    .A(net156),
    .B(_0710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2048_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net91),
    .A2(\daisychain[125] ),
    .Y(_0712_),
    .B1(net46));
 sg13g2_o21ai_1 _2049_ (.B1(net178),
    .VDD(VPWR),
    .Y(_0713_),
    .VSS(VGND),
    .A1(\daisychain[126] ),
    .A2(net23));
 sg13g2_a21oi_1 _2050_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0711_),
    .A2(_0712_),
    .Y(_0254_),
    .B1(_0713_));
 sg13g2_mux2_1 _2051_ (.A0(\state[127] ),
    .A1(\daisychain[127] ),
    .S(net133),
    .X(_0714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2052_ (.Y(_0715_),
    .A(net156),
    .B(_0714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2053_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net91),
    .A2(\daisychain[126] ),
    .Y(_0716_),
    .B1(net46));
 sg13g2_o21ai_1 _2054_ (.B1(net178),
    .VDD(VPWR),
    .Y(_0717_),
    .VSS(VGND),
    .A1(\daisychain[127] ),
    .A2(net23));
 sg13g2_a21oi_1 _2055_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0715_),
    .A2(_0716_),
    .Y(_0255_),
    .B1(_0717_));
 sg13g2_nand2_1 _2056_ (.Y(_0718_),
    .A(net92),
    .B(\state[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2057_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0849_),
    .A2(_0718_),
    .Y(_0256_),
    .B1(net69));
 sg13g2_nand2_1 _2058_ (.Y(_0719_),
    .A(net92),
    .B(\state[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2059_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0855_),
    .A2(_0719_),
    .Y(_0257_),
    .B1(net69));
 sg13g2_nand2_1 _2060_ (.Y(_0720_),
    .A(net92),
    .B(\state[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2061_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0859_),
    .A2(_0720_),
    .Y(_0258_),
    .B1(net69));
 sg13g2_nand2_1 _2062_ (.Y(_0721_),
    .A(net94),
    .B(\state[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2063_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0863_),
    .A2(_0721_),
    .Y(_0259_),
    .B1(net70));
 sg13g2_nand2_1 _2064_ (.Y(_0722_),
    .A(net95),
    .B(\state[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2065_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0867_),
    .A2(_0722_),
    .Y(_0260_),
    .B1(net70));
 sg13g2_nand2_1 _2066_ (.Y(_0723_),
    .A(net95),
    .B(\state[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2067_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0871_),
    .A2(_0723_),
    .Y(_0261_),
    .B1(net70));
 sg13g2_nand2_1 _2068_ (.Y(_0724_),
    .A(net99),
    .B(\state[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2069_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0875_),
    .A2(_0724_),
    .Y(_0262_),
    .B1(net72));
 sg13g2_nand2_1 _2070_ (.Y(_0725_),
    .A(net100),
    .B(\state[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2071_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0879_),
    .A2(_0725_),
    .Y(_0263_),
    .B1(net72));
 sg13g2_nand2_1 _2072_ (.Y(_0726_),
    .A(net99),
    .B(\state[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2073_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0883_),
    .A2(_0726_),
    .Y(_0264_),
    .B1(net72));
 sg13g2_nand2_1 _2074_ (.Y(_0727_),
    .A(net95),
    .B(\state[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2075_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0887_),
    .A2(_0727_),
    .Y(_0265_),
    .B1(net70));
 sg13g2_nand2_1 _2076_ (.Y(_0728_),
    .A(net96),
    .B(\state[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2077_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0891_),
    .A2(_0728_),
    .Y(_0266_),
    .B1(net70));
 sg13g2_nand2_1 _2078_ (.Y(_0729_),
    .A(net96),
    .B(\state[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2079_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0895_),
    .A2(_0729_),
    .Y(_0267_),
    .B1(net70));
 sg13g2_nand2_1 _2080_ (.Y(_0730_),
    .A(net96),
    .B(\state[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2081_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0899_),
    .A2(_0730_),
    .Y(_0268_),
    .B1(net69));
 sg13g2_nand2_1 _2082_ (.Y(_0731_),
    .A(net94),
    .B(\state[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2083_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0903_),
    .A2(_0731_),
    .Y(_0269_),
    .B1(net70));
 sg13g2_nand2_1 _2084_ (.Y(_0732_),
    .A(net95),
    .B(\state[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2085_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0907_),
    .A2(_0732_),
    .Y(_0270_),
    .B1(net70));
 sg13g2_nand2_1 _2086_ (.Y(_0733_),
    .A(net95),
    .B(\state[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2087_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0911_),
    .A2(_0733_),
    .Y(_0271_),
    .B1(net73));
 sg13g2_nand2_1 _2088_ (.Y(_0734_),
    .A(net99),
    .B(\state[16] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2089_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0915_),
    .A2(_0734_),
    .Y(_0272_),
    .B1(net73));
 sg13g2_nand2_1 _2090_ (.Y(_0735_),
    .A(net98),
    .B(\state[17] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2091_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0919_),
    .A2(_0735_),
    .Y(_0273_),
    .B1(net71));
 sg13g2_nand2_1 _2092_ (.Y(_0736_),
    .A(net98),
    .B(\state[18] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2093_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0923_),
    .A2(_0736_),
    .Y(_0274_),
    .B1(net71));
 sg13g2_nand2_1 _2094_ (.Y(_0737_),
    .A(net98),
    .B(\state[19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2095_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0927_),
    .A2(_0737_),
    .Y(_0275_),
    .B1(net71));
 sg13g2_nand2_1 _2096_ (.Y(_0738_),
    .A(net97),
    .B(\state[20] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2097_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0931_),
    .A2(_0738_),
    .Y(_0276_),
    .B1(net71));
 sg13g2_nand2_1 _2098_ (.Y(_0739_),
    .A(net97),
    .B(\state[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2099_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0935_),
    .A2(_0739_),
    .Y(_0277_),
    .B1(net71));
 sg13g2_nand2_1 _2100_ (.Y(_0740_),
    .A(net97),
    .B(\state[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2101_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0939_),
    .A2(_0740_),
    .Y(_0278_),
    .B1(net71));
 sg13g2_nand2_1 _2102_ (.Y(_0741_),
    .A(net101),
    .B(\state[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2103_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0943_),
    .A2(_0741_),
    .Y(_0279_),
    .B1(net71));
 sg13g2_nand2_1 _2104_ (.Y(_0742_),
    .A(net100),
    .B(\state[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2105_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0947_),
    .A2(_0742_),
    .Y(_0280_),
    .B1(net71));
 sg13g2_nand2_1 _2106_ (.Y(_0743_),
    .A(net100),
    .B(\state[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2107_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0951_),
    .A2(_0743_),
    .Y(_0281_),
    .B1(net72));
 sg13g2_nand2_1 _2108_ (.Y(_0744_),
    .A(net99),
    .B(\state[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2109_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0955_),
    .A2(_0744_),
    .Y(_0282_),
    .B1(net72));
 sg13g2_nand2_1 _2110_ (.Y(_0745_),
    .A(net101),
    .B(\state[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2111_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0959_),
    .A2(_0745_),
    .Y(_0283_),
    .B1(net72));
 sg13g2_nand2_1 _2112_ (.Y(_0746_),
    .A(net100),
    .B(\state[28] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2113_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0963_),
    .A2(_0746_),
    .Y(_0284_),
    .B1(net72));
 sg13g2_nand2_1 _2114_ (.Y(_0747_),
    .A(net101),
    .B(\state[29] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2115_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0967_),
    .A2(_0747_),
    .Y(_0285_),
    .B1(net72));
 sg13g2_nand2_1 _2116_ (.Y(_0748_),
    .A(net113),
    .B(\state[30] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2117_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0971_),
    .A2(_0748_),
    .Y(_0286_),
    .B1(net79));
 sg13g2_nand2_1 _2118_ (.Y(_0749_),
    .A(net113),
    .B(\state[31] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2119_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0975_),
    .A2(_0749_),
    .Y(_0287_),
    .B1(net79));
 sg13g2_nand2_1 _2120_ (.Y(_0750_),
    .A(net113),
    .B(\state[32] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2121_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0979_),
    .A2(_0750_),
    .Y(_0288_),
    .B1(net78));
 sg13g2_nand2_1 _2122_ (.Y(_0751_),
    .A(net112),
    .B(\state[33] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2123_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0983_),
    .A2(_0751_),
    .Y(_0289_),
    .B1(net78));
 sg13g2_nand2_1 _2124_ (.Y(_0752_),
    .A(net112),
    .B(\state[34] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2125_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0987_),
    .A2(_0752_),
    .Y(_0290_),
    .B1(net78));
 sg13g2_nand2_1 _2126_ (.Y(_0753_),
    .A(net111),
    .B(\state[35] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2127_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0991_),
    .A2(_0753_),
    .Y(_0291_),
    .B1(net78));
 sg13g2_nand2_1 _2128_ (.Y(_0754_),
    .A(net110),
    .B(\state[36] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2129_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0995_),
    .A2(_0754_),
    .Y(_0292_),
    .B1(net78));
 sg13g2_nand2_1 _2130_ (.Y(_0755_),
    .A(net110),
    .B(\state[37] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2131_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0999_),
    .A2(_0755_),
    .Y(_0293_),
    .B1(net78));
 sg13g2_nand2_1 _2132_ (.Y(_0756_),
    .A(net110),
    .B(\state[38] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2133_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1003_),
    .A2(_0756_),
    .Y(_0294_),
    .B1(net78));
 sg13g2_nand2_1 _2134_ (.Y(_0757_),
    .A(net111),
    .B(\state[39] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2135_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1007_),
    .A2(_0757_),
    .Y(_0295_),
    .B1(net78));
 sg13g2_nand2_1 _2136_ (.Y(_0758_),
    .A(net111),
    .B(\state[40] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2137_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1011_),
    .A2(_0758_),
    .Y(_0296_),
    .B1(net79));
 sg13g2_nand2_1 _2138_ (.Y(_0759_),
    .A(net115),
    .B(\state[41] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2139_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1015_),
    .A2(_0759_),
    .Y(_0297_),
    .B1(net80));
 sg13g2_nand2_1 _2140_ (.Y(_0760_),
    .A(net118),
    .B(\state[42] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2141_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1019_),
    .A2(_0760_),
    .Y(_0298_),
    .B1(net79));
 sg13g2_nand2_1 _2142_ (.Y(_0761_),
    .A(net112),
    .B(\state[43] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2143_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1023_),
    .A2(_0761_),
    .Y(_0299_),
    .B1(net79));
 sg13g2_nand2_1 _2144_ (.Y(_0762_),
    .A(net113),
    .B(\state[44] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2145_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1027_),
    .A2(_0762_),
    .Y(_0300_),
    .B1(net79));
 sg13g2_nand2_1 _2146_ (.Y(_0763_),
    .A(net114),
    .B(\state[45] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2147_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0387_),
    .A2(_0763_),
    .Y(_0301_),
    .B1(net79));
 sg13g2_nand2_1 _2148_ (.Y(_0764_),
    .A(net114),
    .B(\state[46] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2149_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0391_),
    .A2(_0764_),
    .Y(_0302_),
    .B1(net88));
 sg13g2_nand2_1 _2150_ (.Y(_0765_),
    .A(net119),
    .B(\state[47] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2151_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0395_),
    .A2(_0765_),
    .Y(_0303_),
    .B1(net82));
 sg13g2_nand2_1 _2152_ (.Y(_0766_),
    .A(net120),
    .B(\state[48] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2153_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0399_),
    .A2(_0766_),
    .Y(_0304_),
    .B1(net82));
 sg13g2_nand2_1 _2154_ (.Y(_0767_),
    .A(net119),
    .B(\state[49] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2155_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0403_),
    .A2(_0767_),
    .Y(_0305_),
    .B1(net82));
 sg13g2_nand2_1 _2156_ (.Y(_0768_),
    .A(net118),
    .B(\state[50] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2157_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0407_),
    .A2(_0768_),
    .Y(_0306_),
    .B1(net80));
 sg13g2_nand2_1 _2158_ (.Y(_0769_),
    .A(net118),
    .B(\state[51] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2159_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0411_),
    .A2(_0769_),
    .Y(_0307_),
    .B1(net80));
 sg13g2_nand2_1 _2160_ (.Y(_0770_),
    .A(net116),
    .B(\state[52] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2161_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0415_),
    .A2(_0770_),
    .Y(_0308_),
    .B1(net80));
 sg13g2_nand2_1 _2162_ (.Y(_0771_),
    .A(net115),
    .B(\state[53] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2163_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0419_),
    .A2(_0771_),
    .Y(_0309_),
    .B1(net80));
 sg13g2_nand2_1 _2164_ (.Y(_0772_),
    .A(net115),
    .B(\state[54] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2165_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0423_),
    .A2(_0772_),
    .Y(_0310_),
    .B1(net80));
 sg13g2_nand2_1 _2166_ (.Y(_0773_),
    .A(net116),
    .B(\state[55] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2167_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0427_),
    .A2(_0773_),
    .Y(_0311_),
    .B1(net80));
 sg13g2_nand2_1 _2168_ (.Y(_0774_),
    .A(net116),
    .B(\state[56] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2169_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0431_),
    .A2(_0774_),
    .Y(_0312_),
    .B1(net80));
 sg13g2_nand2_1 _2170_ (.Y(_0775_),
    .A(net116),
    .B(\state[57] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2171_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0435_),
    .A2(_0775_),
    .Y(_0313_),
    .B1(net81));
 sg13g2_nand2_1 _2172_ (.Y(_0776_),
    .A(net117),
    .B(\state[58] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2173_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0439_),
    .A2(_0776_),
    .Y(_0314_),
    .B1(net81));
 sg13g2_nand2_1 _2174_ (.Y(_0777_),
    .A(net117),
    .B(\state[59] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2175_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0443_),
    .A2(_0777_),
    .Y(_0315_),
    .B1(net81));
 sg13g2_nand2_1 _2176_ (.Y(_0778_),
    .A(net117),
    .B(\state[60] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2177_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0447_),
    .A2(_0778_),
    .Y(_0316_),
    .B1(net81));
 sg13g2_nand2_1 _2178_ (.Y(_0779_),
    .A(net120),
    .B(\state[61] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2179_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0451_),
    .A2(_0779_),
    .Y(_0317_),
    .B1(net82));
 sg13g2_nand2_1 _2180_ (.Y(_0780_),
    .A(net120),
    .B(\state[62] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2181_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0455_),
    .A2(_0780_),
    .Y(_0318_),
    .B1(net82));
 sg13g2_nand2_1 _2182_ (.Y(_0781_),
    .A(net120),
    .B(\state[63] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2183_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0459_),
    .A2(_0781_),
    .Y(_0319_),
    .B1(net82));
 sg13g2_nand2_1 _2184_ (.Y(_0782_),
    .A(net126),
    .B(\state[64] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2185_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0463_),
    .A2(_0782_),
    .Y(_0320_),
    .B1(net87));
 sg13g2_nand2_1 _2186_ (.Y(_0783_),
    .A(net126),
    .B(\state[65] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2187_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0467_),
    .A2(_0783_),
    .Y(_0321_),
    .B1(net87));
 sg13g2_nand2_1 _2188_ (.Y(_0784_),
    .A(net130),
    .B(\state[66] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2189_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0471_),
    .A2(_0784_),
    .Y(_0322_),
    .B1(net87));
 sg13g2_nand2_1 _2190_ (.Y(_0785_),
    .A(net129),
    .B(\state[67] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2191_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0475_),
    .A2(_0785_),
    .Y(_0323_),
    .B1(net85));
 sg13g2_nand2_1 _2192_ (.Y(_0786_),
    .A(net129),
    .B(\state[68] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2193_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0479_),
    .A2(_0786_),
    .Y(_0324_),
    .B1(net85));
 sg13g2_nand2_1 _2194_ (.Y(_0787_),
    .A(net129),
    .B(\state[69] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2195_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0483_),
    .A2(_0787_),
    .Y(_0325_),
    .B1(net85));
 sg13g2_nand2_1 _2196_ (.Y(_0788_),
    .A(net128),
    .B(\state[70] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2197_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0487_),
    .A2(_0788_),
    .Y(_0326_),
    .B1(net86));
 sg13g2_nand2_1 _2198_ (.Y(_0789_),
    .A(net129),
    .B(\state[71] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2199_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0491_),
    .A2(_0789_),
    .Y(_0327_),
    .B1(net86));
 sg13g2_nand2_1 _2200_ (.Y(_0790_),
    .A(net128),
    .B(\state[72] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2201_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0495_),
    .A2(_0790_),
    .Y(_0328_),
    .B1(net86));
 sg13g2_nand2_1 _2202_ (.Y(_0791_),
    .A(net128),
    .B(\state[73] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2203_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0499_),
    .A2(_0791_),
    .Y(_0329_),
    .B1(net86));
 sg13g2_nand2_1 _2204_ (.Y(_0792_),
    .A(net127),
    .B(\state[74] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2205_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0503_),
    .A2(_0792_),
    .Y(_0330_),
    .B1(net85));
 sg13g2_nand2_1 _2206_ (.Y(_0793_),
    .A(net130),
    .B(\state[75] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2207_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0507_),
    .A2(_0793_),
    .Y(_0331_),
    .B1(net85));
 sg13g2_nand2_1 _2208_ (.Y(_0794_),
    .A(net127),
    .B(\state[76] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2209_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0511_),
    .A2(_0794_),
    .Y(_0332_),
    .B1(net85));
 sg13g2_nand2_1 _2210_ (.Y(_0795_),
    .A(net127),
    .B(\state[77] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2211_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0515_),
    .A2(_0795_),
    .Y(_0333_),
    .B1(net85));
 sg13g2_nand2_1 _2212_ (.Y(_0796_),
    .A(net129),
    .B(\state[78] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2213_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0519_),
    .A2(_0796_),
    .Y(_0334_),
    .B1(net85));
 sg13g2_nand2_1 _2214_ (.Y(_0797_),
    .A(net130),
    .B(\state[79] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2215_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0523_),
    .A2(_0797_),
    .Y(_0335_),
    .B1(net87));
 sg13g2_nand2_1 _2216_ (.Y(_0798_),
    .A(net126),
    .B(\state[80] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2217_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0527_),
    .A2(_0798_),
    .Y(_0336_),
    .B1(net87));
 sg13g2_nand2_1 _2218_ (.Y(_0799_),
    .A(net122),
    .B(\state[81] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2219_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0531_),
    .A2(_0799_),
    .Y(_0337_),
    .B1(net84));
 sg13g2_nand2_1 _2220_ (.Y(_0800_),
    .A(net131),
    .B(\state[82] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2221_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0535_),
    .A2(_0800_),
    .Y(_0338_),
    .B1(net84));
 sg13g2_nand2_1 _2222_ (.Y(_0801_),
    .A(net122),
    .B(\state[83] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2223_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0539_),
    .A2(_0801_),
    .Y(_0339_),
    .B1(net84));
 sg13g2_nand2_1 _2224_ (.Y(_0802_),
    .A(net122),
    .B(\state[84] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2225_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0543_),
    .A2(_0802_),
    .Y(_0340_),
    .B1(net84));
 sg13g2_nand2_1 _2226_ (.Y(_0803_),
    .A(net122),
    .B(\state[85] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2227_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0547_),
    .A2(_0803_),
    .Y(_0341_),
    .B1(net84));
 sg13g2_nand2_1 _2228_ (.Y(_0804_),
    .A(net123),
    .B(\state[86] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2229_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0551_),
    .A2(_0804_),
    .Y(_0342_),
    .B1(net83));
 sg13g2_nand2_1 _2230_ (.Y(_0805_),
    .A(net124),
    .B(\state[87] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2231_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0555_),
    .A2(_0805_),
    .Y(_0343_),
    .B1(net83));
 sg13g2_nand2_1 _2232_ (.Y(_0806_),
    .A(net124),
    .B(\state[88] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2233_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0559_),
    .A2(_0806_),
    .Y(_0344_),
    .B1(net83));
 sg13g2_nand2_1 _2234_ (.Y(_0807_),
    .A(net124),
    .B(\state[89] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2235_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0563_),
    .A2(_0807_),
    .Y(_0345_),
    .B1(net88));
 sg13g2_nand2_1 _2236_ (.Y(_0808_),
    .A(net125),
    .B(\state[90] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2237_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0567_),
    .A2(_0808_),
    .Y(_0346_),
    .B1(net84));
 sg13g2_nand2_1 _2238_ (.Y(_0809_),
    .A(net125),
    .B(\state[91] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2239_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0571_),
    .A2(_0809_),
    .Y(_0347_),
    .B1(net84));
 sg13g2_nand2_1 _2240_ (.Y(_0810_),
    .A(net125),
    .B(\state[92] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2241_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0575_),
    .A2(_0810_),
    .Y(_0348_),
    .B1(net83));
 sg13g2_nand2_1 _2242_ (.Y(_0811_),
    .A(net125),
    .B(\state[93] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2243_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0579_),
    .A2(_0811_),
    .Y(_0349_),
    .B1(net83));
 sg13g2_nand2_1 _2244_ (.Y(_0812_),
    .A(net125),
    .B(\state[94] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2245_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0583_),
    .A2(_0812_),
    .Y(_0350_),
    .B1(net83));
 sg13g2_nand2_1 _2246_ (.Y(_0813_),
    .A(net107),
    .B(\state[95] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2247_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0587_),
    .A2(_0813_),
    .Y(_0351_),
    .B1(net74));
 sg13g2_nand2_1 _2248_ (.Y(_0814_),
    .A(net106),
    .B(\state[96] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2249_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0591_),
    .A2(_0814_),
    .Y(_0352_),
    .B1(net75));
 sg13g2_nand2_1 _2250_ (.Y(_0815_),
    .A(net106),
    .B(\state[97] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2251_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0595_),
    .A2(_0815_),
    .Y(_0353_),
    .B1(net75));
 sg13g2_nand2_1 _2252_ (.Y(_0816_),
    .A(net123),
    .B(\state[98] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2253_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0599_),
    .A2(_0816_),
    .Y(_0354_),
    .B1(net83));
 sg13g2_nand2_1 _2254_ (.Y(_0817_),
    .A(net123),
    .B(\state[99] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2255_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0603_),
    .A2(_0817_),
    .Y(_0355_),
    .B1(net83));
 sg13g2_nand2_1 _2256_ (.Y(_0818_),
    .A(net105),
    .B(\state[100] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2257_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0607_),
    .A2(_0818_),
    .Y(_0356_),
    .B1(net74));
 sg13g2_nand2_1 _2258_ (.Y(_0819_),
    .A(net105),
    .B(\state[101] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2259_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0611_),
    .A2(_0819_),
    .Y(_0357_),
    .B1(net74));
 sg13g2_nand2_1 _2260_ (.Y(_0820_),
    .A(net105),
    .B(\state[102] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2261_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0615_),
    .A2(_0820_),
    .Y(_0358_),
    .B1(net74));
 sg13g2_nand2_1 _2262_ (.Y(_0821_),
    .A(net108),
    .B(\state[103] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2263_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0619_),
    .A2(_0821_),
    .Y(_0359_),
    .B1(net74));
 sg13g2_nand2_1 _2264_ (.Y(_0822_),
    .A(net104),
    .B(\state[104] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2265_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0623_),
    .A2(_0822_),
    .Y(_0360_),
    .B1(net74));
 sg13g2_nand2_1 _2266_ (.Y(_0823_),
    .A(net104),
    .B(\state[105] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2267_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0627_),
    .A2(_0823_),
    .Y(_0361_),
    .B1(net74));
 sg13g2_nand2_1 _2268_ (.Y(_0824_),
    .A(net104),
    .B(\state[106] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2269_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0631_),
    .A2(_0824_),
    .Y(_0362_),
    .B1(net74));
 sg13g2_nand2_1 _2270_ (.Y(_0825_),
    .A(net106),
    .B(\state[107] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2271_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0635_),
    .A2(_0825_),
    .Y(_0363_),
    .B1(net75));
 sg13g2_nand2_1 _2272_ (.Y(_0826_),
    .A(net106),
    .B(\state[108] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2273_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0639_),
    .A2(_0826_),
    .Y(_0364_),
    .B1(net75));
 sg13g2_nand2_1 _2274_ (.Y(_0827_),
    .A(net107),
    .B(\state[109] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2275_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0643_),
    .A2(_0827_),
    .Y(_0365_),
    .B1(net75));
 sg13g2_nand2_1 _2276_ (.Y(_0828_),
    .A(net107),
    .B(\state[110] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2277_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0647_),
    .A2(_0828_),
    .Y(_0366_),
    .B1(net75));
 sg13g2_nand2_1 _2278_ (.Y(_0829_),
    .A(net105),
    .B(\state[111] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2279_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0651_),
    .A2(_0829_),
    .Y(_0367_),
    .B1(net76));
 sg13g2_nand2_1 _2280_ (.Y(_0830_),
    .A(net103),
    .B(\state[112] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2281_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0655_),
    .A2(_0830_),
    .Y(_0368_),
    .B1(net76));
 sg13g2_nand2_1 _2282_ (.Y(_0831_),
    .A(net103),
    .B(\state[113] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2283_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0659_),
    .A2(_0831_),
    .Y(_0369_),
    .B1(net76));
 sg13g2_nand2_1 _2284_ (.Y(_0832_),
    .A(net102),
    .B(\state[114] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2285_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0663_),
    .A2(_0832_),
    .Y(_0370_),
    .B1(net76));
 sg13g2_nand2_1 _2286_ (.Y(_0833_),
    .A(net102),
    .B(\state[115] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2287_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0667_),
    .A2(_0833_),
    .Y(_0371_),
    .B1(net76));
 sg13g2_nand2_1 _2288_ (.Y(_0834_),
    .A(net103),
    .B(\state[116] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2289_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0671_),
    .A2(_0834_),
    .Y(_0372_),
    .B1(net76));
 sg13g2_nand2_1 _2290_ (.Y(_0835_),
    .A(net103),
    .B(\state[117] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2291_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0675_),
    .A2(_0835_),
    .Y(_0373_),
    .B1(net76));
 sg13g2_nand2_1 _2292_ (.Y(_0836_),
    .A(net103),
    .B(\state[118] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2293_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0679_),
    .A2(_0836_),
    .Y(_0374_),
    .B1(net76));
 sg13g2_nand2_1 _2294_ (.Y(_0837_),
    .A(net93),
    .B(\state[119] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2295_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0683_),
    .A2(_0837_),
    .Y(_0375_),
    .B1(net69));
 sg13g2_nand2_1 _2296_ (.Y(_0838_),
    .A(net93),
    .B(\state[120] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2297_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0687_),
    .A2(_0838_),
    .Y(_0376_),
    .B1(net68));
 sg13g2_nand2_1 _2298_ (.Y(_0839_),
    .A(net90),
    .B(\state[121] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2299_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0691_),
    .A2(_0839_),
    .Y(_0377_),
    .B1(net68));
 sg13g2_nand2_1 _2300_ (.Y(_0840_),
    .A(net90),
    .B(\state[122] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2301_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0695_),
    .A2(_0840_),
    .Y(_0378_),
    .B1(net68));
 sg13g2_nand2_1 _2302_ (.Y(_0841_),
    .A(net90),
    .B(\state[123] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2303_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0699_),
    .A2(_0841_),
    .Y(_0379_),
    .B1(net68));
 sg13g2_nand2_1 _2304_ (.Y(_0842_),
    .A(net91),
    .B(\state[124] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2305_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0703_),
    .A2(_0842_),
    .Y(_0380_),
    .B1(net68));
 sg13g2_nand2_1 _2306_ (.Y(_0843_),
    .A(net91),
    .B(\state[125] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2307_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0707_),
    .A2(_0843_),
    .Y(_0381_),
    .B1(net68));
 sg13g2_nand2_1 _2308_ (.Y(_0844_),
    .A(net91),
    .B(\state[126] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2309_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0711_),
    .A2(_0844_),
    .Y(_0382_),
    .B1(net68));
 sg13g2_nand2_1 _2310_ (.Y(_0845_),
    .A(\state[127] ),
    .B(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2311_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0715_),
    .A2(_0845_),
    .Y(_0383_),
    .B1(net68));
 sg13g2_dfrbpq_1 _2312_ (.RESET_B(net326),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0128_),
    .Q(\daisychain[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2313_ (.RESET_B(net325),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0129_),
    .Q(\daisychain[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2314_ (.RESET_B(net323),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0130_),
    .Q(\daisychain[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2315_ (.RESET_B(net321),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0131_),
    .Q(\daisychain[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2316_ (.RESET_B(net319),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0132_),
    .Q(\daisychain[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2317_ (.RESET_B(net317),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0133_),
    .Q(\daisychain[5] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2318_ (.RESET_B(net315),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0134_),
    .Q(\daisychain[6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2319_ (.RESET_B(net313),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0135_),
    .Q(\daisychain[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2320_ (.RESET_B(net311),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0136_),
    .Q(\daisychain[8] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2321_ (.RESET_B(net309),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0137_),
    .Q(\daisychain[9] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2322_ (.RESET_B(net307),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0138_),
    .Q(\daisychain[10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2323_ (.RESET_B(net305),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0139_),
    .Q(\daisychain[11] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2324_ (.RESET_B(net303),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0140_),
    .Q(\daisychain[12] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2325_ (.RESET_B(net301),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0141_),
    .Q(\daisychain[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2326_ (.RESET_B(net299),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0142_),
    .Q(\daisychain[14] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2327_ (.RESET_B(net297),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0143_),
    .Q(\daisychain[15] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2328_ (.RESET_B(net295),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0144_),
    .Q(\daisychain[16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2329_ (.RESET_B(net293),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0145_),
    .Q(\daisychain[17] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2330_ (.RESET_B(net291),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0146_),
    .Q(\daisychain[18] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2331_ (.RESET_B(net289),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0147_),
    .Q(\daisychain[19] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2332_ (.RESET_B(net287),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0148_),
    .Q(\daisychain[20] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2333_ (.RESET_B(net285),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0149_),
    .Q(\daisychain[21] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2334_ (.RESET_B(net283),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0150_),
    .Q(\daisychain[22] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2335_ (.RESET_B(net281),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0151_),
    .Q(\daisychain[23] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2336_ (.RESET_B(net279),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0152_),
    .Q(\daisychain[24] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2337_ (.RESET_B(net277),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0153_),
    .Q(\daisychain[25] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2338_ (.RESET_B(net275),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0154_),
    .Q(\daisychain[26] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2339_ (.RESET_B(net273),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0155_),
    .Q(\daisychain[27] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2340_ (.RESET_B(net271),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0156_),
    .Q(\daisychain[28] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2341_ (.RESET_B(net269),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0157_),
    .Q(\daisychain[29] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2342_ (.RESET_B(net267),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0158_),
    .Q(\daisychain[30] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2343_ (.RESET_B(net265),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0159_),
    .Q(\daisychain[31] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2344_ (.RESET_B(net263),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0160_),
    .Q(\daisychain[32] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2345_ (.RESET_B(net261),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0161_),
    .Q(\daisychain[33] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2346_ (.RESET_B(net259),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0162_),
    .Q(\daisychain[34] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2347_ (.RESET_B(net257),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0163_),
    .Q(\daisychain[35] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2348_ (.RESET_B(net255),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0164_),
    .Q(\daisychain[36] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2349_ (.RESET_B(net253),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0165_),
    .Q(\daisychain[37] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2350_ (.RESET_B(net251),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0166_),
    .Q(\daisychain[38] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2351_ (.RESET_B(net249),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0167_),
    .Q(\daisychain[39] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2352_ (.RESET_B(net247),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0168_),
    .Q(\daisychain[40] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2353_ (.RESET_B(net245),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0169_),
    .Q(\daisychain[41] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2354_ (.RESET_B(net243),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0170_),
    .Q(\daisychain[42] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2355_ (.RESET_B(net241),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0171_),
    .Q(\daisychain[43] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2356_ (.RESET_B(net239),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0172_),
    .Q(\daisychain[44] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2357_ (.RESET_B(net237),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0173_),
    .Q(\daisychain[45] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2358_ (.RESET_B(net235),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0174_),
    .Q(\daisychain[46] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2359_ (.RESET_B(net233),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0175_),
    .Q(\daisychain[47] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2360_ (.RESET_B(net231),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0176_),
    .Q(\daisychain[48] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2361_ (.RESET_B(net229),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0177_),
    .Q(\daisychain[49] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2362_ (.RESET_B(net227),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0178_),
    .Q(\daisychain[50] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2363_ (.RESET_B(net225),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0179_),
    .Q(\daisychain[51] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2364_ (.RESET_B(net223),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0180_),
    .Q(\daisychain[52] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2365_ (.RESET_B(net221),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0181_),
    .Q(\daisychain[53] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2366_ (.RESET_B(net219),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0182_),
    .Q(\daisychain[54] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2367_ (.RESET_B(net217),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0183_),
    .Q(\daisychain[55] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2368_ (.RESET_B(net215),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0184_),
    .Q(\daisychain[56] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2369_ (.RESET_B(net213),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0185_),
    .Q(\daisychain[57] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2370_ (.RESET_B(net211),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0186_),
    .Q(\daisychain[58] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2371_ (.RESET_B(net209),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0187_),
    .Q(\daisychain[59] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2372_ (.RESET_B(net207),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0188_),
    .Q(\daisychain[60] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2373_ (.RESET_B(net205),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0189_),
    .Q(\daisychain[61] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2374_ (.RESET_B(net203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0190_),
    .Q(\daisychain[62] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2375_ (.RESET_B(net201),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0191_),
    .Q(\daisychain[63] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2376_ (.RESET_B(net455),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0192_),
    .Q(\daisychain[64] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2377_ (.RESET_B(net453),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0193_),
    .Q(\daisychain[65] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2378_ (.RESET_B(net451),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0194_),
    .Q(\daisychain[66] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2379_ (.RESET_B(net449),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0195_),
    .Q(\daisychain[67] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2380_ (.RESET_B(net447),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0196_),
    .Q(\daisychain[68] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2381_ (.RESET_B(net445),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0197_),
    .Q(\daisychain[69] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2382_ (.RESET_B(net443),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0198_),
    .Q(\daisychain[70] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2383_ (.RESET_B(net441),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0199_),
    .Q(\daisychain[71] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2384_ (.RESET_B(net439),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0200_),
    .Q(\daisychain[72] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2385_ (.RESET_B(net437),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0201_),
    .Q(\daisychain[73] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2386_ (.RESET_B(net435),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0202_),
    .Q(\daisychain[74] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2387_ (.RESET_B(net433),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0203_),
    .Q(\daisychain[75] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2388_ (.RESET_B(net431),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0204_),
    .Q(\daisychain[76] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2389_ (.RESET_B(net429),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0205_),
    .Q(\daisychain[77] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2390_ (.RESET_B(net427),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0206_),
    .Q(\daisychain[78] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2391_ (.RESET_B(net425),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0207_),
    .Q(\daisychain[79] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2392_ (.RESET_B(net423),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0208_),
    .Q(\daisychain[80] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2393_ (.RESET_B(net421),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0209_),
    .Q(\daisychain[81] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2394_ (.RESET_B(net419),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0210_),
    .Q(\daisychain[82] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2395_ (.RESET_B(net417),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0211_),
    .Q(\daisychain[83] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2396_ (.RESET_B(net415),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0212_),
    .Q(\daisychain[84] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2397_ (.RESET_B(net413),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0213_),
    .Q(\daisychain[85] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2398_ (.RESET_B(net411),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0214_),
    .Q(\daisychain[86] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2399_ (.RESET_B(net409),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0215_),
    .Q(\daisychain[87] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2400_ (.RESET_B(net407),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0216_),
    .Q(\daisychain[88] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2401_ (.RESET_B(net405),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0217_),
    .Q(\daisychain[89] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2402_ (.RESET_B(net403),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0218_),
    .Q(\daisychain[90] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2403_ (.RESET_B(net401),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0219_),
    .Q(\daisychain[91] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2404_ (.RESET_B(net399),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0220_),
    .Q(\daisychain[92] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2405_ (.RESET_B(net397),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0221_),
    .Q(\daisychain[93] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2406_ (.RESET_B(net395),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0222_),
    .Q(\daisychain[94] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2407_ (.RESET_B(net393),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0223_),
    .Q(\daisychain[95] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2408_ (.RESET_B(net391),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0224_),
    .Q(\daisychain[96] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2409_ (.RESET_B(net389),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0225_),
    .Q(\daisychain[97] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2410_ (.RESET_B(net387),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0226_),
    .Q(\daisychain[98] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2411_ (.RESET_B(net385),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0227_),
    .Q(\daisychain[99] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2412_ (.RESET_B(net383),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0228_),
    .Q(\daisychain[100] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2413_ (.RESET_B(net381),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0229_),
    .Q(\daisychain[101] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2414_ (.RESET_B(net379),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0230_),
    .Q(\daisychain[102] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2415_ (.RESET_B(net377),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0231_),
    .Q(\daisychain[103] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2416_ (.RESET_B(net375),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0232_),
    .Q(\daisychain[104] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2417_ (.RESET_B(net373),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0233_),
    .Q(\daisychain[105] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2418_ (.RESET_B(net371),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0234_),
    .Q(\daisychain[106] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2419_ (.RESET_B(net369),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0235_),
    .Q(\daisychain[107] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2420_ (.RESET_B(net367),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0236_),
    .Q(\daisychain[108] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2421_ (.RESET_B(net365),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0237_),
    .Q(\daisychain[109] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2422_ (.RESET_B(net363),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0238_),
    .Q(\daisychain[110] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2423_ (.RESET_B(net361),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0239_),
    .Q(\daisychain[111] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2424_ (.RESET_B(net359),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0240_),
    .Q(\daisychain[112] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2425_ (.RESET_B(net357),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0241_),
    .Q(\daisychain[113] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2426_ (.RESET_B(net355),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0242_),
    .Q(\daisychain[114] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2427_ (.RESET_B(net353),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0243_),
    .Q(\daisychain[115] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2428_ (.RESET_B(net351),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0244_),
    .Q(\daisychain[116] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2429_ (.RESET_B(net349),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0245_),
    .Q(\daisychain[117] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2430_ (.RESET_B(net347),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0246_),
    .Q(\daisychain[118] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2431_ (.RESET_B(net345),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0247_),
    .Q(\daisychain[119] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2432_ (.RESET_B(net343),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0248_),
    .Q(\daisychain[120] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2433_ (.RESET_B(net341),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0249_),
    .Q(\daisychain[121] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2434_ (.RESET_B(net339),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0250_),
    .Q(\daisychain[122] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2435_ (.RESET_B(net337),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0251_),
    .Q(\daisychain[123] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2436_ (.RESET_B(net335),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0252_),
    .Q(\daisychain[124] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2437_ (.RESET_B(net333),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0253_),
    .Q(\daisychain[125] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2438_ (.RESET_B(net331),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0254_),
    .Q(\daisychain[126] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2439_ (.RESET_B(net329),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0255_),
    .Q(\daisychain[127] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2440_ (.RESET_B(net327),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0256_),
    .Q(\state[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2441_ (.RESET_B(net324),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0257_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2442_ (.RESET_B(net320),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0258_),
    .Q(\state[2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2443_ (.RESET_B(net316),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0259_),
    .Q(\state[3] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2444_ (.RESET_B(net312),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0260_),
    .Q(\state[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2445_ (.RESET_B(net308),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0261_),
    .Q(\state[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2446_ (.RESET_B(net304),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0262_),
    .Q(\state[6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2447_ (.RESET_B(net300),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0263_),
    .Q(\state[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2448_ (.RESET_B(net296),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0264_),
    .Q(\state[8] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2449_ (.RESET_B(net292),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0265_),
    .Q(\state[9] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2450_ (.RESET_B(net288),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0266_),
    .Q(\state[10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2451_ (.RESET_B(net284),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0267_),
    .Q(\state[11] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2452_ (.RESET_B(net280),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0268_),
    .Q(\state[12] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2453_ (.RESET_B(net276),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0269_),
    .Q(\state[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2454_ (.RESET_B(net272),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0270_),
    .Q(\state[14] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2455_ (.RESET_B(net268),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0271_),
    .Q(\state[15] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2456_ (.RESET_B(net264),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0272_),
    .Q(\state[16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2457_ (.RESET_B(net260),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0273_),
    .Q(\state[17] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2458_ (.RESET_B(net256),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0274_),
    .Q(\state[18] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2459_ (.RESET_B(net252),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0275_),
    .Q(\state[19] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2460_ (.RESET_B(net248),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0276_),
    .Q(\state[20] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2461_ (.RESET_B(net244),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0277_),
    .Q(\state[21] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2462_ (.RESET_B(net240),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0278_),
    .Q(\state[22] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2463_ (.RESET_B(net236),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0279_),
    .Q(\state[23] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2464_ (.RESET_B(net232),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0280_),
    .Q(\state[24] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2465_ (.RESET_B(net228),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0281_),
    .Q(\state[25] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2466_ (.RESET_B(net224),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0282_),
    .Q(\state[26] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2467_ (.RESET_B(net220),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0283_),
    .Q(\state[27] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2468_ (.RESET_B(net216),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0284_),
    .Q(\state[28] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2469_ (.RESET_B(net212),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0285_),
    .Q(\state[29] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2470_ (.RESET_B(net208),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0286_),
    .Q(\state[30] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2471_ (.RESET_B(net204),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0287_),
    .Q(\state[31] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2472_ (.RESET_B(net),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0288_),
    .Q(\state[32] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2473_ (.RESET_B(net452),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0289_),
    .Q(\state[33] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2474_ (.RESET_B(net448),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0290_),
    .Q(\state[34] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2475_ (.RESET_B(net444),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0291_),
    .Q(\state[35] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2476_ (.RESET_B(net440),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0292_),
    .Q(\state[36] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2477_ (.RESET_B(net436),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0293_),
    .Q(\state[37] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2478_ (.RESET_B(net432),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0294_),
    .Q(\state[38] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2479_ (.RESET_B(net428),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0295_),
    .Q(\state[39] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2480_ (.RESET_B(net424),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0296_),
    .Q(\state[40] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2481_ (.RESET_B(net420),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0297_),
    .Q(\state[41] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2482_ (.RESET_B(net416),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0298_),
    .Q(\state[42] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2483_ (.RESET_B(net412),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0299_),
    .Q(\state[43] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2484_ (.RESET_B(net408),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0300_),
    .Q(\state[44] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2485_ (.RESET_B(net404),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0301_),
    .Q(\state[45] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2486_ (.RESET_B(net400),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0302_),
    .Q(\state[46] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2487_ (.RESET_B(net396),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0303_),
    .Q(\state[47] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2488_ (.RESET_B(net392),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0304_),
    .Q(\state[48] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2489_ (.RESET_B(net388),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0305_),
    .Q(\state[49] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2490_ (.RESET_B(net384),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0306_),
    .Q(\state[50] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2491_ (.RESET_B(net380),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0307_),
    .Q(\state[51] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2492_ (.RESET_B(net376),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0308_),
    .Q(\state[52] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2493_ (.RESET_B(net372),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0309_),
    .Q(\state[53] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2494_ (.RESET_B(net368),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0310_),
    .Q(\state[54] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2495_ (.RESET_B(net364),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0311_),
    .Q(\state[55] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2496_ (.RESET_B(net360),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0312_),
    .Q(\state[56] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2497_ (.RESET_B(net356),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0313_),
    .Q(\state[57] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2498_ (.RESET_B(net352),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0314_),
    .Q(\state[58] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2499_ (.RESET_B(net348),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0315_),
    .Q(\state[59] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2500_ (.RESET_B(net344),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0316_),
    .Q(\state[60] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2501_ (.RESET_B(net340),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0317_),
    .Q(\state[61] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2502_ (.RESET_B(net336),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0318_),
    .Q(\state[62] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2503_ (.RESET_B(net332),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0319_),
    .Q(\state[63] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2504_ (.RESET_B(net328),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0320_),
    .Q(\state[64] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2505_ (.RESET_B(net322),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0321_),
    .Q(\state[65] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2506_ (.RESET_B(net314),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0322_),
    .Q(\state[66] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2507_ (.RESET_B(net306),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0323_),
    .Q(\state[67] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2508_ (.RESET_B(net298),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0324_),
    .Q(\state[68] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2509_ (.RESET_B(net290),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0325_),
    .Q(\state[69] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2510_ (.RESET_B(net282),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0326_),
    .Q(\state[70] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2511_ (.RESET_B(net274),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0327_),
    .Q(\state[71] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2512_ (.RESET_B(net266),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0328_),
    .Q(\state[72] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2513_ (.RESET_B(net258),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0329_),
    .Q(\state[73] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2514_ (.RESET_B(net250),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0330_),
    .Q(\state[74] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2515_ (.RESET_B(net242),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0331_),
    .Q(\state[75] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2516_ (.RESET_B(net234),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0332_),
    .Q(\state[76] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2517_ (.RESET_B(net226),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0333_),
    .Q(\state[77] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2518_ (.RESET_B(net218),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0334_),
    .Q(\state[78] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2519_ (.RESET_B(net210),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0335_),
    .Q(\state[79] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2520_ (.RESET_B(net202),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0336_),
    .Q(\state[80] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2521_ (.RESET_B(net450),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0337_),
    .Q(\state[81] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2522_ (.RESET_B(net442),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0338_),
    .Q(\state[82] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2523_ (.RESET_B(net434),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0339_),
    .Q(\state[83] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2524_ (.RESET_B(net426),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0340_),
    .Q(\state[84] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2525_ (.RESET_B(net418),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0341_),
    .Q(\state[85] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2526_ (.RESET_B(net410),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0342_),
    .Q(\state[86] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2527_ (.RESET_B(net402),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0343_),
    .Q(\state[87] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2528_ (.RESET_B(net394),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0344_),
    .Q(\state[88] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2529_ (.RESET_B(net386),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0345_),
    .Q(\state[89] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2530_ (.RESET_B(net378),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0346_),
    .Q(\state[90] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2531_ (.RESET_B(net370),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0347_),
    .Q(\state[91] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2532_ (.RESET_B(net362),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0348_),
    .Q(\state[92] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2533_ (.RESET_B(net354),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0349_),
    .Q(\state[93] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2534_ (.RESET_B(net346),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0350_),
    .Q(\state[94] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2535_ (.RESET_B(net338),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0351_),
    .Q(\state[95] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2536_ (.RESET_B(net330),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0352_),
    .Q(\state[96] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2537_ (.RESET_B(net318),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0353_),
    .Q(\state[97] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2538_ (.RESET_B(net302),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0354_),
    .Q(\state[98] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2539_ (.RESET_B(net286),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0355_),
    .Q(\state[99] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2540_ (.RESET_B(net270),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0356_),
    .Q(\state[100] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2541_ (.RESET_B(net254),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0357_),
    .Q(\state[101] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2542_ (.RESET_B(net238),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0358_),
    .Q(\state[102] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2543_ (.RESET_B(net222),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0359_),
    .Q(\state[103] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2544_ (.RESET_B(net206),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0360_),
    .Q(\state[104] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2545_ (.RESET_B(net446),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0361_),
    .Q(\state[105] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2546_ (.RESET_B(net430),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0362_),
    .Q(\state[106] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2547_ (.RESET_B(net414),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0363_),
    .Q(\state[107] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2548_ (.RESET_B(net398),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0364_),
    .Q(\state[108] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2549_ (.RESET_B(net382),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0365_),
    .Q(\state[109] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2550_ (.RESET_B(net366),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0366_),
    .Q(\state[110] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2551_ (.RESET_B(net350),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0367_),
    .Q(\state[111] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2552_ (.RESET_B(net334),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0368_),
    .Q(\state[112] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2553_ (.RESET_B(net310),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0369_),
    .Q(\state[113] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2554_ (.RESET_B(net278),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0370_),
    .Q(\state[114] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2555_ (.RESET_B(net246),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0371_),
    .Q(\state[115] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2556_ (.RESET_B(net214),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0372_),
    .Q(\state[116] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2557_ (.RESET_B(net438),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0373_),
    .Q(\state[117] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2558_ (.RESET_B(net406),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0374_),
    .Q(\state[118] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2559_ (.RESET_B(net374),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0375_),
    .Q(\state[119] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2560_ (.RESET_B(net342),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0376_),
    .Q(\state[120] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2561_ (.RESET_B(net294),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0377_),
    .Q(\state[121] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2562_ (.RESET_B(net230),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0378_),
    .Q(\state[122] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2563_ (.RESET_B(net422),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0379_),
    .Q(\state[123] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2564_ (.RESET_B(net358),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0380_),
    .Q(\state[124] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2565_ (.RESET_B(net262),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0381_),
    .Q(\state[125] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2566_ (.RESET_B(net390),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0382_),
    .Q(\state[126] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2567_ (.RESET_B(net454),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0383_),
    .Q(\state[127] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_tiehi _2375__202 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net201));
 sg13g2_tiehi _2520__203 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net202));
 sg13g2_tiehi _2374__204 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net203));
 sg13g2_tiehi _2471__205 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net204));
 sg13g2_tiehi _2373__206 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net205));
 sg13g2_tiehi _2544__207 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net206));
 sg13g2_tiehi _2372__208 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net207));
 sg13g2_tiehi _2470__209 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net208));
 sg13g2_tiehi _2371__210 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net209));
 sg13g2_tiehi _2519__211 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net210));
 sg13g2_tiehi _2370__212 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net211));
 sg13g2_tiehi _2469__213 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net212));
 sg13g2_tiehi _2369__214 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net213));
 sg13g2_tiehi _2556__215 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net214));
 sg13g2_tiehi _2368__216 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net215));
 sg13g2_tiehi _2468__217 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net216));
 sg13g2_tiehi _2367__218 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net217));
 sg13g2_tiehi _2518__219 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net218));
 sg13g2_tiehi _2366__220 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net219));
 sg13g2_tiehi _2467__221 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net220));
 sg13g2_tiehi _2365__222 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net221));
 sg13g2_tiehi _2543__223 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net222));
 sg13g2_tiehi _2364__224 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net223));
 sg13g2_tiehi _2466__225 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net224));
 sg13g2_tiehi _2363__226 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net225));
 sg13g2_tiehi _2517__227 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net226));
 sg13g2_tiehi _2362__228 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net227));
 sg13g2_tiehi _2465__229 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net228));
 sg13g2_tiehi _2361__230 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net229));
 sg13g2_tiehi _2562__231 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net230));
 sg13g2_tiehi _2360__232 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net231));
 sg13g2_tiehi _2464__233 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net232));
 sg13g2_tiehi _2359__234 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net233));
 sg13g2_tiehi _2516__235 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net234));
 sg13g2_tiehi _2358__236 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net235));
 sg13g2_tiehi _2463__237 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net236));
 sg13g2_tiehi _2357__238 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net237));
 sg13g2_tiehi _2542__239 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net238));
 sg13g2_tiehi _2356__240 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net239));
 sg13g2_tiehi _2462__241 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net240));
 sg13g2_tiehi _2355__242 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net241));
 sg13g2_tiehi _2515__243 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net242));
 sg13g2_tiehi _2354__244 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net243));
 sg13g2_tiehi _2461__245 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net244));
 sg13g2_tiehi _2353__246 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net245));
 sg13g2_tiehi _2555__247 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net246));
 sg13g2_tiehi _2352__248 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net247));
 sg13g2_tiehi _2460__249 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net248));
 sg13g2_tiehi _2351__250 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net249));
 sg13g2_tiehi _2514__251 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net250));
 sg13g2_tiehi _2350__252 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net251));
 sg13g2_tiehi _2459__253 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net252));
 sg13g2_tiehi _2349__254 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net253));
 sg13g2_tiehi _2541__255 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net254));
 sg13g2_tiehi _2348__256 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net255));
 sg13g2_tiehi _2458__257 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net256));
 sg13g2_tiehi _2347__258 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net257));
 sg13g2_tiehi _2513__259 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net258));
 sg13g2_tiehi _2346__260 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net259));
 sg13g2_tiehi _2457__261 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net260));
 sg13g2_tiehi _2345__262 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net261));
 sg13g2_tiehi _2565__263 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net262));
 sg13g2_tiehi _2344__264 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net263));
 sg13g2_tiehi _2456__265 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net264));
 sg13g2_tiehi _2343__266 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net265));
 sg13g2_tiehi _2512__267 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net266));
 sg13g2_tiehi _2342__268 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net267));
 sg13g2_tiehi _2455__269 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net268));
 sg13g2_tiehi _2341__270 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net269));
 sg13g2_tiehi _2540__271 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net270));
 sg13g2_tiehi _2340__272 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net271));
 sg13g2_tiehi _2454__273 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net272));
 sg13g2_tiehi _2339__274 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net273));
 sg13g2_tiehi _2511__275 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net274));
 sg13g2_tiehi _2338__276 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net275));
 sg13g2_tiehi _2453__277 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net276));
 sg13g2_tiehi _2337__278 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net277));
 sg13g2_tiehi _2554__279 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net278));
 sg13g2_tiehi _2336__280 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net279));
 sg13g2_tiehi _2452__281 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net280));
 sg13g2_tiehi _2335__282 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net281));
 sg13g2_tiehi _2510__283 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net282));
 sg13g2_tiehi _2334__284 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net283));
 sg13g2_tiehi _2451__285 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net284));
 sg13g2_tiehi _2333__286 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net285));
 sg13g2_tiehi _2539__287 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net286));
 sg13g2_tiehi _2332__288 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net287));
 sg13g2_tiehi _2450__289 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net288));
 sg13g2_tiehi _2331__290 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net289));
 sg13g2_tiehi _2509__291 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net290));
 sg13g2_tiehi _2330__292 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net291));
 sg13g2_tiehi _2449__293 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net292));
 sg13g2_tiehi _2329__294 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net293));
 sg13g2_tiehi _2561__295 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net294));
 sg13g2_tiehi _2328__296 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net295));
 sg13g2_tiehi _2448__297 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net296));
 sg13g2_tiehi _2327__298 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net297));
 sg13g2_tiehi _2508__299 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net298));
 sg13g2_tiehi _2326__300 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net299));
 sg13g2_tiehi _2447__301 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net300));
 sg13g2_tiehi _2325__302 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net301));
 sg13g2_tiehi _2538__303 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net302));
 sg13g2_tiehi _2324__304 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net303));
 sg13g2_tiehi _2446__305 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net304));
 sg13g2_tiehi _2323__306 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net305));
 sg13g2_tiehi _2507__307 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net306));
 sg13g2_tiehi _2322__308 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net307));
 sg13g2_tiehi _2445__309 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net308));
 sg13g2_tiehi _2321__310 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net309));
 sg13g2_tiehi _2553__311 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net310));
 sg13g2_tiehi _2320__312 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net311));
 sg13g2_tiehi _2444__313 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net312));
 sg13g2_tiehi _2319__314 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net313));
 sg13g2_tiehi _2506__315 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net314));
 sg13g2_tiehi _2318__316 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net315));
 sg13g2_tiehi _2443__317 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net316));
 sg13g2_tiehi _2317__318 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net317));
 sg13g2_tiehi _2537__319 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net318));
 sg13g2_tiehi _2316__320 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net319));
 sg13g2_tiehi _2442__321 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net320));
 sg13g2_tiehi _2315__322 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net321));
 sg13g2_tiehi _2505__323 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net322));
 sg13g2_tiehi _2314__324 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net323));
 sg13g2_tiehi _2441__325 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net324));
 sg13g2_tiehi _2313__326 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net325));
 sg13g2_tiehi _2312__327 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net326));
 sg13g2_tiehi _2440__328 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net327));
 sg13g2_tiehi _2504__329 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net328));
 sg13g2_tiehi _2439__330 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net329));
 sg13g2_tiehi _2536__331 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net330));
 sg13g2_tiehi _2438__332 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net331));
 sg13g2_tiehi _2503__333 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net332));
 sg13g2_tiehi _2437__334 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net333));
 sg13g2_tiehi _2552__335 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net334));
 sg13g2_tiehi _2436__336 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net335));
 sg13g2_tiehi _2502__337 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net336));
 sg13g2_tiehi _2435__338 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net337));
 sg13g2_tiehi _2535__339 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net338));
 sg13g2_tiehi _2434__340 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net339));
 sg13g2_tiehi _2501__341 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net340));
 sg13g2_tiehi _2433__342 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net341));
 sg13g2_tiehi _2560__343 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net342));
 sg13g2_tiehi _2432__344 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net343));
 sg13g2_tiehi _2500__345 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net344));
 sg13g2_tiehi _2431__346 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net345));
 sg13g2_tiehi _2534__347 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net346));
 sg13g2_tiehi _2430__348 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net347));
 sg13g2_tiehi _2499__349 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net348));
 sg13g2_tiehi _2429__350 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net349));
 sg13g2_tiehi _2551__351 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net350));
 sg13g2_tiehi _2428__352 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net351));
 sg13g2_tiehi _2498__353 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net352));
 sg13g2_tiehi _2427__354 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net353));
 sg13g2_tiehi _2533__355 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net354));
 sg13g2_tiehi _2426__356 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net355));
 sg13g2_tiehi _2497__357 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net356));
 sg13g2_tiehi _2425__358 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net357));
 sg13g2_tiehi _2564__359 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net358));
 sg13g2_tiehi _2424__360 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net359));
 sg13g2_tiehi _2496__361 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net360));
 sg13g2_tiehi _2423__362 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net361));
 sg13g2_tiehi _2532__363 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net362));
 sg13g2_tiehi _2422__364 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net363));
 sg13g2_tiehi _2495__365 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net364));
 sg13g2_tiehi _2421__366 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net365));
 sg13g2_tiehi _2550__367 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net366));
 sg13g2_tiehi _2420__368 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net367));
 sg13g2_tiehi _2494__369 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net368));
 sg13g2_tiehi _2419__370 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net369));
 sg13g2_tiehi _2531__371 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net370));
 sg13g2_tiehi _2418__372 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net371));
 sg13g2_tiehi _2493__373 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net372));
 sg13g2_tiehi _2417__374 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net373));
 sg13g2_tiehi _2559__375 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net374));
 sg13g2_tiehi _2416__376 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net375));
 sg13g2_tiehi _2492__377 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net376));
 sg13g2_tiehi _2415__378 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net377));
 sg13g2_tiehi _2530__379 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net378));
 sg13g2_tiehi _2414__380 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net379));
 sg13g2_tiehi _2491__381 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net380));
 sg13g2_tiehi _2413__382 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net381));
 sg13g2_tiehi _2549__383 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net382));
 sg13g2_tiehi _2412__384 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net383));
 sg13g2_tiehi _2490__385 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net384));
 sg13g2_tiehi _2411__386 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net385));
 sg13g2_tiehi _2529__387 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net386));
 sg13g2_tiehi _2410__388 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net387));
 sg13g2_tiehi _2489__389 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net388));
 sg13g2_tiehi _2409__390 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net389));
 sg13g2_tiehi _2566__391 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net390));
 sg13g2_tiehi _2408__392 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net391));
 sg13g2_tiehi _2488__393 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net392));
 sg13g2_tiehi _2407__394 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net393));
 sg13g2_tiehi _2528__395 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net394));
 sg13g2_tiehi _2406__396 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net395));
 sg13g2_tiehi _2487__397 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net396));
 sg13g2_tiehi _2405__398 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net397));
 sg13g2_tiehi _2548__399 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net398));
 sg13g2_tiehi _2404__400 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net399));
 sg13g2_tiehi _2486__401 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net400));
 sg13g2_tiehi _2403__402 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net401));
 sg13g2_tiehi _2527__403 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net402));
 sg13g2_tiehi _2402__404 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net403));
 sg13g2_tiehi _2485__405 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net404));
 sg13g2_tiehi _2401__406 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net405));
 sg13g2_tiehi _2558__407 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net406));
 sg13g2_tiehi _2400__408 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net407));
 sg13g2_tiehi _2484__409 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net408));
 sg13g2_tiehi _2399__410 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net409));
 sg13g2_tiehi _2526__411 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net410));
 sg13g2_tiehi _2398__412 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net411));
 sg13g2_tiehi _2483__413 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net412));
 sg13g2_tiehi _2397__414 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net413));
 sg13g2_tiehi _2547__415 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net414));
 sg13g2_tiehi _2396__416 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net415));
 sg13g2_tiehi _2482__417 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net416));
 sg13g2_tiehi _2395__418 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net417));
 sg13g2_tiehi _2525__419 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net418));
 sg13g2_tiehi _2394__420 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net419));
 sg13g2_tiehi _2481__421 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net420));
 sg13g2_tiehi _2393__422 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net421));
 sg13g2_tiehi _2563__423 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net422));
 sg13g2_tiehi _2392__424 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net423));
 sg13g2_tiehi _2480__425 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net424));
 sg13g2_tiehi _2391__426 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net425));
 sg13g2_tiehi _2524__427 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net426));
 sg13g2_tiehi _2390__428 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net427));
 sg13g2_tiehi _2479__429 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net428));
 sg13g2_tiehi _2389__430 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net429));
 sg13g2_tiehi _2546__431 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net430));
 sg13g2_tiehi _2388__432 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net431));
 sg13g2_tiehi _2478__433 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net432));
 sg13g2_tiehi _2387__434 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net433));
 sg13g2_tiehi _2523__435 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net434));
 sg13g2_tiehi _2386__436 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net435));
 sg13g2_tiehi _2477__437 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net436));
 sg13g2_tiehi _2385__438 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net437));
 sg13g2_tiehi _2557__439 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net438));
 sg13g2_tiehi _2384__440 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net439));
 sg13g2_tiehi _2476__441 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net440));
 sg13g2_tiehi _2383__442 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net441));
 sg13g2_tiehi _2522__443 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net442));
 sg13g2_tiehi _2382__444 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net443));
 sg13g2_tiehi _2475__445 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net444));
 sg13g2_tiehi _2381__446 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net445));
 sg13g2_tiehi _2545__447 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net446));
 sg13g2_tiehi _2380__448 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net447));
 sg13g2_tiehi _2474__449 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net448));
 sg13g2_tiehi _2379__450 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net449));
 sg13g2_tiehi _2521__451 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net450));
 sg13g2_tiehi _2378__452 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net451));
 sg13g2_tiehi _2473__453 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net452));
 sg13g2_tiehi _2377__454 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net453));
 sg13g2_tiehi _2567__455 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net454));
 sg13g2_tiehi _2376__456 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net455));
 sg13g2_tiehi heichips25_pudding (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net456));
 sg13g2_tiehi heichips25_pudding_457 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net457));
 sg13g2_tiehi heichips25_pudding_458 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net458));
 sg13g2_tiehi heichips25_pudding_459 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net459));
 sg13g2_tiehi heichips25_pudding_460 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net460));
 sg13g2_tiehi heichips25_pudding_461 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net461));
 sg13g2_tiehi heichips25_pudding_462 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net462));
 sg13g2_tiehi heichips25_pudding_463 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net463));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2832_ (.A(\state[120] ),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2833_ (.A(\state[121] ),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2834_ (.A(\state[122] ),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2835_ (.A(\state[123] ),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2836_ (.A(\state[124] ),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2837_ (.A(\state[125] ),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2838_ (.A(\state[126] ),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2839_ (.A(\state[127] ),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2840_ (.A(\daisychain[120] ),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2841_ (.A(\daisychain[121] ),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2842_ (.A(\daisychain[122] ),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2843_ (.A(\daisychain[123] ),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2844_ (.A(\daisychain[124] ),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2845_ (.A(\daisychain[125] ),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2846_ (.A(\daisychain[126] ),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _2847_ (.A(\daisychain[127] ),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 dac128module dac (.IOUT(i_out),
    .VSS(VGND),
    .VDD(VPWR),
    .EN({\digitalen.g[3].u.OUTP ,
    \digitalen.g[2].u.OUTP ,
    \digitalen.g[1].u.OUTP ,
    \digitalen.g[0].u.OUTP }),
    .ENB({\digitalen.g[3].u.OUTN ,
    \digitalen.g[2].u.OUTN ,
    \digitalen.g[1].u.OUTN ,
    \digitalen.g[0].u.OUTN }),
    .ON({\state[127] ,
    \state[126] ,
    \state[125] ,
    \state[124] ,
    \state[123] ,
    \state[122] ,
    \state[121] ,
    \state[120] ,
    \state[119] ,
    \state[118] ,
    \state[117] ,
    \state[116] ,
    \state[115] ,
    \state[114] ,
    \state[113] ,
    \state[112] ,
    \state[111] ,
    \state[110] ,
    \state[109] ,
    \state[108] ,
    \state[107] ,
    \state[106] ,
    \state[105] ,
    \state[104] ,
    \state[103] ,
    \state[102] ,
    \state[101] ,
    \state[100] ,
    \state[99] ,
    \state[98] ,
    \state[97] ,
    \state[96] ,
    \state[95] ,
    \state[94] ,
    \state[93] ,
    \state[92] ,
    \state[91] ,
    \state[90] ,
    \state[89] ,
    \state[88] ,
    \state[87] ,
    \state[86] ,
    \state[85] ,
    \state[84] ,
    \state[83] ,
    \state[82] ,
    \state[81] ,
    \state[80] ,
    \state[79] ,
    \state[78] ,
    \state[77] ,
    \state[76] ,
    \state[75] ,
    \state[74] ,
    \state[73] ,
    \state[72] ,
    \state[71] ,
    \state[70] ,
    \state[69] ,
    \state[68] ,
    \state[67] ,
    \state[66] ,
    \state[65] ,
    \state[64] ,
    \state[63] ,
    \state[62] ,
    \state[61] ,
    \state[60] ,
    \state[59] ,
    \state[58] ,
    \state[57] ,
    \state[56] ,
    \state[55] ,
    \state[54] ,
    \state[53] ,
    \state[52] ,
    \state[51] ,
    \state[50] ,
    \state[49] ,
    \state[48] ,
    \state[47] ,
    \state[46] ,
    \state[45] ,
    \state[44] ,
    \state[43] ,
    \state[42] ,
    \state[41] ,
    \state[40] ,
    \state[39] ,
    \state[38] ,
    \state[37] ,
    \state[36] ,
    \state[35] ,
    \state[34] ,
    \state[33] ,
    \state[32] ,
    \state[31] ,
    \state[30] ,
    \state[29] ,
    \state[28] ,
    \state[27] ,
    \state[26] ,
    \state[25] ,
    \state[24] ,
    \state[23] ,
    \state[22] ,
    \state[21] ,
    \state[20] ,
    \state[19] ,
    \state[18] ,
    \state[17] ,
    \state[16] ,
    \state[15] ,
    \state[14] ,
    \state[13] ,
    \state[12] ,
    \state[11] ,
    \state[10] ,
    \state[9] ,
    \state[8] ,
    \state[7] ,
    \state[6] ,
    \state[5] ,
    \state[4] ,
    \state[3] ,
    \state[2] ,
    \state[1] ,
    \state[0] }),
    .ONB({_0030_,
    _0029_,
    _0028_,
    _0027_,
    _0026_,
    _0025_,
    _0024_,
    _0023_,
    _0021_,
    _0020_,
    _0019_,
    _0018_,
    _0017_,
    _0016_,
    _0015_,
    _0014_,
    _0013_,
    _0012_,
    _0010_,
    _0009_,
    _0008_,
    _0007_,
    _0006_,
    _0005_,
    _0004_,
    _0003_,
    _0002_,
    _0001_,
    _0126_,
    _0125_,
    _0124_,
    _0123_,
    _0122_,
    _0121_,
    _0120_,
    _0119_,
    _0118_,
    _0117_,
    _0115_,
    _0114_,
    _0113_,
    _0112_,
    _0111_,
    _0110_,
    _0109_,
    _0108_,
    _0107_,
    _0106_,
    _0104_,
    _0103_,
    _0102_,
    _0101_,
    _0100_,
    _0099_,
    _0098_,
    _0097_,
    _0096_,
    _0095_,
    _0093_,
    _0092_,
    _0091_,
    _0090_,
    _0089_,
    _0088_,
    _0087_,
    _0086_,
    _0085_,
    _0084_,
    _0082_,
    _0081_,
    _0080_,
    _0079_,
    _0078_,
    _0077_,
    _0076_,
    _0075_,
    _0074_,
    _0073_,
    _0071_,
    _0070_,
    _0069_,
    _0068_,
    _0067_,
    _0066_,
    _0065_,
    _0064_,
    _0063_,
    _0062_,
    _0060_,
    _0059_,
    _0058_,
    _0057_,
    _0056_,
    _0055_,
    _0054_,
    _0053_,
    _0052_,
    _0051_,
    _0049_,
    _0048_,
    _0047_,
    _0046_,
    _0045_,
    _0044_,
    _0043_,
    _0042_,
    _0041_,
    _0040_,
    _0038_,
    _0037_,
    _0036_,
    _0035_,
    _0034_,
    _0033_,
    _0032_,
    _0031_,
    _0022_,
    _0011_,
    _0127_,
    _0116_,
    _0105_,
    _0094_,
    _0083_,
    _0072_,
    _0061_,
    _0050_,
    _0039_,
    _0000_}),
    .VbiasP({\bias[1] ,
    \bias[0] }),
    .VcascP({i_in,
    i_in}));
 sg13g2_inv_1 \digitalen.g[0].u.inv1  (.VDD(VPWR),
    .Y(\digitalen.g[0].u.OUTN ),
    .A(net6),
    .VSS(VGND));
 sg13g2_inv_1 \digitalen.g[0].u.inv2  (.VDD(VPWR),
    .Y(\digitalen.g[0].u.OUTP ),
    .A(\digitalen.g[0].u.OUTN ),
    .VSS(VGND));
 sg13g2_inv_1 \digitalen.g[1].u.inv1  (.VDD(VPWR),
    .Y(\digitalen.g[1].u.OUTN ),
    .A(net6),
    .VSS(VGND));
 sg13g2_inv_1 \digitalen.g[1].u.inv2  (.VDD(VPWR),
    .Y(\digitalen.g[1].u.OUTP ),
    .A(\digitalen.g[1].u.OUTN ),
    .VSS(VGND));
 sg13g2_inv_1 \digitalen.g[2].u.inv1  (.VDD(VPWR),
    .Y(\digitalen.g[2].u.OUTN ),
    .A(net6),
    .VSS(VGND));
 sg13g2_inv_1 \digitalen.g[2].u.inv2  (.VDD(VPWR),
    .Y(\digitalen.g[2].u.OUTP ),
    .A(\digitalen.g[2].u.OUTN ),
    .VSS(VGND));
 sg13g2_inv_1 \digitalen.g[3].u.inv1  (.VDD(VPWR),
    .Y(\digitalen.g[3].u.OUTN ),
    .A(net6),
    .VSS(VGND));
 sg13g2_inv_1 \digitalen.g[3].u.inv2  (.VDD(VPWR),
    .Y(\digitalen.g[3].u.OUTP ),
    .A(\digitalen.g[3].u.OUTN ),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout23 (.A(net45),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout24 (.A(net45),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout25 (.A(net28),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout26 (.A(net27),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout27 (.A(net28),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout28 (.A(net45),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout29 (.A(net32),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout30 (.A(net32),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout31 (.A(net32),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout32 (.A(net45),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout33 (.A(net34),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout34 (.A(net44),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout35 (.A(net37),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout36 (.A(net37),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout37 (.A(net44),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout38 (.A(net40),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout39 (.A(net40),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout40 (.A(net44),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout41 (.A(net43),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout42 (.A(net43),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout43 (.A(net44),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout44 (.A(net45),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout45 (.A(_0851_),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout46 (.A(net67),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout47 (.A(net50),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout48 (.A(net49),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout49 (.A(net50),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout50 (.A(net67),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout51 (.A(net54),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout52 (.A(net54),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout53 (.A(net54),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout54 (.A(net67),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout55 (.A(net57),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout56 (.A(net57),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout57 (.A(net66),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout58 (.A(net60),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout59 (.A(net60),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout60 (.A(net66),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout61 (.A(net62),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout62 (.A(net66),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout63 (.A(net65),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout64 (.A(net65),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout65 (.A(net66),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout66 (.A(net67),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout67 (.A(_0850_),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout68 (.A(net89),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout69 (.A(net89),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout70 (.A(net73),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout71 (.A(net73),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout72 (.A(net73),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout73 (.A(net77),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout74 (.A(net77),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout75 (.A(net77),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout76 (.A(net77),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout77 (.A(net89),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout78 (.A(net79),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout79 (.A(net88),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout80 (.A(net82),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout81 (.A(net82),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout82 (.A(net88),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout83 (.A(net84),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout84 (.A(net88),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout85 (.A(net87),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout86 (.A(net87),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout87 (.A(net88),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout88 (.A(net89),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout89 (.A(_0847_),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout90 (.A(net91),
    .X(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout91 (.A(net93),
    .X(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout92 (.A(net93),
    .X(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout93 (.A(net132),
    .X(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout94 (.A(net96),
    .X(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout95 (.A(net96),
    .X(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout96 (.A(net109),
    .X(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout97 (.A(net98),
    .X(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout98 (.A(net101),
    .X(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout99 (.A(net100),
    .X(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout100 (.A(net101),
    .X(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout101 (.A(net109),
    .X(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout102 (.A(net103),
    .X(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout103 (.A(net108),
    .X(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout104 (.A(net105),
    .X(net104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout105 (.A(net108),
    .X(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout106 (.A(net107),
    .X(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout107 (.A(net108),
    .X(net107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout108 (.A(net109),
    .X(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout109 (.A(net132),
    .X(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout110 (.A(net112),
    .X(net110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout111 (.A(net112),
    .X(net111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout112 (.A(net114),
    .X(net112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout113 (.A(net114),
    .X(net113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout114 (.A(net121),
    .X(net114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout115 (.A(net118),
    .X(net115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout116 (.A(net118),
    .X(net116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout117 (.A(net118),
    .X(net117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout118 (.A(net121),
    .X(net118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout119 (.A(net121),
    .X(net119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout120 (.A(net121),
    .X(net120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout121 (.A(net132),
    .X(net121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout122 (.A(net131),
    .X(net122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout123 (.A(net125),
    .X(net123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout124 (.A(net125),
    .X(net124),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout125 (.A(net131),
    .X(net125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout126 (.A(net130),
    .X(net126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout127 (.A(net130),
    .X(net127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout128 (.A(net129),
    .X(net128),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout129 (.A(net130),
    .X(net129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout130 (.A(net131),
    .X(net130),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout131 (.A(net132),
    .X(net131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout132 (.A(_0846_),
    .X(net132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout133 (.A(net155),
    .X(net133),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout134 (.A(net155),
    .X(net134),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout135 (.A(net138),
    .X(net135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout136 (.A(net137),
    .X(net136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout137 (.A(net138),
    .X(net137),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout138 (.A(net142),
    .X(net138),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout139 (.A(net142),
    .X(net139),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout140 (.A(net142),
    .X(net140),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout141 (.A(net142),
    .X(net141),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout142 (.A(net155),
    .X(net142),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout143 (.A(net144),
    .X(net143),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout144 (.A(net154),
    .X(net144),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout145 (.A(net147),
    .X(net145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout146 (.A(net147),
    .X(net146),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout147 (.A(net154),
    .X(net147),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout148 (.A(net150),
    .X(net148),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout149 (.A(net150),
    .X(net149),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout150 (.A(net154),
    .X(net150),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout151 (.A(net153),
    .X(net151),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout152 (.A(net153),
    .X(net152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout153 (.A(net154),
    .X(net153),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout154 (.A(net155),
    .X(net154),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout155 (.A(net5),
    .X(net155),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout156 (.A(net157),
    .X(net156),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout157 (.A(net177),
    .X(net157),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout158 (.A(net161),
    .X(net158),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout159 (.A(net160),
    .X(net159),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout160 (.A(net161),
    .X(net160),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout161 (.A(net177),
    .X(net161),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout162 (.A(net163),
    .X(net162),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout163 (.A(net164),
    .X(net163),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout164 (.A(net177),
    .X(net164),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout165 (.A(net166),
    .X(net165),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout166 (.A(net176),
    .X(net166),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout167 (.A(net169),
    .X(net167),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout168 (.A(net169),
    .X(net168),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout169 (.A(net176),
    .X(net169),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout170 (.A(net172),
    .X(net170),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout171 (.A(net172),
    .X(net171),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout172 (.A(net176),
    .X(net172),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout173 (.A(net175),
    .X(net173),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout174 (.A(net175),
    .X(net174),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout175 (.A(net176),
    .X(net175),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout176 (.A(net177),
    .X(net176),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout177 (.A(net4),
    .X(net177),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout178 (.A(net179),
    .X(net178),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout179 (.A(net200),
    .X(net179),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout180 (.A(net183),
    .X(net180),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout181 (.A(net182),
    .X(net181),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout182 (.A(net183),
    .X(net182),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout183 (.A(net200),
    .X(net183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout184 (.A(net187),
    .X(net184),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout185 (.A(net187),
    .X(net185),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout186 (.A(net187),
    .X(net186),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout187 (.A(net200),
    .X(net187),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout188 (.A(net189),
    .X(net188),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout189 (.A(net199),
    .X(net189),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout190 (.A(net192),
    .X(net190),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout191 (.A(net192),
    .X(net191),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout192 (.A(net199),
    .X(net192),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout193 (.A(net195),
    .X(net193),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout194 (.A(net195),
    .X(net194),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout195 (.A(net199),
    .X(net195),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout196 (.A(net198),
    .X(net196),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout197 (.A(net198),
    .X(net197),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout198 (.A(net199),
    .X(net198),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout199 (.A(net200),
    .X(net199),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout200 (.A(net1),
    .X(net200),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi _2472__201 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_14_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_16 clkbuf_2_0__f_clk (.X(clknet_2_0__leaf_clk),
    .A(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_16 clkbuf_2_1__f_clk (.X(clknet_2_1__leaf_clk),
    .A(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_16 clkbuf_2_2__f_clk (.X(clknet_2_2__leaf_clk),
    .A(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_16 clkbuf_2_3__f_clk (.X(clknet_2_3__leaf_clk),
    .A(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload0 (.A(clknet_2_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload1 (.A(clknet_2_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload2 (.A(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload3 (.A(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload5 (.A(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload7 (.A(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload11 (.VDD(VPWR),
    .A(clknet_leaf_12_clk),
    .VSS(VGND));
 sg13g2_buf_8 clkload12 (.A(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net456;
 assign uio_oe[1] = net457;
 assign uio_oe[2] = net458;
 assign uio_oe[3] = net459;
 assign uio_oe[4] = net460;
 assign uio_oe[5] = net461;
 assign uio_oe[6] = net462;
 assign uio_oe[7] = net463;
endmodule
