// SPDX-FileCopyrightText: © 2025 XXX Authors
// SPDX-License-Identifier: Apache-2.0

// Adapted from the Tiny Tapeout template

`default_nettype none

module heichips25_template (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    // List all unused inputs to prevent warnings
    wire _unused = &{ena, ui_in[7:1], uio_in[7:0]};

    logic [7:0] count;
    logic dir_up = 1;
    
	reg [255:0] thermo;

    always_ff @(posedge clk) begin
        if (!rst_n) begin
            count <= '0;
        end else begin
            if (ui_in[0]) begin
                if (dir_up) begin 
                	count <= count + 1;
                	if (count == 254) begin
                		dir_up <= 0;
                	end
                end else begin
                	count <= count - 1;
                	if (count == 1) begin
                		dir_up <= 1;
                	end
                end                
            end
        end
    end
    
	thermometer_encoder #(
		.IN_WIDTH (8),
		.OUT_WIDTH (256))
	te_inst(
		.din (count),
		.thermo (thermo)
	);
    
    assign uo_out  = thermo[7:0];
    assign uio_out = thermo[15:8];
    assign uio_oe  = thermo[23:16];

endmodule
