module non_overlap (VPWR,
    VGND,
    ON,
    ON_N,
    thermo);
 inout VPWR;
 inout VGND;
 output [31:0] ON;
 output [31:0] ON_N;
 input [31:0] thermo;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire \comb_logic[0].delayed[0] ;
 wire \comb_logic[0].pulse_out_n ;
 wire \comb_logic[10].delayed[0] ;
 wire \comb_logic[10].pulse_out_n ;
 wire \comb_logic[11].delayed[0] ;
 wire \comb_logic[11].pulse_out_n ;
 wire \comb_logic[12].delayed[0] ;
 wire \comb_logic[12].pulse_out_n ;
 wire \comb_logic[13].delayed[0] ;
 wire \comb_logic[13].pulse_out_n ;
 wire \comb_logic[14].delayed[0] ;
 wire \comb_logic[14].pulse_out_n ;
 wire \comb_logic[15].delayed[0] ;
 wire \comb_logic[15].pulse_out_n ;
 wire \comb_logic[16].delayed[0] ;
 wire \comb_logic[16].pulse_out_n ;
 wire \comb_logic[17].delayed[0] ;
 wire \comb_logic[17].pulse_out_n ;
 wire \comb_logic[18].delayed[0] ;
 wire \comb_logic[18].pulse_out_n ;
 wire \comb_logic[19].delayed[0] ;
 wire \comb_logic[19].pulse_out_n ;
 wire \comb_logic[1].delayed[0] ;
 wire \comb_logic[1].pulse_out_n ;
 wire \comb_logic[20].delayed[0] ;
 wire \comb_logic[20].pulse_out_n ;
 wire \comb_logic[21].delayed[0] ;
 wire \comb_logic[21].pulse_out_n ;
 wire \comb_logic[22].delayed[0] ;
 wire \comb_logic[22].pulse_out_n ;
 wire \comb_logic[23].delayed[0] ;
 wire \comb_logic[23].pulse_out_n ;
 wire \comb_logic[24].delayed[0] ;
 wire \comb_logic[24].pulse_out_n ;
 wire \comb_logic[25].delayed[0] ;
 wire \comb_logic[25].pulse_out_n ;
 wire \comb_logic[26].delayed[0] ;
 wire \comb_logic[26].pulse_out_n ;
 wire \comb_logic[27].delayed[0] ;
 wire \comb_logic[27].pulse_out_n ;
 wire \comb_logic[28].delayed[0] ;
 wire \comb_logic[28].pulse_out_n ;
 wire \comb_logic[29].delayed[0] ;
 wire \comb_logic[29].pulse_out_n ;
 wire \comb_logic[2].delayed[0] ;
 wire \comb_logic[2].pulse_out_n ;
 wire \comb_logic[30].delayed[0] ;
 wire \comb_logic[30].pulse_out_n ;
 wire \comb_logic[31].delayed[0] ;
 wire \comb_logic[31].pulse_out_n ;
 wire \comb_logic[3].delayed[0] ;
 wire \comb_logic[3].pulse_out_n ;
 wire \comb_logic[4].delayed[0] ;
 wire \comb_logic[4].pulse_out_n ;
 wire \comb_logic[5].delayed[0] ;
 wire \comb_logic[5].pulse_out_n ;
 wire \comb_logic[6].delayed[0] ;
 wire \comb_logic[6].pulse_out_n ;
 wire \comb_logic[7].delayed[0] ;
 wire \comb_logic[7].pulse_out_n ;
 wire \comb_logic[8].delayed[0] ;
 wire \comb_logic[8].pulse_out_n ;
 wire \comb_logic[9].delayed[0] ;
 wire \comb_logic[9].pulse_out_n ;

 sg13g2_tielo _224_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_000_));
 sg13g2_tielo _225_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_001_));
 sg13g2_tielo _226_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_002_));
 sg13g2_tielo _227_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_003_));
 sg13g2_tielo _228_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_004_));
 sg13g2_tielo _229_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_005_));
 sg13g2_tielo _230_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_006_));
 sg13g2_tielo _231_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_007_));
 sg13g2_tielo _232_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_008_));
 sg13g2_tielo _233_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_009_));
 sg13g2_tielo _234_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_010_));
 sg13g2_tielo _235_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_011_));
 sg13g2_tielo _236_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_012_));
 sg13g2_tielo _237_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_013_));
 sg13g2_tielo _238_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_014_));
 sg13g2_tielo _239_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_015_));
 sg13g2_tielo _240_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_016_));
 sg13g2_tielo _241_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_017_));
 sg13g2_tielo _242_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_018_));
 sg13g2_tielo _243_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_019_));
 sg13g2_tielo _244_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_020_));
 sg13g2_tielo _245_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_021_));
 sg13g2_tielo _246_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_022_));
 sg13g2_tielo _247_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_023_));
 sg13g2_tielo _248_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_024_));
 sg13g2_tielo _249_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_025_));
 sg13g2_tielo _250_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_026_));
 sg13g2_tielo _251_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_027_));
 sg13g2_tielo _252_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_028_));
 sg13g2_tielo _253_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_029_));
 sg13g2_tielo _254_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_030_));
 sg13g2_tielo _255_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_031_));
 sg13g2_tielo _256_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_032_));
 sg13g2_tielo _257_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_033_));
 sg13g2_tielo _258_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_034_));
 sg13g2_tielo _259_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_035_));
 sg13g2_tielo _260_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_036_));
 sg13g2_tielo _261_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_037_));
 sg13g2_tielo _262_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_038_));
 sg13g2_tielo _263_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_039_));
 sg13g2_tielo _264_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_040_));
 sg13g2_tielo _265_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_041_));
 sg13g2_tielo _266_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_042_));
 sg13g2_tielo _267_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_043_));
 sg13g2_tielo _268_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_044_));
 sg13g2_tielo _269_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_045_));
 sg13g2_tielo _270_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_046_));
 sg13g2_tielo _271_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_047_));
 sg13g2_tielo _272_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_048_));
 sg13g2_tielo _273_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_049_));
 sg13g2_tielo _274_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_050_));
 sg13g2_tielo _275_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_051_));
 sg13g2_tielo _276_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_052_));
 sg13g2_tielo _277_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_053_));
 sg13g2_tielo _278_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_054_));
 sg13g2_tielo _279_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_055_));
 sg13g2_tielo _280_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_056_));
 sg13g2_tielo _281_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_057_));
 sg13g2_tielo _282_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_058_));
 sg13g2_tielo _283_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_059_));
 sg13g2_tielo _284_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_060_));
 sg13g2_tielo _285_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_061_));
 sg13g2_tielo _286_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_062_));
 sg13g2_tielo _287_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_063_));
 sg13g2_tielo _288_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_064_));
 sg13g2_tielo _289_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_065_));
 sg13g2_tielo _290_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_066_));
 sg13g2_tielo _291_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_067_));
 sg13g2_tielo _292_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_068_));
 sg13g2_tielo _293_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_069_));
 sg13g2_tielo _294_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_070_));
 sg13g2_tielo _295_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_071_));
 sg13g2_tielo _296_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_072_));
 sg13g2_tielo _297_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_073_));
 sg13g2_tielo _298_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_074_));
 sg13g2_tielo _299_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_075_));
 sg13g2_tielo _300_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_076_));
 sg13g2_tielo _301_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_077_));
 sg13g2_tielo _302_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_078_));
 sg13g2_tielo _303_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_079_));
 sg13g2_tielo _304_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_080_));
 sg13g2_tielo _305_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_081_));
 sg13g2_tielo _306_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_082_));
 sg13g2_tielo _307_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_083_));
 sg13g2_tielo _308_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_084_));
 sg13g2_tielo _309_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_085_));
 sg13g2_tielo _310_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_086_));
 sg13g2_tielo _311_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_087_));
 sg13g2_tielo _312_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_088_));
 sg13g2_tielo _313_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_089_));
 sg13g2_tielo _314_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_090_));
 sg13g2_tielo _315_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_091_));
 sg13g2_tielo _316_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_092_));
 sg13g2_tielo _317_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_093_));
 sg13g2_tielo _318_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_094_));
 sg13g2_tielo _319_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_095_));
 sg13g2_tielo _320_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_096_));
 sg13g2_tielo _321_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_097_));
 sg13g2_tielo _322_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_098_));
 sg13g2_tielo _323_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_099_));
 sg13g2_tielo _324_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_100_));
 sg13g2_tielo _325_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_101_));
 sg13g2_tielo _326_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_102_));
 sg13g2_tielo _327_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_103_));
 sg13g2_tielo _328_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_104_));
 sg13g2_tielo _329_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_105_));
 sg13g2_tielo _330_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_106_));
 sg13g2_tielo _331_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_107_));
 sg13g2_tielo _332_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_108_));
 sg13g2_tielo _333_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_109_));
 sg13g2_tielo _334_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_110_));
 sg13g2_tielo _335_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_111_));
 sg13g2_tielo _336_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_112_));
 sg13g2_tielo _337_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_113_));
 sg13g2_tielo _338_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_114_));
 sg13g2_tielo _339_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_115_));
 sg13g2_tielo _340_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_116_));
 sg13g2_tielo _341_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_117_));
 sg13g2_tielo _342_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_118_));
 sg13g2_tielo _343_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_119_));
 sg13g2_tielo _344_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_120_));
 sg13g2_tielo _345_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_121_));
 sg13g2_tielo _346_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_122_));
 sg13g2_tielo _347_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_123_));
 sg13g2_tielo _348_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_124_));
 sg13g2_tielo _349_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_125_));
 sg13g2_tielo _350_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_126_));
 sg13g2_tielo _351_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_127_));
 sg13g2_tielo _352_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_128_));
 sg13g2_tielo _353_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_129_));
 sg13g2_tielo _354_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_130_));
 sg13g2_tielo _355_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_131_));
 sg13g2_tielo _356_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_132_));
 sg13g2_tielo _357_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_133_));
 sg13g2_tielo _358_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_134_));
 sg13g2_tielo _359_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_135_));
 sg13g2_tielo _360_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_136_));
 sg13g2_tielo _361_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_137_));
 sg13g2_tielo _362_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_138_));
 sg13g2_tielo _363_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_139_));
 sg13g2_tielo _364_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_140_));
 sg13g2_tielo _365_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_141_));
 sg13g2_tielo _366_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_142_));
 sg13g2_tielo _367_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_143_));
 sg13g2_tielo _368_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_144_));
 sg13g2_tielo _369_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_145_));
 sg13g2_tielo _370_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_146_));
 sg13g2_tielo _371_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_147_));
 sg13g2_tielo _372_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_148_));
 sg13g2_tielo _373_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_149_));
 sg13g2_tielo _374_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_150_));
 sg13g2_tielo _375_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_151_));
 sg13g2_tielo _376_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_152_));
 sg13g2_tielo _377_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_153_));
 sg13g2_tielo _378_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_154_));
 sg13g2_tielo _379_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_155_));
 sg13g2_tielo _380_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_156_));
 sg13g2_tielo _381_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_157_));
 sg13g2_tielo _382_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_158_));
 sg13g2_tielo _383_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(_159_));
 sg13g2_tielo _384_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[0]));
 sg13g2_tielo _385_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[1]));
 sg13g2_tielo _386_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[2]));
 sg13g2_tielo _387_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[3]));
 sg13g2_tielo _388_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[4]));
 sg13g2_tielo _389_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[5]));
 sg13g2_tielo _390_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[6]));
 sg13g2_tielo _391_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[7]));
 sg13g2_tielo _392_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[8]));
 sg13g2_tielo _393_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[9]));
 sg13g2_tielo _394_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[10]));
 sg13g2_tielo _395_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[11]));
 sg13g2_tielo _396_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[12]));
 sg13g2_tielo _397_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[13]));
 sg13g2_tielo _398_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[14]));
 sg13g2_tielo _399_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[15]));
 sg13g2_tielo _400_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[16]));
 sg13g2_tielo _401_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[17]));
 sg13g2_tielo _402_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[18]));
 sg13g2_tielo _403_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[19]));
 sg13g2_tielo _404_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[20]));
 sg13g2_tielo _405_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[21]));
 sg13g2_tielo _406_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[22]));
 sg13g2_tielo _407_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[23]));
 sg13g2_tielo _408_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[24]));
 sg13g2_tielo _409_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[25]));
 sg13g2_tielo _410_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[26]));
 sg13g2_tielo _411_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[27]));
 sg13g2_tielo _412_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[28]));
 sg13g2_tielo _413_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[29]));
 sg13g2_tielo _414_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[30]));
 sg13g2_tielo _415_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON[31]));
 sg13g2_tielo _416_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[0]));
 sg13g2_tielo _417_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[1]));
 sg13g2_tielo _418_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[2]));
 sg13g2_tielo _419_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[3]));
 sg13g2_tielo _420_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[4]));
 sg13g2_tielo _421_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[5]));
 sg13g2_tielo _422_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[6]));
 sg13g2_tielo _423_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[7]));
 sg13g2_tielo _424_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[8]));
 sg13g2_tielo _425_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[9]));
 sg13g2_tielo _426_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[10]));
 sg13g2_tielo _427_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[11]));
 sg13g2_tielo _428_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[12]));
 sg13g2_tielo _429_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[13]));
 sg13g2_tielo _430_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[14]));
 sg13g2_tielo _431_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[15]));
 sg13g2_tielo _432_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[16]));
 sg13g2_tielo _433_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[17]));
 sg13g2_tielo _434_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[18]));
 sg13g2_tielo _435_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[19]));
 sg13g2_tielo _436_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[20]));
 sg13g2_tielo _437_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[21]));
 sg13g2_tielo _438_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[22]));
 sg13g2_tielo _439_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[23]));
 sg13g2_tielo _440_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[24]));
 sg13g2_tielo _441_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[25]));
 sg13g2_tielo _442_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[26]));
 sg13g2_tielo _443_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[27]));
 sg13g2_tielo _444_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[28]));
 sg13g2_tielo _445_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[29]));
 sg13g2_tielo _446_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[30]));
 sg13g2_tielo _447_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(ON_N[31]));
 sg13g2_tielo _448_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[0].pulse_out_n ));
 sg13g2_tielo _449_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[10].pulse_out_n ));
 sg13g2_tielo _450_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[11].pulse_out_n ));
 sg13g2_tielo _451_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[12].pulse_out_n ));
 sg13g2_tielo _452_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[13].pulse_out_n ));
 sg13g2_tielo _453_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[14].pulse_out_n ));
 sg13g2_tielo _454_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[15].pulse_out_n ));
 sg13g2_tielo _455_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[16].pulse_out_n ));
 sg13g2_tielo _456_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[17].pulse_out_n ));
 sg13g2_tielo _457_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[18].pulse_out_n ));
 sg13g2_tielo _458_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[19].pulse_out_n ));
 sg13g2_tielo _459_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[1].pulse_out_n ));
 sg13g2_tielo _460_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[20].pulse_out_n ));
 sg13g2_tielo _461_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[21].pulse_out_n ));
 sg13g2_tielo _462_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[22].pulse_out_n ));
 sg13g2_tielo _463_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[23].pulse_out_n ));
 sg13g2_tielo _464_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[24].pulse_out_n ));
 sg13g2_tielo _465_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[25].pulse_out_n ));
 sg13g2_tielo _466_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[26].pulse_out_n ));
 sg13g2_tielo _467_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[27].pulse_out_n ));
 sg13g2_tielo _468_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[28].pulse_out_n ));
 sg13g2_tielo _469_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[29].pulse_out_n ));
 sg13g2_tielo _470_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[2].pulse_out_n ));
 sg13g2_tielo _471_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[30].pulse_out_n ));
 sg13g2_tielo _472_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[31].pulse_out_n ));
 sg13g2_tielo _473_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[3].pulse_out_n ));
 sg13g2_tielo _474_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[4].pulse_out_n ));
 sg13g2_tielo _475_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[5].pulse_out_n ));
 sg13g2_tielo _476_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[6].pulse_out_n ));
 sg13g2_tielo _477_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[7].pulse_out_n ));
 sg13g2_tielo _478_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[8].pulse_out_n ));
 sg13g2_tielo _479_ (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(\comb_logic[9].pulse_out_n ));
 sg13g2_dlygate4sd1_1 \comb_logic[0].delay1_I  (.A(thermo[0]),
    .X(_172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[0].nand_on_I  (.Y(_192_),
    .A(_000_),
    .B(_001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[0].nand_on_n_I  (.Y(thermo[0]),
    .A(_002_),
    .B(_003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[0].xor_pulse_I  (.Y(\comb_logic[0].delayed[0] ),
    .A(_004_),
    .B(thermo[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[10].delay1_I  (.A(thermo[10]),
    .X(_176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[10].nand_on_I  (.Y(_202_),
    .A(_005_),
    .B(_006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[10].nand_on_n_I  (.Y(thermo[10]),
    .A(_007_),
    .B(_008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[10].xor_pulse_I  (.Y(\comb_logic[10].delayed[0] ),
    .A(_009_),
    .B(thermo[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[11].delay1_I  (.A(thermo[11]),
    .X(_177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[11].nand_on_I  (.Y(_203_),
    .A(_010_),
    .B(_011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[11].nand_on_n_I  (.Y(thermo[11]),
    .A(_012_),
    .B(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[11].xor_pulse_I  (.Y(\comb_logic[11].delayed[0] ),
    .A(_014_),
    .B(thermo[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[12].delay1_I  (.A(thermo[12]),
    .X(_178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[12].nand_on_I  (.Y(_204_),
    .A(_015_),
    .B(_016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[12].nand_on_n_I  (.Y(thermo[12]),
    .A(_017_),
    .B(_018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[12].xor_pulse_I  (.Y(\comb_logic[12].delayed[0] ),
    .A(_019_),
    .B(thermo[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[13].delay1_I  (.A(thermo[13]),
    .X(_179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[13].nand_on_I  (.Y(_205_),
    .A(_020_),
    .B(_021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[13].nand_on_n_I  (.Y(thermo[13]),
    .A(_022_),
    .B(_023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[13].xor_pulse_I  (.Y(\comb_logic[13].delayed[0] ),
    .A(_024_),
    .B(thermo[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[14].delay1_I  (.A(thermo[14]),
    .X(_180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[14].nand_on_I  (.Y(_206_),
    .A(_025_),
    .B(_026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[14].nand_on_n_I  (.Y(thermo[14]),
    .A(_027_),
    .B(_028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[14].xor_pulse_I  (.Y(\comb_logic[14].delayed[0] ),
    .A(_029_),
    .B(thermo[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[15].delay1_I  (.A(thermo[15]),
    .X(_181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[15].nand_on_I  (.Y(_207_),
    .A(_030_),
    .B(_031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[15].nand_on_n_I  (.Y(thermo[15]),
    .A(_032_),
    .B(_033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[15].xor_pulse_I  (.Y(\comb_logic[15].delayed[0] ),
    .A(_034_),
    .B(thermo[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[16].delay1_I  (.A(thermo[16]),
    .X(_182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[16].nand_on_I  (.Y(_208_),
    .A(_035_),
    .B(_036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[16].nand_on_n_I  (.Y(thermo[16]),
    .A(_037_),
    .B(_038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[16].xor_pulse_I  (.Y(\comb_logic[16].delayed[0] ),
    .A(_039_),
    .B(thermo[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[17].delay1_I  (.A(thermo[17]),
    .X(_184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[17].nand_on_I  (.Y(_209_),
    .A(_040_),
    .B(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[17].nand_on_n_I  (.Y(thermo[17]),
    .A(_042_),
    .B(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[17].xor_pulse_I  (.Y(\comb_logic[17].delayed[0] ),
    .A(_044_),
    .B(thermo[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[18].delay1_I  (.A(thermo[18]),
    .X(_185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[18].nand_on_I  (.Y(_210_),
    .A(_045_),
    .B(_046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[18].nand_on_n_I  (.Y(thermo[18]),
    .A(_047_),
    .B(_048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[18].xor_pulse_I  (.Y(\comb_logic[18].delayed[0] ),
    .A(_049_),
    .B(thermo[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[19].delay1_I  (.A(thermo[19]),
    .X(_186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[19].nand_on_I  (.Y(_211_),
    .A(_050_),
    .B(_051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[19].nand_on_n_I  (.Y(thermo[19]),
    .A(_052_),
    .B(_053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[19].xor_pulse_I  (.Y(\comb_logic[19].delayed[0] ),
    .A(_054_),
    .B(thermo[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[1].delay1_I  (.A(thermo[1]),
    .X(_183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[1].nand_on_I  (.Y(_193_),
    .A(_055_),
    .B(_056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[1].nand_on_n_I  (.Y(thermo[1]),
    .A(_057_),
    .B(_058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[1].xor_pulse_I  (.Y(\comb_logic[1].delayed[0] ),
    .A(_059_),
    .B(thermo[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[20].delay1_I  (.A(thermo[20]),
    .X(_187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[20].nand_on_I  (.Y(_212_),
    .A(_060_),
    .B(_061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[20].nand_on_n_I  (.Y(thermo[20]),
    .A(_062_),
    .B(_063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[20].xor_pulse_I  (.Y(\comb_logic[20].delayed[0] ),
    .A(_064_),
    .B(thermo[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[21].delay1_I  (.A(thermo[21]),
    .X(_188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[21].nand_on_I  (.Y(_213_),
    .A(_065_),
    .B(_066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[21].nand_on_n_I  (.Y(thermo[21]),
    .A(_067_),
    .B(_068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[21].xor_pulse_I  (.Y(\comb_logic[21].delayed[0] ),
    .A(_069_),
    .B(thermo[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[22].delay1_I  (.A(thermo[22]),
    .X(_189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[22].nand_on_I  (.Y(_214_),
    .A(_070_),
    .B(_071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[22].nand_on_n_I  (.Y(thermo[22]),
    .A(_072_),
    .B(_073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[22].xor_pulse_I  (.Y(\comb_logic[22].delayed[0] ),
    .A(_074_),
    .B(thermo[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[23].delay1_I  (.A(thermo[23]),
    .X(_190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[23].nand_on_I  (.Y(_215_),
    .A(_075_),
    .B(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[23].nand_on_n_I  (.Y(thermo[23]),
    .A(_077_),
    .B(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[23].xor_pulse_I  (.Y(\comb_logic[23].delayed[0] ),
    .A(_079_),
    .B(thermo[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[24].delay1_I  (.A(thermo[24]),
    .X(_191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[24].nand_on_I  (.Y(_216_),
    .A(_080_),
    .B(_081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[24].nand_on_n_I  (.Y(thermo[24]),
    .A(_082_),
    .B(_083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[24].xor_pulse_I  (.Y(\comb_logic[24].delayed[0] ),
    .A(_084_),
    .B(thermo[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[25].delay1_I  (.A(thermo[25]),
    .X(_160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[25].nand_on_I  (.Y(_217_),
    .A(_085_),
    .B(_086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[25].nand_on_n_I  (.Y(thermo[25]),
    .A(_087_),
    .B(_088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[25].xor_pulse_I  (.Y(\comb_logic[25].delayed[0] ),
    .A(_089_),
    .B(thermo[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[26].delay1_I  (.A(thermo[26]),
    .X(_161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[26].nand_on_I  (.Y(_218_),
    .A(_090_),
    .B(_091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[26].nand_on_n_I  (.Y(thermo[26]),
    .A(_092_),
    .B(_093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[26].xor_pulse_I  (.Y(\comb_logic[26].delayed[0] ),
    .A(_094_),
    .B(thermo[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[27].delay1_I  (.A(thermo[27]),
    .X(_163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[27].nand_on_I  (.Y(_219_),
    .A(_095_),
    .B(_096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[27].nand_on_n_I  (.Y(thermo[27]),
    .A(_097_),
    .B(_098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[27].xor_pulse_I  (.Y(\comb_logic[27].delayed[0] ),
    .A(_099_),
    .B(thermo[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[28].delay1_I  (.A(thermo[28]),
    .X(_164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[28].nand_on_I  (.Y(_220_),
    .A(_100_),
    .B(_101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[28].nand_on_n_I  (.Y(thermo[28]),
    .A(_102_),
    .B(_103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[28].xor_pulse_I  (.Y(\comb_logic[28].delayed[0] ),
    .A(_104_),
    .B(thermo[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[29].delay1_I  (.A(thermo[29]),
    .X(_165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[29].nand_on_I  (.Y(_221_),
    .A(_105_),
    .B(_106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[29].nand_on_n_I  (.Y(thermo[29]),
    .A(_107_),
    .B(_108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[29].xor_pulse_I  (.Y(\comb_logic[29].delayed[0] ),
    .A(_109_),
    .B(thermo[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[2].delay1_I  (.A(thermo[2]),
    .X(_162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[2].nand_on_I  (.Y(_194_),
    .A(_110_),
    .B(_111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[2].nand_on_n_I  (.Y(thermo[2]),
    .A(_112_),
    .B(_113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[2].xor_pulse_I  (.Y(\comb_logic[2].delayed[0] ),
    .A(_114_),
    .B(thermo[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[30].delay1_I  (.A(thermo[30]),
    .X(_166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[30].nand_on_I  (.Y(_222_),
    .A(_115_),
    .B(_116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[30].nand_on_n_I  (.Y(thermo[30]),
    .A(_117_),
    .B(_118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[30].xor_pulse_I  (.Y(\comb_logic[30].delayed[0] ),
    .A(_119_),
    .B(thermo[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[31].delay1_I  (.A(thermo[31]),
    .X(_167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[31].nand_on_I  (.Y(_223_),
    .A(_120_),
    .B(_121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[31].nand_on_n_I  (.Y(thermo[31]),
    .A(_122_),
    .B(_123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[31].xor_pulse_I  (.Y(\comb_logic[31].delayed[0] ),
    .A(_124_),
    .B(thermo[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[3].delay1_I  (.A(thermo[3]),
    .X(_168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[3].nand_on_I  (.Y(_195_),
    .A(_125_),
    .B(_126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[3].nand_on_n_I  (.Y(thermo[3]),
    .A(_127_),
    .B(_128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[3].xor_pulse_I  (.Y(\comb_logic[3].delayed[0] ),
    .A(_129_),
    .B(thermo[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[4].delay1_I  (.A(thermo[4]),
    .X(_169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[4].nand_on_I  (.Y(_196_),
    .A(_130_),
    .B(_131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[4].nand_on_n_I  (.Y(thermo[4]),
    .A(_132_),
    .B(_133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[4].xor_pulse_I  (.Y(\comb_logic[4].delayed[0] ),
    .A(_134_),
    .B(thermo[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[5].delay1_I  (.A(thermo[5]),
    .X(_170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[5].nand_on_I  (.Y(_197_),
    .A(_135_),
    .B(_136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[5].nand_on_n_I  (.Y(thermo[5]),
    .A(_137_),
    .B(_138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[5].xor_pulse_I  (.Y(\comb_logic[5].delayed[0] ),
    .A(_139_),
    .B(thermo[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[6].delay1_I  (.A(thermo[6]),
    .X(_171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[6].nand_on_I  (.Y(_198_),
    .A(_140_),
    .B(_141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[6].nand_on_n_I  (.Y(thermo[6]),
    .A(_142_),
    .B(_143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[6].xor_pulse_I  (.Y(\comb_logic[6].delayed[0] ),
    .A(_144_),
    .B(thermo[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[7].delay1_I  (.A(thermo[7]),
    .X(_173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[7].nand_on_I  (.Y(_199_),
    .A(_145_),
    .B(_146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[7].nand_on_n_I  (.Y(thermo[7]),
    .A(_147_),
    .B(_148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[7].xor_pulse_I  (.Y(\comb_logic[7].delayed[0] ),
    .A(_149_),
    .B(thermo[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[8].delay1_I  (.A(thermo[8]),
    .X(_174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[8].nand_on_I  (.Y(_200_),
    .A(_150_),
    .B(_151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[8].nand_on_n_I  (.Y(thermo[8]),
    .A(_152_),
    .B(_153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[8].xor_pulse_I  (.Y(\comb_logic[8].delayed[0] ),
    .A(_154_),
    .B(thermo[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd1_1 \comb_logic[9].delay1_I  (.A(thermo[9]),
    .X(_175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[9].nand_on_I  (.Y(_201_),
    .A(_155_),
    .B(_156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 \comb_logic[9].nand_on_n_I  (.Y(thermo[9]),
    .A(_157_),
    .B(_158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 \comb_logic[9].xor_pulse_I  (.Y(\comb_logic[9].delayed[0] ),
    .A(_159_),
    .B(thermo[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_153 (.VDD(VPWR),
    .VSS(VGND));
endmodule
