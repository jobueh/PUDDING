magic
tech ihp-sg13g2
magscale 1 2
timestamp 1756158664
<< metal1 >>
rect 576 12872 15360 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 15360 12872
rect 576 12808 15360 12832
rect 1123 12704 1181 12705
rect 1123 12664 1132 12704
rect 1172 12664 1181 12704
rect 1123 12663 1181 12664
rect 3043 12704 3101 12705
rect 3043 12664 3052 12704
rect 3092 12664 3101 12704
rect 3043 12663 3101 12664
rect 3235 12704 3293 12705
rect 3235 12664 3244 12704
rect 3284 12664 3293 12704
rect 3235 12663 3293 12664
rect 3811 12704 3869 12705
rect 3811 12664 3820 12704
rect 3860 12664 3869 12704
rect 3811 12663 3869 12664
rect 4003 12704 4061 12705
rect 4003 12664 4012 12704
rect 4052 12664 4061 12704
rect 4003 12663 4061 12664
rect 4579 12704 4637 12705
rect 4579 12664 4588 12704
rect 4628 12664 4637 12704
rect 4579 12663 4637 12664
rect 5827 12704 5885 12705
rect 5827 12664 5836 12704
rect 5876 12664 5885 12704
rect 5827 12663 5885 12664
rect 6787 12704 6845 12705
rect 6787 12664 6796 12704
rect 6836 12664 6845 12704
rect 6787 12663 6845 12664
rect 9571 12704 9629 12705
rect 9571 12664 9580 12704
rect 9620 12664 9629 12704
rect 9571 12663 9629 12664
rect 9763 12704 9821 12705
rect 9763 12664 9772 12704
rect 9812 12664 9821 12704
rect 9763 12663 9821 12664
rect 11587 12704 11645 12705
rect 11587 12664 11596 12704
rect 11636 12664 11645 12704
rect 11587 12663 11645 12664
rect 11779 12704 11837 12705
rect 11779 12664 11788 12704
rect 11828 12664 11837 12704
rect 11779 12663 11837 12664
rect 13987 12704 14045 12705
rect 13987 12664 13996 12704
rect 14036 12664 14045 12704
rect 13987 12663 14045 12664
rect 14371 12704 14429 12705
rect 14371 12664 14380 12704
rect 14420 12664 14429 12704
rect 14371 12663 14429 12664
rect 14755 12704 14813 12705
rect 14755 12664 14764 12704
rect 14804 12664 14813 12704
rect 14755 12663 14813 12664
rect 15139 12704 15197 12705
rect 15139 12664 15148 12704
rect 15188 12664 15197 12704
rect 15139 12663 15197 12664
rect 1611 12620 1653 12629
rect 1611 12580 1612 12620
rect 1652 12580 1653 12620
rect 1611 12571 1653 12580
rect 1419 12536 1461 12545
rect 1419 12496 1420 12536
rect 1460 12496 1461 12536
rect 1419 12487 1461 12496
rect 1891 12536 1949 12537
rect 1891 12496 1900 12536
rect 1940 12496 1949 12536
rect 1891 12495 1949 12496
rect 5059 12536 5117 12537
rect 5059 12496 5068 12536
rect 5108 12496 5117 12536
rect 5059 12495 5117 12496
rect 5155 12536 5213 12537
rect 5155 12496 5164 12536
rect 5204 12496 5213 12536
rect 5155 12495 5213 12496
rect 6019 12536 6077 12537
rect 6019 12496 6028 12536
rect 6068 12496 6077 12536
rect 6019 12495 6077 12496
rect 1611 12452 1653 12461
rect 1611 12412 1612 12452
rect 1652 12412 1653 12452
rect 1611 12403 1653 12412
rect 1419 12284 1461 12293
rect 1419 12244 1420 12284
rect 1460 12244 1461 12284
rect 1419 12235 1461 12244
rect 576 12116 15360 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 15360 12116
rect 576 12052 15360 12076
rect 6027 11864 6069 11873
rect 6027 11824 6028 11864
rect 6068 11824 6069 11864
rect 6027 11815 6069 11824
rect 5931 11780 5973 11789
rect 5931 11740 5932 11780
rect 5972 11740 5973 11780
rect 5931 11731 5973 11740
rect 7467 11780 7509 11789
rect 7467 11740 7468 11780
rect 7508 11740 7509 11780
rect 7467 11731 7509 11740
rect 9771 11780 9813 11789
rect 9771 11740 9772 11780
rect 9812 11740 9813 11780
rect 9771 11731 9813 11740
rect 11787 11780 11829 11789
rect 11787 11740 11788 11780
rect 11828 11740 11829 11780
rect 11787 11731 11829 11740
rect 1123 11696 1181 11697
rect 1123 11656 1132 11696
rect 1172 11656 1181 11696
rect 1123 11655 1181 11656
rect 1219 11696 1277 11697
rect 1219 11656 1228 11696
rect 1268 11656 1277 11696
rect 1219 11655 1277 11656
rect 3043 11696 3101 11697
rect 3043 11656 3052 11696
rect 3092 11656 3101 11696
rect 3043 11655 3101 11656
rect 3139 11696 3197 11697
rect 3139 11656 3148 11696
rect 3188 11656 3197 11696
rect 3139 11655 3197 11656
rect 3619 11696 3677 11697
rect 3619 11656 3628 11696
rect 3668 11656 3677 11696
rect 3619 11655 3677 11656
rect 6123 11696 6165 11705
rect 6123 11656 6124 11696
rect 6164 11656 6165 11696
rect 6123 11647 6165 11656
rect 7275 11696 7317 11705
rect 7275 11656 7276 11696
rect 7316 11656 7317 11696
rect 7275 11647 7317 11656
rect 7371 11696 7413 11705
rect 7371 11656 7372 11696
rect 7412 11656 7413 11696
rect 7371 11647 7413 11656
rect 9579 11696 9621 11705
rect 9579 11656 9580 11696
rect 9620 11656 9621 11696
rect 9579 11647 9621 11656
rect 11595 11696 11637 11705
rect 11595 11656 11596 11696
rect 11636 11656 11637 11696
rect 11595 11647 11637 11656
rect 1987 11528 2045 11529
rect 1987 11488 1996 11528
rect 2036 11488 2045 11528
rect 1987 11487 2045 11488
rect 2179 11528 2237 11529
rect 2179 11488 2188 11528
rect 2228 11488 2237 11528
rect 2179 11487 2237 11488
rect 5155 11528 5213 11529
rect 5155 11488 5164 11528
rect 5204 11488 5213 11528
rect 5155 11487 5213 11488
rect 6979 11528 7037 11529
rect 6979 11488 6988 11528
rect 7028 11488 7037 11528
rect 6979 11487 7037 11488
rect 7747 11528 7805 11529
rect 7747 11488 7756 11528
rect 7796 11488 7805 11528
rect 7747 11487 7805 11488
rect 9283 11528 9341 11529
rect 9283 11488 9292 11528
rect 9332 11488 9341 11528
rect 9283 11487 9341 11488
rect 10051 11528 10109 11529
rect 10051 11488 10060 11528
rect 10100 11488 10109 11528
rect 10051 11487 10109 11488
rect 10915 11528 10973 11529
rect 10915 11488 10924 11528
rect 10964 11488 10973 11528
rect 10915 11487 10973 11488
rect 13603 11528 13661 11529
rect 13603 11488 13612 11528
rect 13652 11488 13661 11528
rect 13603 11487 13661 11488
rect 13987 11528 14045 11529
rect 13987 11488 13996 11528
rect 14036 11488 14045 11528
rect 13987 11487 14045 11488
rect 14371 11528 14429 11529
rect 14371 11488 14380 11528
rect 14420 11488 14429 11528
rect 14371 11487 14429 11488
rect 14755 11528 14813 11529
rect 14755 11488 14764 11528
rect 14804 11488 14813 11528
rect 14755 11487 14813 11488
rect 15139 11528 15197 11529
rect 15139 11488 15148 11528
rect 15188 11488 15197 11528
rect 15139 11487 15197 11488
rect 576 11360 15360 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 15360 11360
rect 576 11296 15360 11320
rect 2659 11192 2717 11193
rect 2659 11152 2668 11192
rect 2708 11152 2717 11192
rect 2659 11151 2717 11152
rect 3235 11192 3293 11193
rect 3235 11152 3244 11192
rect 3284 11152 3293 11192
rect 3235 11151 3293 11152
rect 4387 11192 4445 11193
rect 4387 11152 4396 11192
rect 4436 11152 4445 11192
rect 4387 11151 4445 11152
rect 7555 11192 7613 11193
rect 7555 11152 7564 11192
rect 7604 11152 7613 11192
rect 7555 11151 7613 11152
rect 10627 11192 10685 11193
rect 10627 11152 10636 11192
rect 10676 11152 10685 11192
rect 10627 11151 10685 11152
rect 11395 11192 11453 11193
rect 11395 11152 11404 11192
rect 11444 11152 11453 11192
rect 11395 11151 11453 11152
rect 12163 11192 12221 11193
rect 12163 11152 12172 11192
rect 12212 11152 12221 11192
rect 12163 11151 12221 11152
rect 12931 11192 12989 11193
rect 12931 11152 12940 11192
rect 12980 11152 12989 11192
rect 12931 11151 12989 11152
rect 13795 11192 13853 11193
rect 13795 11152 13804 11192
rect 13844 11152 13853 11192
rect 13795 11151 13853 11152
rect 14179 11192 14237 11193
rect 14179 11152 14188 11192
rect 14228 11152 14237 11192
rect 14179 11151 14237 11152
rect 14563 11192 14621 11193
rect 14563 11152 14572 11192
rect 14612 11152 14621 11192
rect 14563 11151 14621 11152
rect 14947 11192 15005 11193
rect 14947 11152 14956 11192
rect 14996 11152 15005 11192
rect 14947 11151 15005 11152
rect 1131 11024 1173 11033
rect 1131 10984 1132 11024
rect 1172 10984 1173 11024
rect 1131 10975 1173 10984
rect 1219 11024 1277 11025
rect 1219 10984 1228 11024
rect 1268 10984 1277 11024
rect 1219 10983 1277 10984
rect 1891 11024 1949 11025
rect 1891 10984 1900 11024
rect 1940 10984 1949 11024
rect 1891 10983 1949 10984
rect 3531 11024 3573 11033
rect 3531 10984 3532 11024
rect 3572 10984 3573 11024
rect 3531 10975 3573 10984
rect 3627 11024 3669 11033
rect 3627 10984 3628 11024
rect 3668 10984 3669 11024
rect 3627 10975 3669 10984
rect 4683 11024 4725 11033
rect 4683 10984 4684 11024
rect 4724 10984 4725 11024
rect 4683 10975 4725 10984
rect 5347 11024 5405 11025
rect 5347 10984 5356 11024
rect 5396 10984 5405 11024
rect 5347 10983 5405 10984
rect 5443 11024 5501 11025
rect 5443 10984 5452 11024
rect 5492 10984 5501 11024
rect 5443 10983 5501 10984
rect 5923 11024 5981 11025
rect 5923 10984 5932 11024
rect 5972 10984 5981 11024
rect 5923 10983 5981 10984
rect 8035 11024 8093 11025
rect 8035 10984 8044 11024
rect 8084 10984 8093 11024
rect 8035 10983 8093 10984
rect 8131 11024 8189 11025
rect 8131 10984 8140 11024
rect 8180 10984 8189 11024
rect 8131 10983 8189 10984
rect 8515 11024 8573 11025
rect 8515 10984 8524 11024
rect 8564 10984 8573 11024
rect 8515 10983 8573 10984
rect 9675 11024 9717 11033
rect 9675 10984 9676 11024
rect 9716 10984 9717 11024
rect 9675 10975 9717 10984
rect 11115 11024 11157 11033
rect 11115 10984 11116 11024
rect 11156 10984 11157 11024
rect 11115 10975 11157 10984
rect 12459 11024 12501 11033
rect 12459 10984 12460 11024
rect 12500 10984 12501 11024
rect 12459 10975 12501 10984
rect 3723 10940 3765 10949
rect 3723 10900 3724 10940
rect 3764 10900 3765 10940
rect 3723 10891 3765 10900
rect 4875 10940 4917 10949
rect 4875 10900 4876 10940
rect 4916 10900 4917 10940
rect 4875 10891 4917 10900
rect 9867 10940 9909 10949
rect 9867 10900 9868 10940
rect 9908 10900 9909 10940
rect 9867 10891 9909 10900
rect 10923 10940 10965 10949
rect 10923 10900 10924 10940
rect 10964 10900 10965 10940
rect 10923 10891 10965 10900
rect 12651 10940 12693 10949
rect 12651 10900 12652 10940
rect 12692 10900 12693 10940
rect 12651 10891 12693 10900
rect 4675 10856 4733 10857
rect 4675 10816 4684 10856
rect 4724 10816 4733 10856
rect 4675 10815 4733 10816
rect 576 10604 15360 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 15360 10604
rect 576 10540 15360 10564
rect 1707 10436 1749 10445
rect 1707 10396 1708 10436
rect 1748 10396 1749 10436
rect 1707 10387 1749 10396
rect 1899 10268 1941 10277
rect 1899 10228 1900 10268
rect 1940 10228 1941 10268
rect 1899 10219 1941 10228
rect 9195 10268 9237 10277
rect 9195 10228 9196 10268
rect 9236 10228 9237 10268
rect 9195 10219 9237 10228
rect 10635 10268 10677 10277
rect 10635 10228 10636 10268
rect 10676 10228 10677 10268
rect 10635 10219 10677 10228
rect 11019 10268 11061 10277
rect 11019 10228 11020 10268
rect 11060 10228 11061 10268
rect 11019 10219 11061 10228
rect 12555 10268 12597 10277
rect 12555 10228 12556 10268
rect 12596 10228 12597 10268
rect 12555 10219 12597 10228
rect 1707 10184 1749 10193
rect 1707 10144 1708 10184
rect 1748 10144 1749 10184
rect 1707 10135 1749 10144
rect 3147 10184 3189 10193
rect 3147 10144 3148 10184
rect 3188 10144 3189 10184
rect 3147 10135 3189 10144
rect 3235 10184 3293 10185
rect 3235 10144 3244 10184
rect 3284 10144 3293 10184
rect 3235 10143 3293 10144
rect 3715 10184 3773 10185
rect 3715 10144 3724 10184
rect 3764 10144 3773 10184
rect 3715 10143 3773 10144
rect 9003 10184 9045 10193
rect 9003 10144 9004 10184
rect 9044 10144 9045 10184
rect 9003 10135 9045 10144
rect 10443 10184 10485 10193
rect 10443 10144 10444 10184
rect 10484 10144 10485 10184
rect 10443 10135 10485 10144
rect 11211 10184 11253 10193
rect 11211 10144 11212 10184
rect 11252 10144 11253 10184
rect 11211 10135 11253 10144
rect 12363 10184 12405 10193
rect 12363 10144 12364 10184
rect 12404 10144 12405 10184
rect 12363 10135 12405 10144
rect 1027 10016 1085 10017
rect 1027 9976 1036 10016
rect 1076 9976 1085 10016
rect 1027 9975 1085 9976
rect 1411 10016 1469 10017
rect 1411 9976 1420 10016
rect 1460 9976 1469 10016
rect 1411 9975 1469 9976
rect 2179 10016 2237 10017
rect 2179 9976 2188 10016
rect 2228 9976 2237 10016
rect 2179 9975 2237 9976
rect 2755 10016 2813 10017
rect 2755 9976 2764 10016
rect 2804 9976 2813 10016
rect 2755 9975 2813 9976
rect 4483 10016 4541 10017
rect 4483 9976 4492 10016
rect 4532 9976 4541 10016
rect 4483 9975 4541 9976
rect 5155 10016 5213 10017
rect 5155 9976 5164 10016
rect 5204 9976 5213 10016
rect 5155 9975 5213 9976
rect 5635 10016 5693 10017
rect 5635 9976 5644 10016
rect 5684 9976 5693 10016
rect 5635 9975 5693 9976
rect 6979 10016 7037 10017
rect 6979 9976 6988 10016
rect 7028 9976 7037 10016
rect 6979 9975 7037 9976
rect 7363 10016 7421 10017
rect 7363 9976 7372 10016
rect 7412 9976 7421 10016
rect 7363 9975 7421 9976
rect 8707 10016 8765 10017
rect 8707 9976 8716 10016
rect 8756 9976 8765 10016
rect 8707 9975 8765 9976
rect 9475 10016 9533 10017
rect 9475 9976 9484 10016
rect 9524 9976 9533 10016
rect 9475 9975 9533 9976
rect 10147 10016 10205 10017
rect 10147 9976 10156 10016
rect 10196 9976 10205 10016
rect 10147 9975 10205 9976
rect 11491 10016 11549 10017
rect 11491 9976 11500 10016
rect 11540 9976 11549 10016
rect 11491 9975 11549 9976
rect 12067 10016 12125 10017
rect 12067 9976 12076 10016
rect 12116 9976 12125 10016
rect 12067 9975 12125 9976
rect 13219 10016 13277 10017
rect 13219 9976 13228 10016
rect 13268 9976 13277 10016
rect 13219 9975 13277 9976
rect 13987 10016 14045 10017
rect 13987 9976 13996 10016
rect 14036 9976 14045 10016
rect 13987 9975 14045 9976
rect 14371 10016 14429 10017
rect 14371 9976 14380 10016
rect 14420 9976 14429 10016
rect 14371 9975 14429 9976
rect 14755 10016 14813 10017
rect 14755 9976 14764 10016
rect 14804 9976 14813 10016
rect 14755 9975 14813 9976
rect 15139 10016 15197 10017
rect 15139 9976 15148 10016
rect 15188 9976 15197 10016
rect 15139 9975 15197 9976
rect 576 9848 15360 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 15360 9848
rect 576 9784 15360 9808
rect 835 9680 893 9681
rect 835 9640 844 9680
rect 884 9640 893 9680
rect 835 9639 893 9640
rect 3235 9680 3293 9681
rect 3235 9640 3244 9680
rect 3284 9640 3293 9680
rect 3235 9639 3293 9640
rect 4387 9680 4445 9681
rect 4387 9640 4396 9680
rect 4436 9640 4445 9680
rect 4387 9639 4445 9640
rect 6211 9680 6269 9681
rect 6211 9640 6220 9680
rect 6260 9640 6269 9680
rect 6211 9639 6269 9640
rect 8515 9680 8573 9681
rect 8515 9640 8524 9680
rect 8564 9640 8573 9680
rect 8515 9639 8573 9640
rect 9283 9680 9341 9681
rect 9283 9640 9292 9680
rect 9332 9640 9341 9680
rect 9283 9639 9341 9640
rect 10819 9680 10877 9681
rect 10819 9640 10828 9680
rect 10868 9640 10877 9680
rect 10819 9639 10877 9640
rect 11011 9680 11069 9681
rect 11011 9640 11020 9680
rect 11060 9640 11069 9680
rect 11011 9639 11069 9640
rect 11971 9680 12029 9681
rect 11971 9640 11980 9680
rect 12020 9640 12029 9680
rect 11971 9639 12029 9640
rect 12739 9680 12797 9681
rect 12739 9640 12748 9680
rect 12788 9640 12797 9680
rect 12739 9639 12797 9640
rect 13603 9680 13661 9681
rect 13603 9640 13612 9680
rect 13652 9640 13661 9680
rect 13603 9639 13661 9640
rect 13987 9680 14045 9681
rect 13987 9640 13996 9680
rect 14036 9640 14045 9680
rect 13987 9639 14045 9640
rect 14371 9680 14429 9681
rect 14371 9640 14380 9680
rect 14420 9640 14429 9680
rect 14371 9639 14429 9640
rect 14755 9680 14813 9681
rect 14755 9640 14764 9680
rect 14804 9640 14813 9680
rect 14755 9639 14813 9640
rect 15139 9680 15197 9681
rect 15139 9640 15148 9680
rect 15188 9640 15197 9680
rect 15139 9639 15197 9640
rect 3531 9596 3573 9605
rect 3531 9556 3532 9596
rect 3572 9556 3573 9596
rect 3531 9547 3573 9556
rect 1315 9512 1373 9513
rect 1315 9472 1324 9512
rect 1364 9472 1373 9512
rect 1315 9471 1373 9472
rect 1411 9512 1469 9513
rect 1411 9472 1420 9512
rect 1460 9472 1469 9512
rect 1411 9471 1469 9472
rect 1891 9512 1949 9513
rect 1891 9472 1900 9512
rect 1940 9472 1949 9512
rect 1891 9471 1949 9472
rect 3723 9512 3765 9521
rect 3723 9472 3724 9512
rect 3764 9472 3765 9512
rect 3723 9463 3765 9472
rect 4683 9512 4725 9521
rect 4683 9472 4684 9512
rect 4724 9472 4725 9512
rect 4683 9463 4725 9472
rect 5155 9512 5213 9513
rect 5155 9472 5164 9512
rect 5204 9472 5213 9512
rect 5155 9471 5213 9472
rect 6691 9512 6749 9513
rect 6691 9472 6700 9512
rect 6740 9472 6749 9512
rect 6691 9471 6749 9472
rect 6787 9512 6845 9513
rect 6787 9472 6796 9512
rect 6836 9472 6845 9512
rect 6787 9471 6845 9472
rect 7171 9512 7229 9513
rect 7171 9472 7180 9512
rect 7220 9472 7229 9512
rect 7171 9471 7229 9472
rect 8811 9512 8853 9521
rect 8811 9472 8812 9512
rect 8852 9472 8853 9512
rect 8811 9463 8853 9472
rect 12267 9512 12309 9521
rect 12267 9472 12268 9512
rect 12308 9472 12309 9512
rect 12267 9463 12309 9472
rect 3531 9428 3573 9437
rect 3531 9388 3532 9428
rect 3572 9388 3573 9428
rect 3531 9379 3573 9388
rect 4779 9428 4821 9437
rect 4779 9388 4780 9428
rect 4820 9388 4821 9428
rect 4779 9379 4821 9388
rect 4875 9428 4917 9437
rect 4875 9388 4876 9428
rect 4916 9388 4917 9428
rect 4875 9379 4917 9388
rect 9003 9428 9045 9437
rect 9003 9388 9004 9428
rect 9044 9388 9045 9428
rect 9003 9379 9045 9388
rect 12459 9428 12501 9437
rect 12459 9388 12460 9428
rect 12500 9388 12501 9428
rect 12459 9379 12501 9388
rect 8907 9344 8949 9353
rect 8907 9304 8908 9344
rect 8948 9304 8949 9344
rect 8907 9295 8949 9304
rect 576 9092 15360 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 15360 9092
rect 576 9028 15360 9052
rect 1515 8840 1557 8849
rect 1515 8800 1516 8840
rect 1556 8800 1557 8840
rect 1515 8791 1557 8800
rect 7179 8840 7221 8849
rect 7179 8800 7180 8840
rect 7220 8800 7221 8840
rect 7179 8791 7221 8800
rect 1419 8756 1461 8765
rect 1419 8716 1420 8756
rect 1460 8716 1461 8756
rect 1419 8707 1461 8716
rect 7275 8756 7317 8765
rect 7275 8716 7276 8756
rect 7316 8716 7317 8756
rect 7275 8707 7317 8716
rect 10731 8756 10773 8765
rect 10731 8716 10732 8756
rect 10772 8716 10773 8756
rect 10731 8707 10773 8716
rect 1611 8672 1653 8681
rect 1611 8632 1612 8672
rect 1652 8632 1653 8672
rect 1611 8623 1653 8632
rect 2859 8672 2901 8681
rect 2859 8632 2860 8672
rect 2900 8632 2901 8672
rect 2859 8623 2901 8632
rect 2947 8672 3005 8673
rect 2947 8632 2956 8672
rect 2996 8632 3005 8672
rect 2947 8631 3005 8632
rect 3907 8672 3965 8673
rect 3907 8632 3916 8672
rect 3956 8632 3965 8672
rect 3907 8631 3965 8632
rect 5155 8672 5213 8673
rect 5155 8632 5164 8672
rect 5204 8632 5213 8672
rect 5155 8631 5213 8632
rect 5251 8672 5309 8673
rect 5251 8632 5260 8672
rect 5300 8632 5309 8672
rect 5251 8631 5309 8632
rect 7083 8672 7125 8681
rect 7083 8632 7084 8672
rect 7124 8632 7125 8672
rect 7083 8623 7125 8632
rect 8803 8672 8861 8673
rect 8803 8632 8812 8672
rect 8852 8632 8861 8672
rect 8803 8631 8861 8632
rect 8899 8672 8957 8673
rect 8899 8632 8908 8672
rect 8948 8632 8957 8672
rect 8899 8631 8957 8632
rect 9283 8672 9341 8673
rect 9283 8632 9292 8672
rect 9332 8632 9341 8672
rect 9283 8631 9341 8632
rect 10539 8672 10581 8681
rect 10539 8632 10540 8672
rect 10580 8632 10581 8672
rect 10539 8623 10581 8632
rect 1123 8504 1181 8505
rect 1123 8464 1132 8504
rect 1172 8464 1181 8504
rect 1123 8463 1181 8464
rect 2467 8504 2525 8505
rect 2467 8464 2476 8504
rect 2516 8464 2525 8504
rect 2467 8463 2525 8464
rect 3715 8504 3773 8505
rect 3715 8464 3724 8504
rect 3764 8464 3773 8504
rect 3715 8463 3773 8464
rect 5731 8504 5789 8505
rect 5731 8464 5740 8504
rect 5780 8464 5789 8504
rect 5731 8463 5789 8464
rect 6787 8504 6845 8505
rect 6787 8464 6796 8504
rect 6836 8464 6845 8504
rect 6787 8463 6845 8464
rect 8323 8504 8381 8505
rect 8323 8464 8332 8504
rect 8372 8464 8381 8504
rect 8323 8463 8381 8464
rect 10243 8504 10301 8505
rect 10243 8464 10252 8504
rect 10292 8464 10301 8504
rect 10243 8463 10301 8464
rect 11011 8504 11069 8505
rect 11011 8464 11020 8504
rect 11060 8464 11069 8504
rect 11011 8463 11069 8464
rect 12259 8504 12317 8505
rect 12259 8464 12268 8504
rect 12308 8464 12317 8504
rect 12259 8463 12317 8464
rect 12643 8504 12701 8505
rect 12643 8464 12652 8504
rect 12692 8464 12701 8504
rect 12643 8463 12701 8464
rect 13987 8504 14045 8505
rect 13987 8464 13996 8504
rect 14036 8464 14045 8504
rect 13987 8463 14045 8464
rect 14371 8504 14429 8505
rect 14371 8464 14380 8504
rect 14420 8464 14429 8504
rect 14371 8463 14429 8464
rect 14755 8504 14813 8505
rect 14755 8464 14764 8504
rect 14804 8464 14813 8504
rect 14755 8463 14813 8464
rect 15139 8504 15197 8505
rect 15139 8464 15148 8504
rect 15188 8464 15197 8504
rect 15139 8463 15197 8464
rect 576 8336 15360 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 15360 8336
rect 576 8272 15360 8296
rect 2563 8168 2621 8169
rect 2563 8128 2572 8168
rect 2612 8128 2621 8168
rect 2563 8127 2621 8128
rect 3427 8168 3485 8169
rect 3427 8128 3436 8168
rect 3476 8128 3485 8168
rect 3427 8127 3485 8128
rect 4195 8168 4253 8169
rect 4195 8128 4204 8168
rect 4244 8128 4253 8168
rect 4195 8127 4253 8128
rect 6019 8168 6077 8169
rect 6019 8128 6028 8168
rect 6068 8128 6077 8168
rect 6019 8127 6077 8128
rect 7747 8168 7805 8169
rect 7747 8128 7756 8168
rect 7796 8128 7805 8168
rect 7747 8127 7805 8128
rect 8515 8168 8573 8169
rect 8515 8128 8524 8168
rect 8564 8128 8573 8168
rect 8515 8127 8573 8128
rect 9283 8168 9341 8169
rect 9283 8128 9292 8168
rect 9332 8128 9341 8168
rect 9283 8127 9341 8128
rect 10435 8168 10493 8169
rect 10435 8128 10444 8168
rect 10484 8128 10493 8168
rect 10435 8127 10493 8128
rect 14371 8168 14429 8169
rect 14371 8128 14380 8168
rect 14420 8128 14429 8168
rect 14371 8127 14429 8128
rect 14755 8168 14813 8169
rect 14755 8128 14764 8168
rect 14804 8128 14813 8168
rect 14755 8127 14813 8128
rect 15139 8168 15197 8169
rect 15139 8128 15148 8168
rect 15188 8128 15197 8168
rect 15139 8127 15197 8128
rect 1131 8000 1173 8009
rect 1131 7960 1132 8000
rect 1172 7960 1173 8000
rect 1131 7951 1173 7960
rect 1219 8000 1277 8001
rect 1219 7960 1228 8000
rect 1268 7960 1277 8000
rect 1219 7959 1277 7960
rect 1795 8000 1853 8001
rect 1795 7960 1804 8000
rect 1844 7960 1853 8000
rect 1795 7959 1853 7960
rect 3915 8000 3957 8009
rect 3915 7960 3916 8000
rect 3956 7960 3957 8000
rect 3915 7951 3957 7960
rect 6499 8000 6557 8001
rect 6499 7960 6508 8000
rect 6548 7960 6557 8000
rect 6499 7959 6557 7960
rect 6595 8000 6653 8001
rect 6595 7960 6604 8000
rect 6644 7960 6653 8000
rect 6595 7959 6653 7960
rect 6979 8000 7037 8001
rect 6979 7960 6988 8000
rect 7028 7960 7037 8000
rect 6979 7959 7037 7960
rect 8811 8000 8853 8009
rect 8811 7960 8812 8000
rect 8852 7960 8853 8000
rect 8811 7951 8853 7960
rect 10731 8000 10773 8009
rect 10731 7960 10732 8000
rect 10772 7960 10773 8000
rect 10731 7951 10773 7960
rect 12363 8000 12405 8009
rect 12363 7960 12364 8000
rect 12404 7960 12405 8000
rect 12363 7951 12405 7960
rect 3723 7916 3765 7925
rect 3723 7876 3724 7916
rect 3764 7876 3765 7916
rect 3723 7867 3765 7876
rect 9003 7916 9045 7925
rect 9003 7876 9004 7916
rect 9044 7876 9045 7916
rect 9003 7867 9045 7876
rect 10923 7916 10965 7925
rect 10923 7876 10924 7916
rect 10964 7876 10965 7916
rect 10923 7867 10965 7876
rect 12555 7916 12597 7925
rect 12555 7876 12556 7916
rect 12596 7876 12597 7916
rect 12555 7867 12597 7876
rect 8907 7832 8949 7841
rect 8907 7792 8908 7832
rect 8948 7792 8949 7832
rect 8907 7783 8949 7792
rect 3915 7748 3957 7757
rect 3915 7708 3916 7748
rect 3956 7708 3957 7748
rect 3915 7699 3957 7708
rect 576 7580 15360 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 15360 7580
rect 576 7516 15360 7540
rect 1515 7412 1557 7421
rect 1515 7372 1516 7412
rect 1556 7372 1557 7412
rect 1515 7363 1557 7372
rect 6987 7412 7029 7421
rect 6987 7372 6988 7412
rect 7028 7372 7029 7412
rect 6987 7363 7029 7372
rect 1707 7244 1749 7253
rect 1707 7204 1708 7244
rect 1748 7204 1749 7244
rect 1707 7195 1749 7204
rect 5355 7244 5397 7253
rect 5355 7204 5356 7244
rect 5396 7204 5397 7244
rect 5355 7195 5397 7204
rect 7179 7244 7221 7253
rect 7179 7204 7180 7244
rect 7220 7204 7221 7244
rect 7179 7195 7221 7204
rect 10923 7244 10965 7253
rect 10923 7204 10924 7244
rect 10964 7204 10965 7244
rect 10923 7195 10965 7204
rect 12555 7244 12597 7253
rect 12555 7204 12556 7244
rect 12596 7204 12597 7244
rect 12555 7195 12597 7204
rect 1515 7160 1557 7169
rect 1515 7120 1516 7160
rect 1556 7120 1557 7160
rect 1515 7111 1557 7120
rect 2859 7160 2901 7169
rect 2859 7120 2860 7160
rect 2900 7120 2901 7160
rect 2859 7111 2901 7120
rect 2947 7160 3005 7161
rect 2947 7120 2956 7160
rect 2996 7120 3005 7160
rect 2947 7119 3005 7120
rect 3715 7160 3773 7161
rect 3715 7120 3724 7160
rect 3764 7120 3773 7160
rect 3715 7119 3773 7120
rect 5547 7160 5589 7169
rect 5547 7120 5548 7160
rect 5588 7120 5589 7160
rect 5547 7111 5589 7120
rect 6987 7160 7029 7169
rect 6987 7120 6988 7160
rect 7028 7120 7029 7160
rect 6987 7111 7029 7120
rect 8803 7160 8861 7161
rect 8803 7120 8812 7160
rect 8852 7120 8861 7160
rect 8803 7119 8861 7120
rect 8899 7160 8957 7161
rect 8899 7120 8908 7160
rect 8948 7120 8957 7160
rect 8899 7119 8957 7120
rect 9283 7160 9341 7161
rect 9283 7120 9292 7160
rect 9332 7120 9341 7160
rect 9283 7119 9341 7120
rect 10731 7160 10773 7169
rect 10731 7120 10732 7160
rect 10772 7120 10773 7160
rect 10731 7111 10773 7120
rect 12363 7160 12405 7169
rect 12363 7120 12364 7160
rect 12404 7120 12405 7160
rect 12363 7111 12405 7120
rect 5355 7076 5397 7085
rect 5355 7036 5356 7076
rect 5396 7036 5397 7076
rect 5355 7027 5397 7036
rect 835 6992 893 6993
rect 835 6952 844 6992
rect 884 6952 893 6992
rect 835 6951 893 6952
rect 1219 6992 1277 6993
rect 1219 6952 1228 6992
rect 1268 6952 1277 6992
rect 1219 6951 1277 6952
rect 2467 6992 2525 6993
rect 2467 6952 2476 6992
rect 2516 6952 2525 6992
rect 2467 6951 2525 6952
rect 4675 6992 4733 6993
rect 4675 6952 4684 6992
rect 4724 6952 4733 6992
rect 4675 6951 4733 6952
rect 5059 6992 5117 6993
rect 5059 6952 5068 6992
rect 5108 6952 5117 6992
rect 5059 6951 5117 6952
rect 7459 6992 7517 6993
rect 7459 6952 7468 6992
rect 7508 6952 7517 6992
rect 7459 6951 7517 6952
rect 8323 6992 8381 6993
rect 8323 6952 8332 6992
rect 8372 6952 8381 6992
rect 8323 6951 8381 6952
rect 10435 6992 10493 6993
rect 10435 6952 10444 6992
rect 10484 6952 10493 6992
rect 10435 6951 10493 6952
rect 11203 6992 11261 6993
rect 11203 6952 11212 6992
rect 11252 6952 11261 6992
rect 11203 6951 11261 6952
rect 12835 6992 12893 6993
rect 12835 6952 12844 6992
rect 12884 6952 12893 6992
rect 12835 6951 12893 6952
rect 13219 6992 13277 6993
rect 13219 6952 13228 6992
rect 13268 6952 13277 6992
rect 13219 6951 13277 6952
rect 13795 6992 13853 6993
rect 13795 6952 13804 6992
rect 13844 6952 13853 6992
rect 13795 6951 13853 6952
rect 14179 6992 14237 6993
rect 14179 6952 14188 6992
rect 14228 6952 14237 6992
rect 14179 6951 14237 6952
rect 14755 6992 14813 6993
rect 14755 6952 14764 6992
rect 14804 6952 14813 6992
rect 14755 6951 14813 6952
rect 15139 6992 15197 6993
rect 15139 6952 15148 6992
rect 15188 6952 15197 6992
rect 15139 6951 15197 6952
rect 576 6824 15360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 15360 6824
rect 576 6760 15360 6784
rect 2371 6656 2429 6657
rect 2371 6616 2380 6656
rect 2420 6616 2429 6656
rect 2371 6615 2429 6616
rect 4579 6656 4637 6657
rect 4579 6616 4588 6656
rect 4628 6616 4637 6656
rect 4579 6615 4637 6616
rect 7843 6656 7901 6657
rect 7843 6616 7852 6656
rect 7892 6616 7901 6656
rect 7843 6615 7901 6616
rect 10147 6656 10205 6657
rect 10147 6616 10156 6656
rect 10196 6616 10205 6656
rect 10147 6615 10205 6616
rect 10915 6656 10973 6657
rect 10915 6616 10924 6656
rect 10964 6616 10973 6656
rect 10915 6615 10973 6616
rect 11875 6656 11933 6657
rect 11875 6616 11884 6656
rect 11924 6616 11933 6656
rect 11875 6615 11933 6616
rect 12643 6656 12701 6657
rect 12643 6616 12652 6656
rect 12692 6616 12701 6656
rect 12643 6615 12701 6616
rect 13507 6656 13565 6657
rect 13507 6616 13516 6656
rect 13556 6616 13565 6656
rect 13507 6615 13565 6616
rect 14371 6656 14429 6657
rect 14371 6616 14380 6656
rect 14420 6616 14429 6656
rect 14371 6615 14429 6616
rect 14755 6656 14813 6657
rect 14755 6616 14764 6656
rect 14804 6616 14813 6656
rect 14755 6615 14813 6616
rect 15139 6656 15197 6657
rect 15139 6616 15148 6656
rect 15188 6616 15197 6656
rect 15139 6615 15197 6616
rect 6795 6572 6837 6581
rect 6795 6532 6796 6572
rect 6836 6532 6837 6572
rect 6795 6523 6837 6532
rect 1035 6488 1077 6497
rect 1035 6448 1036 6488
rect 1076 6448 1077 6488
rect 1035 6439 1077 6448
rect 1123 6488 1181 6489
rect 1123 6448 1132 6488
rect 1172 6448 1181 6488
rect 1123 6447 1181 6448
rect 1603 6488 1661 6489
rect 1603 6448 1612 6488
rect 1652 6448 1661 6488
rect 1603 6447 1661 6448
rect 3627 6488 3669 6497
rect 3627 6448 3628 6488
rect 3668 6448 3669 6488
rect 3627 6439 3669 6448
rect 3723 6488 3765 6497
rect 3723 6448 3724 6488
rect 3764 6448 3765 6488
rect 3723 6439 3765 6448
rect 5059 6488 5117 6489
rect 5059 6448 5068 6488
rect 5108 6448 5117 6488
rect 5059 6447 5117 6448
rect 5155 6488 5213 6489
rect 5155 6448 5164 6488
rect 5204 6448 5213 6488
rect 5155 6447 5213 6448
rect 5539 6488 5597 6489
rect 5539 6448 5548 6488
rect 5588 6448 5597 6488
rect 5539 6447 5597 6448
rect 6603 6488 6645 6497
rect 6603 6448 6604 6488
rect 6644 6448 6645 6488
rect 6603 6439 6645 6448
rect 7267 6488 7325 6489
rect 7267 6448 7276 6488
rect 7316 6448 7325 6488
rect 7267 6447 7325 6448
rect 7363 6488 7421 6489
rect 7363 6448 7372 6488
rect 7412 6448 7421 6488
rect 7363 6447 7421 6448
rect 8323 6488 8381 6489
rect 8323 6448 8332 6488
rect 8372 6448 8381 6488
rect 8323 6447 8381 6448
rect 10443 6488 10485 6497
rect 10443 6448 10444 6488
rect 10484 6448 10485 6488
rect 10443 6439 10485 6448
rect 12171 6488 12213 6497
rect 12171 6448 12172 6488
rect 12212 6448 12213 6488
rect 12171 6439 12213 6448
rect 3819 6404 3861 6413
rect 3819 6364 3820 6404
rect 3860 6364 3861 6404
rect 3819 6355 3861 6364
rect 6795 6404 6837 6413
rect 6795 6364 6796 6404
rect 6836 6364 6837 6404
rect 6795 6355 6837 6364
rect 10635 6404 10677 6413
rect 10635 6364 10636 6404
rect 10676 6364 10677 6404
rect 10635 6355 10677 6364
rect 12363 6404 12405 6413
rect 12363 6364 12364 6404
rect 12404 6364 12405 6404
rect 12363 6355 12405 6364
rect 576 6068 15360 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 15360 6068
rect 576 6004 15360 6028
rect 1419 5900 1461 5909
rect 1419 5860 1420 5900
rect 1460 5860 1461 5900
rect 1419 5851 1461 5860
rect 8035 5816 8093 5817
rect 8035 5776 8044 5816
rect 8084 5776 8093 5816
rect 8035 5775 8093 5776
rect 1611 5732 1653 5741
rect 1611 5692 1612 5732
rect 1652 5692 1653 5732
rect 1611 5683 1653 5692
rect 8235 5732 8277 5741
rect 8235 5692 8236 5732
rect 8276 5692 8277 5732
rect 8235 5683 8277 5692
rect 10635 5732 10677 5741
rect 10635 5692 10636 5732
rect 10676 5692 10677 5732
rect 10635 5683 10677 5692
rect 12555 5732 12597 5741
rect 12555 5692 12556 5732
rect 12596 5692 12597 5732
rect 12555 5683 12597 5692
rect 1419 5648 1461 5657
rect 1419 5608 1420 5648
rect 1460 5608 1461 5648
rect 1419 5599 1461 5608
rect 2859 5648 2901 5657
rect 2859 5608 2860 5648
rect 2900 5608 2901 5648
rect 2859 5599 2901 5608
rect 2947 5648 3005 5649
rect 2947 5608 2956 5648
rect 2996 5608 3005 5648
rect 2947 5607 3005 5608
rect 3811 5648 3869 5649
rect 3811 5608 3820 5648
rect 3860 5608 3869 5648
rect 3811 5607 3869 5608
rect 6211 5648 6269 5649
rect 6211 5608 6220 5648
rect 6260 5608 6269 5648
rect 6211 5607 6269 5608
rect 8043 5648 8085 5657
rect 8043 5608 8044 5648
rect 8084 5608 8085 5648
rect 8043 5599 8085 5608
rect 8515 5648 8573 5649
rect 8515 5608 8524 5648
rect 8564 5608 8573 5648
rect 8515 5607 8573 5608
rect 10443 5648 10485 5657
rect 10443 5608 10444 5648
rect 10484 5608 10485 5648
rect 10443 5599 10485 5608
rect 12363 5648 12405 5657
rect 12363 5608 12364 5648
rect 12404 5608 12405 5648
rect 12363 5599 12405 5608
rect 1123 5480 1181 5481
rect 1123 5440 1132 5480
rect 1172 5440 1181 5480
rect 1123 5439 1181 5440
rect 2467 5480 2525 5481
rect 2467 5440 2476 5480
rect 2516 5440 2525 5480
rect 2467 5439 2525 5440
rect 3619 5480 3677 5481
rect 3619 5440 3628 5480
rect 3668 5440 3677 5480
rect 3619 5439 3677 5440
rect 4579 5480 4637 5481
rect 4579 5440 4588 5480
rect 4628 5440 4637 5480
rect 4579 5439 4637 5440
rect 5251 5480 5309 5481
rect 5251 5440 5260 5480
rect 5300 5440 5309 5480
rect 5251 5439 5309 5440
rect 5635 5480 5693 5481
rect 5635 5440 5644 5480
rect 5684 5440 5693 5480
rect 5635 5439 5693 5440
rect 6019 5480 6077 5481
rect 6019 5440 6028 5480
rect 6068 5440 6077 5480
rect 6019 5439 6077 5440
rect 7075 5480 7133 5481
rect 7075 5440 7084 5480
rect 7124 5440 7133 5480
rect 7075 5439 7133 5440
rect 7459 5480 7517 5481
rect 7459 5440 7468 5480
rect 7508 5440 7517 5480
rect 7459 5439 7517 5440
rect 9283 5480 9341 5481
rect 9283 5440 9292 5480
rect 9332 5440 9341 5480
rect 9283 5439 9341 5440
rect 10147 5480 10205 5481
rect 10147 5440 10156 5480
rect 10196 5440 10205 5480
rect 10147 5439 10205 5440
rect 10915 5480 10973 5481
rect 10915 5440 10924 5480
rect 10964 5440 10973 5480
rect 10915 5439 10973 5440
rect 12067 5480 12125 5481
rect 12067 5440 12076 5480
rect 12116 5440 12125 5480
rect 12067 5439 12125 5440
rect 12835 5480 12893 5481
rect 12835 5440 12844 5480
rect 12884 5440 12893 5480
rect 12835 5439 12893 5440
rect 13987 5480 14045 5481
rect 13987 5440 13996 5480
rect 14036 5440 14045 5480
rect 13987 5439 14045 5440
rect 14371 5480 14429 5481
rect 14371 5440 14380 5480
rect 14420 5440 14429 5480
rect 14371 5439 14429 5440
rect 14755 5480 14813 5481
rect 14755 5440 14764 5480
rect 14804 5440 14813 5480
rect 14755 5439 14813 5440
rect 15139 5480 15197 5481
rect 15139 5440 15148 5480
rect 15188 5440 15197 5480
rect 15139 5439 15197 5440
rect 576 5312 15360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 15360 5312
rect 576 5248 15360 5272
rect 2563 5144 2621 5145
rect 2563 5104 2572 5144
rect 2612 5104 2621 5144
rect 2563 5103 2621 5104
rect 4291 5144 4349 5145
rect 4291 5104 4300 5144
rect 4340 5104 4349 5144
rect 4291 5103 4349 5104
rect 8035 5144 8093 5145
rect 8035 5104 8044 5144
rect 8084 5104 8093 5144
rect 8035 5103 8093 5104
rect 8419 5144 8477 5145
rect 8419 5104 8428 5144
rect 8468 5104 8477 5144
rect 8419 5103 8477 5104
rect 10051 5144 10109 5145
rect 10051 5104 10060 5144
rect 10100 5104 10109 5144
rect 10051 5103 10109 5104
rect 11011 5144 11069 5145
rect 11011 5104 11020 5144
rect 11060 5104 11069 5144
rect 11011 5103 11069 5104
rect 11203 5144 11261 5145
rect 11203 5104 11212 5144
rect 11252 5104 11261 5144
rect 11203 5103 11261 5104
rect 13987 5144 14045 5145
rect 13987 5104 13996 5144
rect 14036 5104 14045 5144
rect 13987 5103 14045 5104
rect 14371 5144 14429 5145
rect 14371 5104 14380 5144
rect 14420 5104 14429 5144
rect 14371 5103 14429 5104
rect 14755 5144 14813 5145
rect 14755 5104 14764 5144
rect 14804 5104 14813 5144
rect 14755 5103 14813 5104
rect 15139 5144 15197 5145
rect 15139 5104 15148 5144
rect 15188 5104 15197 5144
rect 15139 5103 15197 5104
rect 6123 5060 6165 5069
rect 6123 5020 6124 5060
rect 6164 5020 6165 5060
rect 6123 5011 6165 5020
rect 1131 4976 1173 4985
rect 1131 4936 1132 4976
rect 1172 4936 1173 4976
rect 1131 4927 1173 4936
rect 1219 4976 1277 4977
rect 1219 4936 1228 4976
rect 1268 4936 1277 4976
rect 1219 4935 1277 4936
rect 1795 4976 1853 4977
rect 1795 4936 1804 4976
rect 1844 4936 1853 4976
rect 1795 4935 1853 4936
rect 3915 4976 3957 4985
rect 3915 4936 3916 4976
rect 3956 4936 3957 4976
rect 3915 4927 3957 4936
rect 4011 4976 4053 4985
rect 4011 4936 4012 4976
rect 4052 4936 4053 4976
rect 4011 4927 4053 4936
rect 5347 4976 5405 4977
rect 5347 4936 5356 4976
rect 5396 4936 5405 4976
rect 5347 4935 5405 4936
rect 5443 4976 5501 4977
rect 5443 4936 5452 4976
rect 5492 4936 5501 4976
rect 5443 4935 5501 4936
rect 5931 4976 5973 4985
rect 5931 4936 5932 4976
rect 5972 4936 5973 4976
rect 5931 4927 5973 4936
rect 7267 4976 7325 4977
rect 7267 4936 7276 4976
rect 7316 4936 7325 4976
rect 7267 4935 7325 4936
rect 7363 4976 7421 4977
rect 7363 4936 7372 4976
rect 7412 4936 7421 4976
rect 7363 4935 7421 4936
rect 3819 4892 3861 4901
rect 3819 4852 3820 4892
rect 3860 4852 3861 4892
rect 3819 4843 3861 4852
rect 6123 4892 6165 4901
rect 6123 4852 6124 4892
rect 6164 4852 6165 4892
rect 6123 4843 6165 4852
rect 576 4556 15360 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 15360 4556
rect 576 4492 15360 4516
rect 1803 4304 1845 4313
rect 1803 4264 1804 4304
rect 1844 4264 1845 4304
rect 1803 4255 1845 4264
rect 1899 4220 1941 4229
rect 1899 4180 1900 4220
rect 1940 4180 1941 4220
rect 1899 4171 1941 4180
rect 9387 4220 9429 4229
rect 9387 4180 9388 4220
rect 9428 4180 9429 4220
rect 9387 4171 9429 4180
rect 10059 4220 10101 4229
rect 10059 4180 10060 4220
rect 10100 4180 10101 4220
rect 10059 4171 10101 4180
rect 11211 4220 11253 4229
rect 11211 4180 11212 4220
rect 11252 4180 11253 4220
rect 11211 4171 11253 4180
rect 12555 4220 12597 4229
rect 12555 4180 12556 4220
rect 12596 4180 12597 4220
rect 12555 4171 12597 4180
rect 1707 4136 1749 4145
rect 1707 4096 1708 4136
rect 1748 4096 1749 4136
rect 1707 4087 1749 4096
rect 2955 4136 2997 4145
rect 2955 4096 2956 4136
rect 2996 4096 2997 4136
rect 2955 4087 2997 4096
rect 3043 4136 3101 4137
rect 3043 4096 3052 4136
rect 3092 4096 3101 4136
rect 3043 4095 3101 4096
rect 3811 4136 3869 4137
rect 3811 4096 3820 4136
rect 3860 4096 3869 4136
rect 3811 4095 3869 4096
rect 6987 4136 7029 4145
rect 6987 4096 6988 4136
rect 7028 4096 7029 4136
rect 6987 4087 7029 4096
rect 7075 4136 7133 4137
rect 7075 4096 7084 4136
rect 7124 4096 7133 4136
rect 7075 4095 7133 4096
rect 7651 4136 7709 4137
rect 7651 4096 7660 4136
rect 7700 4096 7709 4136
rect 7651 4095 7709 4096
rect 9195 4136 9237 4145
rect 9195 4096 9196 4136
rect 9236 4096 9237 4136
rect 9195 4087 9237 4096
rect 10251 4136 10293 4145
rect 10251 4096 10252 4136
rect 10292 4096 10293 4136
rect 10251 4087 10293 4096
rect 11019 4136 11061 4145
rect 11019 4096 11020 4136
rect 11060 4096 11061 4136
rect 11019 4087 11061 4096
rect 12363 4136 12405 4145
rect 12363 4096 12364 4136
rect 12404 4096 12405 4136
rect 12363 4087 12405 4096
rect 1027 3968 1085 3969
rect 1027 3928 1036 3968
rect 1076 3928 1085 3968
rect 1027 3927 1085 3928
rect 1411 3968 1469 3969
rect 1411 3928 1420 3968
rect 1460 3928 1469 3968
rect 1411 3927 1469 3928
rect 2563 3968 2621 3969
rect 2563 3928 2572 3968
rect 2612 3928 2621 3968
rect 2563 3927 2621 3928
rect 4579 3968 4637 3969
rect 4579 3928 4588 3968
rect 4628 3928 4637 3968
rect 4579 3927 4637 3928
rect 5347 3968 5405 3969
rect 5347 3928 5356 3968
rect 5396 3928 5405 3968
rect 5347 3927 5405 3928
rect 5539 3968 5597 3969
rect 5539 3928 5548 3968
rect 5588 3928 5597 3968
rect 5539 3927 5597 3928
rect 6595 3968 6653 3969
rect 6595 3928 6604 3968
rect 6644 3928 6653 3968
rect 6595 3927 6653 3928
rect 8899 3968 8957 3969
rect 8899 3928 8908 3968
rect 8948 3928 8957 3968
rect 8899 3927 8957 3928
rect 10531 3968 10589 3969
rect 10531 3928 10540 3968
rect 10580 3928 10589 3968
rect 10531 3927 10589 3928
rect 12067 3968 12125 3969
rect 12067 3928 12076 3968
rect 12116 3928 12125 3968
rect 12067 3927 12125 3928
rect 12835 3968 12893 3969
rect 12835 3928 12844 3968
rect 12884 3928 12893 3968
rect 12835 3927 12893 3928
rect 13987 3968 14045 3969
rect 13987 3928 13996 3968
rect 14036 3928 14045 3968
rect 13987 3927 14045 3928
rect 14371 3968 14429 3969
rect 14371 3928 14380 3968
rect 14420 3928 14429 3968
rect 14371 3927 14429 3928
rect 14755 3968 14813 3969
rect 14755 3928 14764 3968
rect 14804 3928 14813 3968
rect 14755 3927 14813 3928
rect 15139 3968 15197 3969
rect 15139 3928 15148 3968
rect 15188 3928 15197 3968
rect 15139 3927 15197 3928
rect 576 3800 15360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 15360 3800
rect 576 3736 15360 3760
rect 835 3632 893 3633
rect 835 3592 844 3632
rect 884 3592 893 3632
rect 835 3591 893 3592
rect 3139 3632 3197 3633
rect 3139 3592 3148 3632
rect 3188 3592 3197 3632
rect 3139 3591 3197 3592
rect 3523 3632 3581 3633
rect 3523 3592 3532 3632
rect 3572 3592 3581 3632
rect 3523 3591 3581 3592
rect 4771 3632 4829 3633
rect 4771 3592 4780 3632
rect 4820 3592 4829 3632
rect 4771 3591 4829 3592
rect 7459 3632 7517 3633
rect 7459 3592 7468 3632
rect 7508 3592 7517 3632
rect 7459 3591 7517 3592
rect 9475 3632 9533 3633
rect 9475 3592 9484 3632
rect 9524 3592 9533 3632
rect 9475 3591 9533 3592
rect 10435 3632 10493 3633
rect 10435 3592 10444 3632
rect 10484 3592 10493 3632
rect 10435 3591 10493 3592
rect 11203 3632 11261 3633
rect 11203 3592 11212 3632
rect 11252 3592 11261 3632
rect 11203 3591 11261 3592
rect 12355 3632 12413 3633
rect 12355 3592 12364 3632
rect 12404 3592 12413 3632
rect 12355 3591 12413 3592
rect 12739 3632 12797 3633
rect 12739 3592 12748 3632
rect 12788 3592 12797 3632
rect 12739 3591 12797 3592
rect 13603 3632 13661 3633
rect 13603 3592 13612 3632
rect 13652 3592 13661 3632
rect 13603 3591 13661 3592
rect 13987 3632 14045 3633
rect 13987 3592 13996 3632
rect 14036 3592 14045 3632
rect 13987 3591 14045 3592
rect 14371 3632 14429 3633
rect 14371 3592 14380 3632
rect 14420 3592 14429 3632
rect 14371 3591 14429 3592
rect 14755 3632 14813 3633
rect 14755 3592 14764 3632
rect 14804 3592 14813 3632
rect 14755 3591 14813 3592
rect 15139 3632 15197 3633
rect 15139 3592 15148 3632
rect 15188 3592 15197 3632
rect 15139 3591 15197 3592
rect 3819 3548 3861 3557
rect 3819 3508 3820 3548
rect 3860 3508 3861 3548
rect 3819 3499 3861 3508
rect 1227 3464 1269 3473
rect 1227 3424 1228 3464
rect 1268 3424 1269 3464
rect 1227 3415 1269 3424
rect 1323 3464 1365 3473
rect 1323 3424 1324 3464
rect 1364 3424 1365 3464
rect 1323 3415 1365 3424
rect 1603 3464 1661 3465
rect 1603 3424 1612 3464
rect 1652 3424 1661 3464
rect 1603 3423 1661 3424
rect 4011 3464 4053 3473
rect 4011 3424 4012 3464
rect 4052 3424 4053 3464
rect 4011 3415 4053 3424
rect 5155 3464 5213 3465
rect 5155 3424 5164 3464
rect 5204 3424 5213 3464
rect 5155 3423 5213 3424
rect 5251 3464 5309 3465
rect 5251 3424 5260 3464
rect 5300 3424 5309 3464
rect 5251 3423 5309 3424
rect 5355 3464 5397 3473
rect 5355 3424 5356 3464
rect 5396 3424 5397 3464
rect 5355 3415 5397 3424
rect 5731 3464 5789 3465
rect 5731 3424 5740 3464
rect 5780 3424 5789 3464
rect 5731 3423 5789 3424
rect 7755 3464 7797 3473
rect 7755 3424 7756 3464
rect 7796 3424 7797 3464
rect 7755 3415 7797 3424
rect 7851 3464 7893 3473
rect 7851 3424 7852 3464
rect 7892 3424 7893 3464
rect 7851 3415 7893 3424
rect 10731 3464 10773 3473
rect 10731 3424 10732 3464
rect 10772 3424 10773 3464
rect 10731 3415 10773 3424
rect 1131 3380 1173 3389
rect 1131 3340 1132 3380
rect 1172 3340 1173 3380
rect 1131 3331 1173 3340
rect 3819 3380 3861 3389
rect 3819 3340 3820 3380
rect 3860 3340 3861 3380
rect 3819 3331 3861 3340
rect 7947 3380 7989 3389
rect 7947 3340 7948 3380
rect 7988 3340 7989 3380
rect 7947 3331 7989 3340
rect 10923 3380 10965 3389
rect 10923 3340 10924 3380
rect 10964 3340 10965 3380
rect 10923 3331 10965 3340
rect 576 3044 15360 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 15360 3044
rect 576 2980 15360 3004
rect 5451 2792 5493 2801
rect 5451 2752 5452 2792
rect 5492 2752 5493 2792
rect 5451 2743 5493 2752
rect 5355 2708 5397 2717
rect 5355 2668 5356 2708
rect 5396 2668 5397 2708
rect 5355 2659 5397 2668
rect 9291 2708 9333 2717
rect 9291 2668 9292 2708
rect 9332 2668 9333 2708
rect 9291 2659 9333 2668
rect 10827 2708 10869 2717
rect 10827 2668 10828 2708
rect 10868 2668 10869 2708
rect 10827 2659 10869 2668
rect 12651 2708 12693 2717
rect 12651 2668 12652 2708
rect 12692 2668 12693 2708
rect 12651 2659 12693 2668
rect 1219 2624 1277 2625
rect 1219 2584 1228 2624
rect 1268 2584 1277 2624
rect 1219 2583 1277 2584
rect 1315 2624 1373 2625
rect 1315 2584 1324 2624
rect 1364 2584 1373 2624
rect 1315 2583 1373 2584
rect 3139 2624 3197 2625
rect 3139 2584 3148 2624
rect 3188 2584 3197 2624
rect 3139 2583 3197 2584
rect 3235 2624 3293 2625
rect 3235 2584 3244 2624
rect 3284 2584 3293 2624
rect 3235 2583 3293 2584
rect 3715 2624 3773 2625
rect 3715 2584 3724 2624
rect 3764 2584 3773 2624
rect 3715 2583 3773 2584
rect 5547 2624 5589 2633
rect 5547 2584 5548 2624
rect 5588 2584 5589 2624
rect 5547 2575 5589 2584
rect 6411 2624 6453 2633
rect 6411 2584 6412 2624
rect 6452 2584 6453 2624
rect 6411 2575 6453 2584
rect 6499 2624 6557 2625
rect 6499 2584 6508 2624
rect 6548 2584 6557 2624
rect 6499 2583 6557 2584
rect 7363 2624 7421 2625
rect 7363 2584 7372 2624
rect 7412 2584 7421 2624
rect 7363 2583 7421 2584
rect 9099 2624 9141 2633
rect 9099 2584 9100 2624
rect 9140 2584 9141 2624
rect 9099 2575 9141 2584
rect 10635 2624 10677 2633
rect 10635 2584 10636 2624
rect 10676 2584 10677 2624
rect 10635 2575 10677 2584
rect 12459 2624 12501 2633
rect 12459 2584 12460 2624
rect 12500 2584 12501 2624
rect 12459 2575 12501 2584
rect 835 2456 893 2457
rect 835 2416 844 2456
rect 884 2416 893 2456
rect 835 2415 893 2416
rect 1795 2456 1853 2457
rect 1795 2416 1804 2456
rect 1844 2416 1853 2456
rect 1795 2415 1853 2416
rect 2659 2456 2717 2457
rect 2659 2416 2668 2456
rect 2708 2416 2717 2456
rect 2659 2415 2717 2416
rect 4867 2456 4925 2457
rect 4867 2416 4876 2456
rect 4916 2416 4925 2456
rect 4867 2415 4925 2416
rect 6019 2456 6077 2457
rect 6019 2416 6028 2456
rect 6068 2416 6077 2456
rect 6019 2415 6077 2416
rect 7171 2456 7229 2457
rect 7171 2416 7180 2456
rect 7220 2416 7229 2456
rect 7171 2415 7229 2416
rect 8131 2456 8189 2457
rect 8131 2416 8140 2456
rect 8180 2416 8189 2456
rect 8131 2415 8189 2416
rect 8803 2456 8861 2457
rect 8803 2416 8812 2456
rect 8852 2416 8861 2456
rect 8803 2415 8861 2416
rect 9571 2456 9629 2457
rect 9571 2416 9580 2456
rect 9620 2416 9629 2456
rect 9571 2415 9629 2416
rect 10339 2456 10397 2457
rect 10339 2416 10348 2456
rect 10388 2416 10397 2456
rect 10339 2415 10397 2416
rect 13795 2456 13853 2457
rect 13795 2416 13804 2456
rect 13844 2416 13853 2456
rect 13795 2415 13853 2416
rect 14179 2456 14237 2457
rect 14179 2416 14188 2456
rect 14228 2416 14237 2456
rect 14179 2415 14237 2416
rect 14563 2456 14621 2457
rect 14563 2416 14572 2456
rect 14612 2416 14621 2456
rect 14563 2415 14621 2416
rect 14947 2456 15005 2457
rect 14947 2416 14956 2456
rect 14996 2416 15005 2456
rect 14947 2415 15005 2416
rect 576 2288 15360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 15360 2288
rect 576 2224 15360 2248
rect 835 2120 893 2121
rect 835 2080 844 2120
rect 884 2080 893 2120
rect 835 2079 893 2080
rect 2851 2120 2909 2121
rect 2851 2080 2860 2120
rect 2900 2080 2909 2120
rect 2851 2079 2909 2080
rect 3235 2120 3293 2121
rect 3235 2080 3244 2120
rect 3284 2080 3293 2120
rect 3235 2079 3293 2080
rect 5827 2120 5885 2121
rect 5827 2080 5836 2120
rect 5876 2080 5885 2120
rect 5827 2079 5885 2080
rect 6211 2120 6269 2121
rect 6211 2080 6220 2120
rect 6260 2080 6269 2120
rect 6211 2079 6269 2080
rect 8227 2120 8285 2121
rect 8227 2080 8236 2120
rect 8276 2080 8285 2120
rect 8227 2079 8285 2080
rect 8899 2120 8957 2121
rect 8899 2080 8908 2120
rect 8948 2080 8957 2120
rect 8899 2079 8957 2080
rect 10819 2120 10877 2121
rect 10819 2080 10828 2120
rect 10868 2080 10877 2120
rect 10819 2079 10877 2080
rect 11011 2120 11069 2121
rect 11011 2080 11020 2120
rect 11060 2080 11069 2120
rect 11011 2079 11069 2080
rect 11395 2120 11453 2121
rect 11395 2080 11404 2120
rect 11444 2080 11453 2120
rect 11395 2079 11453 2080
rect 11971 2120 12029 2121
rect 11971 2080 11980 2120
rect 12020 2080 12029 2120
rect 11971 2079 12029 2080
rect 13123 2120 13181 2121
rect 13123 2080 13132 2120
rect 13172 2080 13181 2120
rect 13123 2079 13181 2080
rect 13987 2120 14045 2121
rect 13987 2080 13996 2120
rect 14036 2080 14045 2120
rect 13987 2079 14045 2080
rect 14371 2120 14429 2121
rect 14371 2080 14380 2120
rect 14420 2080 14429 2120
rect 14371 2079 14429 2080
rect 14755 2120 14813 2121
rect 14755 2080 14764 2120
rect 14804 2080 14813 2120
rect 14755 2079 14813 2080
rect 15139 2120 15197 2121
rect 15139 2080 15148 2120
rect 15188 2080 15197 2120
rect 15139 2079 15197 2080
rect 1323 1952 1365 1961
rect 1323 1912 1324 1952
rect 1364 1912 1365 1952
rect 1323 1903 1365 1912
rect 1603 1952 1661 1953
rect 1603 1912 1612 1952
rect 1652 1912 1661 1952
rect 1603 1911 1661 1912
rect 3627 1952 3669 1961
rect 3627 1912 3628 1952
rect 3668 1912 3669 1952
rect 3627 1903 3669 1912
rect 3723 1952 3765 1961
rect 3723 1912 3724 1952
rect 3764 1912 3765 1952
rect 3723 1903 3765 1912
rect 4483 1952 4541 1953
rect 4483 1912 4492 1952
rect 4532 1912 4541 1952
rect 4483 1911 4541 1912
rect 4579 1952 4637 1953
rect 4579 1912 4588 1952
rect 4628 1912 4637 1952
rect 4579 1911 4637 1912
rect 5059 1952 5117 1953
rect 5059 1912 5068 1952
rect 5108 1912 5117 1952
rect 5059 1911 5117 1912
rect 7467 1952 7509 1961
rect 7467 1912 7468 1952
rect 7508 1912 7509 1952
rect 7467 1903 7509 1912
rect 7563 1952 7605 1961
rect 7563 1912 7564 1952
rect 7604 1912 7605 1952
rect 7563 1903 7605 1912
rect 12651 1952 12693 1961
rect 12651 1912 12652 1952
rect 12692 1912 12693 1952
rect 12651 1903 12693 1912
rect 1131 1868 1173 1877
rect 1131 1828 1132 1868
rect 1172 1828 1173 1868
rect 1131 1819 1173 1828
rect 3531 1868 3573 1877
rect 3531 1828 3532 1868
rect 3572 1828 3573 1868
rect 3531 1819 3573 1828
rect 7371 1868 7413 1877
rect 7371 1828 7372 1868
rect 7412 1828 7413 1868
rect 7371 1819 7413 1828
rect 12843 1868 12885 1877
rect 12843 1828 12844 1868
rect 12884 1828 12885 1868
rect 12843 1819 12885 1828
rect 1227 1784 1269 1793
rect 1227 1744 1228 1784
rect 1268 1744 1269 1784
rect 1227 1735 1269 1744
rect 576 1532 15360 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 15360 1532
rect 576 1468 15360 1492
rect 4491 1280 4533 1289
rect 4491 1240 4492 1280
rect 4532 1240 4533 1280
rect 4491 1231 4533 1240
rect 5355 1280 5397 1289
rect 5355 1240 5356 1280
rect 5396 1240 5397 1280
rect 5355 1231 5397 1240
rect 4395 1196 4437 1205
rect 4395 1156 4396 1196
rect 4436 1156 4437 1196
rect 4395 1147 4437 1156
rect 5259 1196 5301 1205
rect 5259 1156 5260 1196
rect 5300 1156 5301 1196
rect 5259 1147 5301 1156
rect 6795 1196 6837 1205
rect 6795 1156 6796 1196
rect 6836 1156 6837 1196
rect 6795 1147 6837 1156
rect 8139 1196 8181 1205
rect 8139 1156 8140 1196
rect 8180 1156 8181 1196
rect 8139 1147 8181 1156
rect 9003 1196 9045 1205
rect 9003 1156 9004 1196
rect 9044 1156 9045 1196
rect 9003 1147 9045 1156
rect 10923 1196 10965 1205
rect 10923 1156 10924 1196
rect 10964 1156 10965 1196
rect 10923 1147 10965 1156
rect 1315 1112 1373 1113
rect 1315 1072 1324 1112
rect 1364 1072 1373 1112
rect 1315 1071 1373 1072
rect 1411 1112 1469 1113
rect 1411 1072 1420 1112
rect 1460 1072 1469 1112
rect 1411 1071 1469 1072
rect 2947 1112 3005 1113
rect 2947 1072 2956 1112
rect 2996 1072 3005 1112
rect 2947 1071 3005 1072
rect 3043 1112 3101 1113
rect 3043 1072 3052 1112
rect 3092 1072 3101 1112
rect 3043 1071 3101 1072
rect 4099 1112 4157 1113
rect 4099 1072 4108 1112
rect 4148 1072 4157 1112
rect 4099 1071 4157 1072
rect 4587 1112 4629 1121
rect 4587 1072 4588 1112
rect 4628 1072 4629 1112
rect 4587 1063 4629 1072
rect 5451 1112 5493 1121
rect 5451 1072 5452 1112
rect 5492 1072 5493 1112
rect 5451 1063 5493 1072
rect 6987 1112 7029 1121
rect 6987 1072 6988 1112
rect 7028 1072 7029 1112
rect 6987 1063 7029 1072
rect 7947 1112 7989 1121
rect 7947 1072 7948 1112
rect 7988 1072 7989 1112
rect 7947 1063 7989 1072
rect 9195 1112 9237 1121
rect 9195 1072 9196 1112
rect 9236 1072 9237 1112
rect 9195 1063 9237 1072
rect 10731 1112 10773 1121
rect 10731 1072 10732 1112
rect 10772 1072 10773 1112
rect 10731 1063 10773 1072
rect 835 944 893 945
rect 835 904 844 944
rect 884 904 893 944
rect 835 903 893 904
rect 1795 944 1853 945
rect 1795 904 1804 944
rect 1844 904 1853 944
rect 1795 903 1853 904
rect 2467 944 2525 945
rect 2467 904 2476 944
rect 2516 904 2525 944
rect 2467 903 2525 904
rect 6115 944 6173 945
rect 6115 904 6124 944
rect 6164 904 6173 944
rect 6115 903 6173 904
rect 6499 944 6557 945
rect 6499 904 6508 944
rect 6548 904 6557 944
rect 6499 903 6557 904
rect 7651 944 7709 945
rect 7651 904 7660 944
rect 7700 904 7709 944
rect 7651 903 7709 904
rect 8707 944 8765 945
rect 8707 904 8716 944
rect 8756 904 8765 944
rect 8707 903 8765 904
rect 14755 944 14813 945
rect 14755 904 14764 944
rect 14804 904 14813 944
rect 14755 903 14813 904
rect 15139 944 15197 945
rect 15139 904 15148 944
rect 15188 904 15197 944
rect 15139 903 15197 904
rect 576 776 15360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 15360 776
rect 576 712 15360 736
<< via1 >>
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 1132 12664 1172 12704
rect 3052 12664 3092 12704
rect 3244 12664 3284 12704
rect 3820 12664 3860 12704
rect 4012 12664 4052 12704
rect 4588 12664 4628 12704
rect 5836 12664 5876 12704
rect 6796 12664 6836 12704
rect 9580 12664 9620 12704
rect 9772 12664 9812 12704
rect 11596 12664 11636 12704
rect 11788 12664 11828 12704
rect 13996 12664 14036 12704
rect 14380 12664 14420 12704
rect 14764 12664 14804 12704
rect 15148 12664 15188 12704
rect 1612 12580 1652 12620
rect 1420 12496 1460 12536
rect 1900 12496 1940 12536
rect 5068 12496 5108 12536
rect 5164 12496 5204 12536
rect 6028 12496 6068 12536
rect 1612 12412 1652 12452
rect 1420 12244 1460 12284
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 6028 11824 6068 11864
rect 5932 11740 5972 11780
rect 7468 11740 7508 11780
rect 9772 11740 9812 11780
rect 11788 11740 11828 11780
rect 1132 11656 1172 11696
rect 1228 11656 1268 11696
rect 3052 11656 3092 11696
rect 3148 11656 3188 11696
rect 3628 11656 3668 11696
rect 6124 11656 6164 11696
rect 7276 11656 7316 11696
rect 7372 11656 7412 11696
rect 9580 11656 9620 11696
rect 11596 11656 11636 11696
rect 1996 11488 2036 11528
rect 2188 11488 2228 11528
rect 5164 11488 5204 11528
rect 6988 11488 7028 11528
rect 7756 11488 7796 11528
rect 9292 11488 9332 11528
rect 10060 11488 10100 11528
rect 10924 11488 10964 11528
rect 13612 11488 13652 11528
rect 13996 11488 14036 11528
rect 14380 11488 14420 11528
rect 14764 11488 14804 11528
rect 15148 11488 15188 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 2668 11152 2708 11192
rect 3244 11152 3284 11192
rect 4396 11152 4436 11192
rect 7564 11152 7604 11192
rect 10636 11152 10676 11192
rect 11404 11152 11444 11192
rect 12172 11152 12212 11192
rect 12940 11152 12980 11192
rect 13804 11152 13844 11192
rect 14188 11152 14228 11192
rect 14572 11152 14612 11192
rect 14956 11152 14996 11192
rect 1132 10984 1172 11024
rect 1228 10984 1268 11024
rect 1900 10984 1940 11024
rect 3532 10984 3572 11024
rect 3628 10984 3668 11024
rect 4684 10984 4724 11024
rect 5356 10984 5396 11024
rect 5452 10984 5492 11024
rect 5932 10984 5972 11024
rect 8044 10984 8084 11024
rect 8140 10984 8180 11024
rect 8524 10984 8564 11024
rect 9676 10984 9716 11024
rect 11116 10984 11156 11024
rect 12460 10984 12500 11024
rect 3724 10900 3764 10940
rect 4876 10900 4916 10940
rect 9868 10900 9908 10940
rect 10924 10900 10964 10940
rect 12652 10900 12692 10940
rect 4684 10816 4724 10856
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 1708 10396 1748 10436
rect 1900 10228 1940 10268
rect 9196 10228 9236 10268
rect 10636 10228 10676 10268
rect 11020 10228 11060 10268
rect 12556 10228 12596 10268
rect 1708 10144 1748 10184
rect 3148 10144 3188 10184
rect 3244 10144 3284 10184
rect 3724 10144 3764 10184
rect 9004 10144 9044 10184
rect 10444 10144 10484 10184
rect 11212 10144 11252 10184
rect 12364 10144 12404 10184
rect 1036 9976 1076 10016
rect 1420 9976 1460 10016
rect 2188 9976 2228 10016
rect 2764 9976 2804 10016
rect 4492 9976 4532 10016
rect 5164 9976 5204 10016
rect 5644 9976 5684 10016
rect 6988 9976 7028 10016
rect 7372 9976 7412 10016
rect 8716 9976 8756 10016
rect 9484 9976 9524 10016
rect 10156 9976 10196 10016
rect 11500 9976 11540 10016
rect 12076 9976 12116 10016
rect 13228 9976 13268 10016
rect 13996 9976 14036 10016
rect 14380 9976 14420 10016
rect 14764 9976 14804 10016
rect 15148 9976 15188 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 844 9640 884 9680
rect 3244 9640 3284 9680
rect 4396 9640 4436 9680
rect 6220 9640 6260 9680
rect 8524 9640 8564 9680
rect 9292 9640 9332 9680
rect 10828 9640 10868 9680
rect 11020 9640 11060 9680
rect 11980 9640 12020 9680
rect 12748 9640 12788 9680
rect 13612 9640 13652 9680
rect 13996 9640 14036 9680
rect 14380 9640 14420 9680
rect 14764 9640 14804 9680
rect 15148 9640 15188 9680
rect 3532 9556 3572 9596
rect 1324 9472 1364 9512
rect 1420 9472 1460 9512
rect 1900 9472 1940 9512
rect 3724 9472 3764 9512
rect 4684 9472 4724 9512
rect 5164 9472 5204 9512
rect 6700 9472 6740 9512
rect 6796 9472 6836 9512
rect 7180 9472 7220 9512
rect 8812 9472 8852 9512
rect 12268 9472 12308 9512
rect 3532 9388 3572 9428
rect 4780 9388 4820 9428
rect 4876 9388 4916 9428
rect 9004 9388 9044 9428
rect 12460 9388 12500 9428
rect 8908 9304 8948 9344
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 1516 8800 1556 8840
rect 7180 8800 7220 8840
rect 1420 8716 1460 8756
rect 7276 8716 7316 8756
rect 10732 8716 10772 8756
rect 1612 8632 1652 8672
rect 2860 8632 2900 8672
rect 2956 8632 2996 8672
rect 3916 8632 3956 8672
rect 5164 8632 5204 8672
rect 5260 8632 5300 8672
rect 7084 8632 7124 8672
rect 8812 8632 8852 8672
rect 8908 8632 8948 8672
rect 9292 8632 9332 8672
rect 10540 8632 10580 8672
rect 1132 8464 1172 8504
rect 2476 8464 2516 8504
rect 3724 8464 3764 8504
rect 5740 8464 5780 8504
rect 6796 8464 6836 8504
rect 8332 8464 8372 8504
rect 10252 8464 10292 8504
rect 11020 8464 11060 8504
rect 12268 8464 12308 8504
rect 12652 8464 12692 8504
rect 13996 8464 14036 8504
rect 14380 8464 14420 8504
rect 14764 8464 14804 8504
rect 15148 8464 15188 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 2572 8128 2612 8168
rect 3436 8128 3476 8168
rect 4204 8128 4244 8168
rect 6028 8128 6068 8168
rect 7756 8128 7796 8168
rect 8524 8128 8564 8168
rect 9292 8128 9332 8168
rect 10444 8128 10484 8168
rect 14380 8128 14420 8168
rect 14764 8128 14804 8168
rect 15148 8128 15188 8168
rect 1132 7960 1172 8000
rect 1228 7960 1268 8000
rect 1804 7960 1844 8000
rect 3916 7960 3956 8000
rect 6508 7960 6548 8000
rect 6604 7960 6644 8000
rect 6988 7960 7028 8000
rect 8812 7960 8852 8000
rect 10732 7960 10772 8000
rect 12364 7960 12404 8000
rect 3724 7876 3764 7916
rect 9004 7876 9044 7916
rect 10924 7876 10964 7916
rect 12556 7876 12596 7916
rect 8908 7792 8948 7832
rect 3916 7708 3956 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 1516 7372 1556 7412
rect 6988 7372 7028 7412
rect 1708 7204 1748 7244
rect 5356 7204 5396 7244
rect 7180 7204 7220 7244
rect 10924 7204 10964 7244
rect 12556 7204 12596 7244
rect 1516 7120 1556 7160
rect 2860 7120 2900 7160
rect 2956 7120 2996 7160
rect 3724 7120 3764 7160
rect 5548 7120 5588 7160
rect 6988 7120 7028 7160
rect 8812 7120 8852 7160
rect 8908 7120 8948 7160
rect 9292 7120 9332 7160
rect 10732 7120 10772 7160
rect 12364 7120 12404 7160
rect 5356 7036 5396 7076
rect 844 6952 884 6992
rect 1228 6952 1268 6992
rect 2476 6952 2516 6992
rect 4684 6952 4724 6992
rect 5068 6952 5108 6992
rect 7468 6952 7508 6992
rect 8332 6952 8372 6992
rect 10444 6952 10484 6992
rect 11212 6952 11252 6992
rect 12844 6952 12884 6992
rect 13228 6952 13268 6992
rect 13804 6952 13844 6992
rect 14188 6952 14228 6992
rect 14764 6952 14804 6992
rect 15148 6952 15188 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 2380 6616 2420 6656
rect 4588 6616 4628 6656
rect 7852 6616 7892 6656
rect 10156 6616 10196 6656
rect 10924 6616 10964 6656
rect 11884 6616 11924 6656
rect 12652 6616 12692 6656
rect 13516 6616 13556 6656
rect 14380 6616 14420 6656
rect 14764 6616 14804 6656
rect 15148 6616 15188 6656
rect 6796 6532 6836 6572
rect 1036 6448 1076 6488
rect 1132 6448 1172 6488
rect 1612 6448 1652 6488
rect 3628 6448 3668 6488
rect 3724 6448 3764 6488
rect 5068 6448 5108 6488
rect 5164 6448 5204 6488
rect 5548 6448 5588 6488
rect 6604 6448 6644 6488
rect 7276 6448 7316 6488
rect 7372 6448 7412 6488
rect 8332 6448 8372 6488
rect 10444 6448 10484 6488
rect 12172 6448 12212 6488
rect 3820 6364 3860 6404
rect 6796 6364 6836 6404
rect 10636 6364 10676 6404
rect 12364 6364 12404 6404
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 1420 5860 1460 5900
rect 8044 5776 8084 5816
rect 1612 5692 1652 5732
rect 8236 5692 8276 5732
rect 10636 5692 10676 5732
rect 12556 5692 12596 5732
rect 1420 5608 1460 5648
rect 2860 5608 2900 5648
rect 2956 5608 2996 5648
rect 3820 5608 3860 5648
rect 6220 5608 6260 5648
rect 8044 5608 8084 5648
rect 8524 5608 8564 5648
rect 10444 5608 10484 5648
rect 12364 5608 12404 5648
rect 1132 5440 1172 5480
rect 2476 5440 2516 5480
rect 3628 5440 3668 5480
rect 4588 5440 4628 5480
rect 5260 5440 5300 5480
rect 5644 5440 5684 5480
rect 6028 5440 6068 5480
rect 7084 5440 7124 5480
rect 7468 5440 7508 5480
rect 9292 5440 9332 5480
rect 10156 5440 10196 5480
rect 10924 5440 10964 5480
rect 12076 5440 12116 5480
rect 12844 5440 12884 5480
rect 13996 5440 14036 5480
rect 14380 5440 14420 5480
rect 14764 5440 14804 5480
rect 15148 5440 15188 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 2572 5104 2612 5144
rect 4300 5104 4340 5144
rect 8044 5104 8084 5144
rect 8428 5104 8468 5144
rect 10060 5104 10100 5144
rect 11020 5104 11060 5144
rect 11212 5104 11252 5144
rect 13996 5104 14036 5144
rect 14380 5104 14420 5144
rect 14764 5104 14804 5144
rect 15148 5104 15188 5144
rect 6124 5020 6164 5060
rect 1132 4936 1172 4976
rect 1228 4936 1268 4976
rect 1804 4936 1844 4976
rect 3916 4936 3956 4976
rect 4012 4936 4052 4976
rect 5356 4936 5396 4976
rect 5452 4936 5492 4976
rect 5932 4936 5972 4976
rect 7276 4936 7316 4976
rect 7372 4936 7412 4976
rect 3820 4852 3860 4892
rect 6124 4852 6164 4892
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 1804 4264 1844 4304
rect 1900 4180 1940 4220
rect 9388 4180 9428 4220
rect 10060 4180 10100 4220
rect 11212 4180 11252 4220
rect 12556 4180 12596 4220
rect 1708 4096 1748 4136
rect 2956 4096 2996 4136
rect 3052 4096 3092 4136
rect 3820 4096 3860 4136
rect 6988 4096 7028 4136
rect 7084 4096 7124 4136
rect 7660 4096 7700 4136
rect 9196 4096 9236 4136
rect 10252 4096 10292 4136
rect 11020 4096 11060 4136
rect 12364 4096 12404 4136
rect 1036 3928 1076 3968
rect 1420 3928 1460 3968
rect 2572 3928 2612 3968
rect 4588 3928 4628 3968
rect 5356 3928 5396 3968
rect 5548 3928 5588 3968
rect 6604 3928 6644 3968
rect 8908 3928 8948 3968
rect 10540 3928 10580 3968
rect 12076 3928 12116 3968
rect 12844 3928 12884 3968
rect 13996 3928 14036 3968
rect 14380 3928 14420 3968
rect 14764 3928 14804 3968
rect 15148 3928 15188 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 844 3592 884 3632
rect 3148 3592 3188 3632
rect 3532 3592 3572 3632
rect 4780 3592 4820 3632
rect 7468 3592 7508 3632
rect 9484 3592 9524 3632
rect 10444 3592 10484 3632
rect 11212 3592 11252 3632
rect 12364 3592 12404 3632
rect 12748 3592 12788 3632
rect 13612 3592 13652 3632
rect 13996 3592 14036 3632
rect 14380 3592 14420 3632
rect 14764 3592 14804 3632
rect 15148 3592 15188 3632
rect 3820 3508 3860 3548
rect 1228 3424 1268 3464
rect 1324 3424 1364 3464
rect 1612 3424 1652 3464
rect 4012 3424 4052 3464
rect 5164 3424 5204 3464
rect 5260 3424 5300 3464
rect 5356 3424 5396 3464
rect 5740 3424 5780 3464
rect 7756 3424 7796 3464
rect 7852 3424 7892 3464
rect 10732 3424 10772 3464
rect 1132 3340 1172 3380
rect 3820 3340 3860 3380
rect 7948 3340 7988 3380
rect 10924 3340 10964 3380
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 5452 2752 5492 2792
rect 5356 2668 5396 2708
rect 9292 2668 9332 2708
rect 10828 2668 10868 2708
rect 12652 2668 12692 2708
rect 1228 2584 1268 2624
rect 1324 2584 1364 2624
rect 3148 2584 3188 2624
rect 3244 2584 3284 2624
rect 3724 2584 3764 2624
rect 5548 2584 5588 2624
rect 6412 2584 6452 2624
rect 6508 2584 6548 2624
rect 7372 2584 7412 2624
rect 9100 2584 9140 2624
rect 10636 2584 10676 2624
rect 12460 2584 12500 2624
rect 844 2416 884 2456
rect 1804 2416 1844 2456
rect 2668 2416 2708 2456
rect 4876 2416 4916 2456
rect 6028 2416 6068 2456
rect 7180 2416 7220 2456
rect 8140 2416 8180 2456
rect 8812 2416 8852 2456
rect 9580 2416 9620 2456
rect 10348 2416 10388 2456
rect 13804 2416 13844 2456
rect 14188 2416 14228 2456
rect 14572 2416 14612 2456
rect 14956 2416 14996 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 844 2080 884 2120
rect 2860 2080 2900 2120
rect 3244 2080 3284 2120
rect 5836 2080 5876 2120
rect 6220 2080 6260 2120
rect 8236 2080 8276 2120
rect 8908 2080 8948 2120
rect 10828 2080 10868 2120
rect 11020 2080 11060 2120
rect 11404 2080 11444 2120
rect 11980 2080 12020 2120
rect 13132 2080 13172 2120
rect 13996 2080 14036 2120
rect 14380 2080 14420 2120
rect 14764 2080 14804 2120
rect 15148 2080 15188 2120
rect 1324 1912 1364 1952
rect 1612 1912 1652 1952
rect 3628 1912 3668 1952
rect 3724 1912 3764 1952
rect 4492 1912 4532 1952
rect 4588 1912 4628 1952
rect 5068 1912 5108 1952
rect 7468 1912 7508 1952
rect 7564 1912 7604 1952
rect 12652 1912 12692 1952
rect 1132 1828 1172 1868
rect 3532 1828 3572 1868
rect 7372 1828 7412 1868
rect 12844 1828 12884 1868
rect 1228 1744 1268 1784
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 4492 1240 4532 1280
rect 5356 1240 5396 1280
rect 4396 1156 4436 1196
rect 5260 1156 5300 1196
rect 6796 1156 6836 1196
rect 8140 1156 8180 1196
rect 9004 1156 9044 1196
rect 10924 1156 10964 1196
rect 1324 1072 1364 1112
rect 1420 1072 1460 1112
rect 2956 1072 2996 1112
rect 3052 1072 3092 1112
rect 4108 1072 4148 1112
rect 4588 1072 4628 1112
rect 5452 1072 5492 1112
rect 6988 1072 7028 1112
rect 7948 1072 7988 1112
rect 9196 1072 9236 1112
rect 10732 1072 10772 1112
rect 844 904 884 944
rect 1804 904 1844 944
rect 2476 904 2516 944
rect 6124 904 6164 944
rect 6508 904 6548 944
rect 7660 904 7700 944
rect 8716 904 8756 944
rect 14764 904 14804 944
rect 15148 904 15188 944
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
<< metal2 >>
rect 4352 12872 4720 12881
rect 3052 12832 3572 12872
rect 1132 12704 1172 12713
rect 1036 12664 1132 12704
rect 1036 11528 1076 12664
rect 1132 12655 1172 12664
rect 3052 12704 3092 12832
rect 3052 12655 3092 12664
rect 3244 12704 3284 12713
rect 1612 12620 1652 12629
rect 1652 12580 1940 12620
rect 1612 12571 1652 12580
rect 1419 12536 1461 12545
rect 1419 12496 1420 12536
rect 1460 12496 1461 12536
rect 1419 12487 1461 12496
rect 1900 12536 1940 12580
rect 1900 12487 1940 12496
rect 1420 12402 1460 12487
rect 1612 12452 1652 12461
rect 1652 12412 1844 12452
rect 1612 12403 1652 12412
rect 1420 12284 1460 12293
rect 1420 11873 1460 12244
rect 1804 12032 1844 12412
rect 3244 12284 3284 12664
rect 2956 12244 3284 12284
rect 1804 11992 2228 12032
rect 1131 11864 1173 11873
rect 1131 11824 1132 11864
rect 1172 11824 1173 11864
rect 1131 11815 1173 11824
rect 1419 11864 1461 11873
rect 1419 11824 1420 11864
rect 1460 11824 1461 11864
rect 1419 11815 1461 11824
rect 1132 11696 1172 11815
rect 1228 11705 1268 11790
rect 1132 11647 1172 11656
rect 1227 11696 1269 11705
rect 1227 11656 1228 11696
rect 1268 11656 1269 11696
rect 1227 11647 1269 11656
rect 2091 11696 2133 11705
rect 2091 11656 2092 11696
rect 2132 11656 2133 11696
rect 2091 11647 2133 11656
rect 1996 11528 2036 11537
rect 1036 11488 1268 11528
rect 1132 11024 1172 11033
rect 1132 10529 1172 10984
rect 1228 11024 1268 11488
rect 1228 10975 1268 10984
rect 1900 11024 1940 11033
rect 1900 10529 1940 10984
rect 1131 10520 1173 10529
rect 1131 10480 1132 10520
rect 1172 10480 1173 10520
rect 1131 10471 1173 10480
rect 1707 10520 1749 10529
rect 1707 10480 1708 10520
rect 1748 10480 1749 10520
rect 1707 10471 1749 10480
rect 1899 10520 1941 10529
rect 1899 10480 1900 10520
rect 1940 10480 1941 10520
rect 1899 10471 1941 10480
rect 1708 10436 1748 10471
rect 1708 10385 1748 10396
rect 1900 10268 1940 10277
rect 1996 10268 2036 11488
rect 1940 10228 2036 10268
rect 1900 10219 1940 10228
rect 1707 10184 1749 10193
rect 1707 10144 1708 10184
rect 1748 10144 1749 10184
rect 1707 10135 1749 10144
rect 1708 10050 1748 10135
rect 1036 10016 1076 10025
rect 1420 10016 1460 10025
rect 2092 10016 2132 11647
rect 2188 11528 2228 11992
rect 2956 11948 2996 12244
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 2956 11908 3188 11948
rect 3052 11696 3092 11705
rect 3052 11537 3092 11656
rect 3148 11696 3188 11908
rect 3148 11647 3188 11656
rect 2188 11479 2228 11488
rect 3051 11528 3093 11537
rect 3051 11488 3052 11528
rect 3092 11488 3093 11528
rect 3051 11479 3093 11488
rect 2668 11192 2708 11201
rect 2668 10193 2708 11152
rect 3244 11192 3284 11201
rect 3244 10781 3284 11152
rect 3532 11024 3572 12832
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 3820 12704 3860 12713
rect 3628 11696 3668 11705
rect 3628 11537 3668 11656
rect 3627 11528 3669 11537
rect 3627 11488 3628 11528
rect 3668 11488 3669 11528
rect 3627 11479 3669 11488
rect 3532 10975 3572 10984
rect 3628 11024 3668 11479
rect 3628 10975 3668 10984
rect 3724 10940 3764 10949
rect 3820 10940 3860 12664
rect 4012 12704 4052 12713
rect 4012 12545 4052 12664
rect 4587 12704 4629 12713
rect 4587 12664 4588 12704
rect 4628 12664 4629 12704
rect 4587 12655 4629 12664
rect 5067 12704 5109 12713
rect 5067 12664 5068 12704
rect 5108 12664 5109 12704
rect 5067 12655 5109 12664
rect 5836 12704 5876 12713
rect 6796 12704 6836 12713
rect 5876 12664 5972 12704
rect 5836 12655 5876 12664
rect 4588 12570 4628 12655
rect 4011 12536 4053 12545
rect 4011 12496 4012 12536
rect 4052 12496 4053 12536
rect 4011 12487 4053 12496
rect 5068 12536 5108 12655
rect 5068 12487 5108 12496
rect 5163 12536 5205 12545
rect 5163 12496 5164 12536
rect 5204 12496 5205 12536
rect 5163 12487 5205 12496
rect 5164 12209 5204 12487
rect 5163 12200 5205 12209
rect 5163 12160 5164 12200
rect 5204 12160 5205 12200
rect 5163 12151 5205 12160
rect 5932 11780 5972 12664
rect 6027 12536 6069 12545
rect 6027 12496 6028 12536
rect 6068 12496 6069 12536
rect 6027 12487 6069 12496
rect 6028 11864 6068 12487
rect 6028 11815 6068 11824
rect 5932 11731 5972 11740
rect 6796 11705 6836 12664
rect 9580 12704 9620 12713
rect 7468 11780 7508 11789
rect 7508 11740 7604 11780
rect 7468 11731 7508 11740
rect 6123 11696 6165 11705
rect 6123 11656 6124 11696
rect 6164 11656 6165 11696
rect 6123 11647 6165 11656
rect 6795 11696 6837 11705
rect 7276 11696 7316 11705
rect 6795 11656 6796 11696
rect 6836 11656 6837 11696
rect 6795 11647 6837 11656
rect 6988 11656 7276 11696
rect 6124 11562 6164 11647
rect 5164 11528 5204 11537
rect 4876 11488 5164 11528
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 4396 11192 4436 11201
rect 4396 11024 4436 11152
rect 4684 11024 4724 11033
rect 4396 10984 4684 11024
rect 4684 10975 4724 10984
rect 3764 10900 3860 10940
rect 4876 10940 4916 11488
rect 5164 11479 5204 11488
rect 6988 11528 7028 11656
rect 7276 11647 7316 11656
rect 7372 11696 7412 11705
rect 6988 11479 7028 11488
rect 7372 11201 7412 11656
rect 7564 11528 7604 11740
rect 9580 11696 9620 12664
rect 9772 12704 9812 12713
rect 9772 11780 9812 12664
rect 9772 11731 9812 11740
rect 11596 12704 11636 12713
rect 9580 11647 9620 11656
rect 11596 11696 11636 12664
rect 11788 12704 11828 12713
rect 11788 11780 11828 12664
rect 13996 12704 14036 12713
rect 13611 12200 13653 12209
rect 13611 12160 13612 12200
rect 13652 12160 13653 12200
rect 13611 12151 13653 12160
rect 11788 11731 11828 11740
rect 11596 11647 11636 11656
rect 7756 11528 7796 11537
rect 7564 11488 7756 11528
rect 7756 11479 7796 11488
rect 9292 11528 9332 11537
rect 10060 11528 10100 11537
rect 7371 11192 7413 11201
rect 7371 11152 7372 11192
rect 7412 11152 7413 11192
rect 7371 11143 7413 11152
rect 7564 11192 7604 11201
rect 8139 11192 8181 11201
rect 7604 11152 8084 11192
rect 7564 11143 7604 11152
rect 3724 10891 3764 10900
rect 4876 10891 4916 10900
rect 5356 11024 5396 11033
rect 5356 10865 5396 10984
rect 5452 11024 5492 11033
rect 4683 10856 4725 10865
rect 4683 10816 4684 10856
rect 4724 10816 4725 10856
rect 4683 10807 4725 10816
rect 5355 10856 5397 10865
rect 5355 10816 5356 10856
rect 5396 10816 5397 10856
rect 5355 10807 5397 10816
rect 3243 10772 3285 10781
rect 3243 10732 3244 10772
rect 3284 10732 3285 10772
rect 3243 10723 3285 10732
rect 3627 10772 3669 10781
rect 3627 10732 3628 10772
rect 3668 10732 3669 10772
rect 3627 10723 3669 10732
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 3147 10268 3189 10277
rect 3147 10228 3148 10268
rect 3188 10228 3189 10268
rect 3147 10219 3189 10228
rect 3531 10268 3573 10277
rect 3531 10228 3532 10268
rect 3572 10228 3573 10268
rect 3531 10219 3573 10228
rect 2667 10184 2709 10193
rect 2667 10144 2668 10184
rect 2708 10144 2709 10184
rect 2667 10135 2709 10144
rect 3148 10184 3188 10219
rect 3148 10133 3188 10144
rect 3244 10184 3284 10193
rect 2188 10016 2228 10025
rect 1076 9976 1364 10016
rect 1036 9967 1076 9976
rect 844 9680 884 9689
rect 844 8765 884 9640
rect 1324 9512 1364 9976
rect 1460 9976 1652 10016
rect 2092 9976 2188 10016
rect 1420 9967 1460 9976
rect 1419 9848 1461 9857
rect 1419 9808 1420 9848
rect 1460 9808 1461 9848
rect 1419 9799 1461 9808
rect 1420 9521 1460 9799
rect 1324 9463 1364 9472
rect 1419 9512 1461 9521
rect 1419 9472 1420 9512
rect 1460 9472 1556 9512
rect 1419 9463 1461 9472
rect 1420 9378 1460 9463
rect 1420 8765 1460 8850
rect 1516 8840 1556 9472
rect 1516 8791 1556 8800
rect 843 8756 885 8765
rect 843 8716 844 8756
rect 884 8716 885 8756
rect 843 8707 885 8716
rect 1419 8756 1461 8765
rect 1419 8716 1420 8756
rect 1460 8716 1461 8756
rect 1419 8707 1461 8716
rect 1612 8672 1652 9976
rect 2188 9967 2228 9976
rect 2764 10016 2804 10025
rect 3244 10016 3284 10144
rect 2804 9976 3284 10016
rect 2764 9967 2804 9976
rect 3243 9680 3285 9689
rect 3243 9640 3244 9680
rect 3284 9640 3285 9680
rect 3243 9631 3285 9640
rect 3244 9546 3284 9631
rect 3532 9596 3572 10219
rect 3532 9547 3572 9556
rect 1899 9512 1941 9521
rect 1899 9472 1900 9512
rect 1940 9472 1941 9512
rect 1899 9463 1941 9472
rect 1900 9378 1940 9463
rect 3532 9428 3572 9437
rect 3628 9428 3668 10723
rect 4684 10722 4724 10807
rect 3724 10277 3764 10279
rect 3723 10268 3765 10277
rect 3723 10228 3724 10268
rect 3764 10228 3765 10268
rect 3723 10219 3765 10228
rect 3724 10184 3764 10219
rect 3724 10135 3764 10144
rect 4492 10025 4532 10110
rect 3723 10016 3765 10025
rect 3723 9976 3724 10016
rect 3764 9976 3765 10016
rect 3723 9967 3765 9976
rect 4491 10016 4533 10025
rect 5164 10016 5204 10025
rect 4491 9976 4492 10016
rect 4532 9976 4533 10016
rect 4491 9967 4533 9976
rect 4876 9976 5164 10016
rect 5452 10016 5492 10984
rect 5932 11024 5972 11033
rect 5932 10865 5972 10984
rect 8044 11024 8084 11152
rect 8139 11152 8140 11192
rect 8180 11152 8181 11192
rect 8139 11143 8181 11152
rect 8523 11192 8565 11201
rect 8523 11152 8524 11192
rect 8564 11152 8565 11192
rect 8523 11143 8565 11152
rect 8044 10975 8084 10984
rect 8140 11024 8180 11143
rect 8140 10975 8180 10984
rect 8524 11024 8564 11143
rect 9292 11024 9332 11488
rect 9868 11488 10060 11528
rect 9676 11024 9716 11033
rect 9292 10984 9676 11024
rect 8524 10975 8564 10984
rect 9676 10975 9716 10984
rect 9868 10940 9908 11488
rect 10060 11479 10100 11488
rect 10924 11528 10964 11537
rect 9868 10891 9908 10900
rect 10636 11192 10676 11201
rect 5931 10856 5973 10865
rect 5931 10816 5932 10856
rect 5972 10816 5973 10856
rect 5931 10807 5973 10816
rect 9196 10268 9236 10277
rect 9004 10184 9044 10193
rect 8716 10144 9004 10184
rect 5644 10016 5684 10025
rect 5452 9976 5644 10016
rect 3724 9512 3764 9967
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 3819 9680 3861 9689
rect 3819 9640 3820 9680
rect 3860 9640 3861 9680
rect 3819 9631 3861 9640
rect 4396 9680 4436 9689
rect 3724 9463 3764 9472
rect 3572 9388 3668 9428
rect 3532 9379 3572 9388
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 1612 8623 1652 8632
rect 2475 8672 2517 8681
rect 2475 8632 2476 8672
rect 2516 8632 2517 8672
rect 2475 8623 2517 8632
rect 2860 8672 2900 8681
rect 1132 8504 1172 8513
rect 2476 8504 2516 8623
rect 2860 8513 2900 8632
rect 2955 8672 2997 8681
rect 2955 8632 2956 8672
rect 2996 8632 2997 8672
rect 2955 8623 2997 8632
rect 2956 8538 2996 8623
rect 3627 8588 3669 8597
rect 3627 8548 3628 8588
rect 3668 8548 3669 8588
rect 3627 8539 3669 8548
rect 1172 8464 1268 8504
rect 1132 8455 1172 8464
rect 1131 8168 1173 8177
rect 1131 8128 1132 8168
rect 1172 8128 1173 8168
rect 1131 8119 1173 8128
rect 1132 8009 1172 8119
rect 1131 8000 1173 8009
rect 1131 7960 1132 8000
rect 1172 7960 1173 8000
rect 1131 7951 1173 7960
rect 1228 8000 1268 8464
rect 2476 8455 2516 8464
rect 2859 8504 2901 8513
rect 2859 8464 2860 8504
rect 2900 8464 2901 8504
rect 2859 8455 2901 8464
rect 1707 8168 1749 8177
rect 1707 8128 1708 8168
rect 1748 8128 1749 8168
rect 1707 8119 1749 8128
rect 2571 8168 2613 8177
rect 2571 8128 2572 8168
rect 2612 8128 2613 8168
rect 2571 8119 2613 8128
rect 3436 8168 3476 8177
rect 3476 8128 3572 8168
rect 3436 8119 3476 8128
rect 1228 7951 1268 7960
rect 1515 8000 1557 8009
rect 1515 7960 1516 8000
rect 1556 7960 1557 8000
rect 1515 7951 1557 7960
rect 1132 7866 1172 7951
rect 1516 7412 1556 7951
rect 1516 7363 1556 7372
rect 1708 7244 1748 8119
rect 2572 8034 2612 8119
rect 1803 8000 1845 8009
rect 1803 7960 1804 8000
rect 1844 7960 1845 8000
rect 1803 7951 1845 7960
rect 1804 7866 1844 7951
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 1708 7195 1748 7204
rect 2859 7244 2901 7253
rect 2859 7204 2860 7244
rect 2900 7204 2901 7244
rect 2859 7195 2901 7204
rect 1516 7160 1556 7169
rect 1228 7120 1516 7160
rect 844 6992 884 7001
rect 1228 6992 1268 7120
rect 1516 7111 1556 7120
rect 2475 7160 2517 7169
rect 2475 7120 2476 7160
rect 2516 7120 2517 7160
rect 2475 7111 2517 7120
rect 2860 7160 2900 7195
rect 884 6952 1172 6992
rect 844 6943 884 6952
rect 1036 6488 1076 6497
rect 1036 6161 1076 6448
rect 1132 6488 1172 6952
rect 1228 6943 1268 6952
rect 2476 6992 2516 7111
rect 2860 7109 2900 7120
rect 2955 7160 2997 7169
rect 2955 7120 2956 7160
rect 2996 7120 2997 7160
rect 2955 7111 2997 7120
rect 2956 7026 2996 7111
rect 2476 6943 2516 6952
rect 2380 6656 2420 6665
rect 1132 6439 1172 6448
rect 1612 6488 1652 6497
rect 1612 6161 1652 6448
rect 1035 6152 1077 6161
rect 1035 6112 1036 6152
rect 1076 6112 1077 6152
rect 1035 6103 1077 6112
rect 1419 6152 1461 6161
rect 1419 6112 1420 6152
rect 1460 6112 1461 6152
rect 1419 6103 1461 6112
rect 1611 6152 1653 6161
rect 1611 6112 1612 6152
rect 1652 6112 1653 6152
rect 1611 6103 1653 6112
rect 1420 5900 1460 6103
rect 1420 5851 1460 5860
rect 1612 5732 1652 5741
rect 2380 5732 2420 6616
rect 3532 6488 3572 8128
rect 3628 7757 3668 8539
rect 3724 8504 3764 8513
rect 3820 8504 3860 9631
rect 4396 9512 4436 9640
rect 4684 9512 4724 9521
rect 4396 9472 4684 9512
rect 4684 9463 4724 9472
rect 4779 9428 4821 9437
rect 4779 9388 4780 9428
rect 4820 9388 4821 9428
rect 4779 9379 4821 9388
rect 4876 9428 4916 9976
rect 5164 9967 5204 9976
rect 5644 9967 5684 9976
rect 6988 10016 7028 10025
rect 7372 10016 7412 10025
rect 6220 9680 6260 9689
rect 5164 9512 5204 9523
rect 6220 9521 6260 9640
rect 5164 9437 5204 9472
rect 6219 9512 6261 9521
rect 6219 9472 6220 9512
rect 6260 9472 6261 9512
rect 6219 9463 6261 9472
rect 6699 9512 6741 9521
rect 6699 9472 6700 9512
rect 6740 9472 6741 9512
rect 6699 9463 6741 9472
rect 6796 9512 6836 9523
rect 4876 9379 4916 9388
rect 5163 9428 5205 9437
rect 5163 9388 5164 9428
rect 5204 9388 5205 9428
rect 5163 9379 5205 9388
rect 4780 9294 4820 9379
rect 3916 8681 3956 8766
rect 3915 8672 3957 8681
rect 3915 8632 3916 8672
rect 3956 8632 3957 8672
rect 3915 8623 3957 8632
rect 5164 8672 5204 9379
rect 6700 9378 6740 9463
rect 6796 9437 6836 9472
rect 6795 9428 6837 9437
rect 6795 9388 6796 9428
rect 6836 9388 6837 9428
rect 6795 9379 6837 9388
rect 6796 9185 6836 9379
rect 6795 9176 6837 9185
rect 6795 9136 6796 9176
rect 6836 9136 6837 9176
rect 6795 9127 6837 9136
rect 5164 8623 5204 8632
rect 5260 8672 5300 8681
rect 6988 8672 7028 9976
rect 7276 9976 7372 10016
rect 7180 9512 7220 9521
rect 7180 9437 7220 9472
rect 7179 9428 7221 9437
rect 7179 9388 7180 9428
rect 7220 9388 7221 9428
rect 7179 9379 7221 9388
rect 7180 8840 7220 9379
rect 7180 8791 7220 8800
rect 7276 8756 7316 9976
rect 7372 9967 7412 9976
rect 8716 10016 8756 10144
rect 9004 10135 9044 10144
rect 9196 10016 9236 10228
rect 10636 10268 10676 11152
rect 10924 10940 10964 11488
rect 13612 11528 13652 12151
rect 13996 12041 14036 12664
rect 14380 12704 14420 12713
rect 13995 12032 14037 12041
rect 13995 11992 13996 12032
rect 14036 11992 14037 12032
rect 13995 11983 14037 11992
rect 14380 11873 14420 12664
rect 14764 12704 14804 12713
rect 15148 12704 15188 12713
rect 14804 12664 14900 12704
rect 14764 12655 14804 12664
rect 14379 11864 14421 11873
rect 14379 11824 14380 11864
rect 14420 11824 14421 11864
rect 14379 11815 14421 11824
rect 13612 11479 13652 11488
rect 13995 11528 14037 11537
rect 13995 11488 13996 11528
rect 14036 11488 14037 11528
rect 13995 11479 14037 11488
rect 14380 11528 14420 11537
rect 13996 11394 14036 11479
rect 11404 11192 11444 11201
rect 11116 11024 11156 11033
rect 11404 11024 11444 11152
rect 11156 10984 11444 11024
rect 12172 11192 12212 11201
rect 12940 11192 12980 11201
rect 12172 11024 12212 11152
rect 12652 11152 12940 11192
rect 12460 11024 12500 11033
rect 12172 10984 12460 11024
rect 11116 10975 11156 10984
rect 12460 10975 12500 10984
rect 10924 10891 10964 10900
rect 12652 10940 12692 11152
rect 12940 11143 12980 11152
rect 13804 11192 13844 11201
rect 12652 10891 12692 10900
rect 13804 10865 13844 11152
rect 14188 11192 14228 11201
rect 13803 10856 13845 10865
rect 13803 10816 13804 10856
rect 13844 10816 13845 10856
rect 13803 10807 13845 10816
rect 14188 10529 14228 11152
rect 14380 11033 14420 11488
rect 14764 11528 14804 11537
rect 14572 11192 14612 11201
rect 14379 11024 14421 11033
rect 14379 10984 14380 11024
rect 14420 10984 14421 11024
rect 14379 10975 14421 10984
rect 14187 10520 14229 10529
rect 14187 10480 14188 10520
rect 14228 10480 14229 10520
rect 14187 10471 14229 10480
rect 10636 10219 10676 10228
rect 11020 10268 11060 10277
rect 10444 10184 10484 10193
rect 10156 10144 10444 10184
rect 9484 10016 9524 10025
rect 9196 9976 9484 10016
rect 8716 9967 8756 9976
rect 9484 9967 9524 9976
rect 10156 10016 10196 10144
rect 10444 10135 10484 10144
rect 10156 9967 10196 9976
rect 8524 9680 8564 9689
rect 9292 9680 9332 9689
rect 10828 9680 10868 9689
rect 8524 9512 8564 9640
rect 9004 9640 9292 9680
rect 8812 9512 8852 9521
rect 8524 9472 8812 9512
rect 8812 9463 8852 9472
rect 9004 9428 9044 9640
rect 9292 9631 9332 9640
rect 10732 9640 10828 9680
rect 9004 9379 9044 9388
rect 8908 9344 8948 9353
rect 8908 8849 8948 9304
rect 8907 8840 8949 8849
rect 8907 8800 8908 8840
rect 8948 8800 8949 8840
rect 8907 8791 8949 8800
rect 9291 8840 9333 8849
rect 9291 8800 9292 8840
rect 9332 8800 9333 8840
rect 9291 8791 9333 8800
rect 7276 8707 7316 8716
rect 7084 8672 7124 8681
rect 6988 8632 7084 8672
rect 5260 8504 5300 8632
rect 7084 8623 7124 8632
rect 8331 8672 8373 8681
rect 8331 8632 8332 8672
rect 8372 8632 8373 8672
rect 8331 8623 8373 8632
rect 8811 8672 8853 8681
rect 8811 8632 8812 8672
rect 8852 8632 8853 8672
rect 8811 8623 8853 8632
rect 8908 8672 8948 8791
rect 8908 8623 8948 8632
rect 9292 8672 9332 8791
rect 10732 8756 10772 9640
rect 10828 9631 10868 9640
rect 11020 9680 11060 10228
rect 12555 10268 12597 10277
rect 12555 10228 12556 10268
rect 12596 10228 12597 10268
rect 12555 10219 12597 10228
rect 13227 10268 13269 10277
rect 13227 10228 13228 10268
rect 13268 10228 13269 10268
rect 13227 10219 13269 10228
rect 11212 10184 11252 10193
rect 12364 10184 12404 10193
rect 11252 10144 11540 10184
rect 11212 10135 11252 10144
rect 11500 10016 11540 10144
rect 11500 9967 11540 9976
rect 12076 10144 12364 10184
rect 12076 10016 12116 10144
rect 12364 10135 12404 10144
rect 12556 10134 12596 10219
rect 12076 9967 12116 9976
rect 13228 10016 13268 10219
rect 14572 10193 14612 11152
rect 14764 10697 14804 11488
rect 14860 11369 14900 12664
rect 15148 11705 15188 12664
rect 15147 11696 15189 11705
rect 15147 11656 15148 11696
rect 15188 11656 15189 11696
rect 15147 11647 15189 11656
rect 15148 11528 15188 11537
rect 14859 11360 14901 11369
rect 14859 11320 14860 11360
rect 14900 11320 14901 11360
rect 14859 11311 14901 11320
rect 15148 11201 15188 11488
rect 14956 11192 14996 11201
rect 14763 10688 14805 10697
rect 14763 10648 14764 10688
rect 14804 10648 14805 10688
rect 14763 10639 14805 10648
rect 14956 10361 14996 11152
rect 15147 11192 15189 11201
rect 15147 11152 15148 11192
rect 15188 11152 15189 11192
rect 15147 11143 15189 11152
rect 14955 10352 14997 10361
rect 14955 10312 14956 10352
rect 14996 10312 14997 10352
rect 14955 10303 14997 10312
rect 14571 10184 14613 10193
rect 14571 10144 14572 10184
rect 14612 10144 14613 10184
rect 14571 10135 14613 10144
rect 13228 9967 13268 9976
rect 13996 10016 14036 10025
rect 13996 9857 14036 9976
rect 14380 10016 14420 10025
rect 14764 10016 14804 10025
rect 15147 10016 15189 10025
rect 14420 9976 14516 10016
rect 14380 9967 14420 9976
rect 13995 9848 14037 9857
rect 13995 9808 13996 9848
rect 14036 9808 14037 9848
rect 13995 9799 14037 9808
rect 14476 9689 14516 9976
rect 14804 9976 14900 10016
rect 14764 9967 14804 9976
rect 11020 9631 11060 9640
rect 11980 9680 12020 9689
rect 12748 9680 12788 9689
rect 11980 9512 12020 9640
rect 12460 9640 12748 9680
rect 12268 9512 12308 9521
rect 11980 9472 12268 9512
rect 12268 9463 12308 9472
rect 12460 9428 12500 9640
rect 12748 9631 12788 9640
rect 13612 9680 13652 9689
rect 13612 9521 13652 9640
rect 13996 9680 14036 9689
rect 13611 9512 13653 9521
rect 13611 9472 13612 9512
rect 13652 9472 13653 9512
rect 13611 9463 13653 9472
rect 12460 9379 12500 9388
rect 13996 9353 14036 9640
rect 14380 9680 14420 9689
rect 13995 9344 14037 9353
rect 13995 9304 13996 9344
rect 14036 9304 14037 9344
rect 13995 9295 14037 9304
rect 10732 8707 10772 8716
rect 14380 8681 14420 9640
rect 14475 9680 14517 9689
rect 14475 9640 14476 9680
rect 14516 9640 14517 9680
rect 14475 9631 14517 9640
rect 14764 9680 14804 9689
rect 14764 8849 14804 9640
rect 14860 9185 14900 9976
rect 15147 9976 15148 10016
rect 15188 9976 15189 10016
rect 15147 9967 15189 9976
rect 15148 9882 15188 9967
rect 15148 9680 15188 9689
rect 14859 9176 14901 9185
rect 14859 9136 14860 9176
rect 14900 9136 14901 9176
rect 14859 9127 14901 9136
rect 15148 9017 15188 9640
rect 15147 9008 15189 9017
rect 15147 8968 15148 9008
rect 15188 8968 15189 9008
rect 15147 8959 15189 8968
rect 14763 8840 14805 8849
rect 14763 8800 14764 8840
rect 14804 8800 14805 8840
rect 14763 8791 14805 8800
rect 10540 8672 10580 8681
rect 9292 8623 9332 8632
rect 10252 8632 10540 8672
rect 5740 8504 5780 8513
rect 3820 8464 3956 8504
rect 5260 8464 5740 8504
rect 3724 7916 3764 8464
rect 3916 8000 3956 8464
rect 5740 8455 5780 8464
rect 6796 8504 6836 8513
rect 8332 8504 8372 8623
rect 8812 8538 8852 8623
rect 6836 8464 6932 8504
rect 6796 8455 6836 8464
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 4204 8168 4244 8177
rect 3916 7951 3956 7960
rect 4012 8128 4204 8168
rect 3724 7867 3764 7876
rect 3627 7748 3669 7757
rect 3627 7708 3628 7748
rect 3668 7708 3669 7748
rect 3627 7699 3669 7708
rect 3915 7748 3957 7757
rect 3915 7708 3916 7748
rect 3956 7708 3957 7748
rect 3915 7699 3957 7708
rect 3916 7614 3956 7699
rect 3723 7244 3765 7253
rect 3723 7204 3724 7244
rect 3764 7204 3765 7244
rect 3723 7195 3765 7204
rect 3724 7160 3764 7195
rect 3628 6488 3668 6497
rect 3532 6448 3628 6488
rect 3628 6439 3668 6448
rect 3724 6488 3764 7120
rect 3724 6439 3764 6448
rect 3820 6404 3860 6413
rect 4012 6404 4052 8128
rect 4204 8119 4244 8128
rect 6028 8168 6068 8177
rect 6028 8009 6068 8128
rect 6027 8000 6069 8009
rect 6027 7960 6028 8000
rect 6068 7960 6069 8000
rect 6027 7951 6069 7960
rect 6507 8000 6549 8009
rect 6507 7960 6508 8000
rect 6548 7960 6549 8000
rect 6507 7951 6549 7960
rect 6604 8000 6644 8011
rect 6508 7866 6548 7951
rect 6604 7925 6644 7960
rect 6603 7916 6645 7925
rect 6603 7876 6604 7916
rect 6644 7876 6645 7916
rect 6603 7867 6645 7876
rect 5356 7244 5396 7253
rect 5164 7204 5356 7244
rect 4684 7001 4724 7086
rect 4683 6992 4725 7001
rect 4683 6952 4684 6992
rect 4724 6952 4725 6992
rect 4683 6943 4725 6952
rect 5068 6992 5108 7001
rect 5164 6992 5204 7204
rect 5356 7195 5396 7204
rect 5548 7160 5588 7169
rect 6892 7160 6932 8464
rect 8332 8455 8372 8464
rect 10252 8504 10292 8632
rect 10540 8623 10580 8632
rect 14379 8672 14421 8681
rect 14379 8632 14380 8672
rect 14420 8632 14421 8672
rect 14379 8623 14421 8632
rect 10252 8455 10292 8464
rect 11020 8504 11060 8513
rect 7179 8168 7221 8177
rect 7179 8128 7180 8168
rect 7220 8128 7221 8168
rect 7179 8119 7221 8128
rect 7755 8168 7797 8177
rect 7755 8128 7756 8168
rect 7796 8128 7797 8168
rect 7755 8119 7797 8128
rect 8524 8168 8564 8177
rect 9292 8168 9332 8177
rect 6988 8000 7028 8009
rect 6988 7925 7028 7960
rect 6987 7916 7029 7925
rect 6987 7876 6988 7916
rect 7028 7876 7029 7916
rect 6987 7867 7029 7876
rect 6988 7412 7028 7867
rect 6988 7363 7028 7372
rect 7180 7244 7220 8119
rect 7756 8034 7796 8119
rect 8524 8000 8564 8128
rect 9004 8128 9292 8168
rect 8812 8000 8852 8009
rect 8524 7960 8812 8000
rect 8812 7951 8852 7960
rect 9004 7916 9044 8128
rect 9292 8119 9332 8128
rect 10444 8168 10484 8177
rect 10444 8000 10484 8128
rect 10732 8000 10772 8009
rect 10444 7960 10732 8000
rect 10732 7951 10772 7960
rect 9004 7867 9044 7876
rect 10924 7916 10964 7925
rect 11020 7916 11060 8464
rect 12268 8504 12308 8513
rect 12268 8000 12308 8464
rect 12652 8504 12692 8513
rect 12364 8000 12404 8009
rect 12268 7960 12364 8000
rect 12364 7951 12404 7960
rect 10964 7876 11060 7916
rect 12556 7916 12596 7925
rect 12652 7916 12692 8464
rect 13995 8504 14037 8513
rect 13995 8464 13996 8504
rect 14036 8464 14037 8504
rect 13995 8455 14037 8464
rect 14380 8504 14420 8513
rect 13996 8370 14036 8455
rect 14380 8345 14420 8464
rect 14764 8504 14804 8513
rect 15148 8504 15188 8513
rect 14804 8464 14996 8504
rect 14764 8455 14804 8464
rect 14379 8336 14421 8345
rect 14379 8296 14380 8336
rect 14420 8296 14421 8336
rect 14379 8287 14421 8296
rect 12596 7876 12692 7916
rect 14380 8168 14420 8177
rect 10924 7867 10964 7876
rect 12556 7867 12596 7876
rect 14380 7841 14420 8128
rect 14764 8168 14804 8177
rect 8908 7832 8948 7841
rect 8908 7505 8948 7792
rect 14379 7832 14421 7841
rect 14379 7792 14380 7832
rect 14420 7792 14421 7832
rect 14379 7783 14421 7792
rect 14764 7673 14804 8128
rect 14859 8000 14901 8009
rect 14859 7960 14860 8000
rect 14900 7960 14901 8000
rect 14859 7951 14901 7960
rect 14763 7664 14805 7673
rect 14763 7624 14764 7664
rect 14804 7624 14805 7664
rect 14763 7615 14805 7624
rect 8907 7496 8949 7505
rect 8907 7456 8908 7496
rect 8948 7456 8949 7496
rect 8907 7447 8949 7456
rect 9291 7496 9333 7505
rect 9291 7456 9292 7496
rect 9332 7456 9333 7496
rect 9291 7447 9333 7456
rect 7180 7195 7220 7204
rect 6988 7160 7028 7169
rect 6892 7120 6988 7160
rect 5108 6952 5204 6992
rect 5356 7076 5396 7085
rect 5068 6943 5108 6952
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 5356 6749 5396 7036
rect 5548 7001 5588 7120
rect 6988 7111 7028 7120
rect 8331 7160 8373 7169
rect 8331 7120 8332 7160
rect 8372 7120 8373 7160
rect 8331 7111 8373 7120
rect 8811 7160 8853 7169
rect 8811 7120 8812 7160
rect 8852 7120 8853 7160
rect 8811 7111 8853 7120
rect 8908 7160 8948 7447
rect 8908 7111 8948 7120
rect 9292 7160 9332 7447
rect 10924 7244 10964 7253
rect 10732 7160 10772 7169
rect 9292 7111 9332 7120
rect 10444 7120 10732 7160
rect 5547 6992 5589 7001
rect 7468 6992 7508 7001
rect 5547 6952 5548 6992
rect 5588 6952 5589 6992
rect 5547 6943 5589 6952
rect 6604 6952 7468 6992
rect 5163 6740 5205 6749
rect 5163 6700 5164 6740
rect 5204 6700 5205 6740
rect 5163 6691 5205 6700
rect 5355 6740 5397 6749
rect 5355 6700 5356 6740
rect 5396 6700 5397 6740
rect 5355 6691 5397 6700
rect 5547 6740 5589 6749
rect 5547 6700 5548 6740
rect 5588 6700 5589 6740
rect 5547 6691 5589 6700
rect 4588 6656 4628 6665
rect 4588 6497 4628 6616
rect 4587 6488 4629 6497
rect 4587 6448 4588 6488
rect 4628 6448 4629 6488
rect 4587 6439 4629 6448
rect 5067 6488 5109 6497
rect 5067 6448 5068 6488
rect 5108 6448 5109 6488
rect 5067 6439 5109 6448
rect 5164 6488 5204 6691
rect 5164 6439 5204 6448
rect 5548 6488 5588 6691
rect 5548 6439 5588 6448
rect 6604 6488 6644 6952
rect 7468 6943 7508 6952
rect 8332 6992 8372 7111
rect 8812 7026 8852 7111
rect 8332 6943 8372 6952
rect 10444 6992 10484 7120
rect 10732 7111 10772 7120
rect 10924 6992 10964 7204
rect 12555 7244 12597 7253
rect 12555 7204 12556 7244
rect 12596 7204 12597 7244
rect 12555 7195 12597 7204
rect 13227 7244 13269 7253
rect 13227 7204 13228 7244
rect 13268 7204 13269 7244
rect 13227 7195 13269 7204
rect 12364 7160 12404 7169
rect 12364 7001 12404 7120
rect 12556 7110 12596 7195
rect 11212 6992 11252 7001
rect 10924 6952 11212 6992
rect 10444 6943 10484 6952
rect 11212 6943 11252 6952
rect 12363 6992 12405 7001
rect 12363 6952 12364 6992
rect 12404 6952 12405 6992
rect 12363 6943 12405 6952
rect 12843 6992 12885 7001
rect 12843 6952 12844 6992
rect 12884 6952 12885 6992
rect 12843 6943 12885 6952
rect 13228 6992 13268 7195
rect 14187 7160 14229 7169
rect 14187 7120 14188 7160
rect 14228 7120 14229 7160
rect 14187 7111 14229 7120
rect 13228 6943 13268 6952
rect 13803 6992 13845 7001
rect 13803 6952 13804 6992
rect 13844 6952 13845 6992
rect 13803 6943 13845 6952
rect 14188 6992 14228 7111
rect 14188 6943 14228 6952
rect 14764 6992 14804 7001
rect 14860 6992 14900 7951
rect 14956 7337 14996 8464
rect 15188 8464 15284 8504
rect 15148 8455 15188 8464
rect 15244 8177 15284 8464
rect 15148 8168 15188 8177
rect 15148 7505 15188 8128
rect 15243 8168 15285 8177
rect 15243 8128 15244 8168
rect 15284 8128 15285 8168
rect 15243 8119 15285 8128
rect 15147 7496 15189 7505
rect 15147 7456 15148 7496
rect 15188 7456 15189 7496
rect 15147 7447 15189 7456
rect 14955 7328 14997 7337
rect 14955 7288 14956 7328
rect 14996 7288 14997 7328
rect 14955 7279 14997 7288
rect 14804 6952 14900 6992
rect 15148 6992 15188 7001
rect 15188 6952 15284 6992
rect 14764 6943 14804 6952
rect 15148 6943 15188 6952
rect 12844 6858 12884 6943
rect 13804 6858 13844 6943
rect 13515 6824 13557 6833
rect 13515 6784 13516 6824
rect 13556 6784 13557 6824
rect 13515 6775 13557 6784
rect 6796 6581 6836 6666
rect 7852 6656 7892 6665
rect 6795 6572 6837 6581
rect 6795 6532 6796 6572
rect 6836 6532 6837 6572
rect 6795 6523 6837 6532
rect 7275 6572 7317 6581
rect 7275 6532 7276 6572
rect 7316 6532 7317 6572
rect 7275 6523 7317 6532
rect 6604 6439 6644 6448
rect 7276 6488 7316 6523
rect 7852 6497 7892 6616
rect 10156 6656 10196 6665
rect 10924 6656 10964 6665
rect 8331 6572 8373 6581
rect 8331 6532 8332 6572
rect 8372 6532 8373 6572
rect 8331 6523 8373 6532
rect 3860 6364 4052 6404
rect 3820 6355 3860 6364
rect 5068 6354 5108 6439
rect 7276 6437 7316 6448
rect 7371 6488 7413 6497
rect 7371 6448 7372 6488
rect 7412 6448 7413 6488
rect 7371 6439 7413 6448
rect 7851 6488 7893 6497
rect 7851 6448 7852 6488
rect 7892 6448 7893 6488
rect 7851 6439 7893 6448
rect 8332 6488 8372 6523
rect 10156 6488 10196 6616
rect 10636 6616 10924 6656
rect 10444 6488 10484 6497
rect 10156 6448 10444 6488
rect 6796 6404 6836 6413
rect 6796 6320 6836 6364
rect 7372 6354 7412 6439
rect 8332 6437 8372 6448
rect 10444 6439 10484 6448
rect 10636 6404 10676 6616
rect 10924 6607 10964 6616
rect 11884 6656 11924 6665
rect 12652 6656 12692 6665
rect 11884 6488 11924 6616
rect 12364 6616 12652 6656
rect 12172 6488 12212 6497
rect 11884 6448 12172 6488
rect 12172 6439 12212 6448
rect 10636 6355 10676 6364
rect 12364 6404 12404 6616
rect 12652 6607 12692 6616
rect 13516 6656 13556 6775
rect 15244 6665 15284 6952
rect 13516 6607 13556 6616
rect 14380 6656 14420 6665
rect 12364 6355 12404 6364
rect 14380 6329 14420 6616
rect 14764 6656 14804 6665
rect 14764 6497 14804 6616
rect 15148 6656 15188 6665
rect 14763 6488 14805 6497
rect 14763 6448 14764 6488
rect 14804 6448 14805 6488
rect 14763 6439 14805 6448
rect 14379 6320 14421 6329
rect 6796 6280 7124 6320
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 2859 5816 2901 5825
rect 2859 5776 2860 5816
rect 2900 5776 2901 5816
rect 2859 5767 2901 5776
rect 3819 5816 3861 5825
rect 3819 5776 3820 5816
rect 3860 5776 3861 5816
rect 3819 5767 3861 5776
rect 1652 5692 2420 5732
rect 1612 5683 1652 5692
rect 1420 5648 1460 5657
rect 1132 5608 1420 5648
rect 1132 5480 1172 5608
rect 1420 5599 1460 5608
rect 2475 5648 2517 5657
rect 2475 5608 2476 5648
rect 2516 5608 2517 5648
rect 2475 5599 2517 5608
rect 2860 5648 2900 5767
rect 2860 5599 2900 5608
rect 2955 5648 2997 5657
rect 2955 5608 2956 5648
rect 2996 5608 2997 5648
rect 2955 5599 2997 5608
rect 3820 5648 3860 5767
rect 6220 5648 6260 5657
rect 3860 5608 3956 5648
rect 3820 5599 3860 5608
rect 1132 5431 1172 5440
rect 2476 5480 2516 5599
rect 2956 5514 2996 5599
rect 2476 5431 2516 5440
rect 3628 5480 3668 5489
rect 3668 5440 3860 5480
rect 3628 5431 3668 5440
rect 1899 5144 1941 5153
rect 1899 5104 1900 5144
rect 1940 5104 1941 5144
rect 1899 5095 1941 5104
rect 2571 5144 2613 5153
rect 2571 5104 2572 5144
rect 2612 5104 2613 5144
rect 2571 5095 2613 5104
rect 1132 4976 1172 4985
rect 1132 4817 1172 4936
rect 1228 4976 1268 4985
rect 1131 4808 1173 4817
rect 1131 4768 1132 4808
rect 1172 4768 1173 4808
rect 1131 4759 1173 4768
rect 1036 3968 1076 3977
rect 1228 3968 1268 4936
rect 1804 4976 1844 4985
rect 1804 4817 1844 4936
rect 1803 4808 1845 4817
rect 1803 4768 1804 4808
rect 1844 4768 1845 4808
rect 1803 4759 1845 4768
rect 1804 4304 1844 4759
rect 1804 4255 1844 4264
rect 1900 4220 1940 5095
rect 2572 5010 2612 5095
rect 3820 4892 3860 5440
rect 3916 4976 3956 5608
rect 6124 5608 6220 5648
rect 4588 5480 4628 5489
rect 4204 5440 4588 5480
rect 3916 4927 3956 4936
rect 4012 4976 4052 4985
rect 4204 4976 4244 5440
rect 4588 5431 4628 5440
rect 5260 5480 5300 5489
rect 5451 5480 5493 5489
rect 5300 5440 5396 5480
rect 5260 5431 5300 5440
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 4052 4936 4244 4976
rect 4300 5144 4340 5153
rect 4012 4927 4052 4936
rect 3820 4843 3860 4852
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 1900 4171 1940 4180
rect 2956 4145 2996 4230
rect 1708 4136 1748 4145
rect 1076 3928 1268 3968
rect 1420 4096 1708 4136
rect 1420 3968 1460 4096
rect 1708 4087 1748 4096
rect 2955 4136 2997 4145
rect 2955 4096 2956 4136
rect 2996 4096 2997 4136
rect 2955 4087 2997 4096
rect 3052 4136 3092 4145
rect 1036 3919 1076 3928
rect 1420 3919 1460 3928
rect 2572 3968 2612 3977
rect 3052 3968 3092 4096
rect 3819 4136 3861 4145
rect 4300 4136 4340 5104
rect 5356 4976 5396 5440
rect 5451 5440 5452 5480
rect 5492 5440 5493 5480
rect 5451 5431 5493 5440
rect 5644 5480 5684 5489
rect 5452 5069 5492 5431
rect 5451 5060 5493 5069
rect 5451 5020 5452 5060
rect 5492 5020 5493 5060
rect 5451 5011 5493 5020
rect 5356 4927 5396 4936
rect 5452 4976 5492 5011
rect 5644 4976 5684 5440
rect 6028 5480 6068 5489
rect 5932 4976 5972 4985
rect 5644 4936 5932 4976
rect 5452 4926 5492 4936
rect 5932 4927 5972 4936
rect 6028 4892 6068 5440
rect 6124 5069 6164 5608
rect 6220 5599 6260 5608
rect 7084 5480 7124 6280
rect 14379 6280 14380 6320
rect 14420 6280 14421 6320
rect 14379 6271 14421 6280
rect 15148 6161 15188 6616
rect 15243 6656 15285 6665
rect 15243 6616 15244 6656
rect 15284 6616 15285 6656
rect 15243 6607 15285 6616
rect 15147 6152 15189 6161
rect 15147 6112 15148 6152
rect 15188 6112 15189 6152
rect 15147 6103 15189 6112
rect 14763 5984 14805 5993
rect 14763 5944 14764 5984
rect 14804 5944 14805 5984
rect 14763 5935 14805 5944
rect 8044 5816 8084 5825
rect 7948 5776 8044 5816
rect 7948 5657 7988 5776
rect 8044 5767 8084 5776
rect 8236 5741 8276 5826
rect 14379 5816 14421 5825
rect 14379 5776 14380 5816
rect 14420 5776 14421 5816
rect 14379 5767 14421 5776
rect 8235 5732 8277 5741
rect 8235 5692 8236 5732
rect 8276 5692 8277 5732
rect 8235 5683 8277 5692
rect 9291 5732 9333 5741
rect 9291 5692 9292 5732
rect 9332 5692 9333 5732
rect 9291 5683 9333 5692
rect 10636 5732 10676 5741
rect 7947 5648 7989 5657
rect 7947 5608 7948 5648
rect 7988 5608 7989 5648
rect 7947 5599 7989 5608
rect 8044 5648 8084 5657
rect 8523 5648 8565 5657
rect 8084 5608 8180 5648
rect 8044 5599 8084 5608
rect 7084 5431 7124 5440
rect 7468 5480 7508 5489
rect 7275 5228 7317 5237
rect 7275 5188 7276 5228
rect 7316 5188 7317 5228
rect 7275 5179 7317 5188
rect 6123 5060 6165 5069
rect 6123 5020 6124 5060
rect 6164 5020 6165 5060
rect 6123 5011 6165 5020
rect 7276 4976 7316 5179
rect 7276 4927 7316 4936
rect 7372 4976 7412 4985
rect 7468 4976 7508 5440
rect 7948 5237 7988 5599
rect 8140 5396 8180 5608
rect 8523 5608 8524 5648
rect 8564 5608 8565 5648
rect 8523 5599 8565 5608
rect 8524 5514 8564 5599
rect 9292 5480 9332 5683
rect 10444 5648 10484 5657
rect 9292 5431 9332 5440
rect 10156 5608 10444 5648
rect 10156 5480 10196 5608
rect 10444 5599 10484 5608
rect 10636 5480 10676 5692
rect 12556 5732 12596 5741
rect 12364 5648 12404 5657
rect 12076 5608 12364 5648
rect 10924 5480 10964 5489
rect 10636 5440 10924 5480
rect 10156 5431 10196 5440
rect 10924 5431 10964 5440
rect 12076 5480 12116 5608
rect 12364 5599 12404 5608
rect 12556 5480 12596 5692
rect 12844 5480 12884 5489
rect 12556 5440 12844 5480
rect 12076 5431 12116 5440
rect 12844 5431 12884 5440
rect 13996 5480 14036 5489
rect 14380 5480 14420 5767
rect 14036 5440 14132 5480
rect 13996 5431 14036 5440
rect 8140 5356 8468 5396
rect 7947 5228 7989 5237
rect 7947 5188 7948 5228
rect 7988 5188 7989 5228
rect 7947 5179 7989 5188
rect 7412 4936 7508 4976
rect 8044 5144 8084 5153
rect 7372 4927 7412 4936
rect 6124 4892 6164 4901
rect 6028 4852 6124 4892
rect 6124 4843 6164 4852
rect 6987 4472 7029 4481
rect 6987 4432 6988 4472
rect 7028 4432 7029 4472
rect 6987 4423 7029 4432
rect 6988 4145 7028 4423
rect 6987 4136 7029 4145
rect 3819 4096 3820 4136
rect 3860 4096 3861 4136
rect 3819 4087 3861 4096
rect 3916 4096 4340 4136
rect 5260 4096 5492 4136
rect 2612 3928 3092 3968
rect 2572 3919 2612 3928
rect 844 3632 884 3641
rect 3148 3632 3188 3641
rect 884 3592 1172 3632
rect 844 3583 884 3592
rect 1132 3380 1172 3592
rect 2956 3592 3148 3632
rect 1227 3464 1269 3473
rect 1227 3424 1228 3464
rect 1268 3424 1269 3464
rect 1227 3415 1269 3424
rect 1324 3464 1364 3473
rect 1611 3464 1653 3473
rect 1364 3424 1460 3464
rect 1324 3415 1364 3424
rect 1132 3331 1172 3340
rect 1228 2624 1268 3415
rect 1420 2633 1460 3424
rect 1611 3424 1612 3464
rect 1652 3424 1653 3464
rect 1611 3415 1653 3424
rect 1612 3330 1652 3415
rect 1228 2575 1268 2584
rect 1324 2624 1364 2633
rect 843 2456 885 2465
rect 843 2416 844 2456
rect 884 2416 885 2456
rect 1324 2456 1364 2584
rect 1419 2624 1461 2633
rect 1419 2584 1420 2624
rect 1460 2584 1461 2624
rect 2956 2624 2996 3592
rect 3148 3583 3188 3592
rect 3532 3632 3572 3641
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 3243 2876 3285 2885
rect 3243 2836 3244 2876
rect 3284 2836 3285 2876
rect 3243 2827 3285 2836
rect 3148 2624 3188 2633
rect 2956 2584 3148 2624
rect 1419 2575 1461 2584
rect 3148 2575 3188 2584
rect 3244 2624 3284 2827
rect 3244 2575 3284 2584
rect 1804 2456 1844 2465
rect 1324 2416 1804 2456
rect 843 2407 885 2416
rect 1804 2407 1844 2416
rect 2667 2456 2709 2465
rect 2667 2416 2668 2456
rect 2708 2416 2709 2456
rect 2667 2407 2709 2416
rect 844 2322 884 2407
rect 2668 2322 2708 2407
rect 844 2120 884 2129
rect 2860 2120 2900 2129
rect 884 2080 1172 2120
rect 844 2071 884 2080
rect 1132 1868 1172 2080
rect 1324 1952 1364 1961
rect 1612 1952 1652 1961
rect 1364 1912 1556 1952
rect 1324 1903 1364 1912
rect 1132 1819 1172 1828
rect 1227 1784 1269 1793
rect 1227 1744 1228 1784
rect 1268 1744 1269 1784
rect 1227 1735 1269 1744
rect 1419 1784 1461 1793
rect 1419 1744 1420 1784
rect 1460 1744 1461 1784
rect 1419 1735 1461 1744
rect 1228 1650 1268 1735
rect 843 1112 885 1121
rect 843 1072 844 1112
rect 884 1072 885 1112
rect 843 1063 885 1072
rect 1323 1112 1365 1121
rect 1323 1072 1324 1112
rect 1364 1072 1365 1112
rect 1323 1063 1365 1072
rect 1420 1112 1460 1735
rect 1420 1063 1460 1072
rect 844 944 884 1063
rect 1324 978 1364 1063
rect 1516 944 1556 1912
rect 1612 1793 1652 1912
rect 1611 1784 1653 1793
rect 1611 1744 1612 1784
rect 1652 1744 1653 1784
rect 1611 1735 1653 1744
rect 2860 1112 2900 2080
rect 2955 2120 2997 2129
rect 2955 2080 2956 2120
rect 2996 2080 2997 2120
rect 2955 2071 2997 2080
rect 3244 2120 3284 2129
rect 2956 1289 2996 2071
rect 3244 1700 3284 2080
rect 3532 1868 3572 3592
rect 3820 3548 3860 4087
rect 3820 3499 3860 3508
rect 3820 3380 3860 3389
rect 3916 3380 3956 4096
rect 4588 3968 4628 3977
rect 4204 3928 4588 3968
rect 4012 3464 4052 3473
rect 4204 3464 4244 3928
rect 4588 3919 4628 3928
rect 5163 3884 5205 3893
rect 5163 3844 5164 3884
rect 5204 3844 5205 3884
rect 5163 3835 5205 3844
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 4052 3424 4244 3464
rect 4780 3632 4820 3641
rect 4012 3415 4052 3424
rect 3860 3340 3956 3380
rect 3820 3331 3860 3340
rect 3723 2876 3765 2885
rect 3723 2836 3724 2876
rect 3764 2836 3765 2876
rect 3723 2827 3765 2836
rect 3724 2624 3764 2827
rect 4780 2717 4820 3592
rect 5164 3464 5204 3835
rect 5164 3415 5204 3424
rect 5260 3464 5300 4096
rect 5356 3968 5396 3977
rect 5452 3968 5492 4096
rect 6987 4096 6988 4136
rect 7028 4096 7029 4136
rect 6987 4087 7029 4096
rect 7084 4136 7124 4145
rect 5548 3968 5588 3977
rect 5452 3928 5548 3968
rect 5356 3800 5396 3928
rect 5548 3919 5588 3928
rect 6604 3968 6644 3977
rect 7084 3968 7124 4096
rect 7659 4136 7701 4145
rect 7659 4096 7660 4136
rect 7700 4096 7701 4136
rect 7659 4087 7701 4096
rect 7851 4136 7893 4145
rect 7851 4096 7852 4136
rect 7892 4096 7893 4136
rect 7851 4087 7893 4096
rect 7660 4002 7700 4087
rect 6644 3928 7124 3968
rect 6604 3919 6644 3928
rect 5739 3884 5781 3893
rect 5739 3844 5740 3884
rect 5780 3844 5781 3884
rect 5739 3835 5781 3844
rect 5356 3760 5588 3800
rect 5260 3415 5300 3424
rect 5356 3464 5396 3473
rect 5396 3424 5492 3464
rect 5356 3415 5396 3424
rect 5356 2717 5396 2802
rect 5452 2792 5492 3424
rect 5452 2743 5492 2752
rect 4779 2708 4821 2717
rect 4779 2668 4780 2708
rect 4820 2668 4821 2708
rect 4779 2659 4821 2668
rect 5355 2708 5397 2717
rect 5355 2668 5356 2708
rect 5396 2668 5397 2708
rect 5355 2659 5397 2668
rect 3628 2584 3724 2624
rect 3628 1952 3668 2584
rect 3724 2575 3764 2584
rect 5548 2624 5588 3760
rect 5740 3464 5780 3835
rect 7468 3632 7508 3641
rect 7468 3464 7508 3592
rect 7756 3464 7796 3473
rect 7468 3424 7756 3464
rect 5740 3415 5780 3424
rect 7756 3415 7796 3424
rect 7852 3464 7892 4087
rect 7852 3415 7892 3424
rect 7948 3380 7988 3389
rect 8044 3380 8084 5104
rect 8428 5144 8468 5356
rect 14092 5153 14132 5440
rect 14380 5431 14420 5440
rect 14764 5480 14804 5935
rect 15147 5648 15189 5657
rect 15147 5608 15148 5648
rect 15188 5608 15189 5648
rect 15147 5599 15189 5608
rect 14764 5431 14804 5440
rect 14859 5480 14901 5489
rect 14859 5440 14860 5480
rect 14900 5440 14901 5480
rect 14859 5431 14901 5440
rect 15148 5480 15188 5599
rect 15148 5431 15188 5440
rect 14379 5312 14421 5321
rect 14379 5272 14380 5312
rect 14420 5272 14421 5312
rect 14379 5263 14421 5272
rect 8428 5095 8468 5104
rect 10060 5144 10100 5153
rect 9388 4220 9428 4229
rect 10060 4220 10100 5104
rect 9428 4180 9524 4220
rect 9388 4171 9428 4180
rect 9196 4136 9236 4145
rect 8908 4096 9196 4136
rect 8908 3968 8948 4096
rect 9196 4087 9236 4096
rect 8908 3919 8948 3928
rect 9484 3632 9524 4180
rect 10060 4171 10100 4180
rect 11020 5144 11060 5153
rect 10252 4136 10292 4145
rect 11020 4136 11060 5104
rect 11212 5144 11252 5153
rect 11212 4220 11252 5104
rect 13996 5144 14036 5153
rect 13996 4985 14036 5104
rect 14091 5144 14133 5153
rect 14091 5104 14092 5144
rect 14132 5104 14133 5144
rect 14091 5095 14133 5104
rect 14380 5144 14420 5263
rect 14380 5095 14420 5104
rect 14764 5144 14804 5153
rect 14860 5144 14900 5431
rect 14804 5104 14900 5144
rect 15148 5144 15188 5153
rect 14764 5095 14804 5104
rect 13995 4976 14037 4985
rect 13995 4936 13996 4976
rect 14036 4936 14037 4976
rect 13995 4927 14037 4936
rect 15148 4817 15188 5104
rect 15147 4808 15189 4817
rect 15147 4768 15148 4808
rect 15188 4768 15189 4808
rect 15147 4759 15189 4768
rect 14763 4640 14805 4649
rect 14763 4600 14764 4640
rect 14804 4600 14805 4640
rect 14763 4591 14805 4600
rect 14379 4304 14421 4313
rect 14379 4264 14380 4304
rect 14420 4264 14421 4304
rect 14379 4255 14421 4264
rect 11212 4171 11252 4180
rect 12556 4220 12596 4229
rect 12364 4136 12404 4145
rect 10292 4096 10580 4136
rect 10252 4087 10292 4096
rect 10540 3968 10580 4096
rect 11020 4087 11060 4096
rect 12076 4096 12364 4136
rect 10540 3919 10580 3928
rect 12076 3968 12116 4096
rect 12364 4087 12404 4096
rect 12556 3968 12596 4180
rect 12844 3968 12884 3977
rect 12556 3928 12844 3968
rect 12076 3919 12116 3928
rect 12844 3919 12884 3928
rect 13996 3968 14036 3977
rect 13996 3809 14036 3928
rect 14380 3968 14420 4255
rect 14380 3919 14420 3928
rect 14764 3968 14804 4591
rect 15147 4472 15189 4481
rect 15147 4432 15148 4472
rect 15188 4432 15189 4472
rect 15147 4423 15189 4432
rect 14859 4136 14901 4145
rect 14859 4096 14860 4136
rect 14900 4096 14901 4136
rect 14859 4087 14901 4096
rect 14764 3919 14804 3928
rect 13995 3800 14037 3809
rect 13995 3760 13996 3800
rect 14036 3760 14037 3800
rect 13995 3751 14037 3760
rect 9484 3583 9524 3592
rect 10444 3632 10484 3641
rect 11212 3632 11252 3641
rect 10444 3464 10484 3592
rect 10924 3592 11212 3632
rect 10732 3464 10772 3473
rect 10444 3424 10732 3464
rect 10732 3415 10772 3424
rect 7988 3340 8084 3380
rect 10924 3380 10964 3592
rect 11212 3583 11252 3592
rect 12364 3632 12404 3641
rect 12748 3632 12788 3641
rect 7948 3331 7988 3340
rect 10924 3331 10964 3340
rect 6411 2792 6453 2801
rect 6411 2752 6412 2792
rect 6452 2752 6453 2792
rect 6411 2743 6453 2752
rect 7371 2792 7413 2801
rect 7371 2752 7372 2792
rect 7412 2752 7413 2792
rect 7371 2743 7413 2752
rect 5548 2575 5588 2584
rect 6027 2624 6069 2633
rect 6027 2584 6028 2624
rect 6068 2584 6069 2624
rect 6027 2575 6069 2584
rect 6412 2624 6452 2743
rect 6412 2575 6452 2584
rect 6507 2624 6549 2633
rect 6507 2584 6508 2624
rect 6548 2584 6549 2624
rect 6507 2575 6549 2584
rect 7372 2624 7412 2743
rect 9292 2708 9332 2717
rect 9100 2624 9140 2633
rect 7412 2584 7508 2624
rect 7372 2575 7412 2584
rect 3723 2456 3765 2465
rect 4876 2456 4916 2465
rect 3723 2416 3724 2456
rect 3764 2416 3765 2456
rect 3723 2407 3765 2416
rect 4780 2416 4876 2456
rect 3628 1903 3668 1912
rect 3724 1952 3764 2407
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 4491 2120 4533 2129
rect 4780 2120 4820 2416
rect 4876 2407 4916 2416
rect 6028 2456 6068 2575
rect 6508 2490 6548 2575
rect 6028 2407 6068 2416
rect 7180 2456 7220 2465
rect 7220 2416 7412 2456
rect 7180 2407 7220 2416
rect 4491 2080 4492 2120
rect 4532 2080 4533 2120
rect 4491 2071 4533 2080
rect 4588 2080 4820 2120
rect 5067 2120 5109 2129
rect 5836 2120 5876 2129
rect 6220 2120 6260 2129
rect 5067 2080 5068 2120
rect 5108 2080 5109 2120
rect 3724 1903 3764 1912
rect 4492 1952 4532 2071
rect 4492 1903 4532 1912
rect 4588 1952 4628 2080
rect 5067 2071 5109 2080
rect 5260 2080 5836 2120
rect 4588 1903 4628 1912
rect 5068 1952 5108 2071
rect 3532 1819 3572 1828
rect 3244 1660 3572 1700
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 2955 1280 2997 1289
rect 2955 1240 2956 1280
rect 2996 1240 3092 1280
rect 2955 1231 2997 1240
rect 2956 1112 2996 1121
rect 2860 1072 2956 1112
rect 2956 1063 2996 1072
rect 3052 1112 3092 1240
rect 3532 1205 3572 1660
rect 4107 1280 4149 1289
rect 4107 1240 4108 1280
rect 4148 1240 4149 1280
rect 4107 1231 4149 1240
rect 3531 1196 3573 1205
rect 3531 1156 3532 1196
rect 3572 1156 3573 1196
rect 3531 1147 3573 1156
rect 3052 1063 3092 1072
rect 4108 1112 4148 1231
rect 4396 1205 4436 1290
rect 5068 1289 5108 1912
rect 4491 1280 4533 1289
rect 4491 1240 4492 1280
rect 4532 1240 4533 1280
rect 4491 1231 4533 1240
rect 5067 1280 5109 1289
rect 5067 1240 5068 1280
rect 5108 1240 5109 1280
rect 5067 1231 5109 1240
rect 4395 1196 4437 1205
rect 4395 1156 4396 1196
rect 4436 1156 4437 1196
rect 4395 1147 4437 1156
rect 4492 1146 4532 1231
rect 5260 1196 5300 2080
rect 5836 2071 5876 2080
rect 5932 2080 6220 2120
rect 5355 1280 5397 1289
rect 5355 1240 5356 1280
rect 5396 1240 5397 1280
rect 5355 1231 5397 1240
rect 5260 1147 5300 1156
rect 5356 1146 5396 1231
rect 4108 1063 4148 1072
rect 4588 1112 4628 1121
rect 4588 953 4628 1072
rect 5452 1112 5492 1121
rect 5932 1112 5972 2080
rect 6220 2071 6260 2080
rect 7372 1868 7412 2416
rect 7468 1952 7508 2584
rect 8812 2584 9100 2624
rect 8140 2456 8180 2465
rect 7948 2416 8140 2456
rect 7468 1903 7508 1912
rect 7564 1952 7604 1961
rect 7948 1952 7988 2416
rect 8140 2407 8180 2416
rect 8812 2456 8852 2584
rect 9100 2575 9140 2584
rect 9292 2456 9332 2668
rect 10828 2708 10868 2717
rect 10636 2624 10676 2633
rect 10348 2584 10636 2624
rect 9580 2456 9620 2465
rect 9292 2416 9580 2456
rect 8812 2407 8852 2416
rect 9580 2407 9620 2416
rect 10348 2456 10388 2584
rect 10636 2575 10676 2584
rect 10348 2407 10388 2416
rect 8236 2120 8276 2129
rect 7604 1912 7988 1952
rect 8140 2080 8236 2120
rect 7564 1903 7604 1912
rect 7372 1819 7412 1828
rect 5492 1072 5972 1112
rect 6796 1196 6836 1205
rect 5452 1063 5492 1072
rect 1804 944 1844 953
rect 1516 904 1804 944
rect 844 895 884 904
rect 1804 895 1844 904
rect 2475 944 2517 953
rect 2475 904 2476 944
rect 2516 904 2517 944
rect 2475 895 2517 904
rect 4587 944 4629 953
rect 4587 904 4588 944
rect 4628 904 4629 944
rect 4587 895 4629 904
rect 6123 944 6165 953
rect 6123 904 6124 944
rect 6164 904 6165 944
rect 6123 895 6165 904
rect 6508 944 6548 953
rect 6796 944 6836 1156
rect 8140 1196 8180 2080
rect 8236 2071 8276 2080
rect 8908 2120 8948 2129
rect 8908 1196 8948 2080
rect 10828 2120 10868 2668
rect 12364 2624 12404 3592
rect 12652 3592 12748 3632
rect 12652 2708 12692 3592
rect 12748 3583 12788 3592
rect 13612 3632 13652 3641
rect 13612 2969 13652 3592
rect 13996 3632 14036 3641
rect 13996 3473 14036 3592
rect 14379 3632 14421 3641
rect 14379 3592 14380 3632
rect 14420 3592 14421 3632
rect 14379 3583 14421 3592
rect 14764 3632 14804 3641
rect 14860 3632 14900 4087
rect 15148 3968 15188 4423
rect 15148 3919 15188 3928
rect 15243 3968 15285 3977
rect 15243 3928 15244 3968
rect 15284 3928 15285 3968
rect 15243 3919 15285 3928
rect 14804 3592 14900 3632
rect 15148 3632 15188 3641
rect 15244 3632 15284 3919
rect 15188 3592 15284 3632
rect 14764 3583 14804 3592
rect 15148 3583 15188 3592
rect 14380 3498 14420 3583
rect 13995 3464 14037 3473
rect 13995 3424 13996 3464
rect 14036 3424 14037 3464
rect 13995 3415 14037 3424
rect 14571 3296 14613 3305
rect 14571 3256 14572 3296
rect 14612 3256 14613 3296
rect 14571 3247 14613 3256
rect 13611 2960 13653 2969
rect 13611 2920 13612 2960
rect 13652 2920 13653 2960
rect 13611 2911 13653 2920
rect 14187 2792 14229 2801
rect 14187 2752 14188 2792
rect 14228 2752 14229 2792
rect 14187 2743 14229 2752
rect 12652 2659 12692 2668
rect 12460 2624 12500 2633
rect 12364 2584 12460 2624
rect 12460 2575 12500 2584
rect 13803 2456 13845 2465
rect 13803 2416 13804 2456
rect 13844 2416 13845 2456
rect 13803 2407 13845 2416
rect 14188 2456 14228 2743
rect 14188 2407 14228 2416
rect 14572 2456 14612 3247
rect 14955 3128 14997 3137
rect 14955 3088 14956 3128
rect 14996 3088 14997 3128
rect 14955 3079 14997 3088
rect 14763 2624 14805 2633
rect 14763 2584 14764 2624
rect 14804 2584 14805 2624
rect 14763 2575 14805 2584
rect 14572 2407 14612 2416
rect 13804 2322 13844 2407
rect 10828 2071 10868 2080
rect 11020 2120 11060 2129
rect 11020 1364 11060 2080
rect 10732 1324 11060 1364
rect 11404 2120 11444 2129
rect 9004 1196 9044 1205
rect 8908 1156 9004 1196
rect 8140 1147 8180 1156
rect 9004 1147 9044 1156
rect 6988 1112 7028 1121
rect 7948 1112 7988 1121
rect 6988 953 7028 1072
rect 7660 1072 7948 1112
rect 6548 904 6836 944
rect 6987 944 7029 953
rect 6987 904 6988 944
rect 7028 904 7029 944
rect 6508 895 6548 904
rect 6987 895 7029 904
rect 7660 944 7700 1072
rect 7948 1063 7988 1072
rect 9196 1112 9236 1121
rect 9196 953 9236 1072
rect 10732 1112 10772 1324
rect 11404 1205 11444 2080
rect 11979 2120 12021 2129
rect 11979 2080 11980 2120
rect 12020 2080 12021 2120
rect 11979 2071 12021 2080
rect 12651 2120 12693 2129
rect 13132 2120 13172 2129
rect 12651 2080 12652 2120
rect 12692 2080 12693 2120
rect 12651 2071 12693 2080
rect 12844 2080 13132 2120
rect 11980 1986 12020 2071
rect 12652 1952 12692 2071
rect 12652 1903 12692 1912
rect 12844 1868 12884 2080
rect 13132 2071 13172 2080
rect 13996 2120 14036 2129
rect 12844 1819 12884 1828
rect 13996 1793 14036 2080
rect 14379 2120 14421 2129
rect 14379 2080 14380 2120
rect 14420 2080 14421 2120
rect 14379 2071 14421 2080
rect 14764 2120 14804 2575
rect 14956 2456 14996 3079
rect 14956 2407 14996 2416
rect 15147 2288 15189 2297
rect 15147 2248 15148 2288
rect 15188 2248 15189 2288
rect 15147 2239 15189 2248
rect 14764 2071 14804 2080
rect 15148 2120 15188 2239
rect 15148 2071 15188 2080
rect 14380 1986 14420 2071
rect 14763 1952 14805 1961
rect 14763 1912 14764 1952
rect 14804 1912 14805 1952
rect 14763 1903 14805 1912
rect 13995 1784 14037 1793
rect 13995 1744 13996 1784
rect 14036 1744 14037 1784
rect 13995 1735 14037 1744
rect 10923 1196 10965 1205
rect 10923 1156 10924 1196
rect 10964 1156 10965 1196
rect 10923 1147 10965 1156
rect 11403 1196 11445 1205
rect 11403 1156 11404 1196
rect 11444 1156 11445 1196
rect 11403 1147 11445 1156
rect 10732 1063 10772 1072
rect 10924 1062 10964 1147
rect 7660 895 7700 904
rect 8715 944 8757 953
rect 8715 904 8716 944
rect 8756 904 8757 944
rect 8715 895 8757 904
rect 9195 944 9237 953
rect 9195 904 9196 944
rect 9236 904 9237 944
rect 9195 895 9237 904
rect 14764 944 14804 1903
rect 15147 1616 15189 1625
rect 15147 1576 15148 1616
rect 15188 1576 15189 1616
rect 15147 1567 15189 1576
rect 14764 895 14804 904
rect 15148 944 15188 1567
rect 15148 895 15188 904
rect 2476 810 2516 895
rect 6124 810 6164 895
rect 8716 810 8756 895
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
<< via2 >>
rect 1420 12496 1460 12536
rect 1132 11824 1172 11864
rect 1420 11824 1460 11864
rect 1228 11656 1268 11696
rect 2092 11656 2132 11696
rect 1132 10480 1172 10520
rect 1708 10480 1748 10520
rect 1900 10480 1940 10520
rect 1708 10144 1748 10184
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 3052 11488 3092 11528
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3628 11488 3668 11528
rect 4588 12664 4628 12704
rect 5068 12664 5108 12704
rect 4012 12496 4052 12536
rect 5164 12496 5204 12536
rect 5164 12160 5204 12200
rect 6028 12496 6068 12536
rect 6124 11656 6164 11696
rect 6796 11656 6836 11696
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 13612 12160 13652 12200
rect 7372 11152 7412 11192
rect 4684 10816 4724 10856
rect 5356 10816 5396 10856
rect 3244 10732 3284 10772
rect 3628 10732 3668 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 3148 10228 3188 10268
rect 3532 10228 3572 10268
rect 2668 10144 2708 10184
rect 1420 9808 1460 9848
rect 1420 9472 1460 9512
rect 844 8716 884 8756
rect 1420 8716 1460 8756
rect 3244 9640 3284 9680
rect 1900 9472 1940 9512
rect 3724 10228 3764 10268
rect 3724 9976 3764 10016
rect 4492 9976 4532 10016
rect 8140 11152 8180 11192
rect 8524 11152 8564 11192
rect 5932 10816 5972 10856
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3820 9640 3860 9680
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 2476 8632 2516 8672
rect 2956 8632 2996 8672
rect 3628 8548 3668 8588
rect 1132 8128 1172 8168
rect 1132 7960 1172 8000
rect 2860 8464 2900 8504
rect 1708 8128 1748 8168
rect 2572 8128 2612 8168
rect 1516 7960 1556 8000
rect 1804 7960 1844 8000
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 2860 7204 2900 7244
rect 2476 7120 2516 7160
rect 2956 7120 2996 7160
rect 1036 6112 1076 6152
rect 1420 6112 1460 6152
rect 1612 6112 1652 6152
rect 4780 9388 4820 9428
rect 6220 9472 6260 9512
rect 6700 9472 6740 9512
rect 5164 9388 5204 9428
rect 3916 8632 3956 8672
rect 6796 9388 6836 9428
rect 6796 9136 6836 9176
rect 7180 9388 7220 9428
rect 13996 11992 14036 12032
rect 14380 11824 14420 11864
rect 13996 11488 14036 11528
rect 13804 10816 13844 10856
rect 14380 10984 14420 11024
rect 14188 10480 14228 10520
rect 8908 8800 8948 8840
rect 9292 8800 9332 8840
rect 8332 8632 8372 8672
rect 8812 8632 8852 8672
rect 12556 10228 12596 10268
rect 13228 10228 13268 10268
rect 15148 11656 15188 11696
rect 14860 11320 14900 11360
rect 14764 10648 14804 10688
rect 15148 11152 15188 11192
rect 14956 10312 14996 10352
rect 14572 10144 14612 10184
rect 13996 9808 14036 9848
rect 13612 9472 13652 9512
rect 13996 9304 14036 9344
rect 14476 9640 14516 9680
rect 15148 9976 15188 10016
rect 14860 9136 14900 9176
rect 15148 8968 15188 9008
rect 14764 8800 14804 8840
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3628 7708 3668 7748
rect 3916 7708 3956 7748
rect 3724 7204 3764 7244
rect 6028 7960 6068 8000
rect 6508 7960 6548 8000
rect 6604 7876 6644 7916
rect 4684 6952 4724 6992
rect 14380 8632 14420 8672
rect 7180 8128 7220 8168
rect 7756 8128 7796 8168
rect 6988 7876 7028 7916
rect 13996 8464 14036 8504
rect 14380 8296 14420 8336
rect 14380 7792 14420 7832
rect 14860 7960 14900 8000
rect 14764 7624 14804 7664
rect 8908 7456 8948 7496
rect 9292 7456 9332 7496
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 8332 7120 8372 7160
rect 8812 7120 8852 7160
rect 5548 6952 5588 6992
rect 5164 6700 5204 6740
rect 5356 6700 5396 6740
rect 5548 6700 5588 6740
rect 4588 6448 4628 6488
rect 5068 6448 5108 6488
rect 12556 7204 12596 7244
rect 13228 7204 13268 7244
rect 12364 6952 12404 6992
rect 12844 6952 12884 6992
rect 14188 7120 14228 7160
rect 13804 6952 13844 6992
rect 15244 8128 15284 8168
rect 15148 7456 15188 7496
rect 14956 7288 14996 7328
rect 13516 6784 13556 6824
rect 6796 6532 6836 6572
rect 7276 6532 7316 6572
rect 8332 6532 8372 6572
rect 7372 6448 7412 6488
rect 7852 6448 7892 6488
rect 14764 6448 14804 6488
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 2860 5776 2900 5816
rect 3820 5776 3860 5816
rect 2476 5608 2516 5648
rect 2956 5608 2996 5648
rect 1900 5104 1940 5144
rect 2572 5104 2612 5144
rect 1132 4768 1172 4808
rect 1804 4768 1844 4808
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 2956 4096 2996 4136
rect 5452 5440 5492 5480
rect 5452 5020 5492 5060
rect 14380 6280 14420 6320
rect 15244 6616 15284 6656
rect 15148 6112 15188 6152
rect 14764 5944 14804 5984
rect 14380 5776 14420 5816
rect 8236 5692 8276 5732
rect 9292 5692 9332 5732
rect 7948 5608 7988 5648
rect 7276 5188 7316 5228
rect 6124 5020 6164 5060
rect 8524 5608 8564 5648
rect 7948 5188 7988 5228
rect 6988 4432 7028 4472
rect 3820 4096 3860 4136
rect 1228 3424 1268 3464
rect 1612 3424 1652 3464
rect 844 2416 884 2456
rect 1420 2584 1460 2624
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 3244 2836 3284 2876
rect 2668 2416 2708 2456
rect 1228 1744 1268 1784
rect 1420 1744 1460 1784
rect 844 1072 884 1112
rect 1324 1072 1364 1112
rect 1612 1744 1652 1784
rect 2956 2080 2996 2120
rect 5164 3844 5204 3884
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 3724 2836 3764 2876
rect 6988 4096 7028 4136
rect 7660 4096 7700 4136
rect 7852 4096 7892 4136
rect 5740 3844 5780 3884
rect 4780 2668 4820 2708
rect 5356 2668 5396 2708
rect 15148 5608 15188 5648
rect 14860 5440 14900 5480
rect 14380 5272 14420 5312
rect 14092 5104 14132 5144
rect 13996 4936 14036 4976
rect 15148 4768 15188 4808
rect 14764 4600 14804 4640
rect 14380 4264 14420 4304
rect 15148 4432 15188 4472
rect 14860 4096 14900 4136
rect 13996 3760 14036 3800
rect 6412 2752 6452 2792
rect 7372 2752 7412 2792
rect 6028 2584 6068 2624
rect 6508 2584 6548 2624
rect 3724 2416 3764 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 4492 2080 4532 2120
rect 5068 2080 5108 2120
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 2956 1240 2996 1280
rect 4108 1240 4148 1280
rect 3532 1156 3572 1196
rect 4492 1240 4532 1280
rect 5068 1240 5108 1280
rect 4396 1156 4436 1196
rect 5356 1240 5396 1280
rect 2476 904 2516 944
rect 4588 904 4628 944
rect 6124 904 6164 944
rect 14380 3592 14420 3632
rect 15244 3928 15284 3968
rect 13996 3424 14036 3464
rect 14572 3256 14612 3296
rect 13612 2920 13652 2960
rect 14188 2752 14228 2792
rect 13804 2416 13844 2456
rect 14956 3088 14996 3128
rect 14764 2584 14804 2624
rect 6988 904 7028 944
rect 11980 2080 12020 2120
rect 12652 2080 12692 2120
rect 14380 2080 14420 2120
rect 15148 2248 15188 2288
rect 14764 1912 14804 1952
rect 13996 1744 14036 1784
rect 10924 1156 10964 1196
rect 11404 1156 11444 1196
rect 8716 904 8756 944
rect 9196 904 9236 944
rect 15148 1576 15188 1616
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
<< metal3 >>
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 4579 12664 4588 12704
rect 4628 12664 5068 12704
rect 5108 12664 5117 12704
rect 1411 12496 1420 12536
rect 1460 12496 4012 12536
rect 4052 12496 4061 12536
rect 5155 12496 5164 12536
rect 5204 12496 6028 12536
rect 6068 12496 6077 12536
rect 0 12200 80 12220
rect 15920 12200 16000 12220
rect 0 12160 5164 12200
rect 5204 12160 5213 12200
rect 13603 12160 13612 12200
rect 13652 12160 16000 12200
rect 0 12140 80 12160
rect 15920 12140 16000 12160
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 15920 12032 16000 12052
rect 13987 11992 13996 12032
rect 14036 11992 16000 12032
rect 15920 11972 16000 11992
rect 0 11864 80 11884
rect 15920 11864 16000 11884
rect 0 11824 1132 11864
rect 1172 11824 1420 11864
rect 1460 11824 1469 11864
rect 14371 11824 14380 11864
rect 14420 11824 16000 11864
rect 0 11804 80 11824
rect 15920 11804 16000 11824
rect 15920 11696 16000 11716
rect 1219 11656 1228 11696
rect 1268 11656 2092 11696
rect 2132 11656 2141 11696
rect 6115 11656 6124 11696
rect 6164 11656 6796 11696
rect 6836 11656 6845 11696
rect 15139 11656 15148 11696
rect 15188 11656 16000 11696
rect 15920 11636 16000 11656
rect 0 11528 80 11548
rect 15920 11528 16000 11548
rect 0 11488 3052 11528
rect 3092 11488 3628 11528
rect 3668 11488 3677 11528
rect 13987 11488 13996 11528
rect 14036 11488 16000 11528
rect 0 11468 80 11488
rect 15920 11468 16000 11488
rect 15920 11360 16000 11380
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 14851 11320 14860 11360
rect 14900 11320 16000 11360
rect 15920 11300 16000 11320
rect 0 11192 80 11212
rect 15920 11192 16000 11212
rect 0 11152 7372 11192
rect 7412 11152 8140 11192
rect 8180 11152 8524 11192
rect 8564 11152 8573 11192
rect 15139 11152 15148 11192
rect 15188 11152 16000 11192
rect 0 11132 80 11152
rect 15920 11132 16000 11152
rect 15920 11024 16000 11044
rect 14371 10984 14380 11024
rect 14420 10984 16000 11024
rect 15920 10964 16000 10984
rect 0 10856 80 10876
rect 15920 10856 16000 10876
rect 0 10816 4684 10856
rect 4724 10816 5356 10856
rect 5396 10816 5932 10856
rect 5972 10816 5981 10856
rect 13795 10816 13804 10856
rect 13844 10816 16000 10856
rect 0 10796 80 10816
rect 15920 10796 16000 10816
rect 3235 10732 3244 10772
rect 3284 10732 3628 10772
rect 3668 10732 3677 10772
rect 15920 10688 16000 10708
rect 14755 10648 14764 10688
rect 14804 10648 16000 10688
rect 15920 10628 16000 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 0 10520 80 10540
rect 15920 10520 16000 10540
rect 0 10480 1132 10520
rect 1172 10480 1708 10520
rect 1748 10480 1900 10520
rect 1940 10480 1949 10520
rect 14179 10480 14188 10520
rect 14228 10480 16000 10520
rect 0 10460 80 10480
rect 15920 10460 16000 10480
rect 15920 10352 16000 10372
rect 14947 10312 14956 10352
rect 14996 10312 16000 10352
rect 15920 10292 16000 10312
rect 1612 10228 3148 10268
rect 3188 10228 3532 10268
rect 3572 10228 3724 10268
rect 3764 10228 3773 10268
rect 12547 10228 12556 10268
rect 12596 10228 13228 10268
rect 13268 10228 13277 10268
rect 0 10184 80 10204
rect 1612 10184 1652 10228
rect 15920 10184 16000 10204
rect 0 10144 1652 10184
rect 1699 10144 1708 10184
rect 1748 10144 2668 10184
rect 2708 10144 2717 10184
rect 14563 10144 14572 10184
rect 14612 10144 16000 10184
rect 0 10124 80 10144
rect 15920 10124 16000 10144
rect 15920 10016 16000 10036
rect 3715 9976 3724 10016
rect 3764 9976 4492 10016
rect 4532 9976 4541 10016
rect 15139 9976 15148 10016
rect 15188 9976 16000 10016
rect 15920 9956 16000 9976
rect 0 9848 80 9868
rect 15920 9848 16000 9868
rect 0 9808 1420 9848
rect 1460 9808 1469 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 13987 9808 13996 9848
rect 14036 9808 16000 9848
rect 0 9788 80 9808
rect 15920 9788 16000 9808
rect 15920 9680 16000 9700
rect 3235 9640 3244 9680
rect 3284 9640 3820 9680
rect 3860 9640 3869 9680
rect 14467 9640 14476 9680
rect 14516 9640 16000 9680
rect 15920 9620 16000 9640
rect 0 9512 80 9532
rect 15920 9512 16000 9532
rect 0 9472 1364 9512
rect 1411 9472 1420 9512
rect 1460 9472 1900 9512
rect 1940 9472 1949 9512
rect 6211 9472 6220 9512
rect 6260 9472 6700 9512
rect 6740 9472 6749 9512
rect 13603 9472 13612 9512
rect 13652 9472 16000 9512
rect 0 9452 80 9472
rect 1324 9428 1364 9472
rect 15920 9452 16000 9472
rect 1324 9388 4780 9428
rect 4820 9388 5164 9428
rect 5204 9388 5213 9428
rect 6787 9388 6796 9428
rect 6836 9388 7180 9428
rect 7220 9388 7229 9428
rect 15920 9344 16000 9364
rect 13987 9304 13996 9344
rect 14036 9304 16000 9344
rect 15920 9284 16000 9304
rect 0 9176 80 9196
rect 15920 9176 16000 9196
rect 0 9136 6796 9176
rect 6836 9136 6845 9176
rect 14851 9136 14860 9176
rect 14900 9136 16000 9176
rect 0 9116 80 9136
rect 15920 9116 16000 9136
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 15920 9008 16000 9028
rect 15139 8968 15148 9008
rect 15188 8968 16000 9008
rect 15920 8948 16000 8968
rect 0 8840 80 8860
rect 15920 8840 16000 8860
rect 0 8800 8908 8840
rect 8948 8800 9292 8840
rect 9332 8800 9341 8840
rect 14755 8800 14764 8840
rect 14804 8800 16000 8840
rect 0 8780 80 8800
rect 15920 8780 16000 8800
rect 835 8716 844 8756
rect 884 8716 1420 8756
rect 1460 8716 1469 8756
rect 15920 8672 16000 8692
rect 2467 8632 2476 8672
rect 2516 8632 2956 8672
rect 2996 8632 3005 8672
rect 3907 8632 3916 8672
rect 3956 8632 3965 8672
rect 8323 8632 8332 8672
rect 8372 8632 8812 8672
rect 8852 8632 8861 8672
rect 14371 8632 14380 8672
rect 14420 8632 16000 8672
rect 3916 8588 3956 8632
rect 15920 8612 16000 8632
rect 2860 8548 3628 8588
rect 3668 8548 3956 8588
rect 0 8504 80 8524
rect 2860 8504 2900 8548
rect 15920 8504 16000 8524
rect 0 8464 2860 8504
rect 2900 8464 2909 8504
rect 13987 8464 13996 8504
rect 14036 8464 16000 8504
rect 0 8444 80 8464
rect 15920 8444 16000 8464
rect 15920 8336 16000 8356
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 14371 8296 14380 8336
rect 14420 8296 16000 8336
rect 15920 8276 16000 8296
rect 0 8168 80 8188
rect 15920 8168 16000 8188
rect 0 8128 1132 8168
rect 1172 8128 1181 8168
rect 1699 8128 1708 8168
rect 1748 8128 2572 8168
rect 2612 8128 2621 8168
rect 7171 8128 7180 8168
rect 7220 8128 7756 8168
rect 7796 8128 7805 8168
rect 15235 8128 15244 8168
rect 15284 8128 16000 8168
rect 0 8108 80 8128
rect 15920 8108 16000 8128
rect 15920 8000 16000 8020
rect 1123 7960 1132 8000
rect 1172 7960 1516 8000
rect 1556 7960 1804 8000
rect 1844 7960 1853 8000
rect 6019 7960 6028 8000
rect 6068 7960 6508 8000
rect 6548 7960 6557 8000
rect 14851 7960 14860 8000
rect 14900 7960 16000 8000
rect 15920 7940 16000 7960
rect 6280 7876 6604 7916
rect 6644 7876 6988 7916
rect 7028 7876 7037 7916
rect 0 7832 80 7852
rect 6280 7832 6320 7876
rect 15920 7832 16000 7852
rect 0 7792 6320 7832
rect 14371 7792 14380 7832
rect 14420 7792 16000 7832
rect 0 7772 80 7792
rect 15920 7772 16000 7792
rect 3619 7708 3628 7748
rect 3668 7708 3916 7748
rect 3956 7708 3965 7748
rect 15920 7664 16000 7684
rect 14755 7624 14764 7664
rect 14804 7624 16000 7664
rect 15920 7604 16000 7624
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 0 7496 80 7516
rect 15920 7496 16000 7516
rect 0 7456 8908 7496
rect 8948 7456 9292 7496
rect 9332 7456 9341 7496
rect 15139 7456 15148 7496
rect 15188 7456 16000 7496
rect 0 7436 80 7456
rect 15920 7436 16000 7456
rect 15920 7328 16000 7348
rect 14947 7288 14956 7328
rect 14996 7288 16000 7328
rect 15920 7268 16000 7288
rect 2380 7204 2860 7244
rect 2900 7204 3724 7244
rect 3764 7204 3773 7244
rect 12547 7204 12556 7244
rect 12596 7204 13228 7244
rect 13268 7204 13277 7244
rect 0 7160 80 7180
rect 2380 7160 2420 7204
rect 15920 7160 16000 7180
rect 0 7120 2420 7160
rect 2467 7120 2476 7160
rect 2516 7120 2956 7160
rect 2996 7120 3005 7160
rect 8323 7120 8332 7160
rect 8372 7120 8812 7160
rect 8852 7120 8861 7160
rect 14179 7120 14188 7160
rect 14228 7120 16000 7160
rect 0 7100 80 7120
rect 15920 7100 16000 7120
rect 15920 6992 16000 7012
rect 4675 6952 4684 6992
rect 4724 6952 5548 6992
rect 5588 6952 5597 6992
rect 12355 6952 12364 6992
rect 12404 6952 12844 6992
rect 12884 6952 12893 6992
rect 13795 6952 13804 6992
rect 13844 6952 16000 6992
rect 15920 6932 16000 6952
rect 0 6824 80 6844
rect 15920 6824 16000 6844
rect 0 6784 4244 6824
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 13507 6784 13516 6824
rect 13556 6784 16000 6824
rect 0 6764 80 6784
rect 4204 6740 4244 6784
rect 15920 6764 16000 6784
rect 4204 6700 5164 6740
rect 5204 6700 5356 6740
rect 5396 6700 5548 6740
rect 5588 6700 5597 6740
rect 15920 6656 16000 6676
rect 15235 6616 15244 6656
rect 15284 6616 16000 6656
rect 15920 6596 16000 6616
rect 2284 6532 6796 6572
rect 6836 6532 7276 6572
rect 7316 6532 8332 6572
rect 8372 6532 8381 6572
rect 0 6488 80 6508
rect 2284 6488 2324 6532
rect 15920 6488 16000 6508
rect 0 6448 2324 6488
rect 4579 6448 4588 6488
rect 4628 6448 5068 6488
rect 5108 6448 5117 6488
rect 7363 6448 7372 6488
rect 7412 6448 7852 6488
rect 7892 6448 7901 6488
rect 14755 6448 14764 6488
rect 14804 6448 16000 6488
rect 0 6428 80 6448
rect 15920 6428 16000 6448
rect 15920 6320 16000 6340
rect 14340 6280 14380 6320
rect 14420 6280 14429 6320
rect 15532 6280 16000 6320
rect 14380 6236 14420 6280
rect 15532 6236 15572 6280
rect 15920 6260 16000 6280
rect 14380 6196 15572 6236
rect 0 6152 80 6172
rect 15920 6152 16000 6172
rect 0 6112 1036 6152
rect 1076 6112 1420 6152
rect 1460 6112 1612 6152
rect 1652 6112 1661 6152
rect 15139 6112 15148 6152
rect 15188 6112 16000 6152
rect 0 6092 80 6112
rect 15920 6092 16000 6112
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 15920 5984 16000 6004
rect 14755 5944 14764 5984
rect 14804 5944 16000 5984
rect 15920 5924 16000 5944
rect 0 5816 80 5836
rect 15920 5816 16000 5836
rect 0 5776 2860 5816
rect 2900 5776 3820 5816
rect 3860 5776 3869 5816
rect 14371 5776 14380 5816
rect 14420 5776 16000 5816
rect 0 5756 80 5776
rect 15920 5756 16000 5776
rect 8227 5692 8236 5732
rect 8276 5692 9292 5732
rect 9332 5692 9341 5732
rect 15920 5648 16000 5668
rect 2467 5608 2476 5648
rect 2516 5608 2956 5648
rect 2996 5608 3005 5648
rect 7939 5608 7948 5648
rect 7988 5608 8524 5648
rect 8564 5608 8573 5648
rect 15139 5608 15148 5648
rect 15188 5608 16000 5648
rect 15920 5588 16000 5608
rect 0 5480 80 5500
rect 15920 5480 16000 5500
rect 0 5440 5452 5480
rect 5492 5440 5501 5480
rect 14851 5440 14860 5480
rect 14900 5440 16000 5480
rect 0 5420 80 5440
rect 15920 5420 16000 5440
rect 15920 5312 16000 5332
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 14371 5272 14380 5312
rect 14420 5272 16000 5312
rect 15920 5252 16000 5272
rect 1804 5188 7276 5228
rect 7316 5188 7948 5228
rect 7988 5188 7997 5228
rect 0 5144 80 5164
rect 1804 5144 1844 5188
rect 15920 5144 16000 5164
rect 0 5104 1844 5144
rect 1891 5104 1900 5144
rect 1940 5104 2572 5144
rect 2612 5104 2621 5144
rect 14083 5104 14092 5144
rect 14132 5104 16000 5144
rect 0 5084 80 5104
rect 15920 5084 16000 5104
rect 5443 5020 5452 5060
rect 5492 5020 6124 5060
rect 6164 5020 6173 5060
rect 15920 4976 16000 4996
rect 13987 4936 13996 4976
rect 14036 4936 16000 4976
rect 15920 4916 16000 4936
rect 0 4808 80 4828
rect 15920 4808 16000 4828
rect 0 4768 1132 4808
rect 1172 4768 1804 4808
rect 1844 4768 1853 4808
rect 15139 4768 15148 4808
rect 15188 4768 16000 4808
rect 0 4748 80 4768
rect 15920 4748 16000 4768
rect 15920 4640 16000 4660
rect 14755 4600 14764 4640
rect 14804 4600 16000 4640
rect 15920 4580 16000 4600
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 0 4472 80 4492
rect 15920 4472 16000 4492
rect 0 4432 6988 4472
rect 7028 4432 7037 4472
rect 15139 4432 15148 4472
rect 15188 4432 16000 4472
rect 0 4412 80 4432
rect 15920 4412 16000 4432
rect 15920 4304 16000 4324
rect 14371 4264 14380 4304
rect 14420 4264 16000 4304
rect 15920 4244 16000 4264
rect 0 4136 80 4156
rect 15920 4136 16000 4156
rect 0 4096 2956 4136
rect 2996 4096 3820 4136
rect 3860 4096 3869 4136
rect 6979 4096 6988 4136
rect 7028 4096 7660 4136
rect 7700 4096 7852 4136
rect 7892 4096 7901 4136
rect 14851 4096 14860 4136
rect 14900 4096 16000 4136
rect 0 4076 80 4096
rect 15920 4076 16000 4096
rect 15920 3968 16000 3988
rect 15235 3928 15244 3968
rect 15284 3928 16000 3968
rect 15920 3908 16000 3928
rect 4204 3844 5164 3884
rect 5204 3844 5740 3884
rect 5780 3844 5789 3884
rect 0 3800 80 3820
rect 4204 3800 4244 3844
rect 15920 3800 16000 3820
rect 0 3760 4244 3800
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 13987 3760 13996 3800
rect 14036 3760 16000 3800
rect 0 3740 80 3760
rect 15920 3740 16000 3760
rect 15920 3632 16000 3652
rect 14371 3592 14380 3632
rect 14420 3592 16000 3632
rect 15920 3572 16000 3592
rect 0 3464 80 3484
rect 15920 3464 16000 3484
rect 0 3424 1228 3464
rect 1268 3424 1612 3464
rect 1652 3424 1661 3464
rect 13987 3424 13996 3464
rect 14036 3424 16000 3464
rect 0 3404 80 3424
rect 15920 3404 16000 3424
rect 15920 3296 16000 3316
rect 14563 3256 14572 3296
rect 14612 3256 16000 3296
rect 15920 3236 16000 3256
rect 0 3128 80 3148
rect 15920 3128 16000 3148
rect 0 3088 2996 3128
rect 14947 3088 14956 3128
rect 14996 3088 16000 3128
rect 0 3068 80 3088
rect 2956 2876 2996 3088
rect 15920 3068 16000 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 15920 2960 16000 2980
rect 13603 2920 13612 2960
rect 13652 2920 16000 2960
rect 15920 2900 16000 2920
rect 2956 2836 3244 2876
rect 3284 2836 3724 2876
rect 3764 2836 3773 2876
rect 0 2792 80 2812
rect 15920 2792 16000 2812
rect 0 2752 6412 2792
rect 6452 2752 7372 2792
rect 7412 2752 7421 2792
rect 14179 2752 14188 2792
rect 14228 2752 16000 2792
rect 0 2732 80 2752
rect 15920 2732 16000 2752
rect 4771 2668 4780 2708
rect 4820 2668 5356 2708
rect 5396 2668 5405 2708
rect 15920 2624 16000 2644
rect 1411 2584 1420 2624
rect 1460 2584 1469 2624
rect 6019 2584 6028 2624
rect 6068 2584 6508 2624
rect 6548 2584 6557 2624
rect 14755 2584 14764 2624
rect 14804 2584 16000 2624
rect 0 2456 80 2476
rect 1420 2456 1460 2584
rect 15920 2564 16000 2584
rect 15920 2456 16000 2476
rect 0 2416 788 2456
rect 835 2416 844 2456
rect 884 2416 1460 2456
rect 2659 2416 2668 2456
rect 2708 2416 3724 2456
rect 3764 2416 3773 2456
rect 13795 2416 13804 2456
rect 13844 2416 16000 2456
rect 0 2396 80 2416
rect 748 2204 788 2416
rect 15920 2396 16000 2416
rect 15920 2288 16000 2308
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 15139 2248 15148 2288
rect 15188 2248 16000 2288
rect 15920 2228 16000 2248
rect 748 2164 4532 2204
rect 0 2120 80 2140
rect 4492 2120 4532 2164
rect 15920 2120 16000 2140
rect 0 2080 2956 2120
rect 2996 2080 3005 2120
rect 4483 2080 4492 2120
rect 4532 2080 5068 2120
rect 5108 2080 5117 2120
rect 11971 2080 11980 2120
rect 12020 2080 12652 2120
rect 12692 2080 12701 2120
rect 14371 2080 14380 2120
rect 14420 2080 16000 2120
rect 0 2060 80 2080
rect 15920 2060 16000 2080
rect 15920 1952 16000 1972
rect 14755 1912 14764 1952
rect 14804 1912 16000 1952
rect 15920 1892 16000 1912
rect 0 1784 80 1804
rect 15920 1784 16000 1804
rect 0 1744 1228 1784
rect 1268 1744 1420 1784
rect 1460 1744 1612 1784
rect 1652 1744 1661 1784
rect 13987 1744 13996 1784
rect 14036 1744 16000 1784
rect 0 1724 80 1744
rect 15920 1724 16000 1744
rect 15920 1616 16000 1636
rect 15139 1576 15148 1616
rect 15188 1576 16000 1616
rect 15920 1556 16000 1576
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 2947 1240 2956 1280
rect 2996 1240 4108 1280
rect 4148 1240 4492 1280
rect 4532 1240 4541 1280
rect 5059 1240 5068 1280
rect 5108 1240 5356 1280
rect 5396 1240 5405 1280
rect 3523 1156 3532 1196
rect 3572 1156 4396 1196
rect 4436 1156 4445 1196
rect 10915 1156 10924 1196
rect 10964 1156 11404 1196
rect 11444 1156 11453 1196
rect 835 1072 844 1112
rect 884 1072 1324 1112
rect 1364 1072 1373 1112
rect 2467 904 2476 944
rect 2516 904 4588 944
rect 4628 904 4637 944
rect 6115 904 6124 944
rect 6164 904 6988 944
rect 7028 904 7037 944
rect 8707 904 8716 944
rect 8756 904 9196 944
rect 9236 904 9245 944
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
<< via3 >>
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
<< metal4 >>
rect 3076 12116 3516 12896
rect 3076 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3516 12116
rect 3076 10604 3516 12076
rect 3076 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3516 10604
rect 3076 9092 3516 10564
rect 3076 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3516 9092
rect 3076 7580 3516 9052
rect 3076 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3516 7580
rect 3076 6068 3516 7540
rect 3076 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3516 6068
rect 3076 4556 3516 6028
rect 3076 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3516 4556
rect 3076 3640 3516 4516
rect 3076 3600 3132 3640
rect 3172 3600 3228 3640
rect 3268 3600 3324 3640
rect 3364 3600 3420 3640
rect 3460 3600 3516 3640
rect 3076 3544 3516 3600
rect 3076 3504 3132 3544
rect 3172 3504 3228 3544
rect 3268 3504 3324 3544
rect 3364 3504 3420 3544
rect 3460 3504 3516 3544
rect 3076 3448 3516 3504
rect 3076 3408 3132 3448
rect 3172 3408 3228 3448
rect 3268 3408 3324 3448
rect 3364 3408 3420 3448
rect 3460 3408 3516 3448
rect 3076 3352 3516 3408
rect 3076 3312 3132 3352
rect 3172 3312 3228 3352
rect 3268 3312 3324 3352
rect 3364 3312 3420 3352
rect 3460 3312 3516 3352
rect 3076 3044 3516 3312
rect 3076 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3516 3044
rect 3076 1532 3516 3004
rect 3076 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3516 1532
rect 3076 712 3516 1492
rect 4316 12872 4756 12896
rect 4316 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4756 12872
rect 4316 11360 4756 12832
rect 4316 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4756 11360
rect 4316 9848 4756 11320
rect 4316 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4756 9848
rect 4316 8336 4756 9808
rect 4316 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4756 8336
rect 4316 6824 4756 8296
rect 4316 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4756 6824
rect 4316 5312 4756 6784
rect 4316 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4756 5312
rect 4316 4880 4756 5272
rect 4316 4840 4372 4880
rect 4412 4840 4468 4880
rect 4508 4840 4564 4880
rect 4604 4840 4660 4880
rect 4700 4840 4756 4880
rect 4316 4784 4756 4840
rect 4316 4744 4372 4784
rect 4412 4744 4468 4784
rect 4508 4744 4564 4784
rect 4604 4744 4660 4784
rect 4700 4744 4756 4784
rect 4316 4688 4756 4744
rect 4316 4648 4372 4688
rect 4412 4648 4468 4688
rect 4508 4648 4564 4688
rect 4604 4648 4660 4688
rect 4700 4648 4756 4688
rect 4316 4592 4756 4648
rect 4316 4552 4372 4592
rect 4412 4552 4468 4592
rect 4508 4552 4564 4592
rect 4604 4552 4660 4592
rect 4700 4552 4756 4592
rect 4316 3800 4756 4552
rect 4316 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4756 3800
rect 4316 2288 4756 3760
rect 4316 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4756 2288
rect 4316 776 4756 2248
rect 4316 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4756 776
rect 4316 712 4756 736
<< via4 >>
rect 3132 3600 3172 3640
rect 3228 3600 3268 3640
rect 3324 3600 3364 3640
rect 3420 3600 3460 3640
rect 3132 3504 3172 3544
rect 3228 3504 3268 3544
rect 3324 3504 3364 3544
rect 3420 3504 3460 3544
rect 3132 3408 3172 3448
rect 3228 3408 3268 3448
rect 3324 3408 3364 3448
rect 3420 3408 3460 3448
rect 3132 3312 3172 3352
rect 3228 3312 3268 3352
rect 3324 3312 3364 3352
rect 3420 3312 3460 3352
rect 4372 4840 4412 4880
rect 4468 4840 4508 4880
rect 4564 4840 4604 4880
rect 4660 4840 4700 4880
rect 4372 4744 4412 4784
rect 4468 4744 4508 4784
rect 4564 4744 4604 4784
rect 4660 4744 4700 4784
rect 4372 4648 4412 4688
rect 4468 4648 4508 4688
rect 4564 4648 4604 4688
rect 4660 4648 4700 4688
rect 4372 4552 4412 4592
rect 4468 4552 4508 4592
rect 4564 4552 4604 4592
rect 4660 4552 4700 4592
<< metal5 >>
rect 532 4880 15404 4936
rect 532 4840 4372 4880
rect 4412 4840 4468 4880
rect 4508 4840 4564 4880
rect 4604 4840 4660 4880
rect 4700 4840 15404 4880
rect 532 4784 15404 4840
rect 532 4744 4372 4784
rect 4412 4744 4468 4784
rect 4508 4744 4564 4784
rect 4604 4744 4660 4784
rect 4700 4744 15404 4784
rect 532 4688 15404 4744
rect 532 4648 4372 4688
rect 4412 4648 4468 4688
rect 4508 4648 4564 4688
rect 4604 4648 4660 4688
rect 4700 4648 15404 4688
rect 532 4592 15404 4648
rect 532 4552 4372 4592
rect 4412 4552 4468 4592
rect 4508 4552 4564 4592
rect 4604 4552 4660 4592
rect 4700 4552 15404 4592
rect 532 4496 15404 4552
rect 532 3640 15404 3696
rect 532 3600 3132 3640
rect 3172 3600 3228 3640
rect 3268 3600 3324 3640
rect 3364 3600 3420 3640
rect 3460 3600 15404 3640
rect 532 3544 15404 3600
rect 532 3504 3132 3544
rect 3172 3504 3228 3544
rect 3268 3504 3324 3544
rect 3364 3504 3420 3544
rect 3460 3504 15404 3544
rect 532 3448 15404 3504
rect 532 3408 3132 3448
rect 3172 3408 3228 3448
rect 3268 3408 3324 3448
rect 3364 3408 3420 3448
rect 3460 3408 15404 3448
rect 532 3352 15404 3408
rect 532 3312 3132 3352
rect 3172 3312 3228 3352
rect 3268 3312 3324 3352
rect 3364 3312 3420 3352
rect 3460 3312 15404 3352
rect 532 3256 15404 3312
use sg13g2_tielo  _224_
timestamp 1584750033
transform -1 0 11328 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _225_
timestamp 1584750033
transform 1 0 10176 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _226_
timestamp 1584750033
transform 1 0 576 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _227_
timestamp 1584750033
transform -1 0 2112 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _228_
timestamp 1584750033
transform 1 0 576 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _229_
timestamp 1584750033
transform -1 0 13056 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _230_
timestamp 1584750033
transform 1 0 11712 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _231_
timestamp 1584750033
transform -1 0 9600 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _232_
timestamp 1584750033
transform -1 0 8736 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _233_
timestamp 1584750033
transform -1 0 7776 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _234_
timestamp 1584750033
transform -1 0 11520 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _235_
timestamp 1584750033
transform 1 0 10176 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _236_
timestamp 1584750033
transform 1 0 5760 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _237_
timestamp 1584750033
transform 1 0 5376 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _238_
timestamp 1584750033
transform 1 0 4992 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _239_
timestamp 1584750033
transform -1 0 11328 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _240_
timestamp 1584750033
transform -1 0 11808 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _241_
timestamp 1584750033
transform 1 0 3360 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _242_
timestamp 1584750033
transform -1 0 4896 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _243_
timestamp 1584750033
transform 1 0 2208 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _244_
timestamp 1584750033
transform -1 0 11232 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _245_
timestamp 1584750033
transform 1 0 9888 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _246_
timestamp 1584750033
transform -1 0 2688 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _247_
timestamp 1584750033
transform 1 0 864 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _248_
timestamp 1584750033
transform 1 0 576 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _249_
timestamp 1584750033
transform -1 0 11232 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _250_
timestamp 1584750033
transform -1 0 11712 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _251_
timestamp 1584750033
transform -1 0 7392 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _252_
timestamp 1584750033
transform -1 0 7776 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _253_
timestamp 1584750033
transform -1 0 8160 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _254_
timestamp 1584750033
transform 1 0 9216 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _255_
timestamp 1584750033
transform 1 0 8640 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _256_
timestamp 1584750033
transform 1 0 4800 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _257_
timestamp 1584750033
transform 1 0 4416 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _258_
timestamp 1584750033
transform 1 0 4320 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _259_
timestamp 1584750033
transform 1 0 7968 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _260_
timestamp 1584750033
transform 1 0 7392 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _261_
timestamp 1584750033
transform -1 0 4512 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _262_
timestamp 1584750033
transform 1 0 3168 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _263_
timestamp 1584750033
transform 1 0 2208 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _264_
timestamp 1584750033
transform 1 0 10368 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _265_
timestamp 1584750033
transform 1 0 9888 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _266_
timestamp 1584750033
transform -1 0 9600 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _267_
timestamp 1584750033
transform 1 0 8256 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _268_
timestamp 1584750033
transform 1 0 8064 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _269_
timestamp 1584750033
transform -1 0 10368 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _270_
timestamp 1584750033
transform 1 0 9024 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _271_
timestamp 1584750033
transform -1 0 8064 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _272_
timestamp 1584750033
transform 1 0 6528 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _273_
timestamp 1584750033
transform 1 0 5760 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _274_
timestamp 1584750033
transform -1 0 13536 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _275_
timestamp 1584750033
transform 1 0 11808 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _276_
timestamp 1584750033
transform -1 0 2880 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _277_
timestamp 1584750033
transform 1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _278_
timestamp 1584750033
transform 1 0 864 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _279_
timestamp 1584750033
transform -1 0 13056 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _280_
timestamp 1584750033
transform -1 0 12672 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _281_
timestamp 1584750033
transform 1 0 2976 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _282_
timestamp 1584750033
transform 1 0 2208 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _283_
timestamp 1584750033
transform 1 0 2592 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _284_
timestamp 1584750033
transform -1 0 11520 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _285_
timestamp 1584750033
transform 1 0 10752 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _286_
timestamp 1584750033
transform 1 0 3456 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _287_
timestamp 1584750033
transform 1 0 2976 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _288_
timestamp 1584750033
transform 1 0 2208 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _289_
timestamp 1584750033
transform -1 0 9792 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _290_
timestamp 1584750033
transform 1 0 8448 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _291_
timestamp 1584750033
transform -1 0 9600 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _292_
timestamp 1584750033
transform 1 0 8256 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _293_
timestamp 1584750033
transform 1 0 8064 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _294_
timestamp 1584750033
transform -1 0 12096 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _295_
timestamp 1584750033
transform 1 0 11328 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _296_
timestamp 1584750033
transform 1 0 7104 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _297_
timestamp 1584750033
transform 1 0 6720 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _298_
timestamp 1584750033
transform 1 0 5952 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _299_
timestamp 1584750033
transform -1 0 11232 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _300_
timestamp 1584750033
transform 1 0 9888 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _301_
timestamp 1584750033
transform -1 0 5472 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _302_
timestamp 1584750033
transform 1 0 4128 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _303_
timestamp 1584750033
transform -1 0 6048 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _304_
timestamp 1584750033
transform 1 0 6240 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _305_
timestamp 1584750033
transform 1 0 5856 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _306_
timestamp 1584750033
transform 1 0 576 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _307_
timestamp 1584750033
transform 1 0 1152 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _308_
timestamp 1584750033
transform 1 0 768 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _309_
timestamp 1584750033
transform -1 0 13536 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _310_
timestamp 1584750033
transform -1 0 13152 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _311_
timestamp 1584750033
transform 1 0 2976 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _312_
timestamp 1584750033
transform -1 0 4800 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _313_
timestamp 1584750033
transform 1 0 2496 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _314_
timestamp 1584750033
transform -1 0 10368 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _315_
timestamp 1584750033
transform -1 0 10848 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _316_
timestamp 1584750033
transform 1 0 1728 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _317_
timestamp 1584750033
transform -1 0 2976 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _318_
timestamp 1584750033
transform 1 0 864 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _319_
timestamp 1584750033
transform 1 0 10560 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _320_
timestamp 1584750033
transform 1 0 10080 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _321_
timestamp 1584750033
transform -1 0 5472 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _322_
timestamp 1584750033
transform 1 0 4128 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _323_
timestamp 1584750033
transform -1 0 5952 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _324_
timestamp 1584750033
transform -1 0 11712 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _325_
timestamp 1584750033
transform -1 0 11328 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _326_
timestamp 1584750033
transform -1 0 8064 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _327_
timestamp 1584750033
transform 1 0 6720 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _328_
timestamp 1584750033
transform 1 0 7296 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _329_
timestamp 1584750033
transform -1 0 13152 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _330_
timestamp 1584750033
transform 1 0 11808 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _331_
timestamp 1584750033
transform 1 0 3552 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _332_
timestamp 1584750033
transform 1 0 2784 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _333_
timestamp 1584750033
transform -1 0 3552 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _334_
timestamp 1584750033
transform -1 0 9888 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _335_
timestamp 1584750033
transform 1 0 8544 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _336_
timestamp 1584750033
transform -1 0 6144 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _337_
timestamp 1584750033
transform -1 0 6528 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _338_
timestamp 1584750033
transform -1 0 5184 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _339_
timestamp 1584750033
transform -1 0 13248 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _340_
timestamp 1584750033
transform 1 0 11904 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _341_
timestamp 1584750033
transform -1 0 2496 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _342_
timestamp 1584750033
transform -1 0 4320 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _343_
timestamp 1584750033
transform -1 0 2496 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _344_
timestamp 1584750033
transform -1 0 11520 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _345_
timestamp 1584750033
transform 1 0 10176 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _346_
timestamp 1584750033
transform 1 0 5568 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _347_
timestamp 1584750033
transform -1 0 7104 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _348_
timestamp 1584750033
transform 1 0 4320 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _349_
timestamp 1584750033
transform -1 0 13440 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _350_
timestamp 1584750033
transform 1 0 11712 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _351_
timestamp 1584750033
transform 1 0 6912 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _352_
timestamp 1584750033
transform -1 0 8448 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _353_
timestamp 1584750033
transform 1 0 5760 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _354_
timestamp 1584750033
transform -1 0 12960 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _355_
timestamp 1584750033
transform -1 0 12576 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _356_
timestamp 1584750033
transform 1 0 3264 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _357_
timestamp 1584750033
transform 1 0 2400 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _358_
timestamp 1584750033
transform 1 0 2880 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _359_
timestamp 1584750033
transform 1 0 10560 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _360_
timestamp 1584750033
transform 1 0 9984 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _361_
timestamp 1584750033
transform 1 0 576 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _362_
timestamp 1584750033
transform 1 0 576 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _363_
timestamp 1584750033
transform -1 0 2112 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _364_
timestamp 1584750033
transform -1 0 12960 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _365_
timestamp 1584750033
transform 1 0 11616 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _366_
timestamp 1584750033
transform 1 0 4512 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _367_
timestamp 1584750033
transform 1 0 5088 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _368_
timestamp 1584750033
transform -1 0 5856 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _369_
timestamp 1584750033
transform -1 0 13152 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _370_
timestamp 1584750033
transform 1 0 11808 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _371_
timestamp 1584750033
transform -1 0 4608 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _372_
timestamp 1584750033
transform -1 0 4896 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _373_
timestamp 1584750033
transform 1 0 2304 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _374_
timestamp 1584750033
transform 1 0 8640 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _375_
timestamp 1584750033
transform 1 0 8448 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _376_
timestamp 1584750033
transform 1 0 7776 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _377_
timestamp 1584750033
transform 1 0 7200 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _378_
timestamp 1584750033
transform 1 0 6336 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _379_
timestamp 1584750033
transform -1 0 10080 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _380_
timestamp 1584750033
transform 1 0 9312 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _381_
timestamp 1584750033
transform -1 0 2880 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _382_
timestamp 1584750033
transform 1 0 1152 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _383_
timestamp 1584750033
transform 1 0 768 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _384_
timestamp 1584750033
transform 1 0 14880 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _385_
timestamp 1584750033
transform 1 0 14496 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _386_
timestamp 1584750033
transform 1 0 14880 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _387_
timestamp 1584750033
transform 1 0 14496 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _388_
timestamp 1584750033
transform 1 0 13344 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _389_
timestamp 1584750033
transform 1 0 14304 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _390_
timestamp 1584750033
transform 1 0 14112 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _391_
timestamp 1584750033
transform 1 0 14880 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _392_
timestamp 1584750033
transform 1 0 14112 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _393_
timestamp 1584750033
transform 1 0 14496 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _394_
timestamp 1584750033
transform 1 0 13728 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _395_
timestamp 1584750033
transform 1 0 14112 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _396_
timestamp 1584750033
transform 1 0 14880 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _397_
timestamp 1584750033
transform 1 0 14496 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _398_
timestamp 1584750033
transform 1 0 14112 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _399_
timestamp 1584750033
transform 1 0 14880 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _400_
timestamp 1584750033
transform 1 0 13536 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _401_
timestamp 1584750033
transform 1 0 14496 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _402_
timestamp 1584750033
transform 1 0 14496 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _403_
timestamp 1584750033
transform 1 0 14496 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _404_
timestamp 1584750033
transform 1 0 14112 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _405_
timestamp 1584750033
transform 1 0 14112 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _406_
timestamp 1584750033
transform 1 0 14880 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _407_
timestamp 1584750033
transform 1 0 13728 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _408_
timestamp 1584750033
transform 1 0 14112 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _409_
timestamp 1584750033
transform 1 0 14880 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _410_
timestamp 1584750033
transform 1 0 14688 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _411_
timestamp 1584750033
transform 1 0 14496 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _412_
timestamp 1584750033
transform 1 0 14112 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _413_
timestamp 1584750033
transform 1 0 14496 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _414_
timestamp 1584750033
transform 1 0 14880 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _415_
timestamp 1584750033
transform 1 0 13728 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _416_
timestamp 1584750033
transform 1 0 13728 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _417_
timestamp 1584750033
transform 1 0 14112 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _418_
timestamp 1584750033
transform 1 0 13536 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _419_
timestamp 1584750033
transform 1 0 13920 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _420_
timestamp 1584750033
transform 1 0 14688 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _421_
timestamp 1584750033
transform 1 0 13728 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _422_
timestamp 1584750033
transform 1 0 13728 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _423_
timestamp 1584750033
transform 1 0 14496 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _424_
timestamp 1584750033
transform 1 0 14880 0 1 3780
box -48 -56 432 834
use sg13g2_tielo  _425_
timestamp 1584750033
transform 1 0 14880 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _426_
timestamp 1584750033
transform 1 0 13728 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _427_
timestamp 1584750033
transform 1 0 14496 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _428_
timestamp 1584750033
transform 1 0 14112 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _429_
timestamp 1584750033
transform 1 0 14880 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _430_
timestamp 1584750033
transform 1 0 14496 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _431_
timestamp 1584750033
transform 1 0 13248 0 -1 6804
box -48 -56 432 834
use sg13g2_tielo  _432_
timestamp 1584750033
transform 1 0 13920 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _433_
timestamp 1584750033
transform 1 0 14880 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _434_
timestamp 1584750033
transform 1 0 14112 0 -1 8316
box -48 -56 432 834
use sg13g2_tielo  _435_
timestamp 1584750033
transform 1 0 14880 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _436_
timestamp 1584750033
transform 1 0 13728 0 1 8316
box -48 -56 432 834
use sg13g2_tielo  _437_
timestamp 1584750033
transform 1 0 14496 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _438_
timestamp 1584750033
transform 1 0 14496 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _439_
timestamp 1584750033
transform 1 0 13344 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _440_
timestamp 1584750033
transform 1 0 13728 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _441_
timestamp 1584750033
transform 1 0 14304 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _442_
timestamp 1584750033
transform 1 0 13920 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _443_
timestamp 1584750033
transform 1 0 13536 0 -1 11340
box -48 -56 432 834
use sg13g2_tielo  _444_
timestamp 1584750033
transform 1 0 14880 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _445_
timestamp 1584750033
transform 1 0 13728 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _446_
timestamp 1584750033
transform 1 0 14112 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _447_
timestamp 1584750033
transform 1 0 13344 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _448_
timestamp 1584750033
transform -1 0 10176 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _449_
timestamp 1584750033
transform -1 0 9408 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _450_
timestamp 1584750033
transform -1 0 12384 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _451_
timestamp 1584750033
transform -1 0 9024 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _452_
timestamp 1584750033
transform -1 0 12768 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _453_
timestamp 1584750033
transform -1 0 13248 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _454_
timestamp 1584750033
transform -1 0 11136 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _455_
timestamp 1584750033
transform -1 0 12384 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _456_
timestamp 1584750033
transform -1 0 10560 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _457_
timestamp 1584750033
transform -1 0 10560 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _458_
timestamp 1584750033
transform -1 0 12480 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _459_
timestamp 1584750033
transform -1 0 7104 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _460_
timestamp 1584750033
transform -1 0 11616 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _461_
timestamp 1584750033
transform -1 0 10176 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _462_
timestamp 1584750033
transform -1 0 13056 0 1 11340
box -48 -56 432 834
use sg13g2_tielo  _463_
timestamp 1584750033
transform -1 0 13536 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _464_
timestamp 1584750033
transform -1 0 13152 0 1 9828
box -48 -56 432 834
use sg13g2_tielo  _465_
timestamp 1584750033
transform -1 0 13920 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _466_
timestamp 1584750033
transform -1 0 7872 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _467_
timestamp 1584750033
transform -1 0 11904 0 1 6804
box -48 -56 432 834
use sg13g2_tielo  _468_
timestamp 1584750033
transform -1 0 14304 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _469_
timestamp 1584750033
transform -1 0 12480 0 -1 2268
box -48 -56 432 834
use sg13g2_tielo  _470_
timestamp 1584750033
transform -1 0 8256 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _471_
timestamp 1584750033
transform -1 0 9216 0 -1 3780
box -48 -56 432 834
use sg13g2_tielo  _472_
timestamp 1584750033
transform -1 0 12288 0 1 2268
box -48 -56 432 834
use sg13g2_tielo  _473_
timestamp 1584750033
transform -1 0 11616 0 1 5292
box -48 -56 432 834
use sg13g2_tielo  _474_
timestamp 1584750033
transform -1 0 8640 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _475_
timestamp 1584750033
transform -1 0 13152 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _476_
timestamp 1584750033
transform -1 0 10656 0 -1 12852
box -48 -56 432 834
use sg13g2_tielo  _477_
timestamp 1584750033
transform -1 0 9792 0 1 756
box -48 -56 432 834
use sg13g2_tielo  _478_
timestamp 1584750033
transform -1 0 12864 0 -1 5292
box -48 -56 432 834
use sg13g2_tielo  _479_
timestamp 1584750033
transform -1 0 11424 0 1 2268
box -48 -56 432 834
use sg13g2_dlygate4sd1_1  comb_logic\[0\].delay1_I
timestamp 1584750033
transform 1 0 1536 0 -1 2268
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[0\].nand_on_I
timestamp 1584750033
transform 1 0 10560 0 -1 8316
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[0\].nand_on_n_I
timestamp 1584750033
transform -1 0 1536 0 -1 2268
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[0\].xor_pulse_I
timestamp 1584750033
transform 1 0 960 0 1 756
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[1\].delay1_I
timestamp 1584750033
transform -1 0 4224 0 1 756
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[1\].nand_on_I
timestamp 1584750033
transform 1 0 12288 0 1 2268
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[1\].nand_on_n_I
timestamp 1584750033
transform -1 0 4800 0 1 756
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[1\].xor_pulse_I
timestamp 1584750033
transform 1 0 2592 0 1 756
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[2\].delay1_I
timestamp 1584750033
transform 1 0 4992 0 -1 2268
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[2\].nand_on_I
timestamp 1584750033
transform 1 0 8928 0 1 2268
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[2\].nand_on_n_I
timestamp 1584750033
transform -1 0 5664 0 1 756
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[2\].xor_pulse_I
timestamp 1584750033
transform -1 0 4992 0 -1 2268
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[3\].delay1_I
timestamp 1584750033
transform 1 0 7296 0 1 2268
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[3\].nand_on_I
timestamp 1584750033
transform 1 0 12480 0 -1 2268
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[3\].nand_on_n_I
timestamp 1584750033
transform -1 0 7776 0 -1 2268
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[3\].xor_pulse_I
timestamp 1584750033
transform 1 0 6144 0 1 2268
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[4\].delay1_I
timestamp 1584750033
transform 1 0 3648 0 1 2268
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[4\].nand_on_I
timestamp 1584750033
transform 1 0 12192 0 -1 8316
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[4\].nand_on_n_I
timestamp 1584750033
transform -1 0 3936 0 -1 2268
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[4\].xor_pulse_I
timestamp 1584750033
transform 1 0 2784 0 1 2268
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[5\].delay1_I
timestamp 1584750033
transform 1 0 1536 0 -1 3780
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[5\].nand_on_I
timestamp 1584750033
transform 1 0 10368 0 1 8316
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[5\].nand_on_n_I
timestamp 1584750033
transform -1 0 1536 0 -1 3780
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[5\].xor_pulse_I
timestamp 1584750033
transform -1 0 1728 0 1 2268
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[6\].delay1_I
timestamp 1584750033
transform 1 0 5664 0 -1 3780
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[6\].nand_on_I
timestamp 1584750033
transform 1 0 12000 0 -1 6804
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[6\].nand_on_n_I
timestamp 1584750033
transform -1 0 5760 0 1 2268
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[6\].xor_pulse_I
timestamp 1584750033
transform -1 0 5664 0 -1 3780
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[7\].delay1_I
timestamp 1584750033
transform 1 0 3744 0 1 3780
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[7\].nand_on_I
timestamp 1584750033
transform 1 0 12192 0 1 5292
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[7\].nand_on_n_I
timestamp 1584750033
transform -1 0 4224 0 -1 3780
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[7\].xor_pulse_I
timestamp 1584750033
transform 1 0 2688 0 1 3780
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[8\].delay1_I
timestamp 1584750033
transform 1 0 7584 0 1 3780
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[8\].nand_on_I
timestamp 1584750033
transform -1 0 9408 0 1 756
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[8\].nand_on_n_I
timestamp 1584750033
transform 1 0 7584 0 -1 3780
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[8\].xor_pulse_I
timestamp 1584750033
transform 1 0 6720 0 1 3780
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[9\].delay1_I
timestamp 1584750033
transform 1 0 1728 0 -1 5292
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[9\].nand_on_I
timestamp 1584750033
transform 1 0 9408 0 1 11340
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[9\].nand_on_n_I
timestamp 1584750033
transform 1 0 1536 0 1 3780
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[9\].xor_pulse_I
timestamp 1584750033
transform 1 0 864 0 -1 5292
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[10\].delay1_I
timestamp 1584750033
transform 1 0 8448 0 1 5292
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[10\].nand_on_I
timestamp 1584750033
transform 1 0 12096 0 -1 9828
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[10\].nand_on_n_I
timestamp 1584750033
transform 1 0 7872 0 1 5292
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[10\].xor_pulse_I
timestamp 1584750033
transform -1 0 7776 0 -1 5292
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[11\].delay1_I
timestamp 1584750033
transform 1 0 6144 0 1 5292
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[11\].nand_on_I
timestamp 1584750033
transform 1 0 10560 0 -1 3780
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[11\].nand_on_n_I
timestamp 1584750033
transform 1 0 5760 0 -1 5292
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[11\].xor_pulse_I
timestamp 1584750033
transform 1 0 4992 0 -1 5292
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[12\].delay1_I
timestamp 1584750033
transform 1 0 3744 0 1 5292
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[12\].nand_on_I
timestamp 1584750033
transform -1 0 11424 0 1 9828
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[12\].nand_on_n_I
timestamp 1584750033
transform -1 0 4224 0 -1 5292
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[12\].xor_pulse_I
timestamp 1584750033
transform 1 0 2592 0 1 5292
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[13\].delay1_I
timestamp 1584750033
transform 1 0 1536 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[13\].nand_on_I
timestamp 1584750033
transform 1 0 10272 0 -1 6804
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[13\].nand_on_n_I
timestamp 1584750033
transform 1 0 1248 0 1 5292
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[13\].xor_pulse_I
timestamp 1584750033
transform 1 0 768 0 -1 6804
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[14\].delay1_I
timestamp 1584750033
transform 1 0 8256 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[14\].nand_on_I
timestamp 1584750033
transform -1 0 11328 0 -1 11340
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[14\].nand_on_n_I
timestamp 1584750033
transform 1 0 6432 0 -1 6804
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[14\].xor_pulse_I
timestamp 1584750033
transform -1 0 7776 0 -1 6804
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[15\].delay1_I
timestamp 1584750033
transform 1 0 5472 0 -1 6804
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[15\].nand_on_I
timestamp 1584750033
transform 1 0 9024 0 1 3780
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[15\].nand_on_n_I
timestamp 1584750033
transform -1 0 5760 0 1 6804
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[15\].xor_pulse_I
timestamp 1584750033
transform 1 0 4704 0 -1 6804
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[16\].delay1_I
timestamp 1584750033
transform 1 0 3648 0 1 6804
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[16\].nand_on_I
timestamp 1584750033
transform 1 0 7776 0 1 756
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[16\].nand_on_n_I
timestamp 1584750033
transform 1 0 3456 0 -1 6804
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[16\].xor_pulse_I
timestamp 1584750033
transform 1 0 2592 0 1 6804
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[17\].delay1_I
timestamp 1584750033
transform 1 0 9216 0 1 6804
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[17\].nand_on_I
timestamp 1584750033
transform 1 0 10272 0 1 9828
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[17\].nand_on_n_I
timestamp 1584750033
transform 1 0 8640 0 -1 8316
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[17\].xor_pulse_I
timestamp 1584750033
transform 1 0 8448 0 1 6804
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[18\].delay1_I
timestamp 1584750033
transform 1 0 6912 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[18\].nand_on_I
timestamp 1584750033
transform 1 0 9504 0 -1 11340
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[18\].nand_on_n_I
timestamp 1584750033
transform 1 0 6816 0 1 6804
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[18\].xor_pulse_I
timestamp 1584750033
transform 1 0 6144 0 -1 8316
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[19\].delay1_I
timestamp 1584750033
transform 1 0 1728 0 -1 8316
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[19\].nand_on_I
timestamp 1584750033
transform 1 0 12192 0 1 9828
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[19\].nand_on_n_I
timestamp 1584750033
transform 1 0 1344 0 1 6804
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[19\].xor_pulse_I
timestamp 1584750033
transform 1 0 864 0 -1 8316
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[20\].delay1_I
timestamp 1584750033
transform 1 0 3840 0 1 8316
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[20\].nand_on_I
timestamp 1584750033
transform 1 0 10848 0 1 3780
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[20\].nand_on_n_I
timestamp 1584750033
transform -1 0 4128 0 -1 8316
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[20\].xor_pulse_I
timestamp 1584750033
transform 1 0 2592 0 1 8316
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[21\].delay1_I
timestamp 1584750033
transform 1 0 9216 0 1 8316
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[21\].nand_on_I
timestamp 1584750033
transform 1 0 8832 0 1 9828
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[21\].nand_on_n_I
timestamp 1584750033
transform 1 0 8640 0 -1 9828
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[21\].xor_pulse_I
timestamp 1584750033
transform 1 0 8448 0 1 8316
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[22\].delay1_I
timestamp 1584750033
transform 1 0 7104 0 -1 9828
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[22\].nand_on_I
timestamp 1584750033
transform 1 0 11424 0 1 11340
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[22\].nand_on_n_I
timestamp 1584750033
transform 1 0 6912 0 1 8316
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[22\].xor_pulse_I
timestamp 1584750033
transform 1 0 6336 0 -1 9828
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[23\].delay1_I
timestamp 1584750033
transform 1 0 5088 0 -1 9828
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[23\].nand_on_I
timestamp 1584750033
transform 1 0 10272 0 1 5292
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[23\].nand_on_n_I
timestamp 1584750033
transform 1 0 4512 0 -1 9828
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[23\].xor_pulse_I
timestamp 1584750033
transform -1 0 5664 0 1 8316
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[24\].delay1_I
timestamp 1584750033
transform 1 0 1824 0 -1 9828
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[24\].nand_on_I
timestamp 1584750033
transform -1 0 7200 0 1 756
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[24\].nand_on_n_I
timestamp 1584750033
transform -1 0 1824 0 1 8316
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[24\].xor_pulse_I
timestamp 1584750033
transform 1 0 960 0 -1 9828
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[25\].delay1_I
timestamp 1584750033
transform 1 0 3648 0 1 9828
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[25\].nand_on_I
timestamp 1584750033
transform 1 0 12192 0 1 6804
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[25\].nand_on_n_I
timestamp 1584750033
transform -1 0 3936 0 -1 9828
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[25\].xor_pulse_I
timestamp 1584750033
transform 1 0 2880 0 1 9828
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[26\].delay1_I
timestamp 1584750033
transform 1 0 1824 0 -1 11340
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[26\].nand_on_I
timestamp 1584750033
transform -1 0 10464 0 1 3780
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[26\].nand_on_n_I
timestamp 1584750033
transform 1 0 1536 0 1 9828
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[26\].xor_pulse_I
timestamp 1584750033
transform 1 0 864 0 -1 11340
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[27\].delay1_I
timestamp 1584750033
transform 1 0 5856 0 -1 11340
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[27\].nand_on_I
timestamp 1584750033
transform 1 0 10464 0 1 2268
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[27\].nand_on_n_I
timestamp 1584750033
transform 1 0 4512 0 -1 11340
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[27\].xor_pulse_I
timestamp 1584750033
transform -1 0 5856 0 -1 11340
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[28\].delay1_I
timestamp 1584750033
transform 1 0 8448 0 -1 11340
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[28\].nand_on_I
timestamp 1584750033
transform 1 0 10560 0 1 756
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[28\].nand_on_n_I
timestamp 1584750033
transform 1 0 7104 0 1 11340
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[28\].xor_pulse_I
timestamp 1584750033
transform 1 0 7680 0 -1 11340
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[29\].delay1_I
timestamp 1584750033
transform 1 0 3552 0 1 11340
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[29\].nand_on_I
timestamp 1584750033
transform 1 0 12192 0 1 3780
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[29\].nand_on_n_I
timestamp 1584750033
transform 1 0 3360 0 -1 11340
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[29\].xor_pulse_I
timestamp 1584750033
transform -1 0 3552 0 1 11340
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[30\].delay1_I
timestamp 1584750033
transform 1 0 1824 0 -1 12852
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[30\].nand_on_I
timestamp 1584750033
transform 1 0 12288 0 -1 11340
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[30\].nand_on_n_I
timestamp 1584750033
transform 1 0 1248 0 -1 12852
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[30\].xor_pulse_I
timestamp 1584750033
transform -1 0 1632 0 1 11340
box -48 -56 816 834
use sg13g2_dlygate4sd1_1  comb_logic\[31\].delay1_I
timestamp 1584750033
transform 1 0 5952 0 -1 12852
box -48 -56 816 834
use sg13g2_nand2_2  comb_logic\[31\].nand_on_I
timestamp 1584750033
transform 1 0 10560 0 1 6804
box -48 -56 624 834
use sg13g2_nand2_2  comb_logic\[31\].nand_on_n_I
timestamp 1584750033
transform -1 0 6336 0 1 11340
box -48 -56 624 834
use sg13g2_xnor2_1  comb_logic\[31\].xor_pulse_I
timestamp 1584750033
transform 1 0 4704 0 -1 12852
box -48 -56 816 834
use sg13g2_fill_1  FILLER_0_16
timestamp 1584750033
transform 1 0 2112 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_29
timestamp 1584750033
transform 1 0 3360 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_44
timestamp 1584750033
transform 1 0 4800 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_46
timestamp 1584750033
transform 1 0 4992 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_53
timestamp 1584750033
transform 1 0 5664 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_69
timestamp 1584750033
transform 1 0 7200 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_81
timestamp 1584750033
transform 1 0 8352 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_110
timestamp 1584750033
transform 1 0 11136 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_115
timestamp 1584750033
transform 1 0 11616 0 1 756
box -48 -56 432 834
use sg13g2_decap_4  FILLER_0_123
timestamp 1584750033
transform 1 0 12384 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_0_127
timestamp 1584750033
transform 1 0 12768 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_132
timestamp 1584750033
transform 1 0 13248 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_134
timestamp 1584750033
transform 1 0 13440 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_143
timestamp 1584750033
transform 1 0 14304 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_153
timestamp 1584750033
transform 1 0 15264 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_18
timestamp 1584750033
transform 1 0 2304 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_20
timestamp 1584750033
transform 1 0 2496 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_35
timestamp 1584750033
transform 1 0 3936 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_37
timestamp 1584750033
transform 1 0 4128 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_62
timestamp 1584750033
transform 1 0 6528 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_68
timestamp 1584750033
transform 1 0 7104 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_75
timestamp 1584750033
transform 1 0 7776 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_81
timestamp 1584750033
transform 1 0 8352 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_83
timestamp 1584750033
transform 1 0 8544 0 -1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_92
timestamp 1584750033
transform 1 0 9408 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_99
timestamp 1584750033
transform 1 0 10080 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_134
timestamp 1584750033
transform 1 0 13440 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_136
timestamp 1584750033
transform 1 0 13632 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_153
timestamp 1584750033
transform 1 0 15264 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_16
timestamp 1584750033
transform 1 0 2112 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_18
timestamp 1584750033
transform 1 0 2304 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_31
timestamp 1584750033
transform 1 0 3552 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_40
timestamp 1584750033
transform 1 0 4416 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_82
timestamp 1584750033
transform 1 0 8448 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_97
timestamp 1584750033
transform 1 0 9888 0 1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_2_113
timestamp 1584750033
transform 1 0 11424 0 1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_2_117
timestamp 1584750033
transform 1 0 11808 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_128
timestamp 1584750033
transform 1 0 12864 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_151
timestamp 1584750033
transform 1 0 15072 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_153
timestamp 1584750033
transform 1 0 15264 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_18
timestamp 1584750033
transform 1 0 2304 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_22
timestamp 1584750033
transform 1 0 2688 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_38
timestamp 1584750033
transform 1 0 4224 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_40
timestamp 1584750033
transform 1 0 4416 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_61
timestamp 1584750033
transform 1 0 6432 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_68
timestamp 1584750033
transform 1 0 7104 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_79
timestamp 1584750033
transform 1 0 8160 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_94
timestamp 1584750033
transform 1 0 9600 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_114
timestamp 1584750033
transform 1 0 11520 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_121
timestamp 1584750033
transform 1 0 12192 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_130
timestamp 1584750033
transform 1 0 13056 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_132
timestamp 1584750033
transform 1 0 13248 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_153
timestamp 1584750033
transform 1 0 15264 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_0
timestamp 1584750033
transform 1 0 576 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_16
timestamp 1584750033
transform 1 0 2112 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_30
timestamp 1584750033
transform 1 0 3456 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_32
timestamp 1584750033
transform 1 0 3648 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_45
timestamp 1584750033
transform 1 0 4896 0 1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_55
timestamp 1584750033
transform 1 0 5856 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_59
timestamp 1584750033
transform 1 0 6240 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_72
timestamp 1584750033
transform 1 0 7488 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_81
timestamp 1584750033
transform 1 0 8352 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_83
timestamp 1584750033
transform 1 0 8544 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_94
timestamp 1584750033
transform 1 0 9600 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_96
timestamp 1584750033
transform 1 0 9792 0 1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_4_113
timestamp 1584750033
transform 1 0 11424 0 1 3780
box -48 -56 432 834
use sg13g2_decap_4  FILLER_4_131
timestamp 1584750033
transform 1 0 13152 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_135
timestamp 1584750033
transform 1 0 13536 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_153
timestamp 1584750033
transform 1 0 15264 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_0
timestamp 1584750033
transform 1 0 576 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_2
timestamp 1584750033
transform 1 0 768 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_11
timestamp 1584750033
transform 1 0 1632 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_24
timestamp 1584750033
transform 1 0 2880 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_31
timestamp 1584750033
transform 1 0 3552 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_42
timestamp 1584750033
transform 1 0 4608 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1584750033
transform 1 0 6336 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_79
timestamp 1584750033
transform 1 0 8160 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_85
timestamp 1584750033
transform 1 0 8736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_92
timestamp 1584750033
transform 1 0 9408 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_96
timestamp 1584750033
transform 1 0 9792 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_102
timestamp 1584750033
transform 1 0 10368 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_4  FILLER_5_114
timestamp 1584750033
transform 1 0 11520 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_118
timestamp 1584750033
transform 1 0 11904 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_128
timestamp 1584750033
transform 1 0 12864 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_135
timestamp 1584750033
transform 1 0 13536 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_153
timestamp 1584750033
transform 1 0 15264 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_0
timestamp 1584750033
transform 1 0 576 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_2
timestamp 1584750033
transform 1 0 768 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_13
timestamp 1584750033
transform 1 0 1824 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_45
timestamp 1584750033
transform 1 0 4896 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_66
timestamp 1584750033
transform 1 0 6912 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_75
timestamp 1584750033
transform 1 0 7776 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_94
timestamp 1584750033
transform 1 0 9600 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_96
timestamp 1584750033
transform 1 0 9792 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_115
timestamp 1584750033
transform 1 0 11616 0 1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_131
timestamp 1584750033
transform 1 0 13152 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_135
timestamp 1584750033
transform 1 0 13536 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_153
timestamp 1584750033
transform 1 0 15264 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_0
timestamp 1584750033
transform 1 0 576 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_22
timestamp 1584750033
transform 1 0 2688 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_29
timestamp 1584750033
transform 1 0 3360 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_36
timestamp 1584750033
transform 1 0 4032 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_38
timestamp 1584750033
transform 1 0 4224 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_59
timestamp 1584750033
transform 1 0 6240 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_79
timestamp 1584750033
transform 1 0 8160 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_88
timestamp 1584750033
transform 1 0 9024 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_95
timestamp 1584750033
transform 1 0 9696 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_111
timestamp 1584750033
transform 1 0 11232 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_129
timestamp 1584750033
transform 1 0 12960 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_131
timestamp 1584750033
transform 1 0 13152 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_136
timestamp 1584750033
transform 1 0 13632 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_140
timestamp 1584750033
transform 1 0 14016 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_153
timestamp 1584750033
transform 1 0 15264 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_14
timestamp 1584750033
transform 1 0 1920 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_16
timestamp 1584750033
transform 1 0 2112 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_29
timestamp 1584750033
transform 1 0 3360 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_31
timestamp 1584750033
transform 1 0 3552 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_54
timestamp 1584750033
transform 1 0 5760 0 1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_8_61
timestamp 1584750033
transform 1 0 6432 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_75
timestamp 1584750033
transform 1 0 7776 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_77
timestamp 1584750033
transform 1 0 7968 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_98
timestamp 1584750033
transform 1 0 9984 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_118
timestamp 1584750033
transform 1 0 11904 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_120
timestamp 1584750033
transform 1 0 12096 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_143
timestamp 1584750033
transform 1 0 14304 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_153
timestamp 1584750033
transform 1 0 15264 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_0
timestamp 1584750033
transform 1 0 576 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_2
timestamp 1584750033
transform 1 0 768 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_11
timestamp 1584750033
transform 1 0 1632 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_24
timestamp 1584750033
transform 1 0 2880 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_26
timestamp 1584750033
transform 1 0 3072 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_41
timestamp 1584750033
transform 1 0 4512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_48
timestamp 1584750033
transform 1 0 5184 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_52
timestamp 1584750033
transform 1 0 5568 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_78
timestamp 1584750033
transform 1 0 8064 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_94
timestamp 1584750033
transform 1 0 9600 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_98
timestamp 1584750033
transform 1 0 9984 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_110
timestamp 1584750033
transform 1 0 11136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_117
timestamp 1584750033
transform 1 0 11808 0 -1 8316
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_127
timestamp 1584750033
transform 1 0 12768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_134
timestamp 1584750033
transform 1 0 13440 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_153
timestamp 1584750033
transform 1 0 15264 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_0
timestamp 1584750033
transform 1 0 576 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_2
timestamp 1584750033
transform 1 0 768 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_13
timestamp 1584750033
transform 1 0 1824 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_29
timestamp 1584750033
transform 1 0 3360 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_42
timestamp 1584750033
transform 1 0 4608 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_44
timestamp 1584750033
transform 1 0 4800 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_57
timestamp 1584750033
transform 1 0 6048 0 1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_61
timestamp 1584750033
transform 1 0 6432 0 1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_72
timestamp 1584750033
transform 1 0 7488 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_76
timestamp 1584750033
transform 1 0 7872 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_112
timestamp 1584750033
transform 1 0 11328 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_119
timestamp 1584750033
transform 1 0 12000 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_129
timestamp 1584750033
transform 1 0 12960 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_136
timestamp 1584750033
transform 1 0 13632 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_153
timestamp 1584750033
transform 1 0 15264 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_12
timestamp 1584750033
transform 1 0 1728 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_21
timestamp 1584750033
transform 1 0 2592 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_35
timestamp 1584750033
transform 1 0 3936 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_55
timestamp 1584750033
transform 1 0 5856 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_76
timestamp 1584750033
transform 1 0 7872 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_94
timestamp 1584750033
transform 1 0 9600 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_101
timestamp 1584750033
transform 1 0 10272 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_103
timestamp 1584750033
transform 1 0 10464 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_112
timestamp 1584750033
transform 1 0 11328 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_130
timestamp 1584750033
transform 1 0 13056 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_132
timestamp 1584750033
transform 1 0 13248 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_153
timestamp 1584750033
transform 1 0 15264 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_0
timestamp 1584750033
transform 1 0 576 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_44
timestamp 1584750033
transform 1 0 4800 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_46
timestamp 1584750033
transform 1 0 4992 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_51
timestamp 1584750033
transform 1 0 5472 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_56
timestamp 1584750033
transform 1 0 5952 0 1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_63
timestamp 1584750033
transform 1 0 6624 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_72
timestamp 1584750033
transform 1 0 7488 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_79
timestamp 1584750033
transform 1 0 8160 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_81
timestamp 1584750033
transform 1 0 8352 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_96
timestamp 1584750033
transform 1 0 9792 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_135
timestamp 1584750033
transform 1 0 13536 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_153
timestamp 1584750033
transform 1 0 15264 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_0
timestamp 1584750033
transform 1 0 576 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_2
timestamp 1584750033
transform 1 0 768 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_11
timestamp 1584750033
transform 1 0 1632 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_35
timestamp 1584750033
transform 1 0 3936 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_63
timestamp 1584750033
transform 1 0 6624 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_13_90
timestamp 1584750033
transform 1 0 9216 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_92
timestamp 1584750033
transform 1 0 9408 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_99
timestamp 1584750033
transform 1 0 10080 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_101
timestamp 1584750033
transform 1 0 10272 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_116
timestamp 1584750033
transform 1 0 11712 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_132
timestamp 1584750033
transform 1 0 13248 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_134
timestamp 1584750033
transform 1 0 13440 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_151
timestamp 1584750033
transform 1 0 15072 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_153
timestamp 1584750033
transform 1 0 15264 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_0
timestamp 1584750033
transform 1 0 576 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_2
timestamp 1584750033
transform 1 0 768 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_11
timestamp 1584750033
transform 1 0 1632 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_20
timestamp 1584750033
transform 1 0 2496 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_22
timestamp 1584750033
transform 1 0 2688 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_39
timestamp 1584750033
transform 1 0 4320 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_46
timestamp 1584750033
transform 1 0 4992 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_51
timestamp 1584750033
transform 1 0 5472 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_53
timestamp 1584750033
transform 1 0 5664 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_60
timestamp 1584750033
transform 1 0 6336 0 1 11340
box -48 -56 432 834
use sg13g2_decap_8  FILLER_14_78
timestamp 1584750033
transform 1 0 8064 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_85
timestamp 1584750033
transform 1 0 8736 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_87
timestamp 1584750033
transform 1 0 8928 0 1 11340
box -48 -56 144 834
use sg13g2_decap_4  FILLER_14_102
timestamp 1584750033
transform 1 0 10368 0 1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_14_106
timestamp 1584750033
transform 1 0 10752 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_111
timestamp 1584750033
transform 1 0 11232 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_14_123
timestamp 1584750033
transform 1 0 12384 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_125
timestamp 1584750033
transform 1 0 12576 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_130
timestamp 1584750033
transform 1 0 13056 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_132
timestamp 1584750033
transform 1 0 13248 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_153
timestamp 1584750033
transform 1 0 15264 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_0
timestamp 1584750033
transform 1 0 576 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_2
timestamp 1584750033
transform 1 0 768 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_21
timestamp 1584750033
transform 1 0 2592 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_51
timestamp 1584750033
transform 1 0 5472 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_68
timestamp 1584750033
transform 1 0 7104 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_88
timestamp 1584750033
transform 1 0 9024 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_90
timestamp 1584750033
transform 1 0 9216 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_99
timestamp 1584750033
transform 1 0 10080 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_105
timestamp 1584750033
transform 1 0 10656 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_110
timestamp 1584750033
transform 1 0 11136 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_120
timestamp 1584750033
transform 1 0 12096 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_122
timestamp 1584750033
transform 1 0 12288 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_135
timestamp 1584750033
transform 1 0 13536 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_153
timestamp 1584750033
transform 1 0 15264 0 -1 12852
box -48 -56 144 834
<< labels >>
flabel metal3 s 15920 1556 16000 1636 0 FreeSans 320 0 0 0 ON[0]
port 0 nsew signal output
flabel metal3 s 15920 4916 16000 4996 0 FreeSans 320 0 0 0 ON[10]
port 1 nsew signal output
flabel metal3 s 15920 5252 16000 5332 0 FreeSans 320 0 0 0 ON[11]
port 2 nsew signal output
flabel metal3 s 15920 5588 16000 5668 0 FreeSans 320 0 0 0 ON[12]
port 3 nsew signal output
flabel metal3 s 15920 5924 16000 6004 0 FreeSans 320 0 0 0 ON[13]
port 4 nsew signal output
flabel metal3 s 15920 6260 16000 6340 0 FreeSans 320 0 0 0 ON[14]
port 5 nsew signal output
flabel metal3 s 15920 6596 16000 6676 0 FreeSans 320 0 0 0 ON[15]
port 6 nsew signal output
flabel metal3 s 15920 6932 16000 7012 0 FreeSans 320 0 0 0 ON[16]
port 7 nsew signal output
flabel metal3 s 15920 7268 16000 7348 0 FreeSans 320 0 0 0 ON[17]
port 8 nsew signal output
flabel metal3 s 15920 7604 16000 7684 0 FreeSans 320 0 0 0 ON[18]
port 9 nsew signal output
flabel metal3 s 15920 7940 16000 8020 0 FreeSans 320 0 0 0 ON[19]
port 10 nsew signal output
flabel metal3 s 15920 1892 16000 1972 0 FreeSans 320 0 0 0 ON[1]
port 11 nsew signal output
flabel metal3 s 15920 8276 16000 8356 0 FreeSans 320 0 0 0 ON[20]
port 12 nsew signal output
flabel metal3 s 15920 8612 16000 8692 0 FreeSans 320 0 0 0 ON[21]
port 13 nsew signal output
flabel metal3 s 15920 8948 16000 9028 0 FreeSans 320 0 0 0 ON[22]
port 14 nsew signal output
flabel metal3 s 15920 9284 16000 9364 0 FreeSans 320 0 0 0 ON[23]
port 15 nsew signal output
flabel metal3 s 15920 9620 16000 9700 0 FreeSans 320 0 0 0 ON[24]
port 16 nsew signal output
flabel metal3 s 15920 9956 16000 10036 0 FreeSans 320 0 0 0 ON[25]
port 17 nsew signal output
flabel metal3 s 15920 10292 16000 10372 0 FreeSans 320 0 0 0 ON[26]
port 18 nsew signal output
flabel metal3 s 15920 10628 16000 10708 0 FreeSans 320 0 0 0 ON[27]
port 19 nsew signal output
flabel metal3 s 15920 10964 16000 11044 0 FreeSans 320 0 0 0 ON[28]
port 20 nsew signal output
flabel metal3 s 15920 11300 16000 11380 0 FreeSans 320 0 0 0 ON[29]
port 21 nsew signal output
flabel metal3 s 15920 2228 16000 2308 0 FreeSans 320 0 0 0 ON[2]
port 22 nsew signal output
flabel metal3 s 15920 11636 16000 11716 0 FreeSans 320 0 0 0 ON[30]
port 23 nsew signal output
flabel metal3 s 15920 11972 16000 12052 0 FreeSans 320 0 0 0 ON[31]
port 24 nsew signal output
flabel metal3 s 15920 2564 16000 2644 0 FreeSans 320 0 0 0 ON[3]
port 25 nsew signal output
flabel metal3 s 15920 2900 16000 2980 0 FreeSans 320 0 0 0 ON[4]
port 26 nsew signal output
flabel metal3 s 15920 3236 16000 3316 0 FreeSans 320 0 0 0 ON[5]
port 27 nsew signal output
flabel metal3 s 15920 3572 16000 3652 0 FreeSans 320 0 0 0 ON[6]
port 28 nsew signal output
flabel metal3 s 15920 3908 16000 3988 0 FreeSans 320 0 0 0 ON[7]
port 29 nsew signal output
flabel metal3 s 15920 4244 16000 4324 0 FreeSans 320 0 0 0 ON[8]
port 30 nsew signal output
flabel metal3 s 15920 4580 16000 4660 0 FreeSans 320 0 0 0 ON[9]
port 31 nsew signal output
flabel metal3 s 15920 1724 16000 1804 0 FreeSans 320 0 0 0 ON_N[0]
port 32 nsew signal output
flabel metal3 s 15920 5084 16000 5164 0 FreeSans 320 0 0 0 ON_N[10]
port 33 nsew signal output
flabel metal3 s 15920 5420 16000 5500 0 FreeSans 320 0 0 0 ON_N[11]
port 34 nsew signal output
flabel metal3 s 15920 5756 16000 5836 0 FreeSans 320 0 0 0 ON_N[12]
port 35 nsew signal output
flabel metal3 s 15920 6092 16000 6172 0 FreeSans 320 0 0 0 ON_N[13]
port 36 nsew signal output
flabel metal3 s 15920 6428 16000 6508 0 FreeSans 320 0 0 0 ON_N[14]
port 37 nsew signal output
flabel metal3 s 15920 6764 16000 6844 0 FreeSans 320 0 0 0 ON_N[15]
port 38 nsew signal output
flabel metal3 s 15920 7100 16000 7180 0 FreeSans 320 0 0 0 ON_N[16]
port 39 nsew signal output
flabel metal3 s 15920 7436 16000 7516 0 FreeSans 320 0 0 0 ON_N[17]
port 40 nsew signal output
flabel metal3 s 15920 7772 16000 7852 0 FreeSans 320 0 0 0 ON_N[18]
port 41 nsew signal output
flabel metal3 s 15920 8108 16000 8188 0 FreeSans 320 0 0 0 ON_N[19]
port 42 nsew signal output
flabel metal3 s 15920 2060 16000 2140 0 FreeSans 320 0 0 0 ON_N[1]
port 43 nsew signal output
flabel metal3 s 15920 8444 16000 8524 0 FreeSans 320 0 0 0 ON_N[20]
port 44 nsew signal output
flabel metal3 s 15920 8780 16000 8860 0 FreeSans 320 0 0 0 ON_N[21]
port 45 nsew signal output
flabel metal3 s 15920 9116 16000 9196 0 FreeSans 320 0 0 0 ON_N[22]
port 46 nsew signal output
flabel metal3 s 15920 9452 16000 9532 0 FreeSans 320 0 0 0 ON_N[23]
port 47 nsew signal output
flabel metal3 s 15920 9788 16000 9868 0 FreeSans 320 0 0 0 ON_N[24]
port 48 nsew signal output
flabel metal3 s 15920 10124 16000 10204 0 FreeSans 320 0 0 0 ON_N[25]
port 49 nsew signal output
flabel metal3 s 15920 10460 16000 10540 0 FreeSans 320 0 0 0 ON_N[26]
port 50 nsew signal output
flabel metal3 s 15920 10796 16000 10876 0 FreeSans 320 0 0 0 ON_N[27]
port 51 nsew signal output
flabel metal3 s 15920 11132 16000 11212 0 FreeSans 320 0 0 0 ON_N[28]
port 52 nsew signal output
flabel metal3 s 15920 11468 16000 11548 0 FreeSans 320 0 0 0 ON_N[29]
port 53 nsew signal output
flabel metal3 s 15920 2396 16000 2476 0 FreeSans 320 0 0 0 ON_N[2]
port 54 nsew signal output
flabel metal3 s 15920 11804 16000 11884 0 FreeSans 320 0 0 0 ON_N[30]
port 55 nsew signal output
flabel metal3 s 15920 12140 16000 12220 0 FreeSans 320 0 0 0 ON_N[31]
port 56 nsew signal output
flabel metal3 s 15920 2732 16000 2812 0 FreeSans 320 0 0 0 ON_N[3]
port 57 nsew signal output
flabel metal3 s 15920 3068 16000 3148 0 FreeSans 320 0 0 0 ON_N[4]
port 58 nsew signal output
flabel metal3 s 15920 3404 16000 3484 0 FreeSans 320 0 0 0 ON_N[5]
port 59 nsew signal output
flabel metal3 s 15920 3740 16000 3820 0 FreeSans 320 0 0 0 ON_N[6]
port 60 nsew signal output
flabel metal3 s 15920 4076 16000 4156 0 FreeSans 320 0 0 0 ON_N[7]
port 61 nsew signal output
flabel metal3 s 15920 4412 16000 4492 0 FreeSans 320 0 0 0 ON_N[8]
port 62 nsew signal output
flabel metal3 s 15920 4748 16000 4828 0 FreeSans 320 0 0 0 ON_N[9]
port 63 nsew signal output
flabel metal4 s 4316 712 4756 12896 0 FreeSans 2560 90 0 0 VGND
port 64 nsew ground bidirectional
flabel metal5 s 532 4496 15404 4936 0 FreeSans 2560 0 0 0 VGND
port 64 nsew ground bidirectional
flabel metal4 s 3076 712 3516 12896 0 FreeSans 2560 90 0 0 VPWR
port 65 nsew power bidirectional
flabel metal5 s 532 3256 15404 3696 0 FreeSans 2560 0 0 0 VPWR
port 65 nsew power bidirectional
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 thermo[0]
port 66 nsew signal input
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 thermo[10]
port 67 nsew signal input
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 thermo[11]
port 68 nsew signal input
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 thermo[12]
port 69 nsew signal input
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 thermo[13]
port 70 nsew signal input
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 thermo[14]
port 71 nsew signal input
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 thermo[15]
port 72 nsew signal input
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 thermo[16]
port 73 nsew signal input
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 thermo[17]
port 74 nsew signal input
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 thermo[18]
port 75 nsew signal input
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 thermo[19]
port 76 nsew signal input
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 thermo[1]
port 77 nsew signal input
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 thermo[20]
port 78 nsew signal input
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 thermo[21]
port 79 nsew signal input
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 thermo[22]
port 80 nsew signal input
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 thermo[23]
port 81 nsew signal input
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 thermo[24]
port 82 nsew signal input
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 thermo[25]
port 83 nsew signal input
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 thermo[26]
port 84 nsew signal input
flabel metal3 s 0 10796 80 10876 0 FreeSans 320 0 0 0 thermo[27]
port 85 nsew signal input
flabel metal3 s 0 11132 80 11212 0 FreeSans 320 0 0 0 thermo[28]
port 86 nsew signal input
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 thermo[29]
port 87 nsew signal input
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 thermo[2]
port 88 nsew signal input
flabel metal3 s 0 11804 80 11884 0 FreeSans 320 0 0 0 thermo[30]
port 89 nsew signal input
flabel metal3 s 0 12140 80 12220 0 FreeSans 320 0 0 0 thermo[31]
port 90 nsew signal input
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 thermo[3]
port 91 nsew signal input
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 thermo[4]
port 92 nsew signal input
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 thermo[5]
port 93 nsew signal input
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 thermo[6]
port 94 nsew signal input
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 thermo[7]
port 95 nsew signal input
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 thermo[8]
port 96 nsew signal input
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 thermo[9]
port 97 nsew signal input
rlabel metal1 7968 12852 7968 12852 0 VGND
rlabel metal1 7968 12096 7968 12096 0 VPWR
rlabel metal3 15554 1596 15554 1596 0 ON[0]
rlabel metal3 14978 4956 14978 4956 0 ON[10]
rlabel metal3 15170 5292 15170 5292 0 ON[11]
rlabel metal3 15554 5628 15554 5628 0 ON[12]
rlabel metal3 15362 5964 15362 5964 0 ON[13]
rlabel metal3 14976 6216 14976 6216 0 ON[14]
rlabel metal3 15602 6636 15602 6636 0 ON[15]
rlabel metal3 14882 6972 14882 6972 0 ON[16]
rlabel metal3 15458 7308 15458 7308 0 ON[17]
rlabel metal3 15362 7644 15362 7644 0 ON[18]
rlabel metal3 15410 7980 15410 7980 0 ON[19]
rlabel metal3 15362 1932 15362 1932 0 ON[1]
rlabel metal3 15170 8316 15170 8316 0 ON[20]
rlabel metal3 15170 8652 15170 8652 0 ON[21]
rlabel metal3 15554 8988 15554 8988 0 ON[22]
rlabel metal3 14978 9324 14978 9324 0 ON[23]
rlabel metal3 15218 9660 15218 9660 0 ON[24]
rlabel metal3 15554 9996 15554 9996 0 ON[25]
rlabel metal3 15458 10332 15458 10332 0 ON[26]
rlabel metal3 15362 10668 15362 10668 0 ON[27]
rlabel metal3 15170 11004 15170 11004 0 ON[28]
rlabel metal3 15410 11340 15410 11340 0 ON[29]
rlabel metal3 15554 2268 15554 2268 0 ON[2]
rlabel metal3 15554 11676 15554 11676 0 ON[30]
rlabel metal3 14978 12012 14978 12012 0 ON[31]
rlabel metal3 15362 2604 15362 2604 0 ON[3]
rlabel metal3 14786 2940 14786 2940 0 ON[4]
rlabel metal3 15266 3276 15266 3276 0 ON[5]
rlabel metal3 15170 3612 15170 3612 0 ON[6]
rlabel metal3 15602 3948 15602 3948 0 ON[7]
rlabel metal3 15170 4284 15170 4284 0 ON[8]
rlabel metal3 15362 4620 15362 4620 0 ON[9]
rlabel metal3 14978 1764 14978 1764 0 ON_N[0]
rlabel metal3 15026 5124 15026 5124 0 ON_N[10]
rlabel metal3 15410 5460 15410 5460 0 ON_N[11]
rlabel metal3 15170 5796 15170 5796 0 ON_N[12]
rlabel metal3 15554 6132 15554 6132 0 ON_N[13]
rlabel metal3 15362 6468 15362 6468 0 ON_N[14]
rlabel metal3 14738 6804 14738 6804 0 ON_N[15]
rlabel metal3 15074 7140 15074 7140 0 ON_N[16]
rlabel metal3 15554 7476 15554 7476 0 ON_N[17]
rlabel metal3 15170 7812 15170 7812 0 ON_N[18]
rlabel metal3 15602 8148 15602 8148 0 ON_N[19]
rlabel metal3 15170 2100 15170 2100 0 ON_N[1]
rlabel metal3 14978 8484 14978 8484 0 ON_N[20]
rlabel metal3 15362 8820 15362 8820 0 ON_N[21]
rlabel metal3 15410 9156 15410 9156 0 ON_N[22]
rlabel metal3 14786 9492 14786 9492 0 ON_N[23]
rlabel metal3 14978 9828 14978 9828 0 ON_N[24]
rlabel metal3 15266 10164 15266 10164 0 ON_N[25]
rlabel metal3 15074 10500 15074 10500 0 ON_N[26]
rlabel metal3 14882 10836 14882 10836 0 ON_N[27]
rlabel metal3 15554 11172 15554 11172 0 ON_N[28]
rlabel metal3 14978 11508 14978 11508 0 ON_N[29]
rlabel metal3 14882 2436 14882 2436 0 ON_N[2]
rlabel metal3 15170 11844 15170 11844 0 ON_N[30]
rlabel metal3 14786 12180 14786 12180 0 ON_N[31]
rlabel metal3 15074 2772 15074 2772 0 ON_N[3]
rlabel metal3 15458 3108 15458 3108 0 ON_N[4]
rlabel metal3 14978 3444 14978 3444 0 ON_N[5]
rlabel metal3 14978 3780 14978 3780 0 ON_N[6]
rlabel metal3 15410 4116 15410 4116 0 ON_N[7]
rlabel metal3 15554 4452 15554 4452 0 ON_N[8]
rlabel metal3 15554 4788 15554 4788 0 ON_N[9]
rlabel metal2 10992 7896 10992 7896 0 _000_
rlabel metal2 10464 8064 10464 8064 0 _001_
rlabel metal2 1152 1974 1152 1974 0 _002_
rlabel metal2 1440 1932 1440 1932 0 _003_
rlabel metal3 1104 1092 1104 1092 0 _004_
rlabel metal2 12480 9534 12480 9534 0 _005_
rlabel metal2 12000 9576 12000 9576 0 _006_
rlabel metal3 8784 5712 8784 5712 0 _007_
rlabel metal2 8448 5250 8448 5250 0 _008_
rlabel metal2 7440 4956 7440 4956 0 _009_
rlabel metal2 10944 3486 10944 3486 0 _010_
rlabel metal2 10464 3528 10464 3528 0 _011_
rlabel metal2 6096 4872 6096 4872 0 _012_
rlabel metal2 5664 5208 5664 5208 0 _013_
rlabel metal2 5376 5208 5376 5208 0 _014_
rlabel metal2 11040 9954 11040 9954 0 _015_
rlabel metal2 11520 10080 11520 10080 0 _016_
rlabel metal2 3840 5166 3840 5166 0 _017_
rlabel metal2 4416 5460 4416 5460 0 _018_
rlabel metal3 2736 5628 2736 5628 0 _019_
rlabel metal2 10656 6510 10656 6510 0 _020_
rlabel metal2 10176 6552 10176 6552 0 _021_
rlabel metal2 2016 5712 2016 5712 0 _022_
rlabel metal2 1152 5544 1152 5544 0 _023_
rlabel metal2 1152 6720 1152 6720 0 _024_
rlabel metal2 10944 11214 10944 11214 0 _025_
rlabel metal2 11424 11088 11424 11088 0 _026_
rlabel metal2 7104 5880 7104 5880 0 _027_
rlabel metal2 7056 6972 7056 6972 0 _028_
rlabel metal3 7632 6468 7632 6468 0 _029_
rlabel metal2 9456 4200 9456 4200 0 _030_
rlabel metal2 8928 4032 8928 4032 0 _031_
rlabel metal2 5280 7224 5280 7224 0 _032_
rlabel metal3 5136 6972 5136 6972 0 _033_
rlabel metal3 4848 6468 4848 6468 0 _034_
rlabel metal2 8208 2100 8208 2100 0 _035_
rlabel metal2 7680 1008 7680 1008 0 _036_
rlabel metal2 3936 6384 3936 6384 0 _037_
rlabel metal2 3504 8148 3504 8148 0 _038_
rlabel metal3 2736 7140 2736 7140 0 _039_
rlabel metal2 10656 10710 10656 10710 0 _040_
rlabel metal2 10176 10080 10176 10080 0 _041_
rlabel metal2 9024 8022 9024 8022 0 _042_
rlabel metal2 8544 8064 8544 8064 0 _043_
rlabel metal3 8592 7140 8592 7140 0 _044_
rlabel metal2 9888 11214 9888 11214 0 _045_
rlabel metal2 9312 11256 9312 11256 0 _046_
rlabel metal3 7488 8148 7488 8148 0 _047_
rlabel metal2 6960 7140 6960 7140 0 _048_
rlabel metal2 6048 8064 6048 8064 0 _049_
rlabel metal3 12912 10248 12912 10248 0 _050_
rlabel metal2 12096 10080 12096 10080 0 _051_
rlabel metal3 2160 8148 2160 8148 0 _052_
rlabel metal2 1248 7056 1248 7056 0 _053_
rlabel metal2 1248 8232 1248 8232 0 _054_
rlabel metal2 12720 3612 12720 3612 0 _055_
rlabel metal2 12432 2604 12432 2604 0 _056_
rlabel metal2 3264 1890 3264 1890 0 _057_
rlabel metal3 3552 924 3552 924 0 _058_
rlabel metal2 2928 1092 2928 1092 0 _059_
rlabel metal2 11232 4662 11232 4662 0 _060_
rlabel metal2 11040 4620 11040 4620 0 _061_
rlabel metal2 3744 8190 3744 8190 0 _062_
rlabel metal3 3552 9660 3552 9660 0 _063_
rlabel metal3 2736 8652 2736 8652 0 _064_
rlabel metal2 9216 10122 9216 10122 0 _065_
rlabel metal2 8736 10080 8736 10080 0 _066_
rlabel metal2 9024 9534 9024 9534 0 _067_
rlabel metal2 8544 9576 8544 9576 0 _068_
rlabel metal3 8592 8652 8592 8652 0 _069_
rlabel metal2 11808 12222 11808 12222 0 _070_
rlabel metal2 11616 12180 11616 12180 0 _071_
rlabel metal2 7344 9996 7344 9996 0 _072_
rlabel metal2 7056 8652 7056 8652 0 _073_
rlabel metal2 6240 9576 6240 9576 0 _074_
rlabel metal2 10656 5586 10656 5586 0 _075_
rlabel metal2 10176 5544 10176 5544 0 _076_
rlabel metal2 4896 9702 4896 9702 0 _077_
rlabel metal2 4416 9576 4416 9576 0 _078_
rlabel metal2 5280 8568 5280 8568 0 _079_
rlabel metal2 6816 1050 6816 1050 0 _080_
rlabel metal2 7008 1008 7008 1008 0 _081_
rlabel metal2 864 9198 864 9198 0 _082_
rlabel metal2 1632 9324 1632 9324 0 _083_
rlabel metal2 1344 9744 1344 9744 0 _084_
rlabel metal3 12912 7224 12912 7224 0 _085_
rlabel metal3 12624 6972 12624 6972 0 _086_
rlabel metal2 3600 9408 3600 9408 0 _087_
rlabel metal3 4128 9996 4128 9996 0 _088_
rlabel metal2 3264 10080 3264 10080 0 _089_
rlabel metal2 10080 4662 10080 4662 0 _090_
rlabel metal2 10560 4032 10560 4032 0 _091_
rlabel metal2 2016 10878 2016 10878 0 _092_
rlabel metal3 2208 10164 2208 10164 0 _093_
rlabel metal2 1248 11256 1248 11256 0 _094_
rlabel metal2 10848 2394 10848 2394 0 _095_
rlabel metal2 10368 2520 10368 2520 0 _096_
rlabel metal2 4896 11214 4896 11214 0 _097_
rlabel metal2 4416 11088 4416 11088 0 _098_
rlabel metal2 5472 10500 5472 10500 0 _099_
rlabel metal2 11424 1638 11424 1638 0 _100_
rlabel metal2 10752 1218 10752 1218 0 _101_
rlabel metal2 7536 11760 7536 11760 0 _102_
rlabel metal2 7008 11592 7008 11592 0 _103_
rlabel metal2 8064 11088 8064 11088 0 _104_
rlabel metal2 12576 4074 12576 4074 0 _105_
rlabel metal2 12096 4032 12096 4032 0 _106_
rlabel metal2 3792 10920 3792 10920 0 _107_
rlabel metal2 3072 12768 3072 12768 0 _108_
rlabel metal2 3168 11802 3168 11802 0 _109_
rlabel metal2 9312 2562 9312 2562 0 _110_
rlabel metal2 8832 2520 8832 2520 0 _111_
rlabel metal2 5568 2100 5568 2100 0 _112_
rlabel metal2 5712 1092 5712 1092 0 _113_
rlabel metal2 4608 2016 4608 2016 0 _114_
rlabel metal2 12672 11046 12672 11046 0 _115_
rlabel metal2 12192 11088 12192 11088 0 _116_
rlabel metal2 2208 11760 2208 11760 0 _117_
rlabel metal2 4032 12600 4032 12600 0 _118_
rlabel metal3 1680 11676 1680 11676 0 _119_
rlabel metal2 10944 7098 10944 7098 0 _120_
rlabel metal2 10464 7056 10464 7056 0 _121_
rlabel metal2 5904 12684 5904 12684 0 _122_
rlabel metal2 6816 12180 6816 12180 0 _123_
rlabel metal2 5088 12600 5088 12600 0 _124_
rlabel metal2 12864 1974 12864 1974 0 _125_
rlabel metal3 12336 2100 12336 2100 0 _126_
rlabel metal2 7392 2142 7392 2142 0 _127_
rlabel metal2 8064 2436 8064 2436 0 _128_
rlabel metal2 6048 2520 6048 2520 0 _129_
rlabel metal2 12624 7896 12624 7896 0 _130_
rlabel metal2 12288 8232 12288 8232 0 _131_
rlabel metal2 3552 2730 3552 2730 0 _132_
rlabel metal3 3216 2436 3216 2436 0 _133_
rlabel metal2 3072 2604 3072 2604 0 _134_
rlabel metal2 10800 9660 10800 9660 0 _135_
rlabel metal2 10272 8568 10272 8568 0 _136_
rlabel metal2 1152 3486 1152 3486 0 _137_
rlabel metal2 1392 3444 1392 3444 0 _138_
rlabel metal2 1344 2520 1344 2520 0 _139_
rlabel metal2 12384 6510 12384 6510 0 _140_
rlabel metal2 11904 6552 11904 6552 0 _141_
rlabel metal2 4800 3150 4800 3150 0 _142_
rlabel metal2 5568 3192 5568 3192 0 _143_
rlabel metal2 5280 3780 5280 3780 0 _144_
rlabel metal2 12576 5586 12576 5586 0 _145_
rlabel metal2 12096 5544 12096 5544 0 _146_
rlabel metal2 3888 3360 3888 3360 0 _147_
rlabel metal2 4416 3948 4416 3948 0 _148_
rlabel metal2 3072 4032 3072 4032 0 _149_
rlabel metal2 8928 1638 8928 1638 0 _150_
rlabel metal3 8976 924 8976 924 0 _151_
rlabel metal2 8016 3360 8016 3360 0 _152_
rlabel metal2 7488 3528 7488 3528 0 _153_
rlabel metal2 7104 4032 7104 4032 0 _154_
rlabel metal2 9792 12222 9792 12222 0 _155_
rlabel metal2 9600 12180 9600 12180 0 _156_
rlabel metal3 2256 5124 2256 5124 0 _157_
rlabel metal2 1440 4032 1440 4032 0 _158_
rlabel metal2 1248 4452 1248 4452 0 _159_
rlabel metal3 654 1764 654 1764 0 thermo[0]
rlabel metal3 942 5124 942 5124 0 thermo[10]
rlabel metal2 5472 5208 5472 5208 0 thermo[11]
rlabel metal2 2880 5712 2880 5712 0 thermo[12]
rlabel metal3 558 6132 558 6132 0 thermo[13]
rlabel metal3 1182 6468 1182 6468 0 thermo[14]
rlabel metal2 5184 6594 5184 6594 0 thermo[15]
rlabel metal2 2880 7182 2880 7182 0 thermo[16]
rlabel metal2 8928 7308 8928 7308 0 thermo[17]
rlabel metal3 3180 7812 3180 7812 0 thermo[18]
rlabel metal2 1152 8064 1152 8064 0 thermo[19]
rlabel metal2 3072 1176 3072 1176 0 thermo[1]
rlabel metal2 2880 8568 2880 8568 0 thermo[20]
rlabel metal2 8928 8736 8928 8736 0 thermo[21]
rlabel metal2 7200 9156 7200 9156 0 thermo[22]
rlabel metal3 3072 9408 3072 9408 0 thermo[23]
rlabel metal2 1440 9660 1440 9660 0 thermo[24]
rlabel metal2 3168 10206 3168 10206 0 thermo[25]
rlabel metal2 1152 10752 1152 10752 0 thermo[26]
rlabel metal3 2382 10836 2382 10836 0 thermo[27]
rlabel metal2 7392 11424 7392 11424 0 thermo[28]
rlabel metal2 3072 11592 3072 11592 0 thermo[29]
rlabel metal2 4512 2016 4512 2016 0 thermo[2]
rlabel metal2 1152 11760 1152 11760 0 thermo[30]
rlabel metal2 5184 12348 5184 12348 0 thermo[31]
rlabel metal2 6432 2688 6432 2688 0 thermo[3]
rlabel metal2 3264 2730 3264 2730 0 thermo[4]
rlabel metal3 654 3444 654 3444 0 thermo[5]
rlabel metal2 5184 3654 5184 3654 0 thermo[6]
rlabel metal3 1518 4116 1518 4116 0 thermo[7]
rlabel metal2 7008 4284 7008 4284 0 thermo[8]
rlabel metal2 1152 4872 1152 4872 0 thermo[9]
<< properties >>
string FIXED_BBOX 0 0 16000 14000
<< end >>
