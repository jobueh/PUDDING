VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO non_overlap
  CLASS BLOCK ;
  FOREIGN non_overlap ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 70.000 ;
  PIN ON[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 7.780 80.000 8.180 ;
    END
  END ON[0]
  PIN ON[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 24.580 80.000 24.980 ;
    END
  END ON[10]
  PIN ON[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 26.260 80.000 26.660 ;
    END
  END ON[11]
  PIN ON[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 27.940 80.000 28.340 ;
    END
  END ON[12]
  PIN ON[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 29.620 80.000 30.020 ;
    END
  END ON[13]
  PIN ON[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 31.300 80.000 31.700 ;
    END
  END ON[14]
  PIN ON[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 32.980 80.000 33.380 ;
    END
  END ON[15]
  PIN ON[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 34.660 80.000 35.060 ;
    END
  END ON[16]
  PIN ON[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 36.340 80.000 36.740 ;
    END
  END ON[17]
  PIN ON[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 38.020 80.000 38.420 ;
    END
  END ON[18]
  PIN ON[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 39.700 80.000 40.100 ;
    END
  END ON[19]
  PIN ON[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 9.460 80.000 9.860 ;
    END
  END ON[1]
  PIN ON[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 41.380 80.000 41.780 ;
    END
  END ON[20]
  PIN ON[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 43.060 80.000 43.460 ;
    END
  END ON[21]
  PIN ON[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 44.740 80.000 45.140 ;
    END
  END ON[22]
  PIN ON[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 46.420 80.000 46.820 ;
    END
  END ON[23]
  PIN ON[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 48.100 80.000 48.500 ;
    END
  END ON[24]
  PIN ON[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 49.780 80.000 50.180 ;
    END
  END ON[25]
  PIN ON[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 51.460 80.000 51.860 ;
    END
  END ON[26]
  PIN ON[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 53.140 80.000 53.540 ;
    END
  END ON[27]
  PIN ON[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 54.820 80.000 55.220 ;
    END
  END ON[28]
  PIN ON[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 56.500 80.000 56.900 ;
    END
  END ON[29]
  PIN ON[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 11.140 80.000 11.540 ;
    END
  END ON[2]
  PIN ON[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 58.180 80.000 58.580 ;
    END
  END ON[30]
  PIN ON[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 59.860 80.000 60.260 ;
    END
  END ON[31]
  PIN ON[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 12.820 80.000 13.220 ;
    END
  END ON[3]
  PIN ON[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 14.500 80.000 14.900 ;
    END
  END ON[4]
  PIN ON[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 16.180 80.000 16.580 ;
    END
  END ON[5]
  PIN ON[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 17.860 80.000 18.260 ;
    END
  END ON[6]
  PIN ON[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 19.540 80.000 19.940 ;
    END
  END ON[7]
  PIN ON[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 21.220 80.000 21.620 ;
    END
  END ON[8]
  PIN ON[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 22.900 80.000 23.300 ;
    END
  END ON[9]
  PIN ON_N[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 8.620 80.000 9.020 ;
    END
  END ON_N[0]
  PIN ON_N[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 25.420 80.000 25.820 ;
    END
  END ON_N[10]
  PIN ON_N[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 27.100 80.000 27.500 ;
    END
  END ON_N[11]
  PIN ON_N[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 28.780 80.000 29.180 ;
    END
  END ON_N[12]
  PIN ON_N[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 30.460 80.000 30.860 ;
    END
  END ON_N[13]
  PIN ON_N[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 32.140 80.000 32.540 ;
    END
  END ON_N[14]
  PIN ON_N[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 33.820 80.000 34.220 ;
    END
  END ON_N[15]
  PIN ON_N[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 35.500 80.000 35.900 ;
    END
  END ON_N[16]
  PIN ON_N[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 37.180 80.000 37.580 ;
    END
  END ON_N[17]
  PIN ON_N[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 38.860 80.000 39.260 ;
    END
  END ON_N[18]
  PIN ON_N[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 40.540 80.000 40.940 ;
    END
  END ON_N[19]
  PIN ON_N[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 10.300 80.000 10.700 ;
    END
  END ON_N[1]
  PIN ON_N[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 42.220 80.000 42.620 ;
    END
  END ON_N[20]
  PIN ON_N[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 43.900 80.000 44.300 ;
    END
  END ON_N[21]
  PIN ON_N[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 45.580 80.000 45.980 ;
    END
  END ON_N[22]
  PIN ON_N[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 47.260 80.000 47.660 ;
    END
  END ON_N[23]
  PIN ON_N[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 48.940 80.000 49.340 ;
    END
  END ON_N[24]
  PIN ON_N[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 50.620 80.000 51.020 ;
    END
  END ON_N[25]
  PIN ON_N[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 52.300 80.000 52.700 ;
    END
  END ON_N[26]
  PIN ON_N[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 53.980 80.000 54.380 ;
    END
  END ON_N[27]
  PIN ON_N[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 55.660 80.000 56.060 ;
    END
  END ON_N[28]
  PIN ON_N[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 57.340 80.000 57.740 ;
    END
  END ON_N[29]
  PIN ON_N[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 11.980 80.000 12.380 ;
    END
  END ON_N[2]
  PIN ON_N[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 59.020 80.000 59.420 ;
    END
  END ON_N[30]
  PIN ON_N[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 60.700 80.000 61.100 ;
    END
  END ON_N[31]
  PIN ON_N[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 13.660 80.000 14.060 ;
    END
  END ON_N[3]
  PIN ON_N[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 15.340 80.000 15.740 ;
    END
  END ON_N[4]
  PIN ON_N[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 17.020 80.000 17.420 ;
    END
  END ON_N[5]
  PIN ON_N[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 18.700 80.000 19.100 ;
    END
  END ON_N[6]
  PIN ON_N[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 20.380 80.000 20.780 ;
    END
  END ON_N[7]
  PIN ON_N[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 22.060 80.000 22.460 ;
    END
  END ON_N[8]
  PIN ON_N[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal3 ;
        RECT 79.600 23.740 80.000 24.140 ;
    END
  END ON_N[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 21.580 3.560 23.780 64.480 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.660 22.480 77.020 24.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 15.380 3.560 17.580 64.480 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.660 16.280 77.020 18.480 ;
    END
  END VPWR
  PIN thermo[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 8.620 0.400 9.020 ;
    END
  END thermo[0]
  PIN thermo[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.420 0.400 25.820 ;
    END
  END thermo[10]
  PIN thermo[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 27.100 0.400 27.500 ;
    END
  END thermo[11]
  PIN thermo[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.780 0.400 29.180 ;
    END
  END thermo[12]
  PIN thermo[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.460 0.400 30.860 ;
    END
  END thermo[13]
  PIN thermo[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.140 0.400 32.540 ;
    END
  END thermo[14]
  PIN thermo[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.820 0.400 34.220 ;
    END
  END thermo[15]
  PIN thermo[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 35.500 0.400 35.900 ;
    END
  END thermo[16]
  PIN thermo[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 37.180 0.400 37.580 ;
    END
  END thermo[17]
  PIN thermo[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.860 0.400 39.260 ;
    END
  END thermo[18]
  PIN thermo[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.540 0.400 40.940 ;
    END
  END thermo[19]
  PIN thermo[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.300 0.400 10.700 ;
    END
  END thermo[1]
  PIN thermo[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.220 0.400 42.620 ;
    END
  END thermo[20]
  PIN thermo[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.900 0.400 44.300 ;
    END
  END thermo[21]
  PIN thermo[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.580 0.400 45.980 ;
    END
  END thermo[22]
  PIN thermo[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.260 0.400 47.660 ;
    END
  END thermo[23]
  PIN thermo[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.940 0.400 49.340 ;
    END
  END thermo[24]
  PIN thermo[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.620 0.400 51.020 ;
    END
  END thermo[25]
  PIN thermo[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.300 0.400 52.700 ;
    END
  END thermo[26]
  PIN thermo[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.980 0.400 54.380 ;
    END
  END thermo[27]
  PIN thermo[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 55.660 0.400 56.060 ;
    END
  END thermo[28]
  PIN thermo[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.340 0.400 57.740 ;
    END
  END thermo[29]
  PIN thermo[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.980 0.400 12.380 ;
    END
  END thermo[2]
  PIN thermo[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.020 0.400 59.420 ;
    END
  END thermo[30]
  PIN thermo[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.700 0.400 61.100 ;
    END
  END thermo[31]
  PIN thermo[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 13.660 0.400 14.060 ;
    END
  END thermo[3]
  PIN thermo[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.340 0.400 15.740 ;
    END
  END thermo[4]
  PIN thermo[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 17.020 0.400 17.420 ;
    END
  END thermo[5]
  PIN thermo[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 18.700 0.400 19.100 ;
    END
  END thermo[6]
  PIN thermo[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.380 0.400 20.780 ;
    END
  END thermo[7]
  PIN thermo[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.060 0.400 22.460 ;
    END
  END thermo[8]
  PIN thermo[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543400 ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.740 0.400 24.140 ;
    END
  END thermo[9]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 76.800 64.410 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 76.800 64.480 ;
      LAYER Metal2 ;
        RECT 4.215 3.635 76.425 64.405 ;
      LAYER Metal3 ;
        RECT 0.400 61.310 79.600 64.360 ;
        RECT 0.610 60.490 79.390 61.310 ;
        RECT 0.400 60.470 79.600 60.490 ;
        RECT 0.400 59.650 79.390 60.470 ;
        RECT 0.400 59.630 79.600 59.650 ;
        RECT 0.610 58.810 79.390 59.630 ;
        RECT 0.400 58.790 79.600 58.810 ;
        RECT 0.400 57.970 79.390 58.790 ;
        RECT 0.400 57.950 79.600 57.970 ;
        RECT 0.610 57.130 79.390 57.950 ;
        RECT 0.400 57.110 79.600 57.130 ;
        RECT 0.400 56.290 79.390 57.110 ;
        RECT 0.400 56.270 79.600 56.290 ;
        RECT 0.610 55.450 79.390 56.270 ;
        RECT 0.400 55.430 79.600 55.450 ;
        RECT 0.400 54.610 79.390 55.430 ;
        RECT 0.400 54.590 79.600 54.610 ;
        RECT 0.610 53.770 79.390 54.590 ;
        RECT 0.400 53.750 79.600 53.770 ;
        RECT 0.400 52.930 79.390 53.750 ;
        RECT 0.400 52.910 79.600 52.930 ;
        RECT 0.610 52.090 79.390 52.910 ;
        RECT 0.400 52.070 79.600 52.090 ;
        RECT 0.400 51.250 79.390 52.070 ;
        RECT 0.400 51.230 79.600 51.250 ;
        RECT 0.610 50.410 79.390 51.230 ;
        RECT 0.400 50.390 79.600 50.410 ;
        RECT 0.400 49.570 79.390 50.390 ;
        RECT 0.400 49.550 79.600 49.570 ;
        RECT 0.610 48.730 79.390 49.550 ;
        RECT 0.400 48.710 79.600 48.730 ;
        RECT 0.400 47.890 79.390 48.710 ;
        RECT 0.400 47.870 79.600 47.890 ;
        RECT 0.610 47.050 79.390 47.870 ;
        RECT 0.400 47.030 79.600 47.050 ;
        RECT 0.400 46.210 79.390 47.030 ;
        RECT 0.400 46.190 79.600 46.210 ;
        RECT 0.610 45.370 79.390 46.190 ;
        RECT 0.400 45.350 79.600 45.370 ;
        RECT 0.400 44.530 79.390 45.350 ;
        RECT 0.400 44.510 79.600 44.530 ;
        RECT 0.610 43.690 79.390 44.510 ;
        RECT 0.400 43.670 79.600 43.690 ;
        RECT 0.400 42.850 79.390 43.670 ;
        RECT 0.400 42.830 79.600 42.850 ;
        RECT 0.610 42.010 79.390 42.830 ;
        RECT 0.400 41.990 79.600 42.010 ;
        RECT 0.400 41.170 79.390 41.990 ;
        RECT 0.400 41.150 79.600 41.170 ;
        RECT 0.610 40.330 79.390 41.150 ;
        RECT 0.400 40.310 79.600 40.330 ;
        RECT 0.400 39.490 79.390 40.310 ;
        RECT 0.400 39.470 79.600 39.490 ;
        RECT 0.610 38.650 79.390 39.470 ;
        RECT 0.400 38.630 79.600 38.650 ;
        RECT 0.400 37.810 79.390 38.630 ;
        RECT 0.400 37.790 79.600 37.810 ;
        RECT 0.610 36.970 79.390 37.790 ;
        RECT 0.400 36.950 79.600 36.970 ;
        RECT 0.400 36.130 79.390 36.950 ;
        RECT 0.400 36.110 79.600 36.130 ;
        RECT 0.610 35.290 79.390 36.110 ;
        RECT 0.400 35.270 79.600 35.290 ;
        RECT 0.400 34.450 79.390 35.270 ;
        RECT 0.400 34.430 79.600 34.450 ;
        RECT 0.610 33.610 79.390 34.430 ;
        RECT 0.400 33.590 79.600 33.610 ;
        RECT 0.400 32.770 79.390 33.590 ;
        RECT 0.400 32.750 79.600 32.770 ;
        RECT 0.610 31.930 79.390 32.750 ;
        RECT 0.400 31.910 79.600 31.930 ;
        RECT 0.400 31.090 79.390 31.910 ;
        RECT 0.400 31.070 79.600 31.090 ;
        RECT 0.610 30.250 79.390 31.070 ;
        RECT 0.400 30.230 79.600 30.250 ;
        RECT 0.400 29.410 79.390 30.230 ;
        RECT 0.400 29.390 79.600 29.410 ;
        RECT 0.610 28.570 79.390 29.390 ;
        RECT 0.400 28.550 79.600 28.570 ;
        RECT 0.400 27.730 79.390 28.550 ;
        RECT 0.400 27.710 79.600 27.730 ;
        RECT 0.610 26.890 79.390 27.710 ;
        RECT 0.400 26.870 79.600 26.890 ;
        RECT 0.400 26.050 79.390 26.870 ;
        RECT 0.400 26.030 79.600 26.050 ;
        RECT 0.610 25.210 79.390 26.030 ;
        RECT 0.400 25.190 79.600 25.210 ;
        RECT 0.400 24.370 79.390 25.190 ;
        RECT 0.400 24.350 79.600 24.370 ;
        RECT 0.610 23.530 79.390 24.350 ;
        RECT 0.400 23.510 79.600 23.530 ;
        RECT 0.400 22.690 79.390 23.510 ;
        RECT 0.400 22.670 79.600 22.690 ;
        RECT 0.610 21.850 79.390 22.670 ;
        RECT 0.400 21.830 79.600 21.850 ;
        RECT 0.400 21.010 79.390 21.830 ;
        RECT 0.400 20.990 79.600 21.010 ;
        RECT 0.610 20.170 79.390 20.990 ;
        RECT 0.400 20.150 79.600 20.170 ;
        RECT 0.400 19.330 79.390 20.150 ;
        RECT 0.400 19.310 79.600 19.330 ;
        RECT 0.610 18.490 79.390 19.310 ;
        RECT 0.400 18.470 79.600 18.490 ;
        RECT 0.400 17.650 79.390 18.470 ;
        RECT 0.400 17.630 79.600 17.650 ;
        RECT 0.610 16.810 79.390 17.630 ;
        RECT 0.400 16.790 79.600 16.810 ;
        RECT 0.400 15.970 79.390 16.790 ;
        RECT 0.400 15.950 79.600 15.970 ;
        RECT 0.610 15.130 79.390 15.950 ;
        RECT 0.400 15.110 79.600 15.130 ;
        RECT 0.400 14.290 79.390 15.110 ;
        RECT 0.400 14.270 79.600 14.290 ;
        RECT 0.610 13.450 79.390 14.270 ;
        RECT 0.400 13.430 79.600 13.450 ;
        RECT 0.400 12.610 79.390 13.430 ;
        RECT 0.400 12.590 79.600 12.610 ;
        RECT 0.610 11.770 79.390 12.590 ;
        RECT 0.400 11.750 79.600 11.770 ;
        RECT 0.400 10.930 79.390 11.750 ;
        RECT 0.400 10.910 79.600 10.930 ;
        RECT 0.610 10.090 79.390 10.910 ;
        RECT 0.400 10.070 79.600 10.090 ;
        RECT 0.400 9.250 79.390 10.070 ;
        RECT 0.400 9.230 79.600 9.250 ;
        RECT 0.610 8.410 79.390 9.230 ;
        RECT 0.400 8.390 79.600 8.410 ;
        RECT 0.400 7.570 79.390 8.390 ;
        RECT 0.400 3.680 79.600 7.570 ;
  END
END non_overlap
END LIBRARY

