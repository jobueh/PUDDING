VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DAC2U128OUT4IN
  CLASS BLOCK ;
  FOREIGN DAC2U128OUT4IN ;
  ORIGIN 2.210 5.110 ;
  SIZE 134.420 BY 26.590 ;
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT -1.900 15.150 131.900 15.820 ;
    END
    PORT
      LAYER Metal1 ;
        RECT -1.900 17.200 131.900 17.700 ;
    END
    PORT
      LAYER Metal1 ;
        RECT -1.900 0.550 131.900 1.220 ;
    END
    PORT
      LAYER Metal1 ;
        RECT -1.900 -1.330 131.900 -0.830 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT -1.900 20.780 131.900 21.280 ;
    END
    PORT
      LAYER Metal1 ;
        RECT -1.900 -4.910 131.900 -4.410 ;
    END
  END VSS
  PIN VbiasP[1]
    ANTENNAGATEAREA 478.500000 ;
    ANTENNADIFFAREA 5.010000 ;
    PORT
      LAYER Metal1 ;
        RECT -1.000 10.040 131.000 14.970 ;
    END
  END VbiasP[1]
  PIN Iout
    ANTENNADIFFAREA 66.047997 ;
    PORT
      LAYER Metal1 ;
        RECT -1.900 7.835 131.900 8.535 ;
    END
  END Iout
  PIN VbiasP[0]
    ANTENNAGATEAREA 478.500000 ;
    ANTENNADIFFAREA 5.010000 ;
    PORT
      LAYER Metal1 ;
        RECT -1.000 1.400 131.000 6.330 ;
    END
  END VbiasP[0]
  PIN ON[64]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 128.130 20.990 128.420 21.280 ;
    END
  END ON[64]
  PIN ONB[64]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 127.580 20.990 127.870 21.280 ;
    END
  END ONB[64]
  PIN ON[65]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 126.130 20.990 126.420 21.280 ;
    END
  END ON[65]
  PIN ONB[65]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 125.580 20.990 125.870 21.280 ;
    END
  END ONB[65]
  PIN ON[66]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 124.130 20.990 124.420 21.280 ;
    END
  END ON[66]
  PIN ONB[66]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 123.580 20.990 123.870 21.280 ;
    END
  END ONB[66]
  PIN ON[67]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 122.130 20.990 122.420 21.280 ;
    END
  END ON[67]
  PIN ONB[67]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 121.580 20.990 121.870 21.280 ;
    END
  END ONB[67]
  PIN ON[68]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 120.130 20.990 120.420 21.280 ;
    END
  END ON[68]
  PIN ONB[68]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 119.580 20.990 119.870 21.280 ;
    END
  END ONB[68]
  PIN ON[69]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.130 20.990 118.420 21.280 ;
    END
  END ON[69]
  PIN ONB[69]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.580 20.990 117.870 21.280 ;
    END
  END ONB[69]
  PIN ON[70]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 116.130 20.990 116.420 21.280 ;
    END
  END ON[70]
  PIN ONB[70]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 115.580 20.990 115.870 21.280 ;
    END
  END ONB[70]
  PIN ON[71]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 114.130 20.990 114.420 21.280 ;
    END
  END ON[71]
  PIN ONB[71]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 113.580 20.990 113.870 21.280 ;
    END
  END ONB[71]
  PIN ON[72]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 112.130 20.990 112.420 21.280 ;
    END
  END ON[72]
  PIN ONB[72]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 111.580 20.990 111.870 21.280 ;
    END
  END ONB[72]
  PIN ON[73]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.130 20.990 110.420 21.280 ;
    END
  END ON[73]
  PIN ONB[73]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 109.580 20.990 109.870 21.280 ;
    END
  END ONB[73]
  PIN ON[74]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 108.130 20.990 108.420 21.280 ;
    END
  END ON[74]
  PIN ONB[74]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 107.580 20.990 107.870 21.280 ;
    END
  END ONB[74]
  PIN ON[75]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 106.130 20.990 106.420 21.280 ;
    END
  END ON[75]
  PIN ONB[75]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 105.580 20.990 105.870 21.280 ;
    END
  END ONB[75]
  PIN ON[76]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 104.130 20.990 104.420 21.280 ;
    END
  END ON[76]
  PIN ONB[76]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 103.580 20.990 103.870 21.280 ;
    END
  END ONB[76]
  PIN ON[77]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 102.130 20.990 102.420 21.280 ;
    END
  END ON[77]
  PIN ONB[77]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 101.580 20.990 101.870 21.280 ;
    END
  END ONB[77]
  PIN ON[78]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 100.130 20.990 100.420 21.280 ;
    END
  END ON[78]
  PIN ONB[78]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 99.580 20.990 99.870 21.280 ;
    END
  END ONB[78]
  PIN ON[79]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 98.130 20.990 98.420 21.280 ;
    END
  END ON[79]
  PIN ONB[79]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 97.580 20.990 97.870 21.280 ;
    END
  END ONB[79]
  PIN ON[80]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 96.130 20.990 96.420 21.280 ;
    END
  END ON[80]
  PIN ONB[80]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 95.580 20.990 95.870 21.280 ;
    END
  END ONB[80]
  PIN ON[81]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 94.130 20.990 94.420 21.280 ;
    END
  END ON[81]
  PIN ONB[81]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 93.580 20.990 93.870 21.280 ;
    END
  END ONB[81]
  PIN ON[82]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 92.130 20.990 92.420 21.280 ;
    END
  END ON[82]
  PIN ONB[82]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 91.580 20.990 91.870 21.280 ;
    END
  END ONB[82]
  PIN ON[83]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 90.130 20.990 90.420 21.280 ;
    END
  END ON[83]
  PIN ONB[83]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 89.580 20.990 89.870 21.280 ;
    END
  END ONB[83]
  PIN ON[84]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 88.130 20.990 88.420 21.280 ;
    END
  END ON[84]
  PIN ONB[84]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 87.580 20.990 87.870 21.280 ;
    END
  END ONB[84]
  PIN ON[85]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 86.130 20.990 86.420 21.280 ;
    END
  END ON[85]
  PIN ONB[85]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 85.580 20.990 85.870 21.280 ;
    END
  END ONB[85]
  PIN ON[86]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 84.130 20.990 84.420 21.280 ;
    END
  END ON[86]
  PIN ONB[86]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 83.580 20.990 83.870 21.280 ;
    END
  END ONB[86]
  PIN ON[87]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 82.130 20.990 82.420 21.280 ;
    END
  END ON[87]
  PIN ONB[87]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 81.580 20.990 81.870 21.280 ;
    END
  END ONB[87]
  PIN ON[88]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 80.130 20.990 80.420 21.280 ;
    END
  END ON[88]
  PIN ONB[88]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 79.580 20.990 79.870 21.280 ;
    END
  END ONB[88]
  PIN ON[89]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 78.130 20.990 78.420 21.280 ;
    END
  END ON[89]
  PIN ONB[89]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.580 20.990 77.870 21.280 ;
    END
  END ONB[89]
  PIN ON[90]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 76.130 20.990 76.420 21.280 ;
    END
  END ON[90]
  PIN ONB[90]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 75.580 20.990 75.870 21.280 ;
    END
  END ONB[90]
  PIN ON[91]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 74.130 20.990 74.420 21.280 ;
    END
  END ON[91]
  PIN ONB[91]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 73.580 20.990 73.870 21.280 ;
    END
  END ONB[91]
  PIN ON[92]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 72.130 20.990 72.420 21.280 ;
    END
  END ON[92]
  PIN ONB[92]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 71.580 20.990 71.870 21.280 ;
    END
  END ONB[92]
  PIN ON[93]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.130 20.990 70.420 21.280 ;
    END
  END ON[93]
  PIN ONB[93]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.580 20.990 69.870 21.280 ;
    END
  END ONB[93]
  PIN ON[94]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.130 20.990 68.420 21.280 ;
    END
  END ON[94]
  PIN ONB[94]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 67.580 20.990 67.870 21.280 ;
    END
  END ONB[94]
  PIN ON[95]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 66.130 20.990 66.420 21.280 ;
    END
  END ON[95]
  PIN ONB[95]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 65.580 20.990 65.870 21.280 ;
    END
  END ONB[95]
  PIN EN[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 130.130 20.990 130.420 21.280 ;
    END
  END EN[2]
  PIN ENB[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 129.580 20.990 129.870 21.280 ;
    END
  END ENB[2]
  PIN ON[97]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 62.130 20.990 62.420 21.280 ;
    END
  END ON[97]
  PIN ONB[97]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 61.580 20.990 61.870 21.280 ;
    END
  END ONB[97]
  PIN ON[98]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 60.130 20.990 60.420 21.280 ;
    END
  END ON[98]
  PIN ONB[98]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 59.580 20.990 59.870 21.280 ;
    END
  END ONB[98]
  PIN ON[99]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 58.130 20.990 58.420 21.280 ;
    END
  END ON[99]
  PIN ONB[99]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.580 20.990 57.870 21.280 ;
    END
  END ONB[99]
  PIN ON[100]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 56.130 20.990 56.420 21.280 ;
    END
  END ON[100]
  PIN ONB[100]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 55.580 20.990 55.870 21.280 ;
    END
  END ONB[100]
  PIN ON[101]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 54.130 20.990 54.420 21.280 ;
    END
  END ON[101]
  PIN ONB[101]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 53.580 20.990 53.870 21.280 ;
    END
  END ONB[101]
  PIN ON[102]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 52.130 20.990 52.420 21.280 ;
    END
  END ON[102]
  PIN ONB[102]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 51.580 20.990 51.870 21.280 ;
    END
  END ONB[102]
  PIN ON[103]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 50.130 20.990 50.420 21.280 ;
    END
  END ON[103]
  PIN ONB[103]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 49.580 20.990 49.870 21.280 ;
    END
  END ONB[103]
  PIN ON[104]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 48.130 20.990 48.420 21.280 ;
    END
  END ON[104]
  PIN ONB[104]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 47.580 20.990 47.870 21.280 ;
    END
  END ONB[104]
  PIN ON[105]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 46.130 20.990 46.420 21.280 ;
    END
  END ON[105]
  PIN ONB[105]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 45.580 20.990 45.870 21.280 ;
    END
  END ONB[105]
  PIN ON[106]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 44.130 20.990 44.420 21.280 ;
    END
  END ON[106]
  PIN ONB[106]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 43.580 20.990 43.870 21.280 ;
    END
  END ONB[106]
  PIN ON[107]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 42.130 20.990 42.420 21.280 ;
    END
  END ON[107]
  PIN ONB[107]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 41.580 20.990 41.870 21.280 ;
    END
  END ONB[107]
  PIN ON[108]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 40.130 20.990 40.420 21.280 ;
    END
  END ON[108]
  PIN ONB[108]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 39.580 20.990 39.870 21.280 ;
    END
  END ONB[108]
  PIN ON[109]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 38.130 20.990 38.420 21.280 ;
    END
  END ON[109]
  PIN ONB[109]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 37.580 20.990 37.870 21.280 ;
    END
  END ONB[109]
  PIN ON[110]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.130 20.990 36.420 21.280 ;
    END
  END ON[110]
  PIN ONB[110]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 35.580 20.990 35.870 21.280 ;
    END
  END ONB[110]
  PIN ON[111]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 34.130 20.990 34.420 21.280 ;
    END
  END ON[111]
  PIN ONB[111]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 33.580 20.990 33.870 21.280 ;
    END
  END ONB[111]
  PIN ON[112]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 32.130 20.990 32.420 21.280 ;
    END
  END ON[112]
  PIN ONB[112]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 31.580 20.990 31.870 21.280 ;
    END
  END ONB[112]
  PIN ON[113]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.130 20.990 30.420 21.280 ;
    END
  END ON[113]
  PIN ONB[113]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 29.580 20.990 29.870 21.280 ;
    END
  END ONB[113]
  PIN ON[114]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.130 20.990 28.420 21.280 ;
    END
  END ON[114]
  PIN ONB[114]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 27.580 20.990 27.870 21.280 ;
    END
  END ONB[114]
  PIN ON[115]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 26.130 20.990 26.420 21.280 ;
    END
  END ON[115]
  PIN ONB[115]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.580 20.990 25.870 21.280 ;
    END
  END ONB[115]
  PIN ON[116]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 24.130 20.990 24.420 21.280 ;
    END
  END ON[116]
  PIN ONB[116]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 23.580 20.990 23.870 21.280 ;
    END
  END ONB[116]
  PIN ON[117]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 22.130 20.990 22.420 21.280 ;
    END
  END ON[117]
  PIN ONB[117]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.580 20.990 21.870 21.280 ;
    END
  END ONB[117]
  PIN ON[118]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 20.130 20.990 20.420 21.280 ;
    END
  END ON[118]
  PIN ONB[118]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 19.580 20.990 19.870 21.280 ;
    END
  END ONB[118]
  PIN ON[119]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 18.130 20.990 18.420 21.280 ;
    END
  END ON[119]
  PIN ONB[119]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.580 20.990 17.870 21.280 ;
    END
  END ONB[119]
  PIN ON[120]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.130 20.990 16.420 21.280 ;
    END
  END ON[120]
  PIN ONB[120]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 15.580 20.990 15.870 21.280 ;
    END
  END ONB[120]
  PIN ON[121]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.130 20.990 14.420 21.280 ;
    END
  END ON[121]
  PIN ONB[121]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.580 20.990 13.870 21.280 ;
    END
  END ONB[121]
  PIN ON[122]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.130 20.990 12.420 21.280 ;
    END
  END ON[122]
  PIN ONB[122]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.580 20.990 11.870 21.280 ;
    END
  END ONB[122]
  PIN ON[123]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.130 20.990 10.420 21.280 ;
    END
  END ON[123]
  PIN ONB[123]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.580 20.990 9.870 21.280 ;
    END
  END ONB[123]
  PIN ON[124]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 8.130 20.990 8.420 21.280 ;
    END
  END ON[124]
  PIN ONB[124]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.580 20.990 7.870 21.280 ;
    END
  END ONB[124]
  PIN ON[125]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 6.130 20.990 6.420 21.280 ;
    END
  END ON[125]
  PIN ONB[125]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.580 20.990 5.870 21.280 ;
    END
  END ONB[125]
  PIN ON[126]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 4.130 20.990 4.420 21.280 ;
    END
  END ON[126]
  PIN ONB[126]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.580 20.990 3.870 21.280 ;
    END
  END ONB[126]
  PIN ON[127]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.130 20.990 2.420 21.280 ;
    END
  END ON[127]
  PIN ONB[127]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.580 20.990 1.870 21.280 ;
    END
  END ONB[127]
  PIN ON[96]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.130 20.990 64.420 21.280 ;
    END
  END ON[96]
  PIN ONB[96]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.580 20.990 63.870 21.280 ;
    END
  END ONB[96]
  PIN EN[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.130 20.990 0.420 21.280 ;
    END
  END EN[3]
  PIN ENB[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT -0.420 20.990 -0.130 21.280 ;
    END
  END ENB[3]
  PIN ON[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.580 -4.910 1.870 -4.620 ;
    END
  END ON[0]
  PIN ONB[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.130 -4.910 2.420 -4.620 ;
    END
  END ONB[0]
  PIN ON[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.580 -4.910 3.870 -4.620 ;
    END
  END ON[1]
  PIN ONB[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 4.130 -4.910 4.420 -4.620 ;
    END
  END ONB[1]
  PIN ON[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.580 -4.910 5.870 -4.620 ;
    END
  END ON[2]
  PIN ONB[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 6.130 -4.910 6.420 -4.620 ;
    END
  END ONB[2]
  PIN ON[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.580 -4.910 7.870 -4.620 ;
    END
  END ON[3]
  PIN ONB[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 8.130 -4.910 8.420 -4.620 ;
    END
  END ONB[3]
  PIN ON[4]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.580 -4.910 9.870 -4.620 ;
    END
  END ON[4]
  PIN ONB[4]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.130 -4.910 10.420 -4.620 ;
    END
  END ONB[4]
  PIN ON[5]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.580 -4.910 11.870 -4.620 ;
    END
  END ON[5]
  PIN ONB[5]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.130 -4.910 12.420 -4.620 ;
    END
  END ONB[5]
  PIN ON[6]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.580 -4.910 13.870 -4.620 ;
    END
  END ON[6]
  PIN ONB[6]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.130 -4.910 14.420 -4.620 ;
    END
  END ONB[6]
  PIN ON[7]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 15.580 -4.910 15.870 -4.620 ;
    END
  END ON[7]
  PIN ONB[7]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.130 -4.910 16.420 -4.620 ;
    END
  END ONB[7]
  PIN ON[8]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.580 -4.910 17.870 -4.620 ;
    END
  END ON[8]
  PIN ONB[8]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 18.130 -4.910 18.420 -4.620 ;
    END
  END ONB[8]
  PIN ON[9]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 19.580 -4.910 19.870 -4.620 ;
    END
  END ON[9]
  PIN ONB[9]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 20.130 -4.910 20.420 -4.620 ;
    END
  END ONB[9]
  PIN ON[10]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.580 -4.910 21.870 -4.620 ;
    END
  END ON[10]
  PIN ONB[10]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 22.130 -4.910 22.420 -4.620 ;
    END
  END ONB[10]
  PIN ON[11]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 23.580 -4.910 23.870 -4.620 ;
    END
  END ON[11]
  PIN ONB[11]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 24.130 -4.910 24.420 -4.620 ;
    END
  END ONB[11]
  PIN ON[12]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.580 -4.910 25.870 -4.620 ;
    END
  END ON[12]
  PIN ONB[12]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 26.130 -4.910 26.420 -4.620 ;
    END
  END ONB[12]
  PIN ON[13]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 27.580 -4.910 27.870 -4.620 ;
    END
  END ON[13]
  PIN ONB[13]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.130 -4.910 28.420 -4.620 ;
    END
  END ONB[13]
  PIN ON[14]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 29.580 -4.910 29.870 -4.620 ;
    END
  END ON[14]
  PIN ONB[14]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.130 -4.910 30.420 -4.620 ;
    END
  END ONB[14]
  PIN ON[15]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 31.580 -4.910 31.870 -4.620 ;
    END
  END ON[15]
  PIN ONB[15]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 32.130 -4.910 32.420 -4.620 ;
    END
  END ONB[15]
  PIN ON[16]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 33.580 -4.910 33.870 -4.620 ;
    END
  END ON[16]
  PIN ONB[16]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 34.130 -4.910 34.420 -4.620 ;
    END
  END ONB[16]
  PIN ON[17]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 35.580 -4.910 35.870 -4.620 ;
    END
  END ON[17]
  PIN ONB[17]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.130 -4.910 36.420 -4.620 ;
    END
  END ONB[17]
  PIN ON[18]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 37.580 -4.910 37.870 -4.620 ;
    END
  END ON[18]
  PIN ONB[18]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 38.130 -4.910 38.420 -4.620 ;
    END
  END ONB[18]
  PIN ON[19]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 39.580 -4.910 39.870 -4.620 ;
    END
  END ON[19]
  PIN ONB[19]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 40.130 -4.910 40.420 -4.620 ;
    END
  END ONB[19]
  PIN ON[20]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 41.580 -4.910 41.870 -4.620 ;
    END
  END ON[20]
  PIN ONB[20]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 42.130 -4.910 42.420 -4.620 ;
    END
  END ONB[20]
  PIN ON[21]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 43.580 -4.910 43.870 -4.620 ;
    END
  END ON[21]
  PIN ONB[21]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 44.130 -4.910 44.420 -4.620 ;
    END
  END ONB[21]
  PIN ON[22]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 45.580 -4.910 45.870 -4.620 ;
    END
  END ON[22]
  PIN ONB[22]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 46.130 -4.910 46.420 -4.620 ;
    END
  END ONB[22]
  PIN ON[23]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 47.580 -4.910 47.870 -4.620 ;
    END
  END ON[23]
  PIN ONB[23]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 48.130 -4.910 48.420 -4.620 ;
    END
  END ONB[23]
  PIN ON[24]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 49.580 -4.910 49.870 -4.620 ;
    END
  END ON[24]
  PIN ONB[24]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 50.130 -4.910 50.420 -4.620 ;
    END
  END ONB[24]
  PIN ON[25]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 51.580 -4.910 51.870 -4.620 ;
    END
  END ON[25]
  PIN ONB[25]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 52.130 -4.910 52.420 -4.620 ;
    END
  END ONB[25]
  PIN ON[26]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 53.580 -4.910 53.870 -4.620 ;
    END
  END ON[26]
  PIN ONB[26]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 54.130 -4.910 54.420 -4.620 ;
    END
  END ONB[26]
  PIN ON[27]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 55.580 -4.910 55.870 -4.620 ;
    END
  END ON[27]
  PIN ONB[27]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 56.130 -4.910 56.420 -4.620 ;
    END
  END ONB[27]
  PIN ON[28]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.580 -4.910 57.870 -4.620 ;
    END
  END ON[28]
  PIN ONB[28]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 58.130 -4.910 58.420 -4.620 ;
    END
  END ONB[28]
  PIN ON[29]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 59.580 -4.910 59.870 -4.620 ;
    END
  END ON[29]
  PIN ONB[29]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 60.130 -4.910 60.420 -4.620 ;
    END
  END ONB[29]
  PIN ON[30]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 61.580 -4.910 61.870 -4.620 ;
    END
  END ON[30]
  PIN ONB[30]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 62.130 -4.910 62.420 -4.620 ;
    END
  END ONB[30]
  PIN ON[31]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.580 -4.910 63.870 -4.620 ;
    END
  END ON[31]
  PIN ONB[31]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.130 -4.910 64.420 -4.620 ;
    END
  END ONB[31]
  PIN EN[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT -0.420 -4.910 -0.130 -4.620 ;
    END
  END EN[0]
  PIN ENB[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 0.130 -4.910 0.420 -4.620 ;
    END
  END ENB[0]
  PIN ON[33]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 67.580 -4.910 67.870 -4.620 ;
    END
  END ON[33]
  PIN ONB[33]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.130 -4.910 68.420 -4.620 ;
    END
  END ONB[33]
  PIN ON[34]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.580 -4.910 69.870 -4.620 ;
    END
  END ON[34]
  PIN ONB[34]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.130 -4.910 70.420 -4.620 ;
    END
  END ONB[34]
  PIN ON[35]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 71.580 -4.910 71.870 -4.620 ;
    END
  END ON[35]
  PIN ONB[35]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 72.130 -4.910 72.420 -4.620 ;
    END
  END ONB[35]
  PIN ON[36]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 73.580 -4.910 73.870 -4.620 ;
    END
  END ON[36]
  PIN ONB[36]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 74.130 -4.910 74.420 -4.620 ;
    END
  END ONB[36]
  PIN ON[37]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 75.580 -4.910 75.870 -4.620 ;
    END
  END ON[37]
  PIN ONB[37]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 76.130 -4.910 76.420 -4.620 ;
    END
  END ONB[37]
  PIN ON[38]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.580 -4.910 77.870 -4.620 ;
    END
  END ON[38]
  PIN ONB[38]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 78.130 -4.910 78.420 -4.620 ;
    END
  END ONB[38]
  PIN ON[39]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 79.580 -4.910 79.870 -4.620 ;
    END
  END ON[39]
  PIN ONB[39]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 80.130 -4.910 80.420 -4.620 ;
    END
  END ONB[39]
  PIN ON[40]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 81.580 -4.910 81.870 -4.620 ;
    END
  END ON[40]
  PIN ONB[40]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 82.130 -4.910 82.420 -4.620 ;
    END
  END ONB[40]
  PIN ON[41]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 83.580 -4.910 83.870 -4.620 ;
    END
  END ON[41]
  PIN ONB[41]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 84.130 -4.910 84.420 -4.620 ;
    END
  END ONB[41]
  PIN ON[42]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 85.580 -4.910 85.870 -4.620 ;
    END
  END ON[42]
  PIN ONB[42]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 86.130 -4.910 86.420 -4.620 ;
    END
  END ONB[42]
  PIN ON[43]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 87.580 -4.910 87.870 -4.620 ;
    END
  END ON[43]
  PIN ONB[43]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 88.130 -4.910 88.420 -4.620 ;
    END
  END ONB[43]
  PIN ON[44]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 89.580 -4.910 89.870 -4.620 ;
    END
  END ON[44]
  PIN ONB[44]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 90.130 -4.910 90.420 -4.620 ;
    END
  END ONB[44]
  PIN ON[45]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 91.580 -4.910 91.870 -4.620 ;
    END
  END ON[45]
  PIN ONB[45]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 92.130 -4.910 92.420 -4.620 ;
    END
  END ONB[45]
  PIN ON[46]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 93.580 -4.910 93.870 -4.620 ;
    END
  END ON[46]
  PIN ONB[46]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 94.130 -4.910 94.420 -4.620 ;
    END
  END ONB[46]
  PIN ON[47]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 95.580 -4.910 95.870 -4.620 ;
    END
  END ON[47]
  PIN ONB[47]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 96.130 -4.910 96.420 -4.620 ;
    END
  END ONB[47]
  PIN ON[48]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 97.580 -4.910 97.870 -4.620 ;
    END
  END ON[48]
  PIN ONB[48]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 98.130 -4.910 98.420 -4.620 ;
    END
  END ONB[48]
  PIN ON[49]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 99.580 -4.910 99.870 -4.620 ;
    END
  END ON[49]
  PIN ONB[49]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 100.130 -4.910 100.420 -4.620 ;
    END
  END ONB[49]
  PIN ON[50]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 101.580 -4.910 101.870 -4.620 ;
    END
  END ON[50]
  PIN ONB[50]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 102.130 -4.910 102.420 -4.620 ;
    END
  END ONB[50]
  PIN ON[51]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 103.580 -4.910 103.870 -4.620 ;
    END
  END ON[51]
  PIN ONB[51]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 104.130 -4.910 104.420 -4.620 ;
    END
  END ONB[51]
  PIN ON[52]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 105.580 -4.910 105.870 -4.620 ;
    END
  END ON[52]
  PIN ONB[52]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 106.130 -4.910 106.420 -4.620 ;
    END
  END ONB[52]
  PIN ON[53]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 107.580 -4.910 107.870 -4.620 ;
    END
  END ON[53]
  PIN ONB[53]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 108.130 -4.910 108.420 -4.620 ;
    END
  END ONB[53]
  PIN ON[54]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 109.580 -4.910 109.870 -4.620 ;
    END
  END ON[54]
  PIN ONB[54]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.130 -4.910 110.420 -4.620 ;
    END
  END ONB[54]
  PIN ON[55]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 111.580 -4.910 111.870 -4.620 ;
    END
  END ON[55]
  PIN ONB[55]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 112.130 -4.910 112.420 -4.620 ;
    END
  END ONB[55]
  PIN ON[56]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 113.580 -4.910 113.870 -4.620 ;
    END
  END ON[56]
  PIN ONB[56]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 114.130 -4.910 114.420 -4.620 ;
    END
  END ONB[56]
  PIN ON[57]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 115.580 -4.910 115.870 -4.620 ;
    END
  END ON[57]
  PIN ONB[57]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 116.130 -4.910 116.420 -4.620 ;
    END
  END ONB[57]
  PIN ON[58]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.580 -4.910 117.870 -4.620 ;
    END
  END ON[58]
  PIN ONB[58]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.130 -4.910 118.420 -4.620 ;
    END
  END ONB[58]
  PIN ON[59]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 119.580 -4.910 119.870 -4.620 ;
    END
  END ON[59]
  PIN ONB[59]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 120.130 -4.910 120.420 -4.620 ;
    END
  END ONB[59]
  PIN ON[60]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 121.580 -4.910 121.870 -4.620 ;
    END
  END ON[60]
  PIN ONB[60]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 122.130 -4.910 122.420 -4.620 ;
    END
  END ONB[60]
  PIN ON[61]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 123.580 -4.910 123.870 -4.620 ;
    END
  END ON[61]
  PIN ONB[61]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 124.130 -4.910 124.420 -4.620 ;
    END
  END ONB[61]
  PIN ON[62]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 125.580 -4.910 125.870 -4.620 ;
    END
  END ON[62]
  PIN ONB[62]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 126.130 -4.910 126.420 -4.620 ;
    END
  END ONB[62]
  PIN ON[63]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 127.580 -4.910 127.870 -4.620 ;
    END
  END ON[63]
  PIN ONB[63]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 128.130 -4.910 128.420 -4.620 ;
    END
  END ONB[63]
  PIN ON[32]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 65.580 -4.910 65.870 -4.620 ;
    END
  END ON[32]
  PIN ONB[32]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 66.130 -4.910 66.420 -4.620 ;
    END
  END ONB[32]
  PIN EN[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 129.580 -4.910 129.870 -4.620 ;
    END
  END EN[1]
  PIN ENB[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 130.130 -4.910 130.420 -4.620 ;
    END
  END ENB[1]
  PIN VcascP[1]
    ANTENNAGATEAREA 1.755000 ;
    ANTENNADIFFAREA 10.710000 ;
    PORT
      LAYER Metal3 ;
        RECT -1.900 16.020 131.900 16.720 ;
    END
  END VcascP[1]
  PIN VcascP[0]
    ANTENNAGATEAREA 1.755000 ;
    ANTENNADIFFAREA 10.710000 ;
    PORT
      LAYER Metal3 ;
        RECT -1.900 -0.350 131.900 0.350 ;
    END
  END VcascP[0]
  OBS
      LAYER GatPoly ;
        RECT -0.665 19.950 -0.145 20.130 ;
        RECT 0.145 19.950 0.665 20.130 ;
        RECT 1.335 19.950 1.855 20.130 ;
        RECT 2.145 19.950 2.665 20.130 ;
        RECT 3.335 19.950 3.855 20.130 ;
        RECT 4.145 19.950 4.665 20.130 ;
        RECT 5.335 19.950 5.855 20.130 ;
        RECT 6.145 19.950 6.665 20.130 ;
        RECT 7.335 19.950 7.855 20.130 ;
        RECT 8.145 19.950 8.665 20.130 ;
        RECT 9.335 19.950 9.855 20.130 ;
        RECT 10.145 19.950 10.665 20.130 ;
        RECT 11.335 19.950 11.855 20.130 ;
        RECT 12.145 19.950 12.665 20.130 ;
        RECT 13.335 19.950 13.855 20.130 ;
        RECT 14.145 19.950 14.665 20.130 ;
        RECT 15.335 19.950 15.855 20.130 ;
        RECT 16.145 19.950 16.665 20.130 ;
        RECT 17.335 19.950 17.855 20.130 ;
        RECT 18.145 19.950 18.665 20.130 ;
        RECT 19.335 19.950 19.855 20.130 ;
        RECT 20.145 19.950 20.665 20.130 ;
        RECT 21.335 19.950 21.855 20.130 ;
        RECT 22.145 19.950 22.665 20.130 ;
        RECT 23.335 19.950 23.855 20.130 ;
        RECT 24.145 19.950 24.665 20.130 ;
        RECT 25.335 19.950 25.855 20.130 ;
        RECT 26.145 19.950 26.665 20.130 ;
        RECT 27.335 19.950 27.855 20.130 ;
        RECT 28.145 19.950 28.665 20.130 ;
        RECT 29.335 19.950 29.855 20.130 ;
        RECT 30.145 19.950 30.665 20.130 ;
        RECT 31.335 19.950 31.855 20.130 ;
        RECT 32.145 19.950 32.665 20.130 ;
        RECT 33.335 19.950 33.855 20.130 ;
        RECT 34.145 19.950 34.665 20.130 ;
        RECT 35.335 19.950 35.855 20.130 ;
        RECT 36.145 19.950 36.665 20.130 ;
        RECT 37.335 19.950 37.855 20.130 ;
        RECT 38.145 19.950 38.665 20.130 ;
        RECT 39.335 19.950 39.855 20.130 ;
        RECT 40.145 19.950 40.665 20.130 ;
        RECT 41.335 19.950 41.855 20.130 ;
        RECT 42.145 19.950 42.665 20.130 ;
        RECT 43.335 19.950 43.855 20.130 ;
        RECT 44.145 19.950 44.665 20.130 ;
        RECT 45.335 19.950 45.855 20.130 ;
        RECT 46.145 19.950 46.665 20.130 ;
        RECT 47.335 19.950 47.855 20.130 ;
        RECT 48.145 19.950 48.665 20.130 ;
        RECT 49.335 19.950 49.855 20.130 ;
        RECT 50.145 19.950 50.665 20.130 ;
        RECT 51.335 19.950 51.855 20.130 ;
        RECT 52.145 19.950 52.665 20.130 ;
        RECT 53.335 19.950 53.855 20.130 ;
        RECT 54.145 19.950 54.665 20.130 ;
        RECT 55.335 19.950 55.855 20.130 ;
        RECT 56.145 19.950 56.665 20.130 ;
        RECT 57.335 19.950 57.855 20.130 ;
        RECT 58.145 19.950 58.665 20.130 ;
        RECT 59.335 19.950 59.855 20.130 ;
        RECT 60.145 19.950 60.665 20.130 ;
        RECT 61.335 19.950 61.855 20.130 ;
        RECT 62.145 19.950 62.665 20.130 ;
        RECT 63.335 19.950 63.855 20.130 ;
        RECT 64.145 19.950 64.665 20.130 ;
        RECT 65.335 19.950 65.855 20.130 ;
        RECT 66.145 19.950 66.665 20.130 ;
        RECT 67.335 19.950 67.855 20.130 ;
        RECT 68.145 19.950 68.665 20.130 ;
        RECT 69.335 19.950 69.855 20.130 ;
        RECT 70.145 19.950 70.665 20.130 ;
        RECT 71.335 19.950 71.855 20.130 ;
        RECT 72.145 19.950 72.665 20.130 ;
        RECT 73.335 19.950 73.855 20.130 ;
        RECT 74.145 19.950 74.665 20.130 ;
        RECT 75.335 19.950 75.855 20.130 ;
        RECT 76.145 19.950 76.665 20.130 ;
        RECT 77.335 19.950 77.855 20.130 ;
        RECT 78.145 19.950 78.665 20.130 ;
        RECT 79.335 19.950 79.855 20.130 ;
        RECT 80.145 19.950 80.665 20.130 ;
        RECT 81.335 19.950 81.855 20.130 ;
        RECT 82.145 19.950 82.665 20.130 ;
        RECT 83.335 19.950 83.855 20.130 ;
        RECT 84.145 19.950 84.665 20.130 ;
        RECT 85.335 19.950 85.855 20.130 ;
        RECT 86.145 19.950 86.665 20.130 ;
        RECT 87.335 19.950 87.855 20.130 ;
        RECT 88.145 19.950 88.665 20.130 ;
        RECT 89.335 19.950 89.855 20.130 ;
        RECT 90.145 19.950 90.665 20.130 ;
        RECT 91.335 19.950 91.855 20.130 ;
        RECT 92.145 19.950 92.665 20.130 ;
        RECT 93.335 19.950 93.855 20.130 ;
        RECT 94.145 19.950 94.665 20.130 ;
        RECT 95.335 19.950 95.855 20.130 ;
        RECT 96.145 19.950 96.665 20.130 ;
        RECT 97.335 19.950 97.855 20.130 ;
        RECT 98.145 19.950 98.665 20.130 ;
        RECT 99.335 19.950 99.855 20.130 ;
        RECT 100.145 19.950 100.665 20.130 ;
        RECT 101.335 19.950 101.855 20.130 ;
        RECT 102.145 19.950 102.665 20.130 ;
        RECT 103.335 19.950 103.855 20.130 ;
        RECT 104.145 19.950 104.665 20.130 ;
        RECT 105.335 19.950 105.855 20.130 ;
        RECT 106.145 19.950 106.665 20.130 ;
        RECT 107.335 19.950 107.855 20.130 ;
        RECT 108.145 19.950 108.665 20.130 ;
        RECT 109.335 19.950 109.855 20.130 ;
        RECT 110.145 19.950 110.665 20.130 ;
        RECT 111.335 19.950 111.855 20.130 ;
        RECT 112.145 19.950 112.665 20.130 ;
        RECT 113.335 19.950 113.855 20.130 ;
        RECT 114.145 19.950 114.665 20.130 ;
        RECT 115.335 19.950 115.855 20.130 ;
        RECT 116.145 19.950 116.665 20.130 ;
        RECT 117.335 19.950 117.855 20.130 ;
        RECT 118.145 19.950 118.665 20.130 ;
        RECT 119.335 19.950 119.855 20.130 ;
        RECT 120.145 19.950 120.665 20.130 ;
        RECT 121.335 19.950 121.855 20.130 ;
        RECT 122.145 19.950 122.665 20.130 ;
        RECT 123.335 19.950 123.855 20.130 ;
        RECT 124.145 19.950 124.665 20.130 ;
        RECT 125.335 19.950 125.855 20.130 ;
        RECT 126.145 19.950 126.665 20.130 ;
        RECT 127.335 19.950 127.855 20.130 ;
        RECT 128.145 19.950 128.665 20.130 ;
        RECT 129.335 19.950 129.855 20.130 ;
        RECT 130.145 19.950 130.665 20.130 ;
        RECT -0.665 19.620 -0.145 19.800 ;
        RECT -0.445 19.430 -0.145 19.620 ;
        RECT 0.145 19.620 0.665 19.800 ;
        RECT 1.335 19.620 1.855 19.800 ;
        RECT 0.145 19.250 0.445 19.620 ;
        RECT 1.555 19.430 1.855 19.620 ;
        RECT 2.145 19.620 2.665 19.800 ;
        RECT 3.335 19.620 3.855 19.800 ;
        RECT 2.145 19.250 2.445 19.620 ;
        RECT 3.555 19.430 3.855 19.620 ;
        RECT 4.145 19.620 4.665 19.800 ;
        RECT 5.335 19.620 5.855 19.800 ;
        RECT 4.145 19.250 4.445 19.620 ;
        RECT 5.555 19.430 5.855 19.620 ;
        RECT 6.145 19.620 6.665 19.800 ;
        RECT 7.335 19.620 7.855 19.800 ;
        RECT 6.145 19.250 6.445 19.620 ;
        RECT 7.555 19.430 7.855 19.620 ;
        RECT 8.145 19.620 8.665 19.800 ;
        RECT 9.335 19.620 9.855 19.800 ;
        RECT 8.145 19.250 8.445 19.620 ;
        RECT 9.555 19.430 9.855 19.620 ;
        RECT 10.145 19.620 10.665 19.800 ;
        RECT 11.335 19.620 11.855 19.800 ;
        RECT 10.145 19.250 10.445 19.620 ;
        RECT 11.555 19.430 11.855 19.620 ;
        RECT 12.145 19.620 12.665 19.800 ;
        RECT 13.335 19.620 13.855 19.800 ;
        RECT 12.145 19.250 12.445 19.620 ;
        RECT 13.555 19.430 13.855 19.620 ;
        RECT 14.145 19.620 14.665 19.800 ;
        RECT 15.335 19.620 15.855 19.800 ;
        RECT 14.145 19.250 14.445 19.620 ;
        RECT 15.555 19.430 15.855 19.620 ;
        RECT 16.145 19.620 16.665 19.800 ;
        RECT 17.335 19.620 17.855 19.800 ;
        RECT 16.145 19.250 16.445 19.620 ;
        RECT 17.555 19.430 17.855 19.620 ;
        RECT 18.145 19.620 18.665 19.800 ;
        RECT 19.335 19.620 19.855 19.800 ;
        RECT 18.145 19.250 18.445 19.620 ;
        RECT 19.555 19.430 19.855 19.620 ;
        RECT 20.145 19.620 20.665 19.800 ;
        RECT 21.335 19.620 21.855 19.800 ;
        RECT 20.145 19.250 20.445 19.620 ;
        RECT 21.555 19.430 21.855 19.620 ;
        RECT 22.145 19.620 22.665 19.800 ;
        RECT 23.335 19.620 23.855 19.800 ;
        RECT 22.145 19.250 22.445 19.620 ;
        RECT 23.555 19.430 23.855 19.620 ;
        RECT 24.145 19.620 24.665 19.800 ;
        RECT 25.335 19.620 25.855 19.800 ;
        RECT 24.145 19.250 24.445 19.620 ;
        RECT 25.555 19.430 25.855 19.620 ;
        RECT 26.145 19.620 26.665 19.800 ;
        RECT 27.335 19.620 27.855 19.800 ;
        RECT 26.145 19.250 26.445 19.620 ;
        RECT 27.555 19.430 27.855 19.620 ;
        RECT 28.145 19.620 28.665 19.800 ;
        RECT 29.335 19.620 29.855 19.800 ;
        RECT 28.145 19.250 28.445 19.620 ;
        RECT 29.555 19.430 29.855 19.620 ;
        RECT 30.145 19.620 30.665 19.800 ;
        RECT 31.335 19.620 31.855 19.800 ;
        RECT 30.145 19.250 30.445 19.620 ;
        RECT 31.555 19.430 31.855 19.620 ;
        RECT 32.145 19.620 32.665 19.800 ;
        RECT 33.335 19.620 33.855 19.800 ;
        RECT 32.145 19.250 32.445 19.620 ;
        RECT 33.555 19.430 33.855 19.620 ;
        RECT 34.145 19.620 34.665 19.800 ;
        RECT 35.335 19.620 35.855 19.800 ;
        RECT 34.145 19.250 34.445 19.620 ;
        RECT 35.555 19.430 35.855 19.620 ;
        RECT 36.145 19.620 36.665 19.800 ;
        RECT 37.335 19.620 37.855 19.800 ;
        RECT 36.145 19.250 36.445 19.620 ;
        RECT 37.555 19.430 37.855 19.620 ;
        RECT 38.145 19.620 38.665 19.800 ;
        RECT 39.335 19.620 39.855 19.800 ;
        RECT 38.145 19.250 38.445 19.620 ;
        RECT 39.555 19.430 39.855 19.620 ;
        RECT 40.145 19.620 40.665 19.800 ;
        RECT 41.335 19.620 41.855 19.800 ;
        RECT 40.145 19.250 40.445 19.620 ;
        RECT 41.555 19.430 41.855 19.620 ;
        RECT 42.145 19.620 42.665 19.800 ;
        RECT 43.335 19.620 43.855 19.800 ;
        RECT 42.145 19.250 42.445 19.620 ;
        RECT 43.555 19.430 43.855 19.620 ;
        RECT 44.145 19.620 44.665 19.800 ;
        RECT 45.335 19.620 45.855 19.800 ;
        RECT 44.145 19.250 44.445 19.620 ;
        RECT 45.555 19.430 45.855 19.620 ;
        RECT 46.145 19.620 46.665 19.800 ;
        RECT 47.335 19.620 47.855 19.800 ;
        RECT 46.145 19.250 46.445 19.620 ;
        RECT 47.555 19.430 47.855 19.620 ;
        RECT 48.145 19.620 48.665 19.800 ;
        RECT 49.335 19.620 49.855 19.800 ;
        RECT 48.145 19.250 48.445 19.620 ;
        RECT 49.555 19.430 49.855 19.620 ;
        RECT 50.145 19.620 50.665 19.800 ;
        RECT 51.335 19.620 51.855 19.800 ;
        RECT 50.145 19.250 50.445 19.620 ;
        RECT 51.555 19.430 51.855 19.620 ;
        RECT 52.145 19.620 52.665 19.800 ;
        RECT 53.335 19.620 53.855 19.800 ;
        RECT 52.145 19.250 52.445 19.620 ;
        RECT 53.555 19.430 53.855 19.620 ;
        RECT 54.145 19.620 54.665 19.800 ;
        RECT 55.335 19.620 55.855 19.800 ;
        RECT 54.145 19.250 54.445 19.620 ;
        RECT 55.555 19.430 55.855 19.620 ;
        RECT 56.145 19.620 56.665 19.800 ;
        RECT 57.335 19.620 57.855 19.800 ;
        RECT 56.145 19.250 56.445 19.620 ;
        RECT 57.555 19.430 57.855 19.620 ;
        RECT 58.145 19.620 58.665 19.800 ;
        RECT 59.335 19.620 59.855 19.800 ;
        RECT 58.145 19.250 58.445 19.620 ;
        RECT 59.555 19.430 59.855 19.620 ;
        RECT 60.145 19.620 60.665 19.800 ;
        RECT 61.335 19.620 61.855 19.800 ;
        RECT 60.145 19.250 60.445 19.620 ;
        RECT 61.555 19.430 61.855 19.620 ;
        RECT 62.145 19.620 62.665 19.800 ;
        RECT 63.335 19.620 63.855 19.800 ;
        RECT 62.145 19.250 62.445 19.620 ;
        RECT 63.555 19.430 63.855 19.620 ;
        RECT 64.145 19.620 64.665 19.800 ;
        RECT 65.335 19.620 65.855 19.800 ;
        RECT 64.145 19.250 64.445 19.620 ;
        RECT 65.555 19.430 65.855 19.620 ;
        RECT 66.145 19.620 66.665 19.800 ;
        RECT 67.335 19.620 67.855 19.800 ;
        RECT 66.145 19.250 66.445 19.620 ;
        RECT 67.555 19.430 67.855 19.620 ;
        RECT 68.145 19.620 68.665 19.800 ;
        RECT 69.335 19.620 69.855 19.800 ;
        RECT 68.145 19.250 68.445 19.620 ;
        RECT 69.555 19.430 69.855 19.620 ;
        RECT 70.145 19.620 70.665 19.800 ;
        RECT 71.335 19.620 71.855 19.800 ;
        RECT 70.145 19.250 70.445 19.620 ;
        RECT 71.555 19.430 71.855 19.620 ;
        RECT 72.145 19.620 72.665 19.800 ;
        RECT 73.335 19.620 73.855 19.800 ;
        RECT 72.145 19.250 72.445 19.620 ;
        RECT 73.555 19.430 73.855 19.620 ;
        RECT 74.145 19.620 74.665 19.800 ;
        RECT 75.335 19.620 75.855 19.800 ;
        RECT 74.145 19.250 74.445 19.620 ;
        RECT 75.555 19.430 75.855 19.620 ;
        RECT 76.145 19.620 76.665 19.800 ;
        RECT 77.335 19.620 77.855 19.800 ;
        RECT 76.145 19.250 76.445 19.620 ;
        RECT 77.555 19.430 77.855 19.620 ;
        RECT 78.145 19.620 78.665 19.800 ;
        RECT 79.335 19.620 79.855 19.800 ;
        RECT 78.145 19.250 78.445 19.620 ;
        RECT 79.555 19.430 79.855 19.620 ;
        RECT 80.145 19.620 80.665 19.800 ;
        RECT 81.335 19.620 81.855 19.800 ;
        RECT 80.145 19.250 80.445 19.620 ;
        RECT 81.555 19.430 81.855 19.620 ;
        RECT 82.145 19.620 82.665 19.800 ;
        RECT 83.335 19.620 83.855 19.800 ;
        RECT 82.145 19.250 82.445 19.620 ;
        RECT 83.555 19.430 83.855 19.620 ;
        RECT 84.145 19.620 84.665 19.800 ;
        RECT 85.335 19.620 85.855 19.800 ;
        RECT 84.145 19.250 84.445 19.620 ;
        RECT 85.555 19.430 85.855 19.620 ;
        RECT 86.145 19.620 86.665 19.800 ;
        RECT 87.335 19.620 87.855 19.800 ;
        RECT 86.145 19.250 86.445 19.620 ;
        RECT 87.555 19.430 87.855 19.620 ;
        RECT 88.145 19.620 88.665 19.800 ;
        RECT 89.335 19.620 89.855 19.800 ;
        RECT 88.145 19.250 88.445 19.620 ;
        RECT 89.555 19.430 89.855 19.620 ;
        RECT 90.145 19.620 90.665 19.800 ;
        RECT 91.335 19.620 91.855 19.800 ;
        RECT 90.145 19.250 90.445 19.620 ;
        RECT 91.555 19.430 91.855 19.620 ;
        RECT 92.145 19.620 92.665 19.800 ;
        RECT 93.335 19.620 93.855 19.800 ;
        RECT 92.145 19.250 92.445 19.620 ;
        RECT 93.555 19.430 93.855 19.620 ;
        RECT 94.145 19.620 94.665 19.800 ;
        RECT 95.335 19.620 95.855 19.800 ;
        RECT 94.145 19.250 94.445 19.620 ;
        RECT 95.555 19.430 95.855 19.620 ;
        RECT 96.145 19.620 96.665 19.800 ;
        RECT 97.335 19.620 97.855 19.800 ;
        RECT 96.145 19.250 96.445 19.620 ;
        RECT 97.555 19.430 97.855 19.620 ;
        RECT 98.145 19.620 98.665 19.800 ;
        RECT 99.335 19.620 99.855 19.800 ;
        RECT 98.145 19.250 98.445 19.620 ;
        RECT 99.555 19.430 99.855 19.620 ;
        RECT 100.145 19.620 100.665 19.800 ;
        RECT 101.335 19.620 101.855 19.800 ;
        RECT 100.145 19.250 100.445 19.620 ;
        RECT 101.555 19.430 101.855 19.620 ;
        RECT 102.145 19.620 102.665 19.800 ;
        RECT 103.335 19.620 103.855 19.800 ;
        RECT 102.145 19.250 102.445 19.620 ;
        RECT 103.555 19.430 103.855 19.620 ;
        RECT 104.145 19.620 104.665 19.800 ;
        RECT 105.335 19.620 105.855 19.800 ;
        RECT 104.145 19.250 104.445 19.620 ;
        RECT 105.555 19.430 105.855 19.620 ;
        RECT 106.145 19.620 106.665 19.800 ;
        RECT 107.335 19.620 107.855 19.800 ;
        RECT 106.145 19.250 106.445 19.620 ;
        RECT 107.555 19.430 107.855 19.620 ;
        RECT 108.145 19.620 108.665 19.800 ;
        RECT 109.335 19.620 109.855 19.800 ;
        RECT 108.145 19.250 108.445 19.620 ;
        RECT 109.555 19.430 109.855 19.620 ;
        RECT 110.145 19.620 110.665 19.800 ;
        RECT 111.335 19.620 111.855 19.800 ;
        RECT 110.145 19.250 110.445 19.620 ;
        RECT 111.555 19.430 111.855 19.620 ;
        RECT 112.145 19.620 112.665 19.800 ;
        RECT 113.335 19.620 113.855 19.800 ;
        RECT 112.145 19.250 112.445 19.620 ;
        RECT 113.555 19.430 113.855 19.620 ;
        RECT 114.145 19.620 114.665 19.800 ;
        RECT 115.335 19.620 115.855 19.800 ;
        RECT 114.145 19.250 114.445 19.620 ;
        RECT 115.555 19.430 115.855 19.620 ;
        RECT 116.145 19.620 116.665 19.800 ;
        RECT 117.335 19.620 117.855 19.800 ;
        RECT 116.145 19.250 116.445 19.620 ;
        RECT 117.555 19.430 117.855 19.620 ;
        RECT 118.145 19.620 118.665 19.800 ;
        RECT 119.335 19.620 119.855 19.800 ;
        RECT 118.145 19.250 118.445 19.620 ;
        RECT 119.555 19.430 119.855 19.620 ;
        RECT 120.145 19.620 120.665 19.800 ;
        RECT 121.335 19.620 121.855 19.800 ;
        RECT 120.145 19.250 120.445 19.620 ;
        RECT 121.555 19.430 121.855 19.620 ;
        RECT 122.145 19.620 122.665 19.800 ;
        RECT 123.335 19.620 123.855 19.800 ;
        RECT 122.145 19.250 122.445 19.620 ;
        RECT 123.555 19.430 123.855 19.620 ;
        RECT 124.145 19.620 124.665 19.800 ;
        RECT 125.335 19.620 125.855 19.800 ;
        RECT 124.145 19.250 124.445 19.620 ;
        RECT 125.555 19.430 125.855 19.620 ;
        RECT 126.145 19.620 126.665 19.800 ;
        RECT 127.335 19.620 127.855 19.800 ;
        RECT 126.145 19.250 126.445 19.620 ;
        RECT 127.555 19.430 127.855 19.620 ;
        RECT 128.145 19.620 128.665 19.800 ;
        RECT 129.335 19.620 129.855 19.800 ;
        RECT 128.145 19.250 128.445 19.620 ;
        RECT 129.555 19.430 129.855 19.620 ;
        RECT 130.145 19.620 130.665 19.800 ;
        RECT 130.145 19.250 130.445 19.620 ;
        RECT -0.895 18.950 0.445 19.250 ;
        RECT 1.105 18.950 2.445 19.250 ;
        RECT 3.105 18.950 4.445 19.250 ;
        RECT 5.105 18.950 6.445 19.250 ;
        RECT 7.105 18.950 8.445 19.250 ;
        RECT 9.105 18.950 10.445 19.250 ;
        RECT 11.105 18.950 12.445 19.250 ;
        RECT 13.105 18.950 14.445 19.250 ;
        RECT 15.105 18.950 16.445 19.250 ;
        RECT 17.105 18.950 18.445 19.250 ;
        RECT 19.105 18.950 20.445 19.250 ;
        RECT 21.105 18.950 22.445 19.250 ;
        RECT 23.105 18.950 24.445 19.250 ;
        RECT 25.105 18.950 26.445 19.250 ;
        RECT 27.105 18.950 28.445 19.250 ;
        RECT 29.105 18.950 30.445 19.250 ;
        RECT 31.105 18.950 32.445 19.250 ;
        RECT 33.105 18.950 34.445 19.250 ;
        RECT 35.105 18.950 36.445 19.250 ;
        RECT 37.105 18.950 38.445 19.250 ;
        RECT 39.105 18.950 40.445 19.250 ;
        RECT 41.105 18.950 42.445 19.250 ;
        RECT 43.105 18.950 44.445 19.250 ;
        RECT 45.105 18.950 46.445 19.250 ;
        RECT 47.105 18.950 48.445 19.250 ;
        RECT 49.105 18.950 50.445 19.250 ;
        RECT 51.105 18.950 52.445 19.250 ;
        RECT 53.105 18.950 54.445 19.250 ;
        RECT 55.105 18.950 56.445 19.250 ;
        RECT 57.105 18.950 58.445 19.250 ;
        RECT 59.105 18.950 60.445 19.250 ;
        RECT 61.105 18.950 62.445 19.250 ;
        RECT 63.105 18.950 64.445 19.250 ;
        RECT 65.105 18.950 66.445 19.250 ;
        RECT 67.105 18.950 68.445 19.250 ;
        RECT 69.105 18.950 70.445 19.250 ;
        RECT 71.105 18.950 72.445 19.250 ;
        RECT 73.105 18.950 74.445 19.250 ;
        RECT 75.105 18.950 76.445 19.250 ;
        RECT 77.105 18.950 78.445 19.250 ;
        RECT 79.105 18.950 80.445 19.250 ;
        RECT 81.105 18.950 82.445 19.250 ;
        RECT 83.105 18.950 84.445 19.250 ;
        RECT 85.105 18.950 86.445 19.250 ;
        RECT 87.105 18.950 88.445 19.250 ;
        RECT 89.105 18.950 90.445 19.250 ;
        RECT 91.105 18.950 92.445 19.250 ;
        RECT 93.105 18.950 94.445 19.250 ;
        RECT 95.105 18.950 96.445 19.250 ;
        RECT 97.105 18.950 98.445 19.250 ;
        RECT 99.105 18.950 100.445 19.250 ;
        RECT 101.105 18.950 102.445 19.250 ;
        RECT 103.105 18.950 104.445 19.250 ;
        RECT 105.105 18.950 106.445 19.250 ;
        RECT 107.105 18.950 108.445 19.250 ;
        RECT 109.105 18.950 110.445 19.250 ;
        RECT 111.105 18.950 112.445 19.250 ;
        RECT 113.105 18.950 114.445 19.250 ;
        RECT 115.105 18.950 116.445 19.250 ;
        RECT 117.105 18.950 118.445 19.250 ;
        RECT 119.105 18.950 120.445 19.250 ;
        RECT 121.105 18.950 122.445 19.250 ;
        RECT 123.105 18.950 124.445 19.250 ;
        RECT 125.105 18.950 126.445 19.250 ;
        RECT 127.105 18.950 128.445 19.250 ;
        RECT 129.105 18.950 130.445 19.250 ;
        RECT -0.490 18.470 -0.190 18.770 ;
        RECT -0.320 18.400 -0.190 18.470 ;
        RECT 0.190 18.470 0.490 18.770 ;
        RECT 1.510 18.470 1.810 18.770 ;
        RECT 0.190 18.400 0.320 18.470 ;
        RECT 1.680 18.400 1.810 18.470 ;
        RECT 2.190 18.470 2.490 18.770 ;
        RECT 3.510 18.470 3.810 18.770 ;
        RECT 2.190 18.400 2.320 18.470 ;
        RECT 3.680 18.400 3.810 18.470 ;
        RECT 4.190 18.470 4.490 18.770 ;
        RECT 5.510 18.470 5.810 18.770 ;
        RECT 4.190 18.400 4.320 18.470 ;
        RECT 5.680 18.400 5.810 18.470 ;
        RECT 6.190 18.470 6.490 18.770 ;
        RECT 7.510 18.470 7.810 18.770 ;
        RECT 6.190 18.400 6.320 18.470 ;
        RECT 7.680 18.400 7.810 18.470 ;
        RECT 8.190 18.470 8.490 18.770 ;
        RECT 9.510 18.470 9.810 18.770 ;
        RECT 8.190 18.400 8.320 18.470 ;
        RECT 9.680 18.400 9.810 18.470 ;
        RECT 10.190 18.470 10.490 18.770 ;
        RECT 11.510 18.470 11.810 18.770 ;
        RECT 10.190 18.400 10.320 18.470 ;
        RECT 11.680 18.400 11.810 18.470 ;
        RECT 12.190 18.470 12.490 18.770 ;
        RECT 13.510 18.470 13.810 18.770 ;
        RECT 12.190 18.400 12.320 18.470 ;
        RECT 13.680 18.400 13.810 18.470 ;
        RECT 14.190 18.470 14.490 18.770 ;
        RECT 15.510 18.470 15.810 18.770 ;
        RECT 14.190 18.400 14.320 18.470 ;
        RECT 15.680 18.400 15.810 18.470 ;
        RECT 16.190 18.470 16.490 18.770 ;
        RECT 17.510 18.470 17.810 18.770 ;
        RECT 16.190 18.400 16.320 18.470 ;
        RECT 17.680 18.400 17.810 18.470 ;
        RECT 18.190 18.470 18.490 18.770 ;
        RECT 19.510 18.470 19.810 18.770 ;
        RECT 18.190 18.400 18.320 18.470 ;
        RECT 19.680 18.400 19.810 18.470 ;
        RECT 20.190 18.470 20.490 18.770 ;
        RECT 21.510 18.470 21.810 18.770 ;
        RECT 20.190 18.400 20.320 18.470 ;
        RECT 21.680 18.400 21.810 18.470 ;
        RECT 22.190 18.470 22.490 18.770 ;
        RECT 23.510 18.470 23.810 18.770 ;
        RECT 22.190 18.400 22.320 18.470 ;
        RECT 23.680 18.400 23.810 18.470 ;
        RECT 24.190 18.470 24.490 18.770 ;
        RECT 25.510 18.470 25.810 18.770 ;
        RECT 24.190 18.400 24.320 18.470 ;
        RECT 25.680 18.400 25.810 18.470 ;
        RECT 26.190 18.470 26.490 18.770 ;
        RECT 27.510 18.470 27.810 18.770 ;
        RECT 26.190 18.400 26.320 18.470 ;
        RECT 27.680 18.400 27.810 18.470 ;
        RECT 28.190 18.470 28.490 18.770 ;
        RECT 29.510 18.470 29.810 18.770 ;
        RECT 28.190 18.400 28.320 18.470 ;
        RECT 29.680 18.400 29.810 18.470 ;
        RECT 30.190 18.470 30.490 18.770 ;
        RECT 31.510 18.470 31.810 18.770 ;
        RECT 30.190 18.400 30.320 18.470 ;
        RECT 31.680 18.400 31.810 18.470 ;
        RECT 32.190 18.470 32.490 18.770 ;
        RECT 33.510 18.470 33.810 18.770 ;
        RECT 32.190 18.400 32.320 18.470 ;
        RECT 33.680 18.400 33.810 18.470 ;
        RECT 34.190 18.470 34.490 18.770 ;
        RECT 35.510 18.470 35.810 18.770 ;
        RECT 34.190 18.400 34.320 18.470 ;
        RECT 35.680 18.400 35.810 18.470 ;
        RECT 36.190 18.470 36.490 18.770 ;
        RECT 37.510 18.470 37.810 18.770 ;
        RECT 36.190 18.400 36.320 18.470 ;
        RECT 37.680 18.400 37.810 18.470 ;
        RECT 38.190 18.470 38.490 18.770 ;
        RECT 39.510 18.470 39.810 18.770 ;
        RECT 38.190 18.400 38.320 18.470 ;
        RECT 39.680 18.400 39.810 18.470 ;
        RECT 40.190 18.470 40.490 18.770 ;
        RECT 41.510 18.470 41.810 18.770 ;
        RECT 40.190 18.400 40.320 18.470 ;
        RECT 41.680 18.400 41.810 18.470 ;
        RECT 42.190 18.470 42.490 18.770 ;
        RECT 43.510 18.470 43.810 18.770 ;
        RECT 42.190 18.400 42.320 18.470 ;
        RECT 43.680 18.400 43.810 18.470 ;
        RECT 44.190 18.470 44.490 18.770 ;
        RECT 45.510 18.470 45.810 18.770 ;
        RECT 44.190 18.400 44.320 18.470 ;
        RECT 45.680 18.400 45.810 18.470 ;
        RECT 46.190 18.470 46.490 18.770 ;
        RECT 47.510 18.470 47.810 18.770 ;
        RECT 46.190 18.400 46.320 18.470 ;
        RECT 47.680 18.400 47.810 18.470 ;
        RECT 48.190 18.470 48.490 18.770 ;
        RECT 49.510 18.470 49.810 18.770 ;
        RECT 48.190 18.400 48.320 18.470 ;
        RECT 49.680 18.400 49.810 18.470 ;
        RECT 50.190 18.470 50.490 18.770 ;
        RECT 51.510 18.470 51.810 18.770 ;
        RECT 50.190 18.400 50.320 18.470 ;
        RECT 51.680 18.400 51.810 18.470 ;
        RECT 52.190 18.470 52.490 18.770 ;
        RECT 53.510 18.470 53.810 18.770 ;
        RECT 52.190 18.400 52.320 18.470 ;
        RECT 53.680 18.400 53.810 18.470 ;
        RECT 54.190 18.470 54.490 18.770 ;
        RECT 55.510 18.470 55.810 18.770 ;
        RECT 54.190 18.400 54.320 18.470 ;
        RECT 55.680 18.400 55.810 18.470 ;
        RECT 56.190 18.470 56.490 18.770 ;
        RECT 57.510 18.470 57.810 18.770 ;
        RECT 56.190 18.400 56.320 18.470 ;
        RECT 57.680 18.400 57.810 18.470 ;
        RECT 58.190 18.470 58.490 18.770 ;
        RECT 59.510 18.470 59.810 18.770 ;
        RECT 58.190 18.400 58.320 18.470 ;
        RECT 59.680 18.400 59.810 18.470 ;
        RECT 60.190 18.470 60.490 18.770 ;
        RECT 61.510 18.470 61.810 18.770 ;
        RECT 60.190 18.400 60.320 18.470 ;
        RECT 61.680 18.400 61.810 18.470 ;
        RECT 62.190 18.470 62.490 18.770 ;
        RECT 63.510 18.470 63.810 18.770 ;
        RECT 62.190 18.400 62.320 18.470 ;
        RECT 63.680 18.400 63.810 18.470 ;
        RECT 64.190 18.470 64.490 18.770 ;
        RECT 65.510 18.470 65.810 18.770 ;
        RECT 64.190 18.400 64.320 18.470 ;
        RECT 65.680 18.400 65.810 18.470 ;
        RECT 66.190 18.470 66.490 18.770 ;
        RECT 67.510 18.470 67.810 18.770 ;
        RECT 66.190 18.400 66.320 18.470 ;
        RECT 67.680 18.400 67.810 18.470 ;
        RECT 68.190 18.470 68.490 18.770 ;
        RECT 69.510 18.470 69.810 18.770 ;
        RECT 68.190 18.400 68.320 18.470 ;
        RECT 69.680 18.400 69.810 18.470 ;
        RECT 70.190 18.470 70.490 18.770 ;
        RECT 71.510 18.470 71.810 18.770 ;
        RECT 70.190 18.400 70.320 18.470 ;
        RECT 71.680 18.400 71.810 18.470 ;
        RECT 72.190 18.470 72.490 18.770 ;
        RECT 73.510 18.470 73.810 18.770 ;
        RECT 72.190 18.400 72.320 18.470 ;
        RECT 73.680 18.400 73.810 18.470 ;
        RECT 74.190 18.470 74.490 18.770 ;
        RECT 75.510 18.470 75.810 18.770 ;
        RECT 74.190 18.400 74.320 18.470 ;
        RECT 75.680 18.400 75.810 18.470 ;
        RECT 76.190 18.470 76.490 18.770 ;
        RECT 77.510 18.470 77.810 18.770 ;
        RECT 76.190 18.400 76.320 18.470 ;
        RECT 77.680 18.400 77.810 18.470 ;
        RECT 78.190 18.470 78.490 18.770 ;
        RECT 79.510 18.470 79.810 18.770 ;
        RECT 78.190 18.400 78.320 18.470 ;
        RECT 79.680 18.400 79.810 18.470 ;
        RECT 80.190 18.470 80.490 18.770 ;
        RECT 81.510 18.470 81.810 18.770 ;
        RECT 80.190 18.400 80.320 18.470 ;
        RECT 81.680 18.400 81.810 18.470 ;
        RECT 82.190 18.470 82.490 18.770 ;
        RECT 83.510 18.470 83.810 18.770 ;
        RECT 82.190 18.400 82.320 18.470 ;
        RECT 83.680 18.400 83.810 18.470 ;
        RECT 84.190 18.470 84.490 18.770 ;
        RECT 85.510 18.470 85.810 18.770 ;
        RECT 84.190 18.400 84.320 18.470 ;
        RECT 85.680 18.400 85.810 18.470 ;
        RECT 86.190 18.470 86.490 18.770 ;
        RECT 87.510 18.470 87.810 18.770 ;
        RECT 86.190 18.400 86.320 18.470 ;
        RECT 87.680 18.400 87.810 18.470 ;
        RECT 88.190 18.470 88.490 18.770 ;
        RECT 89.510 18.470 89.810 18.770 ;
        RECT 88.190 18.400 88.320 18.470 ;
        RECT 89.680 18.400 89.810 18.470 ;
        RECT 90.190 18.470 90.490 18.770 ;
        RECT 91.510 18.470 91.810 18.770 ;
        RECT 90.190 18.400 90.320 18.470 ;
        RECT 91.680 18.400 91.810 18.470 ;
        RECT 92.190 18.470 92.490 18.770 ;
        RECT 93.510 18.470 93.810 18.770 ;
        RECT 92.190 18.400 92.320 18.470 ;
        RECT 93.680 18.400 93.810 18.470 ;
        RECT 94.190 18.470 94.490 18.770 ;
        RECT 95.510 18.470 95.810 18.770 ;
        RECT 94.190 18.400 94.320 18.470 ;
        RECT 95.680 18.400 95.810 18.470 ;
        RECT 96.190 18.470 96.490 18.770 ;
        RECT 97.510 18.470 97.810 18.770 ;
        RECT 96.190 18.400 96.320 18.470 ;
        RECT 97.680 18.400 97.810 18.470 ;
        RECT 98.190 18.470 98.490 18.770 ;
        RECT 99.510 18.470 99.810 18.770 ;
        RECT 98.190 18.400 98.320 18.470 ;
        RECT 99.680 18.400 99.810 18.470 ;
        RECT 100.190 18.470 100.490 18.770 ;
        RECT 101.510 18.470 101.810 18.770 ;
        RECT 100.190 18.400 100.320 18.470 ;
        RECT 101.680 18.400 101.810 18.470 ;
        RECT 102.190 18.470 102.490 18.770 ;
        RECT 103.510 18.470 103.810 18.770 ;
        RECT 102.190 18.400 102.320 18.470 ;
        RECT 103.680 18.400 103.810 18.470 ;
        RECT 104.190 18.470 104.490 18.770 ;
        RECT 105.510 18.470 105.810 18.770 ;
        RECT 104.190 18.400 104.320 18.470 ;
        RECT 105.680 18.400 105.810 18.470 ;
        RECT 106.190 18.470 106.490 18.770 ;
        RECT 107.510 18.470 107.810 18.770 ;
        RECT 106.190 18.400 106.320 18.470 ;
        RECT 107.680 18.400 107.810 18.470 ;
        RECT 108.190 18.470 108.490 18.770 ;
        RECT 109.510 18.470 109.810 18.770 ;
        RECT 108.190 18.400 108.320 18.470 ;
        RECT 109.680 18.400 109.810 18.470 ;
        RECT 110.190 18.470 110.490 18.770 ;
        RECT 111.510 18.470 111.810 18.770 ;
        RECT 110.190 18.400 110.320 18.470 ;
        RECT 111.680 18.400 111.810 18.470 ;
        RECT 112.190 18.470 112.490 18.770 ;
        RECT 113.510 18.470 113.810 18.770 ;
        RECT 112.190 18.400 112.320 18.470 ;
        RECT 113.680 18.400 113.810 18.470 ;
        RECT 114.190 18.470 114.490 18.770 ;
        RECT 115.510 18.470 115.810 18.770 ;
        RECT 114.190 18.400 114.320 18.470 ;
        RECT 115.680 18.400 115.810 18.470 ;
        RECT 116.190 18.470 116.490 18.770 ;
        RECT 117.510 18.470 117.810 18.770 ;
        RECT 116.190 18.400 116.320 18.470 ;
        RECT 117.680 18.400 117.810 18.470 ;
        RECT 118.190 18.470 118.490 18.770 ;
        RECT 119.510 18.470 119.810 18.770 ;
        RECT 118.190 18.400 118.320 18.470 ;
        RECT 119.680 18.400 119.810 18.470 ;
        RECT 120.190 18.470 120.490 18.770 ;
        RECT 121.510 18.470 121.810 18.770 ;
        RECT 120.190 18.400 120.320 18.470 ;
        RECT 121.680 18.400 121.810 18.470 ;
        RECT 122.190 18.470 122.490 18.770 ;
        RECT 123.510 18.470 123.810 18.770 ;
        RECT 122.190 18.400 122.320 18.470 ;
        RECT 123.680 18.400 123.810 18.470 ;
        RECT 124.190 18.470 124.490 18.770 ;
        RECT 125.510 18.470 125.810 18.770 ;
        RECT 124.190 18.400 124.320 18.470 ;
        RECT 125.680 18.400 125.810 18.470 ;
        RECT 126.190 18.470 126.490 18.770 ;
        RECT 127.510 18.470 127.810 18.770 ;
        RECT 126.190 18.400 126.320 18.470 ;
        RECT 127.680 18.400 127.810 18.470 ;
        RECT 128.190 18.470 128.490 18.770 ;
        RECT 129.510 18.470 129.810 18.770 ;
        RECT 128.190 18.400 128.320 18.470 ;
        RECT 129.680 18.400 129.810 18.470 ;
        RECT 130.190 18.470 130.490 18.770 ;
        RECT 130.190 18.400 130.320 18.470 ;
        RECT -0.320 17.920 -0.190 18.100 ;
        RECT 0.190 17.920 0.320 18.100 ;
        RECT 1.680 17.920 1.810 18.100 ;
        RECT 2.190 17.920 2.320 18.100 ;
        RECT 3.680 17.920 3.810 18.100 ;
        RECT 4.190 17.920 4.320 18.100 ;
        RECT 5.680 17.920 5.810 18.100 ;
        RECT 6.190 17.920 6.320 18.100 ;
        RECT 7.680 17.920 7.810 18.100 ;
        RECT 8.190 17.920 8.320 18.100 ;
        RECT 9.680 17.920 9.810 18.100 ;
        RECT 10.190 17.920 10.320 18.100 ;
        RECT 11.680 17.920 11.810 18.100 ;
        RECT 12.190 17.920 12.320 18.100 ;
        RECT 13.680 17.920 13.810 18.100 ;
        RECT 14.190 17.920 14.320 18.100 ;
        RECT 15.680 17.920 15.810 18.100 ;
        RECT 16.190 17.920 16.320 18.100 ;
        RECT 17.680 17.920 17.810 18.100 ;
        RECT 18.190 17.920 18.320 18.100 ;
        RECT 19.680 17.920 19.810 18.100 ;
        RECT 20.190 17.920 20.320 18.100 ;
        RECT 21.680 17.920 21.810 18.100 ;
        RECT 22.190 17.920 22.320 18.100 ;
        RECT 23.680 17.920 23.810 18.100 ;
        RECT 24.190 17.920 24.320 18.100 ;
        RECT 25.680 17.920 25.810 18.100 ;
        RECT 26.190 17.920 26.320 18.100 ;
        RECT 27.680 17.920 27.810 18.100 ;
        RECT 28.190 17.920 28.320 18.100 ;
        RECT 29.680 17.920 29.810 18.100 ;
        RECT 30.190 17.920 30.320 18.100 ;
        RECT 31.680 17.920 31.810 18.100 ;
        RECT 32.190 17.920 32.320 18.100 ;
        RECT 33.680 17.920 33.810 18.100 ;
        RECT 34.190 17.920 34.320 18.100 ;
        RECT 35.680 17.920 35.810 18.100 ;
        RECT 36.190 17.920 36.320 18.100 ;
        RECT 37.680 17.920 37.810 18.100 ;
        RECT 38.190 17.920 38.320 18.100 ;
        RECT 39.680 17.920 39.810 18.100 ;
        RECT 40.190 17.920 40.320 18.100 ;
        RECT 41.680 17.920 41.810 18.100 ;
        RECT 42.190 17.920 42.320 18.100 ;
        RECT 43.680 17.920 43.810 18.100 ;
        RECT 44.190 17.920 44.320 18.100 ;
        RECT 45.680 17.920 45.810 18.100 ;
        RECT 46.190 17.920 46.320 18.100 ;
        RECT 47.680 17.920 47.810 18.100 ;
        RECT 48.190 17.920 48.320 18.100 ;
        RECT 49.680 17.920 49.810 18.100 ;
        RECT 50.190 17.920 50.320 18.100 ;
        RECT 51.680 17.920 51.810 18.100 ;
        RECT 52.190 17.920 52.320 18.100 ;
        RECT 53.680 17.920 53.810 18.100 ;
        RECT 54.190 17.920 54.320 18.100 ;
        RECT 55.680 17.920 55.810 18.100 ;
        RECT 56.190 17.920 56.320 18.100 ;
        RECT 57.680 17.920 57.810 18.100 ;
        RECT 58.190 17.920 58.320 18.100 ;
        RECT 59.680 17.920 59.810 18.100 ;
        RECT 60.190 17.920 60.320 18.100 ;
        RECT 61.680 17.920 61.810 18.100 ;
        RECT 62.190 17.920 62.320 18.100 ;
        RECT 63.680 17.920 63.810 18.100 ;
        RECT 64.190 17.920 64.320 18.100 ;
        RECT 65.680 17.920 65.810 18.100 ;
        RECT 66.190 17.920 66.320 18.100 ;
        RECT 67.680 17.920 67.810 18.100 ;
        RECT 68.190 17.920 68.320 18.100 ;
        RECT 69.680 17.920 69.810 18.100 ;
        RECT 70.190 17.920 70.320 18.100 ;
        RECT 71.680 17.920 71.810 18.100 ;
        RECT 72.190 17.920 72.320 18.100 ;
        RECT 73.680 17.920 73.810 18.100 ;
        RECT 74.190 17.920 74.320 18.100 ;
        RECT 75.680 17.920 75.810 18.100 ;
        RECT 76.190 17.920 76.320 18.100 ;
        RECT 77.680 17.920 77.810 18.100 ;
        RECT 78.190 17.920 78.320 18.100 ;
        RECT 79.680 17.920 79.810 18.100 ;
        RECT 80.190 17.920 80.320 18.100 ;
        RECT 81.680 17.920 81.810 18.100 ;
        RECT 82.190 17.920 82.320 18.100 ;
        RECT 83.680 17.920 83.810 18.100 ;
        RECT 84.190 17.920 84.320 18.100 ;
        RECT 85.680 17.920 85.810 18.100 ;
        RECT 86.190 17.920 86.320 18.100 ;
        RECT 87.680 17.920 87.810 18.100 ;
        RECT 88.190 17.920 88.320 18.100 ;
        RECT 89.680 17.920 89.810 18.100 ;
        RECT 90.190 17.920 90.320 18.100 ;
        RECT 91.680 17.920 91.810 18.100 ;
        RECT 92.190 17.920 92.320 18.100 ;
        RECT 93.680 17.920 93.810 18.100 ;
        RECT 94.190 17.920 94.320 18.100 ;
        RECT 95.680 17.920 95.810 18.100 ;
        RECT 96.190 17.920 96.320 18.100 ;
        RECT 97.680 17.920 97.810 18.100 ;
        RECT 98.190 17.920 98.320 18.100 ;
        RECT 99.680 17.920 99.810 18.100 ;
        RECT 100.190 17.920 100.320 18.100 ;
        RECT 101.680 17.920 101.810 18.100 ;
        RECT 102.190 17.920 102.320 18.100 ;
        RECT 103.680 17.920 103.810 18.100 ;
        RECT 104.190 17.920 104.320 18.100 ;
        RECT 105.680 17.920 105.810 18.100 ;
        RECT 106.190 17.920 106.320 18.100 ;
        RECT 107.680 17.920 107.810 18.100 ;
        RECT 108.190 17.920 108.320 18.100 ;
        RECT 109.680 17.920 109.810 18.100 ;
        RECT 110.190 17.920 110.320 18.100 ;
        RECT 111.680 17.920 111.810 18.100 ;
        RECT 112.190 17.920 112.320 18.100 ;
        RECT 113.680 17.920 113.810 18.100 ;
        RECT 114.190 17.920 114.320 18.100 ;
        RECT 115.680 17.920 115.810 18.100 ;
        RECT 116.190 17.920 116.320 18.100 ;
        RECT 117.680 17.920 117.810 18.100 ;
        RECT 118.190 17.920 118.320 18.100 ;
        RECT 119.680 17.920 119.810 18.100 ;
        RECT 120.190 17.920 120.320 18.100 ;
        RECT 121.680 17.920 121.810 18.100 ;
        RECT 122.190 17.920 122.320 18.100 ;
        RECT 123.680 17.920 123.810 18.100 ;
        RECT 124.190 17.920 124.320 18.100 ;
        RECT 125.680 17.920 125.810 18.100 ;
        RECT 126.190 17.920 126.320 18.100 ;
        RECT 127.680 17.920 127.810 18.100 ;
        RECT 128.190 17.920 128.320 18.100 ;
        RECT 129.680 17.920 129.810 18.100 ;
        RECT 130.190 17.920 130.320 18.100 ;
        RECT -0.490 16.720 -0.190 17.020 ;
        RECT -0.320 16.520 -0.190 16.720 ;
        RECT 0.190 16.720 0.490 17.020 ;
        RECT 1.510 16.720 1.810 17.020 ;
        RECT 0.190 16.520 0.320 16.720 ;
        RECT 1.680 16.520 1.810 16.720 ;
        RECT 2.190 16.720 2.490 17.020 ;
        RECT 3.510 16.720 3.810 17.020 ;
        RECT 2.190 16.520 2.320 16.720 ;
        RECT 3.680 16.520 3.810 16.720 ;
        RECT 4.190 16.720 4.490 17.020 ;
        RECT 5.510 16.720 5.810 17.020 ;
        RECT 4.190 16.520 4.320 16.720 ;
        RECT 5.680 16.520 5.810 16.720 ;
        RECT 6.190 16.720 6.490 17.020 ;
        RECT 7.510 16.720 7.810 17.020 ;
        RECT 6.190 16.520 6.320 16.720 ;
        RECT 7.680 16.520 7.810 16.720 ;
        RECT 8.190 16.720 8.490 17.020 ;
        RECT 9.510 16.720 9.810 17.020 ;
        RECT 8.190 16.520 8.320 16.720 ;
        RECT 9.680 16.520 9.810 16.720 ;
        RECT 10.190 16.720 10.490 17.020 ;
        RECT 11.510 16.720 11.810 17.020 ;
        RECT 10.190 16.520 10.320 16.720 ;
        RECT 11.680 16.520 11.810 16.720 ;
        RECT 12.190 16.720 12.490 17.020 ;
        RECT 13.510 16.720 13.810 17.020 ;
        RECT 12.190 16.520 12.320 16.720 ;
        RECT 13.680 16.520 13.810 16.720 ;
        RECT 14.190 16.720 14.490 17.020 ;
        RECT 15.510 16.720 15.810 17.020 ;
        RECT 14.190 16.520 14.320 16.720 ;
        RECT 15.680 16.520 15.810 16.720 ;
        RECT 16.190 16.720 16.490 17.020 ;
        RECT 17.510 16.720 17.810 17.020 ;
        RECT 16.190 16.520 16.320 16.720 ;
        RECT 17.680 16.520 17.810 16.720 ;
        RECT 18.190 16.720 18.490 17.020 ;
        RECT 19.510 16.720 19.810 17.020 ;
        RECT 18.190 16.520 18.320 16.720 ;
        RECT 19.680 16.520 19.810 16.720 ;
        RECT 20.190 16.720 20.490 17.020 ;
        RECT 21.510 16.720 21.810 17.020 ;
        RECT 20.190 16.520 20.320 16.720 ;
        RECT 21.680 16.520 21.810 16.720 ;
        RECT 22.190 16.720 22.490 17.020 ;
        RECT 23.510 16.720 23.810 17.020 ;
        RECT 22.190 16.520 22.320 16.720 ;
        RECT 23.680 16.520 23.810 16.720 ;
        RECT 24.190 16.720 24.490 17.020 ;
        RECT 25.510 16.720 25.810 17.020 ;
        RECT 24.190 16.520 24.320 16.720 ;
        RECT 25.680 16.520 25.810 16.720 ;
        RECT 26.190 16.720 26.490 17.020 ;
        RECT 27.510 16.720 27.810 17.020 ;
        RECT 26.190 16.520 26.320 16.720 ;
        RECT 27.680 16.520 27.810 16.720 ;
        RECT 28.190 16.720 28.490 17.020 ;
        RECT 29.510 16.720 29.810 17.020 ;
        RECT 28.190 16.520 28.320 16.720 ;
        RECT 29.680 16.520 29.810 16.720 ;
        RECT 30.190 16.720 30.490 17.020 ;
        RECT 31.510 16.720 31.810 17.020 ;
        RECT 30.190 16.520 30.320 16.720 ;
        RECT 31.680 16.520 31.810 16.720 ;
        RECT 32.190 16.720 32.490 17.020 ;
        RECT 33.510 16.720 33.810 17.020 ;
        RECT 32.190 16.520 32.320 16.720 ;
        RECT 33.680 16.520 33.810 16.720 ;
        RECT 34.190 16.720 34.490 17.020 ;
        RECT 35.510 16.720 35.810 17.020 ;
        RECT 34.190 16.520 34.320 16.720 ;
        RECT 35.680 16.520 35.810 16.720 ;
        RECT 36.190 16.720 36.490 17.020 ;
        RECT 37.510 16.720 37.810 17.020 ;
        RECT 36.190 16.520 36.320 16.720 ;
        RECT 37.680 16.520 37.810 16.720 ;
        RECT 38.190 16.720 38.490 17.020 ;
        RECT 39.510 16.720 39.810 17.020 ;
        RECT 38.190 16.520 38.320 16.720 ;
        RECT 39.680 16.520 39.810 16.720 ;
        RECT 40.190 16.720 40.490 17.020 ;
        RECT 41.510 16.720 41.810 17.020 ;
        RECT 40.190 16.520 40.320 16.720 ;
        RECT 41.680 16.520 41.810 16.720 ;
        RECT 42.190 16.720 42.490 17.020 ;
        RECT 43.510 16.720 43.810 17.020 ;
        RECT 42.190 16.520 42.320 16.720 ;
        RECT 43.680 16.520 43.810 16.720 ;
        RECT 44.190 16.720 44.490 17.020 ;
        RECT 45.510 16.720 45.810 17.020 ;
        RECT 44.190 16.520 44.320 16.720 ;
        RECT 45.680 16.520 45.810 16.720 ;
        RECT 46.190 16.720 46.490 17.020 ;
        RECT 47.510 16.720 47.810 17.020 ;
        RECT 46.190 16.520 46.320 16.720 ;
        RECT 47.680 16.520 47.810 16.720 ;
        RECT 48.190 16.720 48.490 17.020 ;
        RECT 49.510 16.720 49.810 17.020 ;
        RECT 48.190 16.520 48.320 16.720 ;
        RECT 49.680 16.520 49.810 16.720 ;
        RECT 50.190 16.720 50.490 17.020 ;
        RECT 51.510 16.720 51.810 17.020 ;
        RECT 50.190 16.520 50.320 16.720 ;
        RECT 51.680 16.520 51.810 16.720 ;
        RECT 52.190 16.720 52.490 17.020 ;
        RECT 53.510 16.720 53.810 17.020 ;
        RECT 52.190 16.520 52.320 16.720 ;
        RECT 53.680 16.520 53.810 16.720 ;
        RECT 54.190 16.720 54.490 17.020 ;
        RECT 55.510 16.720 55.810 17.020 ;
        RECT 54.190 16.520 54.320 16.720 ;
        RECT 55.680 16.520 55.810 16.720 ;
        RECT 56.190 16.720 56.490 17.020 ;
        RECT 57.510 16.720 57.810 17.020 ;
        RECT 56.190 16.520 56.320 16.720 ;
        RECT 57.680 16.520 57.810 16.720 ;
        RECT 58.190 16.720 58.490 17.020 ;
        RECT 59.510 16.720 59.810 17.020 ;
        RECT 58.190 16.520 58.320 16.720 ;
        RECT 59.680 16.520 59.810 16.720 ;
        RECT 60.190 16.720 60.490 17.020 ;
        RECT 61.510 16.720 61.810 17.020 ;
        RECT 60.190 16.520 60.320 16.720 ;
        RECT 61.680 16.520 61.810 16.720 ;
        RECT 62.190 16.720 62.490 17.020 ;
        RECT 63.510 16.720 63.810 17.020 ;
        RECT 62.190 16.520 62.320 16.720 ;
        RECT 63.680 16.520 63.810 16.720 ;
        RECT 64.190 16.720 64.490 17.020 ;
        RECT 65.510 16.720 65.810 17.020 ;
        RECT 64.190 16.520 64.320 16.720 ;
        RECT 65.680 16.520 65.810 16.720 ;
        RECT 66.190 16.720 66.490 17.020 ;
        RECT 67.510 16.720 67.810 17.020 ;
        RECT 66.190 16.520 66.320 16.720 ;
        RECT 67.680 16.520 67.810 16.720 ;
        RECT 68.190 16.720 68.490 17.020 ;
        RECT 69.510 16.720 69.810 17.020 ;
        RECT 68.190 16.520 68.320 16.720 ;
        RECT 69.680 16.520 69.810 16.720 ;
        RECT 70.190 16.720 70.490 17.020 ;
        RECT 71.510 16.720 71.810 17.020 ;
        RECT 70.190 16.520 70.320 16.720 ;
        RECT 71.680 16.520 71.810 16.720 ;
        RECT 72.190 16.720 72.490 17.020 ;
        RECT 73.510 16.720 73.810 17.020 ;
        RECT 72.190 16.520 72.320 16.720 ;
        RECT 73.680 16.520 73.810 16.720 ;
        RECT 74.190 16.720 74.490 17.020 ;
        RECT 75.510 16.720 75.810 17.020 ;
        RECT 74.190 16.520 74.320 16.720 ;
        RECT 75.680 16.520 75.810 16.720 ;
        RECT 76.190 16.720 76.490 17.020 ;
        RECT 77.510 16.720 77.810 17.020 ;
        RECT 76.190 16.520 76.320 16.720 ;
        RECT 77.680 16.520 77.810 16.720 ;
        RECT 78.190 16.720 78.490 17.020 ;
        RECT 79.510 16.720 79.810 17.020 ;
        RECT 78.190 16.520 78.320 16.720 ;
        RECT 79.680 16.520 79.810 16.720 ;
        RECT 80.190 16.720 80.490 17.020 ;
        RECT 81.510 16.720 81.810 17.020 ;
        RECT 80.190 16.520 80.320 16.720 ;
        RECT 81.680 16.520 81.810 16.720 ;
        RECT 82.190 16.720 82.490 17.020 ;
        RECT 83.510 16.720 83.810 17.020 ;
        RECT 82.190 16.520 82.320 16.720 ;
        RECT 83.680 16.520 83.810 16.720 ;
        RECT 84.190 16.720 84.490 17.020 ;
        RECT 85.510 16.720 85.810 17.020 ;
        RECT 84.190 16.520 84.320 16.720 ;
        RECT 85.680 16.520 85.810 16.720 ;
        RECT 86.190 16.720 86.490 17.020 ;
        RECT 87.510 16.720 87.810 17.020 ;
        RECT 86.190 16.520 86.320 16.720 ;
        RECT 87.680 16.520 87.810 16.720 ;
        RECT 88.190 16.720 88.490 17.020 ;
        RECT 89.510 16.720 89.810 17.020 ;
        RECT 88.190 16.520 88.320 16.720 ;
        RECT 89.680 16.520 89.810 16.720 ;
        RECT 90.190 16.720 90.490 17.020 ;
        RECT 91.510 16.720 91.810 17.020 ;
        RECT 90.190 16.520 90.320 16.720 ;
        RECT 91.680 16.520 91.810 16.720 ;
        RECT 92.190 16.720 92.490 17.020 ;
        RECT 93.510 16.720 93.810 17.020 ;
        RECT 92.190 16.520 92.320 16.720 ;
        RECT 93.680 16.520 93.810 16.720 ;
        RECT 94.190 16.720 94.490 17.020 ;
        RECT 95.510 16.720 95.810 17.020 ;
        RECT 94.190 16.520 94.320 16.720 ;
        RECT 95.680 16.520 95.810 16.720 ;
        RECT 96.190 16.720 96.490 17.020 ;
        RECT 97.510 16.720 97.810 17.020 ;
        RECT 96.190 16.520 96.320 16.720 ;
        RECT 97.680 16.520 97.810 16.720 ;
        RECT 98.190 16.720 98.490 17.020 ;
        RECT 99.510 16.720 99.810 17.020 ;
        RECT 98.190 16.520 98.320 16.720 ;
        RECT 99.680 16.520 99.810 16.720 ;
        RECT 100.190 16.720 100.490 17.020 ;
        RECT 101.510 16.720 101.810 17.020 ;
        RECT 100.190 16.520 100.320 16.720 ;
        RECT 101.680 16.520 101.810 16.720 ;
        RECT 102.190 16.720 102.490 17.020 ;
        RECT 103.510 16.720 103.810 17.020 ;
        RECT 102.190 16.520 102.320 16.720 ;
        RECT 103.680 16.520 103.810 16.720 ;
        RECT 104.190 16.720 104.490 17.020 ;
        RECT 105.510 16.720 105.810 17.020 ;
        RECT 104.190 16.520 104.320 16.720 ;
        RECT 105.680 16.520 105.810 16.720 ;
        RECT 106.190 16.720 106.490 17.020 ;
        RECT 107.510 16.720 107.810 17.020 ;
        RECT 106.190 16.520 106.320 16.720 ;
        RECT 107.680 16.520 107.810 16.720 ;
        RECT 108.190 16.720 108.490 17.020 ;
        RECT 109.510 16.720 109.810 17.020 ;
        RECT 108.190 16.520 108.320 16.720 ;
        RECT 109.680 16.520 109.810 16.720 ;
        RECT 110.190 16.720 110.490 17.020 ;
        RECT 111.510 16.720 111.810 17.020 ;
        RECT 110.190 16.520 110.320 16.720 ;
        RECT 111.680 16.520 111.810 16.720 ;
        RECT 112.190 16.720 112.490 17.020 ;
        RECT 113.510 16.720 113.810 17.020 ;
        RECT 112.190 16.520 112.320 16.720 ;
        RECT 113.680 16.520 113.810 16.720 ;
        RECT 114.190 16.720 114.490 17.020 ;
        RECT 115.510 16.720 115.810 17.020 ;
        RECT 114.190 16.520 114.320 16.720 ;
        RECT 115.680 16.520 115.810 16.720 ;
        RECT 116.190 16.720 116.490 17.020 ;
        RECT 117.510 16.720 117.810 17.020 ;
        RECT 116.190 16.520 116.320 16.720 ;
        RECT 117.680 16.520 117.810 16.720 ;
        RECT 118.190 16.720 118.490 17.020 ;
        RECT 119.510 16.720 119.810 17.020 ;
        RECT 118.190 16.520 118.320 16.720 ;
        RECT 119.680 16.520 119.810 16.720 ;
        RECT 120.190 16.720 120.490 17.020 ;
        RECT 121.510 16.720 121.810 17.020 ;
        RECT 120.190 16.520 120.320 16.720 ;
        RECT 121.680 16.520 121.810 16.720 ;
        RECT 122.190 16.720 122.490 17.020 ;
        RECT 123.510 16.720 123.810 17.020 ;
        RECT 122.190 16.520 122.320 16.720 ;
        RECT 123.680 16.520 123.810 16.720 ;
        RECT 124.190 16.720 124.490 17.020 ;
        RECT 125.510 16.720 125.810 17.020 ;
        RECT 124.190 16.520 124.320 16.720 ;
        RECT 125.680 16.520 125.810 16.720 ;
        RECT 126.190 16.720 126.490 17.020 ;
        RECT 127.510 16.720 127.810 17.020 ;
        RECT 126.190 16.520 126.320 16.720 ;
        RECT 127.680 16.520 127.810 16.720 ;
        RECT 128.190 16.720 128.490 17.020 ;
        RECT 129.510 16.720 129.810 17.020 ;
        RECT 128.190 16.520 128.320 16.720 ;
        RECT 129.680 16.520 129.810 16.720 ;
        RECT 130.190 16.720 130.490 17.020 ;
        RECT 130.190 16.520 130.320 16.720 ;
        RECT -0.320 16.040 -0.190 16.220 ;
        RECT 0.190 16.040 0.320 16.220 ;
        RECT 1.680 16.040 1.810 16.220 ;
        RECT 2.190 16.040 2.320 16.220 ;
        RECT 3.680 16.040 3.810 16.220 ;
        RECT 4.190 16.040 4.320 16.220 ;
        RECT 5.680 16.040 5.810 16.220 ;
        RECT 6.190 16.040 6.320 16.220 ;
        RECT 7.680 16.040 7.810 16.220 ;
        RECT 8.190 16.040 8.320 16.220 ;
        RECT 9.680 16.040 9.810 16.220 ;
        RECT 10.190 16.040 10.320 16.220 ;
        RECT 11.680 16.040 11.810 16.220 ;
        RECT 12.190 16.040 12.320 16.220 ;
        RECT 13.680 16.040 13.810 16.220 ;
        RECT 14.190 16.040 14.320 16.220 ;
        RECT 15.680 16.040 15.810 16.220 ;
        RECT 16.190 16.040 16.320 16.220 ;
        RECT 17.680 16.040 17.810 16.220 ;
        RECT 18.190 16.040 18.320 16.220 ;
        RECT 19.680 16.040 19.810 16.220 ;
        RECT 20.190 16.040 20.320 16.220 ;
        RECT 21.680 16.040 21.810 16.220 ;
        RECT 22.190 16.040 22.320 16.220 ;
        RECT 23.680 16.040 23.810 16.220 ;
        RECT 24.190 16.040 24.320 16.220 ;
        RECT 25.680 16.040 25.810 16.220 ;
        RECT 26.190 16.040 26.320 16.220 ;
        RECT 27.680 16.040 27.810 16.220 ;
        RECT 28.190 16.040 28.320 16.220 ;
        RECT 29.680 16.040 29.810 16.220 ;
        RECT 30.190 16.040 30.320 16.220 ;
        RECT 31.680 16.040 31.810 16.220 ;
        RECT 32.190 16.040 32.320 16.220 ;
        RECT 33.680 16.040 33.810 16.220 ;
        RECT 34.190 16.040 34.320 16.220 ;
        RECT 35.680 16.040 35.810 16.220 ;
        RECT 36.190 16.040 36.320 16.220 ;
        RECT 37.680 16.040 37.810 16.220 ;
        RECT 38.190 16.040 38.320 16.220 ;
        RECT 39.680 16.040 39.810 16.220 ;
        RECT 40.190 16.040 40.320 16.220 ;
        RECT 41.680 16.040 41.810 16.220 ;
        RECT 42.190 16.040 42.320 16.220 ;
        RECT 43.680 16.040 43.810 16.220 ;
        RECT 44.190 16.040 44.320 16.220 ;
        RECT 45.680 16.040 45.810 16.220 ;
        RECT 46.190 16.040 46.320 16.220 ;
        RECT 47.680 16.040 47.810 16.220 ;
        RECT 48.190 16.040 48.320 16.220 ;
        RECT 49.680 16.040 49.810 16.220 ;
        RECT 50.190 16.040 50.320 16.220 ;
        RECT 51.680 16.040 51.810 16.220 ;
        RECT 52.190 16.040 52.320 16.220 ;
        RECT 53.680 16.040 53.810 16.220 ;
        RECT 54.190 16.040 54.320 16.220 ;
        RECT 55.680 16.040 55.810 16.220 ;
        RECT 56.190 16.040 56.320 16.220 ;
        RECT 57.680 16.040 57.810 16.220 ;
        RECT 58.190 16.040 58.320 16.220 ;
        RECT 59.680 16.040 59.810 16.220 ;
        RECT 60.190 16.040 60.320 16.220 ;
        RECT 61.680 16.040 61.810 16.220 ;
        RECT 62.190 16.040 62.320 16.220 ;
        RECT 63.680 16.040 63.810 16.220 ;
        RECT 64.190 16.040 64.320 16.220 ;
        RECT 65.680 16.040 65.810 16.220 ;
        RECT 66.190 16.040 66.320 16.220 ;
        RECT 67.680 16.040 67.810 16.220 ;
        RECT 68.190 16.040 68.320 16.220 ;
        RECT 69.680 16.040 69.810 16.220 ;
        RECT 70.190 16.040 70.320 16.220 ;
        RECT 71.680 16.040 71.810 16.220 ;
        RECT 72.190 16.040 72.320 16.220 ;
        RECT 73.680 16.040 73.810 16.220 ;
        RECT 74.190 16.040 74.320 16.220 ;
        RECT 75.680 16.040 75.810 16.220 ;
        RECT 76.190 16.040 76.320 16.220 ;
        RECT 77.680 16.040 77.810 16.220 ;
        RECT 78.190 16.040 78.320 16.220 ;
        RECT 79.680 16.040 79.810 16.220 ;
        RECT 80.190 16.040 80.320 16.220 ;
        RECT 81.680 16.040 81.810 16.220 ;
        RECT 82.190 16.040 82.320 16.220 ;
        RECT 83.680 16.040 83.810 16.220 ;
        RECT 84.190 16.040 84.320 16.220 ;
        RECT 85.680 16.040 85.810 16.220 ;
        RECT 86.190 16.040 86.320 16.220 ;
        RECT 87.680 16.040 87.810 16.220 ;
        RECT 88.190 16.040 88.320 16.220 ;
        RECT 89.680 16.040 89.810 16.220 ;
        RECT 90.190 16.040 90.320 16.220 ;
        RECT 91.680 16.040 91.810 16.220 ;
        RECT 92.190 16.040 92.320 16.220 ;
        RECT 93.680 16.040 93.810 16.220 ;
        RECT 94.190 16.040 94.320 16.220 ;
        RECT 95.680 16.040 95.810 16.220 ;
        RECT 96.190 16.040 96.320 16.220 ;
        RECT 97.680 16.040 97.810 16.220 ;
        RECT 98.190 16.040 98.320 16.220 ;
        RECT 99.680 16.040 99.810 16.220 ;
        RECT 100.190 16.040 100.320 16.220 ;
        RECT 101.680 16.040 101.810 16.220 ;
        RECT 102.190 16.040 102.320 16.220 ;
        RECT 103.680 16.040 103.810 16.220 ;
        RECT 104.190 16.040 104.320 16.220 ;
        RECT 105.680 16.040 105.810 16.220 ;
        RECT 106.190 16.040 106.320 16.220 ;
        RECT 107.680 16.040 107.810 16.220 ;
        RECT 108.190 16.040 108.320 16.220 ;
        RECT 109.680 16.040 109.810 16.220 ;
        RECT 110.190 16.040 110.320 16.220 ;
        RECT 111.680 16.040 111.810 16.220 ;
        RECT 112.190 16.040 112.320 16.220 ;
        RECT 113.680 16.040 113.810 16.220 ;
        RECT 114.190 16.040 114.320 16.220 ;
        RECT 115.680 16.040 115.810 16.220 ;
        RECT 116.190 16.040 116.320 16.220 ;
        RECT 117.680 16.040 117.810 16.220 ;
        RECT 118.190 16.040 118.320 16.220 ;
        RECT 119.680 16.040 119.810 16.220 ;
        RECT 120.190 16.040 120.320 16.220 ;
        RECT 121.680 16.040 121.810 16.220 ;
        RECT 122.190 16.040 122.320 16.220 ;
        RECT 123.680 16.040 123.810 16.220 ;
        RECT 124.190 16.040 124.320 16.220 ;
        RECT 125.680 16.040 125.810 16.220 ;
        RECT 126.190 16.040 126.320 16.220 ;
        RECT 127.680 16.040 127.810 16.220 ;
        RECT 128.190 16.040 128.320 16.220 ;
        RECT 129.680 16.040 129.810 16.220 ;
        RECT 130.190 16.040 130.320 16.220 ;
        RECT -1.900 14.690 -1.410 14.990 ;
        RECT -1.560 14.610 -1.410 14.690 ;
        RECT -1.000 10.040 -0.820 15.040 ;
        RECT 0.630 10.040 1.180 15.040 ;
        RECT 2.630 10.040 3.180 15.040 ;
        RECT 4.630 10.040 5.180 15.040 ;
        RECT 6.630 10.040 7.180 15.040 ;
        RECT 8.630 10.040 9.180 15.040 ;
        RECT 10.630 10.040 11.180 15.040 ;
        RECT 12.630 10.040 13.180 15.040 ;
        RECT 14.630 10.040 15.180 15.040 ;
        RECT 16.630 10.040 17.180 15.040 ;
        RECT 18.630 10.040 19.180 15.040 ;
        RECT 20.630 10.040 21.180 15.040 ;
        RECT 22.630 10.040 23.180 15.040 ;
        RECT 24.630 10.040 25.180 15.040 ;
        RECT 26.630 10.040 27.180 15.040 ;
        RECT 28.630 10.040 29.180 15.040 ;
        RECT 30.630 10.040 31.180 15.040 ;
        RECT 32.630 10.040 33.180 15.040 ;
        RECT 34.630 10.040 35.180 15.040 ;
        RECT 36.630 10.040 37.180 15.040 ;
        RECT 38.630 10.040 39.180 15.040 ;
        RECT 40.630 10.040 41.180 15.040 ;
        RECT 42.630 10.040 43.180 15.040 ;
        RECT 44.630 10.040 45.180 15.040 ;
        RECT 46.630 10.040 47.180 15.040 ;
        RECT 48.630 10.040 49.180 15.040 ;
        RECT 50.630 10.040 51.180 15.040 ;
        RECT 52.630 10.040 53.180 15.040 ;
        RECT 54.630 10.040 55.180 15.040 ;
        RECT 56.630 10.040 57.180 15.040 ;
        RECT 58.630 10.040 59.180 15.040 ;
        RECT 60.630 10.040 61.180 15.040 ;
        RECT 62.630 10.040 63.180 15.040 ;
        RECT 64.630 10.040 65.180 15.040 ;
        RECT 66.630 10.040 67.180 15.040 ;
        RECT 68.630 10.040 69.180 15.040 ;
        RECT 70.630 10.040 71.180 15.040 ;
        RECT 72.630 10.040 73.180 15.040 ;
        RECT 74.630 10.040 75.180 15.040 ;
        RECT 76.630 10.040 77.180 15.040 ;
        RECT 78.630 10.040 79.180 15.040 ;
        RECT 80.630 10.040 81.180 15.040 ;
        RECT 82.630 10.040 83.180 15.040 ;
        RECT 84.630 10.040 85.180 15.040 ;
        RECT 86.630 10.040 87.180 15.040 ;
        RECT 88.630 10.040 89.180 15.040 ;
        RECT 90.630 10.040 91.180 15.040 ;
        RECT 92.630 10.040 93.180 15.040 ;
        RECT 94.630 10.040 95.180 15.040 ;
        RECT 96.630 10.040 97.180 15.040 ;
        RECT 98.630 10.040 99.180 15.040 ;
        RECT 100.630 10.040 101.180 15.040 ;
        RECT 102.630 10.040 103.180 15.040 ;
        RECT 104.630 10.040 105.180 15.040 ;
        RECT 106.630 10.040 107.180 15.040 ;
        RECT 108.630 10.040 109.180 15.040 ;
        RECT 110.630 10.040 111.180 15.040 ;
        RECT 112.630 10.040 113.180 15.040 ;
        RECT 114.630 10.040 115.180 15.040 ;
        RECT 116.630 10.040 117.180 15.040 ;
        RECT 118.630 10.040 119.180 15.040 ;
        RECT 120.630 10.040 121.180 15.040 ;
        RECT 122.630 10.040 123.180 15.040 ;
        RECT 124.630 10.040 125.180 15.040 ;
        RECT 126.630 10.040 127.180 15.040 ;
        RECT 128.630 10.040 129.180 15.040 ;
        RECT 130.630 10.040 131.000 15.040 ;
        RECT 131.410 14.690 131.900 14.990 ;
        RECT 131.410 14.610 131.560 14.690 ;
        RECT -1.000 9.140 -0.820 9.740 ;
        RECT 0.380 9.140 0.820 9.740 ;
        RECT 1.000 9.140 1.180 9.740 ;
        RECT 2.380 9.140 2.820 9.740 ;
        RECT 3.000 9.140 3.180 9.740 ;
        RECT 4.380 9.140 4.820 9.740 ;
        RECT 5.000 9.140 5.180 9.740 ;
        RECT 6.380 9.140 6.820 9.740 ;
        RECT 7.000 9.140 7.180 9.740 ;
        RECT 8.380 9.140 8.820 9.740 ;
        RECT 9.000 9.140 9.180 9.740 ;
        RECT 10.380 9.140 10.820 9.740 ;
        RECT 11.000 9.140 11.180 9.740 ;
        RECT 12.380 9.140 12.820 9.740 ;
        RECT 13.000 9.140 13.180 9.740 ;
        RECT 14.380 9.140 14.820 9.740 ;
        RECT 15.000 9.140 15.180 9.740 ;
        RECT 16.380 9.140 16.820 9.740 ;
        RECT 17.000 9.140 17.180 9.740 ;
        RECT 18.380 9.140 18.820 9.740 ;
        RECT 19.000 9.140 19.180 9.740 ;
        RECT 20.380 9.140 20.820 9.740 ;
        RECT 21.000 9.140 21.180 9.740 ;
        RECT 22.380 9.140 22.820 9.740 ;
        RECT 23.000 9.140 23.180 9.740 ;
        RECT 24.380 9.140 24.820 9.740 ;
        RECT 25.000 9.140 25.180 9.740 ;
        RECT 26.380 9.140 26.820 9.740 ;
        RECT 27.000 9.140 27.180 9.740 ;
        RECT 28.380 9.140 28.820 9.740 ;
        RECT 29.000 9.140 29.180 9.740 ;
        RECT 30.380 9.140 30.820 9.740 ;
        RECT 31.000 9.140 31.180 9.740 ;
        RECT 32.380 9.140 32.820 9.740 ;
        RECT 33.000 9.140 33.180 9.740 ;
        RECT 34.380 9.140 34.820 9.740 ;
        RECT 35.000 9.140 35.180 9.740 ;
        RECT 36.380 9.140 36.820 9.740 ;
        RECT 37.000 9.140 37.180 9.740 ;
        RECT 38.380 9.140 38.820 9.740 ;
        RECT 39.000 9.140 39.180 9.740 ;
        RECT 40.380 9.140 40.820 9.740 ;
        RECT 41.000 9.140 41.180 9.740 ;
        RECT 42.380 9.140 42.820 9.740 ;
        RECT 43.000 9.140 43.180 9.740 ;
        RECT 44.380 9.140 44.820 9.740 ;
        RECT 45.000 9.140 45.180 9.740 ;
        RECT 46.380 9.140 46.820 9.740 ;
        RECT 47.000 9.140 47.180 9.740 ;
        RECT 48.380 9.140 48.820 9.740 ;
        RECT 49.000 9.140 49.180 9.740 ;
        RECT 50.380 9.140 50.820 9.740 ;
        RECT 51.000 9.140 51.180 9.740 ;
        RECT 52.380 9.140 52.820 9.740 ;
        RECT 53.000 9.140 53.180 9.740 ;
        RECT 54.380 9.140 54.820 9.740 ;
        RECT 55.000 9.140 55.180 9.740 ;
        RECT 56.380 9.140 56.820 9.740 ;
        RECT 57.000 9.140 57.180 9.740 ;
        RECT 58.380 9.140 58.820 9.740 ;
        RECT 59.000 9.140 59.180 9.740 ;
        RECT 60.380 9.140 60.820 9.740 ;
        RECT 61.000 9.140 61.180 9.740 ;
        RECT 62.380 9.140 62.820 9.740 ;
        RECT 63.000 9.140 63.180 9.740 ;
        RECT 64.380 9.140 64.820 9.740 ;
        RECT 65.000 9.140 65.180 9.740 ;
        RECT 66.380 9.140 66.820 9.740 ;
        RECT 67.000 9.140 67.180 9.740 ;
        RECT 68.380 9.140 68.820 9.740 ;
        RECT 69.000 9.140 69.180 9.740 ;
        RECT 70.380 9.140 70.820 9.740 ;
        RECT 71.000 9.140 71.180 9.740 ;
        RECT 72.380 9.140 72.820 9.740 ;
        RECT 73.000 9.140 73.180 9.740 ;
        RECT 74.380 9.140 74.820 9.740 ;
        RECT 75.000 9.140 75.180 9.740 ;
        RECT 76.380 9.140 76.820 9.740 ;
        RECT 77.000 9.140 77.180 9.740 ;
        RECT 78.380 9.140 78.820 9.740 ;
        RECT 79.000 9.140 79.180 9.740 ;
        RECT 80.380 9.140 80.820 9.740 ;
        RECT 81.000 9.140 81.180 9.740 ;
        RECT 82.380 9.140 82.820 9.740 ;
        RECT 83.000 9.140 83.180 9.740 ;
        RECT 84.380 9.140 84.820 9.740 ;
        RECT 85.000 9.140 85.180 9.740 ;
        RECT 86.380 9.140 86.820 9.740 ;
        RECT 87.000 9.140 87.180 9.740 ;
        RECT 88.380 9.140 88.820 9.740 ;
        RECT 89.000 9.140 89.180 9.740 ;
        RECT 90.380 9.140 90.820 9.740 ;
        RECT 91.000 9.140 91.180 9.740 ;
        RECT 92.380 9.140 92.820 9.740 ;
        RECT 93.000 9.140 93.180 9.740 ;
        RECT 94.380 9.140 94.820 9.740 ;
        RECT 95.000 9.140 95.180 9.740 ;
        RECT 96.380 9.140 96.820 9.740 ;
        RECT 97.000 9.140 97.180 9.740 ;
        RECT 98.380 9.140 98.820 9.740 ;
        RECT 99.000 9.140 99.180 9.740 ;
        RECT 100.380 9.140 100.820 9.740 ;
        RECT 101.000 9.140 101.180 9.740 ;
        RECT 102.380 9.140 102.820 9.740 ;
        RECT 103.000 9.140 103.180 9.740 ;
        RECT 104.380 9.140 104.820 9.740 ;
        RECT 105.000 9.140 105.180 9.740 ;
        RECT 106.380 9.140 106.820 9.740 ;
        RECT 107.000 9.140 107.180 9.740 ;
        RECT 108.380 9.140 108.820 9.740 ;
        RECT 109.000 9.140 109.180 9.740 ;
        RECT 110.380 9.140 110.820 9.740 ;
        RECT 111.000 9.140 111.180 9.740 ;
        RECT 112.380 9.140 112.820 9.740 ;
        RECT 113.000 9.140 113.180 9.740 ;
        RECT 114.380 9.140 114.820 9.740 ;
        RECT 115.000 9.140 115.180 9.740 ;
        RECT 116.380 9.140 116.820 9.740 ;
        RECT 117.000 9.140 117.180 9.740 ;
        RECT 118.380 9.140 118.820 9.740 ;
        RECT 119.000 9.140 119.180 9.740 ;
        RECT 120.380 9.140 120.820 9.740 ;
        RECT 121.000 9.140 121.180 9.740 ;
        RECT 122.380 9.140 122.820 9.740 ;
        RECT 123.000 9.140 123.180 9.740 ;
        RECT 124.380 9.140 124.820 9.740 ;
        RECT 125.000 9.140 125.180 9.740 ;
        RECT 126.380 9.140 126.820 9.740 ;
        RECT 127.000 9.140 127.180 9.740 ;
        RECT 128.380 9.140 128.820 9.740 ;
        RECT 129.000 9.140 129.180 9.740 ;
        RECT 130.380 9.140 130.820 9.740 ;
        RECT -1.560 8.580 -1.410 8.760 ;
        RECT 131.410 8.580 131.560 8.760 ;
        RECT -1.560 7.610 -1.410 7.790 ;
        RECT 131.410 7.610 131.560 7.790 ;
        RECT -0.820 6.630 -0.380 7.230 ;
        RECT 0.820 6.630 1.000 7.230 ;
        RECT 1.180 6.630 1.620 7.230 ;
        RECT 2.820 6.630 3.000 7.230 ;
        RECT 3.180 6.630 3.620 7.230 ;
        RECT 4.820 6.630 5.000 7.230 ;
        RECT 5.180 6.630 5.620 7.230 ;
        RECT 6.820 6.630 7.000 7.230 ;
        RECT 7.180 6.630 7.620 7.230 ;
        RECT 8.820 6.630 9.000 7.230 ;
        RECT 9.180 6.630 9.620 7.230 ;
        RECT 10.820 6.630 11.000 7.230 ;
        RECT 11.180 6.630 11.620 7.230 ;
        RECT 12.820 6.630 13.000 7.230 ;
        RECT 13.180 6.630 13.620 7.230 ;
        RECT 14.820 6.630 15.000 7.230 ;
        RECT 15.180 6.630 15.620 7.230 ;
        RECT 16.820 6.630 17.000 7.230 ;
        RECT 17.180 6.630 17.620 7.230 ;
        RECT 18.820 6.630 19.000 7.230 ;
        RECT 19.180 6.630 19.620 7.230 ;
        RECT 20.820 6.630 21.000 7.230 ;
        RECT 21.180 6.630 21.620 7.230 ;
        RECT 22.820 6.630 23.000 7.230 ;
        RECT 23.180 6.630 23.620 7.230 ;
        RECT 24.820 6.630 25.000 7.230 ;
        RECT 25.180 6.630 25.620 7.230 ;
        RECT 26.820 6.630 27.000 7.230 ;
        RECT 27.180 6.630 27.620 7.230 ;
        RECT 28.820 6.630 29.000 7.230 ;
        RECT 29.180 6.630 29.620 7.230 ;
        RECT 30.820 6.630 31.000 7.230 ;
        RECT 31.180 6.630 31.620 7.230 ;
        RECT 32.820 6.630 33.000 7.230 ;
        RECT 33.180 6.630 33.620 7.230 ;
        RECT 34.820 6.630 35.000 7.230 ;
        RECT 35.180 6.630 35.620 7.230 ;
        RECT 36.820 6.630 37.000 7.230 ;
        RECT 37.180 6.630 37.620 7.230 ;
        RECT 38.820 6.630 39.000 7.230 ;
        RECT 39.180 6.630 39.620 7.230 ;
        RECT 40.820 6.630 41.000 7.230 ;
        RECT 41.180 6.630 41.620 7.230 ;
        RECT 42.820 6.630 43.000 7.230 ;
        RECT 43.180 6.630 43.620 7.230 ;
        RECT 44.820 6.630 45.000 7.230 ;
        RECT 45.180 6.630 45.620 7.230 ;
        RECT 46.820 6.630 47.000 7.230 ;
        RECT 47.180 6.630 47.620 7.230 ;
        RECT 48.820 6.630 49.000 7.230 ;
        RECT 49.180 6.630 49.620 7.230 ;
        RECT 50.820 6.630 51.000 7.230 ;
        RECT 51.180 6.630 51.620 7.230 ;
        RECT 52.820 6.630 53.000 7.230 ;
        RECT 53.180 6.630 53.620 7.230 ;
        RECT 54.820 6.630 55.000 7.230 ;
        RECT 55.180 6.630 55.620 7.230 ;
        RECT 56.820 6.630 57.000 7.230 ;
        RECT 57.180 6.630 57.620 7.230 ;
        RECT 58.820 6.630 59.000 7.230 ;
        RECT 59.180 6.630 59.620 7.230 ;
        RECT 60.820 6.630 61.000 7.230 ;
        RECT 61.180 6.630 61.620 7.230 ;
        RECT 62.820 6.630 63.000 7.230 ;
        RECT 63.180 6.630 63.620 7.230 ;
        RECT 64.820 6.630 65.000 7.230 ;
        RECT 65.180 6.630 65.620 7.230 ;
        RECT 66.820 6.630 67.000 7.230 ;
        RECT 67.180 6.630 67.620 7.230 ;
        RECT 68.820 6.630 69.000 7.230 ;
        RECT 69.180 6.630 69.620 7.230 ;
        RECT 70.820 6.630 71.000 7.230 ;
        RECT 71.180 6.630 71.620 7.230 ;
        RECT 72.820 6.630 73.000 7.230 ;
        RECT 73.180 6.630 73.620 7.230 ;
        RECT 74.820 6.630 75.000 7.230 ;
        RECT 75.180 6.630 75.620 7.230 ;
        RECT 76.820 6.630 77.000 7.230 ;
        RECT 77.180 6.630 77.620 7.230 ;
        RECT 78.820 6.630 79.000 7.230 ;
        RECT 79.180 6.630 79.620 7.230 ;
        RECT 80.820 6.630 81.000 7.230 ;
        RECT 81.180 6.630 81.620 7.230 ;
        RECT 82.820 6.630 83.000 7.230 ;
        RECT 83.180 6.630 83.620 7.230 ;
        RECT 84.820 6.630 85.000 7.230 ;
        RECT 85.180 6.630 85.620 7.230 ;
        RECT 86.820 6.630 87.000 7.230 ;
        RECT 87.180 6.630 87.620 7.230 ;
        RECT 88.820 6.630 89.000 7.230 ;
        RECT 89.180 6.630 89.620 7.230 ;
        RECT 90.820 6.630 91.000 7.230 ;
        RECT 91.180 6.630 91.620 7.230 ;
        RECT 92.820 6.630 93.000 7.230 ;
        RECT 93.180 6.630 93.620 7.230 ;
        RECT 94.820 6.630 95.000 7.230 ;
        RECT 95.180 6.630 95.620 7.230 ;
        RECT 96.820 6.630 97.000 7.230 ;
        RECT 97.180 6.630 97.620 7.230 ;
        RECT 98.820 6.630 99.000 7.230 ;
        RECT 99.180 6.630 99.620 7.230 ;
        RECT 100.820 6.630 101.000 7.230 ;
        RECT 101.180 6.630 101.620 7.230 ;
        RECT 102.820 6.630 103.000 7.230 ;
        RECT 103.180 6.630 103.620 7.230 ;
        RECT 104.820 6.630 105.000 7.230 ;
        RECT 105.180 6.630 105.620 7.230 ;
        RECT 106.820 6.630 107.000 7.230 ;
        RECT 107.180 6.630 107.620 7.230 ;
        RECT 108.820 6.630 109.000 7.230 ;
        RECT 109.180 6.630 109.620 7.230 ;
        RECT 110.820 6.630 111.000 7.230 ;
        RECT 111.180 6.630 111.620 7.230 ;
        RECT 112.820 6.630 113.000 7.230 ;
        RECT 113.180 6.630 113.620 7.230 ;
        RECT 114.820 6.630 115.000 7.230 ;
        RECT 115.180 6.630 115.620 7.230 ;
        RECT 116.820 6.630 117.000 7.230 ;
        RECT 117.180 6.630 117.620 7.230 ;
        RECT 118.820 6.630 119.000 7.230 ;
        RECT 119.180 6.630 119.620 7.230 ;
        RECT 120.820 6.630 121.000 7.230 ;
        RECT 121.180 6.630 121.620 7.230 ;
        RECT 122.820 6.630 123.000 7.230 ;
        RECT 123.180 6.630 123.620 7.230 ;
        RECT 124.820 6.630 125.000 7.230 ;
        RECT 125.180 6.630 125.620 7.230 ;
        RECT 126.820 6.630 127.000 7.230 ;
        RECT 127.180 6.630 127.620 7.230 ;
        RECT 128.820 6.630 129.000 7.230 ;
        RECT 129.180 6.630 129.620 7.230 ;
        RECT 130.820 6.630 131.000 7.230 ;
        RECT -1.560 1.680 -1.410 1.760 ;
        RECT -1.900 1.380 -1.410 1.680 ;
        RECT -1.000 1.330 -0.630 6.330 ;
        RECT 0.820 1.330 1.370 6.330 ;
        RECT 2.820 1.330 3.370 6.330 ;
        RECT 4.820 1.330 5.370 6.330 ;
        RECT 6.820 1.330 7.370 6.330 ;
        RECT 8.820 1.330 9.370 6.330 ;
        RECT 10.820 1.330 11.370 6.330 ;
        RECT 12.820 1.330 13.370 6.330 ;
        RECT 14.820 1.330 15.370 6.330 ;
        RECT 16.820 1.330 17.370 6.330 ;
        RECT 18.820 1.330 19.370 6.330 ;
        RECT 20.820 1.330 21.370 6.330 ;
        RECT 22.820 1.330 23.370 6.330 ;
        RECT 24.820 1.330 25.370 6.330 ;
        RECT 26.820 1.330 27.370 6.330 ;
        RECT 28.820 1.330 29.370 6.330 ;
        RECT 30.820 1.330 31.370 6.330 ;
        RECT 32.820 1.330 33.370 6.330 ;
        RECT 34.820 1.330 35.370 6.330 ;
        RECT 36.820 1.330 37.370 6.330 ;
        RECT 38.820 1.330 39.370 6.330 ;
        RECT 40.820 1.330 41.370 6.330 ;
        RECT 42.820 1.330 43.370 6.330 ;
        RECT 44.820 1.330 45.370 6.330 ;
        RECT 46.820 1.330 47.370 6.330 ;
        RECT 48.820 1.330 49.370 6.330 ;
        RECT 50.820 1.330 51.370 6.330 ;
        RECT 52.820 1.330 53.370 6.330 ;
        RECT 54.820 1.330 55.370 6.330 ;
        RECT 56.820 1.330 57.370 6.330 ;
        RECT 58.820 1.330 59.370 6.330 ;
        RECT 60.820 1.330 61.370 6.330 ;
        RECT 62.820 1.330 63.370 6.330 ;
        RECT 64.820 1.330 65.370 6.330 ;
        RECT 66.820 1.330 67.370 6.330 ;
        RECT 68.820 1.330 69.370 6.330 ;
        RECT 70.820 1.330 71.370 6.330 ;
        RECT 72.820 1.330 73.370 6.330 ;
        RECT 74.820 1.330 75.370 6.330 ;
        RECT 76.820 1.330 77.370 6.330 ;
        RECT 78.820 1.330 79.370 6.330 ;
        RECT 80.820 1.330 81.370 6.330 ;
        RECT 82.820 1.330 83.370 6.330 ;
        RECT 84.820 1.330 85.370 6.330 ;
        RECT 86.820 1.330 87.370 6.330 ;
        RECT 88.820 1.330 89.370 6.330 ;
        RECT 90.820 1.330 91.370 6.330 ;
        RECT 92.820 1.330 93.370 6.330 ;
        RECT 94.820 1.330 95.370 6.330 ;
        RECT 96.820 1.330 97.370 6.330 ;
        RECT 98.820 1.330 99.370 6.330 ;
        RECT 100.820 1.330 101.370 6.330 ;
        RECT 102.820 1.330 103.370 6.330 ;
        RECT 104.820 1.330 105.370 6.330 ;
        RECT 106.820 1.330 107.370 6.330 ;
        RECT 108.820 1.330 109.370 6.330 ;
        RECT 110.820 1.330 111.370 6.330 ;
        RECT 112.820 1.330 113.370 6.330 ;
        RECT 114.820 1.330 115.370 6.330 ;
        RECT 116.820 1.330 117.370 6.330 ;
        RECT 118.820 1.330 119.370 6.330 ;
        RECT 120.820 1.330 121.370 6.330 ;
        RECT 122.820 1.330 123.370 6.330 ;
        RECT 124.820 1.330 125.370 6.330 ;
        RECT 126.820 1.330 127.370 6.330 ;
        RECT 128.820 1.330 129.370 6.330 ;
        RECT 130.820 1.330 131.000 6.330 ;
        RECT 131.410 1.680 131.560 1.760 ;
        RECT 131.410 1.380 131.900 1.680 ;
        RECT -0.320 0.150 -0.190 0.330 ;
        RECT 0.190 0.150 0.320 0.330 ;
        RECT 1.680 0.150 1.810 0.330 ;
        RECT 2.190 0.150 2.320 0.330 ;
        RECT 3.680 0.150 3.810 0.330 ;
        RECT 4.190 0.150 4.320 0.330 ;
        RECT 5.680 0.150 5.810 0.330 ;
        RECT 6.190 0.150 6.320 0.330 ;
        RECT 7.680 0.150 7.810 0.330 ;
        RECT 8.190 0.150 8.320 0.330 ;
        RECT 9.680 0.150 9.810 0.330 ;
        RECT 10.190 0.150 10.320 0.330 ;
        RECT 11.680 0.150 11.810 0.330 ;
        RECT 12.190 0.150 12.320 0.330 ;
        RECT 13.680 0.150 13.810 0.330 ;
        RECT 14.190 0.150 14.320 0.330 ;
        RECT 15.680 0.150 15.810 0.330 ;
        RECT 16.190 0.150 16.320 0.330 ;
        RECT 17.680 0.150 17.810 0.330 ;
        RECT 18.190 0.150 18.320 0.330 ;
        RECT 19.680 0.150 19.810 0.330 ;
        RECT 20.190 0.150 20.320 0.330 ;
        RECT 21.680 0.150 21.810 0.330 ;
        RECT 22.190 0.150 22.320 0.330 ;
        RECT 23.680 0.150 23.810 0.330 ;
        RECT 24.190 0.150 24.320 0.330 ;
        RECT 25.680 0.150 25.810 0.330 ;
        RECT 26.190 0.150 26.320 0.330 ;
        RECT 27.680 0.150 27.810 0.330 ;
        RECT 28.190 0.150 28.320 0.330 ;
        RECT 29.680 0.150 29.810 0.330 ;
        RECT 30.190 0.150 30.320 0.330 ;
        RECT 31.680 0.150 31.810 0.330 ;
        RECT 32.190 0.150 32.320 0.330 ;
        RECT 33.680 0.150 33.810 0.330 ;
        RECT 34.190 0.150 34.320 0.330 ;
        RECT 35.680 0.150 35.810 0.330 ;
        RECT 36.190 0.150 36.320 0.330 ;
        RECT 37.680 0.150 37.810 0.330 ;
        RECT 38.190 0.150 38.320 0.330 ;
        RECT 39.680 0.150 39.810 0.330 ;
        RECT 40.190 0.150 40.320 0.330 ;
        RECT 41.680 0.150 41.810 0.330 ;
        RECT 42.190 0.150 42.320 0.330 ;
        RECT 43.680 0.150 43.810 0.330 ;
        RECT 44.190 0.150 44.320 0.330 ;
        RECT 45.680 0.150 45.810 0.330 ;
        RECT 46.190 0.150 46.320 0.330 ;
        RECT 47.680 0.150 47.810 0.330 ;
        RECT 48.190 0.150 48.320 0.330 ;
        RECT 49.680 0.150 49.810 0.330 ;
        RECT 50.190 0.150 50.320 0.330 ;
        RECT 51.680 0.150 51.810 0.330 ;
        RECT 52.190 0.150 52.320 0.330 ;
        RECT 53.680 0.150 53.810 0.330 ;
        RECT 54.190 0.150 54.320 0.330 ;
        RECT 55.680 0.150 55.810 0.330 ;
        RECT 56.190 0.150 56.320 0.330 ;
        RECT 57.680 0.150 57.810 0.330 ;
        RECT 58.190 0.150 58.320 0.330 ;
        RECT 59.680 0.150 59.810 0.330 ;
        RECT 60.190 0.150 60.320 0.330 ;
        RECT 61.680 0.150 61.810 0.330 ;
        RECT 62.190 0.150 62.320 0.330 ;
        RECT 63.680 0.150 63.810 0.330 ;
        RECT 64.190 0.150 64.320 0.330 ;
        RECT 65.680 0.150 65.810 0.330 ;
        RECT 66.190 0.150 66.320 0.330 ;
        RECT 67.680 0.150 67.810 0.330 ;
        RECT 68.190 0.150 68.320 0.330 ;
        RECT 69.680 0.150 69.810 0.330 ;
        RECT 70.190 0.150 70.320 0.330 ;
        RECT 71.680 0.150 71.810 0.330 ;
        RECT 72.190 0.150 72.320 0.330 ;
        RECT 73.680 0.150 73.810 0.330 ;
        RECT 74.190 0.150 74.320 0.330 ;
        RECT 75.680 0.150 75.810 0.330 ;
        RECT 76.190 0.150 76.320 0.330 ;
        RECT 77.680 0.150 77.810 0.330 ;
        RECT 78.190 0.150 78.320 0.330 ;
        RECT 79.680 0.150 79.810 0.330 ;
        RECT 80.190 0.150 80.320 0.330 ;
        RECT 81.680 0.150 81.810 0.330 ;
        RECT 82.190 0.150 82.320 0.330 ;
        RECT 83.680 0.150 83.810 0.330 ;
        RECT 84.190 0.150 84.320 0.330 ;
        RECT 85.680 0.150 85.810 0.330 ;
        RECT 86.190 0.150 86.320 0.330 ;
        RECT 87.680 0.150 87.810 0.330 ;
        RECT 88.190 0.150 88.320 0.330 ;
        RECT 89.680 0.150 89.810 0.330 ;
        RECT 90.190 0.150 90.320 0.330 ;
        RECT 91.680 0.150 91.810 0.330 ;
        RECT 92.190 0.150 92.320 0.330 ;
        RECT 93.680 0.150 93.810 0.330 ;
        RECT 94.190 0.150 94.320 0.330 ;
        RECT 95.680 0.150 95.810 0.330 ;
        RECT 96.190 0.150 96.320 0.330 ;
        RECT 97.680 0.150 97.810 0.330 ;
        RECT 98.190 0.150 98.320 0.330 ;
        RECT 99.680 0.150 99.810 0.330 ;
        RECT 100.190 0.150 100.320 0.330 ;
        RECT 101.680 0.150 101.810 0.330 ;
        RECT 102.190 0.150 102.320 0.330 ;
        RECT 103.680 0.150 103.810 0.330 ;
        RECT 104.190 0.150 104.320 0.330 ;
        RECT 105.680 0.150 105.810 0.330 ;
        RECT 106.190 0.150 106.320 0.330 ;
        RECT 107.680 0.150 107.810 0.330 ;
        RECT 108.190 0.150 108.320 0.330 ;
        RECT 109.680 0.150 109.810 0.330 ;
        RECT 110.190 0.150 110.320 0.330 ;
        RECT 111.680 0.150 111.810 0.330 ;
        RECT 112.190 0.150 112.320 0.330 ;
        RECT 113.680 0.150 113.810 0.330 ;
        RECT 114.190 0.150 114.320 0.330 ;
        RECT 115.680 0.150 115.810 0.330 ;
        RECT 116.190 0.150 116.320 0.330 ;
        RECT 117.680 0.150 117.810 0.330 ;
        RECT 118.190 0.150 118.320 0.330 ;
        RECT 119.680 0.150 119.810 0.330 ;
        RECT 120.190 0.150 120.320 0.330 ;
        RECT 121.680 0.150 121.810 0.330 ;
        RECT 122.190 0.150 122.320 0.330 ;
        RECT 123.680 0.150 123.810 0.330 ;
        RECT 124.190 0.150 124.320 0.330 ;
        RECT 125.680 0.150 125.810 0.330 ;
        RECT 126.190 0.150 126.320 0.330 ;
        RECT 127.680 0.150 127.810 0.330 ;
        RECT 128.190 0.150 128.320 0.330 ;
        RECT 129.680 0.150 129.810 0.330 ;
        RECT 130.190 0.150 130.320 0.330 ;
        RECT -0.320 -0.350 -0.190 -0.150 ;
        RECT -0.490 -0.650 -0.190 -0.350 ;
        RECT 0.190 -0.350 0.320 -0.150 ;
        RECT 1.680 -0.350 1.810 -0.150 ;
        RECT 0.190 -0.650 0.490 -0.350 ;
        RECT 1.510 -0.650 1.810 -0.350 ;
        RECT 2.190 -0.350 2.320 -0.150 ;
        RECT 3.680 -0.350 3.810 -0.150 ;
        RECT 2.190 -0.650 2.490 -0.350 ;
        RECT 3.510 -0.650 3.810 -0.350 ;
        RECT 4.190 -0.350 4.320 -0.150 ;
        RECT 5.680 -0.350 5.810 -0.150 ;
        RECT 4.190 -0.650 4.490 -0.350 ;
        RECT 5.510 -0.650 5.810 -0.350 ;
        RECT 6.190 -0.350 6.320 -0.150 ;
        RECT 7.680 -0.350 7.810 -0.150 ;
        RECT 6.190 -0.650 6.490 -0.350 ;
        RECT 7.510 -0.650 7.810 -0.350 ;
        RECT 8.190 -0.350 8.320 -0.150 ;
        RECT 9.680 -0.350 9.810 -0.150 ;
        RECT 8.190 -0.650 8.490 -0.350 ;
        RECT 9.510 -0.650 9.810 -0.350 ;
        RECT 10.190 -0.350 10.320 -0.150 ;
        RECT 11.680 -0.350 11.810 -0.150 ;
        RECT 10.190 -0.650 10.490 -0.350 ;
        RECT 11.510 -0.650 11.810 -0.350 ;
        RECT 12.190 -0.350 12.320 -0.150 ;
        RECT 13.680 -0.350 13.810 -0.150 ;
        RECT 12.190 -0.650 12.490 -0.350 ;
        RECT 13.510 -0.650 13.810 -0.350 ;
        RECT 14.190 -0.350 14.320 -0.150 ;
        RECT 15.680 -0.350 15.810 -0.150 ;
        RECT 14.190 -0.650 14.490 -0.350 ;
        RECT 15.510 -0.650 15.810 -0.350 ;
        RECT 16.190 -0.350 16.320 -0.150 ;
        RECT 17.680 -0.350 17.810 -0.150 ;
        RECT 16.190 -0.650 16.490 -0.350 ;
        RECT 17.510 -0.650 17.810 -0.350 ;
        RECT 18.190 -0.350 18.320 -0.150 ;
        RECT 19.680 -0.350 19.810 -0.150 ;
        RECT 18.190 -0.650 18.490 -0.350 ;
        RECT 19.510 -0.650 19.810 -0.350 ;
        RECT 20.190 -0.350 20.320 -0.150 ;
        RECT 21.680 -0.350 21.810 -0.150 ;
        RECT 20.190 -0.650 20.490 -0.350 ;
        RECT 21.510 -0.650 21.810 -0.350 ;
        RECT 22.190 -0.350 22.320 -0.150 ;
        RECT 23.680 -0.350 23.810 -0.150 ;
        RECT 22.190 -0.650 22.490 -0.350 ;
        RECT 23.510 -0.650 23.810 -0.350 ;
        RECT 24.190 -0.350 24.320 -0.150 ;
        RECT 25.680 -0.350 25.810 -0.150 ;
        RECT 24.190 -0.650 24.490 -0.350 ;
        RECT 25.510 -0.650 25.810 -0.350 ;
        RECT 26.190 -0.350 26.320 -0.150 ;
        RECT 27.680 -0.350 27.810 -0.150 ;
        RECT 26.190 -0.650 26.490 -0.350 ;
        RECT 27.510 -0.650 27.810 -0.350 ;
        RECT 28.190 -0.350 28.320 -0.150 ;
        RECT 29.680 -0.350 29.810 -0.150 ;
        RECT 28.190 -0.650 28.490 -0.350 ;
        RECT 29.510 -0.650 29.810 -0.350 ;
        RECT 30.190 -0.350 30.320 -0.150 ;
        RECT 31.680 -0.350 31.810 -0.150 ;
        RECT 30.190 -0.650 30.490 -0.350 ;
        RECT 31.510 -0.650 31.810 -0.350 ;
        RECT 32.190 -0.350 32.320 -0.150 ;
        RECT 33.680 -0.350 33.810 -0.150 ;
        RECT 32.190 -0.650 32.490 -0.350 ;
        RECT 33.510 -0.650 33.810 -0.350 ;
        RECT 34.190 -0.350 34.320 -0.150 ;
        RECT 35.680 -0.350 35.810 -0.150 ;
        RECT 34.190 -0.650 34.490 -0.350 ;
        RECT 35.510 -0.650 35.810 -0.350 ;
        RECT 36.190 -0.350 36.320 -0.150 ;
        RECT 37.680 -0.350 37.810 -0.150 ;
        RECT 36.190 -0.650 36.490 -0.350 ;
        RECT 37.510 -0.650 37.810 -0.350 ;
        RECT 38.190 -0.350 38.320 -0.150 ;
        RECT 39.680 -0.350 39.810 -0.150 ;
        RECT 38.190 -0.650 38.490 -0.350 ;
        RECT 39.510 -0.650 39.810 -0.350 ;
        RECT 40.190 -0.350 40.320 -0.150 ;
        RECT 41.680 -0.350 41.810 -0.150 ;
        RECT 40.190 -0.650 40.490 -0.350 ;
        RECT 41.510 -0.650 41.810 -0.350 ;
        RECT 42.190 -0.350 42.320 -0.150 ;
        RECT 43.680 -0.350 43.810 -0.150 ;
        RECT 42.190 -0.650 42.490 -0.350 ;
        RECT 43.510 -0.650 43.810 -0.350 ;
        RECT 44.190 -0.350 44.320 -0.150 ;
        RECT 45.680 -0.350 45.810 -0.150 ;
        RECT 44.190 -0.650 44.490 -0.350 ;
        RECT 45.510 -0.650 45.810 -0.350 ;
        RECT 46.190 -0.350 46.320 -0.150 ;
        RECT 47.680 -0.350 47.810 -0.150 ;
        RECT 46.190 -0.650 46.490 -0.350 ;
        RECT 47.510 -0.650 47.810 -0.350 ;
        RECT 48.190 -0.350 48.320 -0.150 ;
        RECT 49.680 -0.350 49.810 -0.150 ;
        RECT 48.190 -0.650 48.490 -0.350 ;
        RECT 49.510 -0.650 49.810 -0.350 ;
        RECT 50.190 -0.350 50.320 -0.150 ;
        RECT 51.680 -0.350 51.810 -0.150 ;
        RECT 50.190 -0.650 50.490 -0.350 ;
        RECT 51.510 -0.650 51.810 -0.350 ;
        RECT 52.190 -0.350 52.320 -0.150 ;
        RECT 53.680 -0.350 53.810 -0.150 ;
        RECT 52.190 -0.650 52.490 -0.350 ;
        RECT 53.510 -0.650 53.810 -0.350 ;
        RECT 54.190 -0.350 54.320 -0.150 ;
        RECT 55.680 -0.350 55.810 -0.150 ;
        RECT 54.190 -0.650 54.490 -0.350 ;
        RECT 55.510 -0.650 55.810 -0.350 ;
        RECT 56.190 -0.350 56.320 -0.150 ;
        RECT 57.680 -0.350 57.810 -0.150 ;
        RECT 56.190 -0.650 56.490 -0.350 ;
        RECT 57.510 -0.650 57.810 -0.350 ;
        RECT 58.190 -0.350 58.320 -0.150 ;
        RECT 59.680 -0.350 59.810 -0.150 ;
        RECT 58.190 -0.650 58.490 -0.350 ;
        RECT 59.510 -0.650 59.810 -0.350 ;
        RECT 60.190 -0.350 60.320 -0.150 ;
        RECT 61.680 -0.350 61.810 -0.150 ;
        RECT 60.190 -0.650 60.490 -0.350 ;
        RECT 61.510 -0.650 61.810 -0.350 ;
        RECT 62.190 -0.350 62.320 -0.150 ;
        RECT 63.680 -0.350 63.810 -0.150 ;
        RECT 62.190 -0.650 62.490 -0.350 ;
        RECT 63.510 -0.650 63.810 -0.350 ;
        RECT 64.190 -0.350 64.320 -0.150 ;
        RECT 65.680 -0.350 65.810 -0.150 ;
        RECT 64.190 -0.650 64.490 -0.350 ;
        RECT 65.510 -0.650 65.810 -0.350 ;
        RECT 66.190 -0.350 66.320 -0.150 ;
        RECT 67.680 -0.350 67.810 -0.150 ;
        RECT 66.190 -0.650 66.490 -0.350 ;
        RECT 67.510 -0.650 67.810 -0.350 ;
        RECT 68.190 -0.350 68.320 -0.150 ;
        RECT 69.680 -0.350 69.810 -0.150 ;
        RECT 68.190 -0.650 68.490 -0.350 ;
        RECT 69.510 -0.650 69.810 -0.350 ;
        RECT 70.190 -0.350 70.320 -0.150 ;
        RECT 71.680 -0.350 71.810 -0.150 ;
        RECT 70.190 -0.650 70.490 -0.350 ;
        RECT 71.510 -0.650 71.810 -0.350 ;
        RECT 72.190 -0.350 72.320 -0.150 ;
        RECT 73.680 -0.350 73.810 -0.150 ;
        RECT 72.190 -0.650 72.490 -0.350 ;
        RECT 73.510 -0.650 73.810 -0.350 ;
        RECT 74.190 -0.350 74.320 -0.150 ;
        RECT 75.680 -0.350 75.810 -0.150 ;
        RECT 74.190 -0.650 74.490 -0.350 ;
        RECT 75.510 -0.650 75.810 -0.350 ;
        RECT 76.190 -0.350 76.320 -0.150 ;
        RECT 77.680 -0.350 77.810 -0.150 ;
        RECT 76.190 -0.650 76.490 -0.350 ;
        RECT 77.510 -0.650 77.810 -0.350 ;
        RECT 78.190 -0.350 78.320 -0.150 ;
        RECT 79.680 -0.350 79.810 -0.150 ;
        RECT 78.190 -0.650 78.490 -0.350 ;
        RECT 79.510 -0.650 79.810 -0.350 ;
        RECT 80.190 -0.350 80.320 -0.150 ;
        RECT 81.680 -0.350 81.810 -0.150 ;
        RECT 80.190 -0.650 80.490 -0.350 ;
        RECT 81.510 -0.650 81.810 -0.350 ;
        RECT 82.190 -0.350 82.320 -0.150 ;
        RECT 83.680 -0.350 83.810 -0.150 ;
        RECT 82.190 -0.650 82.490 -0.350 ;
        RECT 83.510 -0.650 83.810 -0.350 ;
        RECT 84.190 -0.350 84.320 -0.150 ;
        RECT 85.680 -0.350 85.810 -0.150 ;
        RECT 84.190 -0.650 84.490 -0.350 ;
        RECT 85.510 -0.650 85.810 -0.350 ;
        RECT 86.190 -0.350 86.320 -0.150 ;
        RECT 87.680 -0.350 87.810 -0.150 ;
        RECT 86.190 -0.650 86.490 -0.350 ;
        RECT 87.510 -0.650 87.810 -0.350 ;
        RECT 88.190 -0.350 88.320 -0.150 ;
        RECT 89.680 -0.350 89.810 -0.150 ;
        RECT 88.190 -0.650 88.490 -0.350 ;
        RECT 89.510 -0.650 89.810 -0.350 ;
        RECT 90.190 -0.350 90.320 -0.150 ;
        RECT 91.680 -0.350 91.810 -0.150 ;
        RECT 90.190 -0.650 90.490 -0.350 ;
        RECT 91.510 -0.650 91.810 -0.350 ;
        RECT 92.190 -0.350 92.320 -0.150 ;
        RECT 93.680 -0.350 93.810 -0.150 ;
        RECT 92.190 -0.650 92.490 -0.350 ;
        RECT 93.510 -0.650 93.810 -0.350 ;
        RECT 94.190 -0.350 94.320 -0.150 ;
        RECT 95.680 -0.350 95.810 -0.150 ;
        RECT 94.190 -0.650 94.490 -0.350 ;
        RECT 95.510 -0.650 95.810 -0.350 ;
        RECT 96.190 -0.350 96.320 -0.150 ;
        RECT 97.680 -0.350 97.810 -0.150 ;
        RECT 96.190 -0.650 96.490 -0.350 ;
        RECT 97.510 -0.650 97.810 -0.350 ;
        RECT 98.190 -0.350 98.320 -0.150 ;
        RECT 99.680 -0.350 99.810 -0.150 ;
        RECT 98.190 -0.650 98.490 -0.350 ;
        RECT 99.510 -0.650 99.810 -0.350 ;
        RECT 100.190 -0.350 100.320 -0.150 ;
        RECT 101.680 -0.350 101.810 -0.150 ;
        RECT 100.190 -0.650 100.490 -0.350 ;
        RECT 101.510 -0.650 101.810 -0.350 ;
        RECT 102.190 -0.350 102.320 -0.150 ;
        RECT 103.680 -0.350 103.810 -0.150 ;
        RECT 102.190 -0.650 102.490 -0.350 ;
        RECT 103.510 -0.650 103.810 -0.350 ;
        RECT 104.190 -0.350 104.320 -0.150 ;
        RECT 105.680 -0.350 105.810 -0.150 ;
        RECT 104.190 -0.650 104.490 -0.350 ;
        RECT 105.510 -0.650 105.810 -0.350 ;
        RECT 106.190 -0.350 106.320 -0.150 ;
        RECT 107.680 -0.350 107.810 -0.150 ;
        RECT 106.190 -0.650 106.490 -0.350 ;
        RECT 107.510 -0.650 107.810 -0.350 ;
        RECT 108.190 -0.350 108.320 -0.150 ;
        RECT 109.680 -0.350 109.810 -0.150 ;
        RECT 108.190 -0.650 108.490 -0.350 ;
        RECT 109.510 -0.650 109.810 -0.350 ;
        RECT 110.190 -0.350 110.320 -0.150 ;
        RECT 111.680 -0.350 111.810 -0.150 ;
        RECT 110.190 -0.650 110.490 -0.350 ;
        RECT 111.510 -0.650 111.810 -0.350 ;
        RECT 112.190 -0.350 112.320 -0.150 ;
        RECT 113.680 -0.350 113.810 -0.150 ;
        RECT 112.190 -0.650 112.490 -0.350 ;
        RECT 113.510 -0.650 113.810 -0.350 ;
        RECT 114.190 -0.350 114.320 -0.150 ;
        RECT 115.680 -0.350 115.810 -0.150 ;
        RECT 114.190 -0.650 114.490 -0.350 ;
        RECT 115.510 -0.650 115.810 -0.350 ;
        RECT 116.190 -0.350 116.320 -0.150 ;
        RECT 117.680 -0.350 117.810 -0.150 ;
        RECT 116.190 -0.650 116.490 -0.350 ;
        RECT 117.510 -0.650 117.810 -0.350 ;
        RECT 118.190 -0.350 118.320 -0.150 ;
        RECT 119.680 -0.350 119.810 -0.150 ;
        RECT 118.190 -0.650 118.490 -0.350 ;
        RECT 119.510 -0.650 119.810 -0.350 ;
        RECT 120.190 -0.350 120.320 -0.150 ;
        RECT 121.680 -0.350 121.810 -0.150 ;
        RECT 120.190 -0.650 120.490 -0.350 ;
        RECT 121.510 -0.650 121.810 -0.350 ;
        RECT 122.190 -0.350 122.320 -0.150 ;
        RECT 123.680 -0.350 123.810 -0.150 ;
        RECT 122.190 -0.650 122.490 -0.350 ;
        RECT 123.510 -0.650 123.810 -0.350 ;
        RECT 124.190 -0.350 124.320 -0.150 ;
        RECT 125.680 -0.350 125.810 -0.150 ;
        RECT 124.190 -0.650 124.490 -0.350 ;
        RECT 125.510 -0.650 125.810 -0.350 ;
        RECT 126.190 -0.350 126.320 -0.150 ;
        RECT 127.680 -0.350 127.810 -0.150 ;
        RECT 126.190 -0.650 126.490 -0.350 ;
        RECT 127.510 -0.650 127.810 -0.350 ;
        RECT 128.190 -0.350 128.320 -0.150 ;
        RECT 129.680 -0.350 129.810 -0.150 ;
        RECT 128.190 -0.650 128.490 -0.350 ;
        RECT 129.510 -0.650 129.810 -0.350 ;
        RECT 130.190 -0.350 130.320 -0.150 ;
        RECT 130.190 -0.650 130.490 -0.350 ;
        RECT -0.320 -1.730 -0.190 -1.550 ;
        RECT 0.190 -1.730 0.320 -1.550 ;
        RECT 1.680 -1.730 1.810 -1.550 ;
        RECT 2.190 -1.730 2.320 -1.550 ;
        RECT 3.680 -1.730 3.810 -1.550 ;
        RECT 4.190 -1.730 4.320 -1.550 ;
        RECT 5.680 -1.730 5.810 -1.550 ;
        RECT 6.190 -1.730 6.320 -1.550 ;
        RECT 7.680 -1.730 7.810 -1.550 ;
        RECT 8.190 -1.730 8.320 -1.550 ;
        RECT 9.680 -1.730 9.810 -1.550 ;
        RECT 10.190 -1.730 10.320 -1.550 ;
        RECT 11.680 -1.730 11.810 -1.550 ;
        RECT 12.190 -1.730 12.320 -1.550 ;
        RECT 13.680 -1.730 13.810 -1.550 ;
        RECT 14.190 -1.730 14.320 -1.550 ;
        RECT 15.680 -1.730 15.810 -1.550 ;
        RECT 16.190 -1.730 16.320 -1.550 ;
        RECT 17.680 -1.730 17.810 -1.550 ;
        RECT 18.190 -1.730 18.320 -1.550 ;
        RECT 19.680 -1.730 19.810 -1.550 ;
        RECT 20.190 -1.730 20.320 -1.550 ;
        RECT 21.680 -1.730 21.810 -1.550 ;
        RECT 22.190 -1.730 22.320 -1.550 ;
        RECT 23.680 -1.730 23.810 -1.550 ;
        RECT 24.190 -1.730 24.320 -1.550 ;
        RECT 25.680 -1.730 25.810 -1.550 ;
        RECT 26.190 -1.730 26.320 -1.550 ;
        RECT 27.680 -1.730 27.810 -1.550 ;
        RECT 28.190 -1.730 28.320 -1.550 ;
        RECT 29.680 -1.730 29.810 -1.550 ;
        RECT 30.190 -1.730 30.320 -1.550 ;
        RECT 31.680 -1.730 31.810 -1.550 ;
        RECT 32.190 -1.730 32.320 -1.550 ;
        RECT 33.680 -1.730 33.810 -1.550 ;
        RECT 34.190 -1.730 34.320 -1.550 ;
        RECT 35.680 -1.730 35.810 -1.550 ;
        RECT 36.190 -1.730 36.320 -1.550 ;
        RECT 37.680 -1.730 37.810 -1.550 ;
        RECT 38.190 -1.730 38.320 -1.550 ;
        RECT 39.680 -1.730 39.810 -1.550 ;
        RECT 40.190 -1.730 40.320 -1.550 ;
        RECT 41.680 -1.730 41.810 -1.550 ;
        RECT 42.190 -1.730 42.320 -1.550 ;
        RECT 43.680 -1.730 43.810 -1.550 ;
        RECT 44.190 -1.730 44.320 -1.550 ;
        RECT 45.680 -1.730 45.810 -1.550 ;
        RECT 46.190 -1.730 46.320 -1.550 ;
        RECT 47.680 -1.730 47.810 -1.550 ;
        RECT 48.190 -1.730 48.320 -1.550 ;
        RECT 49.680 -1.730 49.810 -1.550 ;
        RECT 50.190 -1.730 50.320 -1.550 ;
        RECT 51.680 -1.730 51.810 -1.550 ;
        RECT 52.190 -1.730 52.320 -1.550 ;
        RECT 53.680 -1.730 53.810 -1.550 ;
        RECT 54.190 -1.730 54.320 -1.550 ;
        RECT 55.680 -1.730 55.810 -1.550 ;
        RECT 56.190 -1.730 56.320 -1.550 ;
        RECT 57.680 -1.730 57.810 -1.550 ;
        RECT 58.190 -1.730 58.320 -1.550 ;
        RECT 59.680 -1.730 59.810 -1.550 ;
        RECT 60.190 -1.730 60.320 -1.550 ;
        RECT 61.680 -1.730 61.810 -1.550 ;
        RECT 62.190 -1.730 62.320 -1.550 ;
        RECT 63.680 -1.730 63.810 -1.550 ;
        RECT 64.190 -1.730 64.320 -1.550 ;
        RECT 65.680 -1.730 65.810 -1.550 ;
        RECT 66.190 -1.730 66.320 -1.550 ;
        RECT 67.680 -1.730 67.810 -1.550 ;
        RECT 68.190 -1.730 68.320 -1.550 ;
        RECT 69.680 -1.730 69.810 -1.550 ;
        RECT 70.190 -1.730 70.320 -1.550 ;
        RECT 71.680 -1.730 71.810 -1.550 ;
        RECT 72.190 -1.730 72.320 -1.550 ;
        RECT 73.680 -1.730 73.810 -1.550 ;
        RECT 74.190 -1.730 74.320 -1.550 ;
        RECT 75.680 -1.730 75.810 -1.550 ;
        RECT 76.190 -1.730 76.320 -1.550 ;
        RECT 77.680 -1.730 77.810 -1.550 ;
        RECT 78.190 -1.730 78.320 -1.550 ;
        RECT 79.680 -1.730 79.810 -1.550 ;
        RECT 80.190 -1.730 80.320 -1.550 ;
        RECT 81.680 -1.730 81.810 -1.550 ;
        RECT 82.190 -1.730 82.320 -1.550 ;
        RECT 83.680 -1.730 83.810 -1.550 ;
        RECT 84.190 -1.730 84.320 -1.550 ;
        RECT 85.680 -1.730 85.810 -1.550 ;
        RECT 86.190 -1.730 86.320 -1.550 ;
        RECT 87.680 -1.730 87.810 -1.550 ;
        RECT 88.190 -1.730 88.320 -1.550 ;
        RECT 89.680 -1.730 89.810 -1.550 ;
        RECT 90.190 -1.730 90.320 -1.550 ;
        RECT 91.680 -1.730 91.810 -1.550 ;
        RECT 92.190 -1.730 92.320 -1.550 ;
        RECT 93.680 -1.730 93.810 -1.550 ;
        RECT 94.190 -1.730 94.320 -1.550 ;
        RECT 95.680 -1.730 95.810 -1.550 ;
        RECT 96.190 -1.730 96.320 -1.550 ;
        RECT 97.680 -1.730 97.810 -1.550 ;
        RECT 98.190 -1.730 98.320 -1.550 ;
        RECT 99.680 -1.730 99.810 -1.550 ;
        RECT 100.190 -1.730 100.320 -1.550 ;
        RECT 101.680 -1.730 101.810 -1.550 ;
        RECT 102.190 -1.730 102.320 -1.550 ;
        RECT 103.680 -1.730 103.810 -1.550 ;
        RECT 104.190 -1.730 104.320 -1.550 ;
        RECT 105.680 -1.730 105.810 -1.550 ;
        RECT 106.190 -1.730 106.320 -1.550 ;
        RECT 107.680 -1.730 107.810 -1.550 ;
        RECT 108.190 -1.730 108.320 -1.550 ;
        RECT 109.680 -1.730 109.810 -1.550 ;
        RECT 110.190 -1.730 110.320 -1.550 ;
        RECT 111.680 -1.730 111.810 -1.550 ;
        RECT 112.190 -1.730 112.320 -1.550 ;
        RECT 113.680 -1.730 113.810 -1.550 ;
        RECT 114.190 -1.730 114.320 -1.550 ;
        RECT 115.680 -1.730 115.810 -1.550 ;
        RECT 116.190 -1.730 116.320 -1.550 ;
        RECT 117.680 -1.730 117.810 -1.550 ;
        RECT 118.190 -1.730 118.320 -1.550 ;
        RECT 119.680 -1.730 119.810 -1.550 ;
        RECT 120.190 -1.730 120.320 -1.550 ;
        RECT 121.680 -1.730 121.810 -1.550 ;
        RECT 122.190 -1.730 122.320 -1.550 ;
        RECT 123.680 -1.730 123.810 -1.550 ;
        RECT 124.190 -1.730 124.320 -1.550 ;
        RECT 125.680 -1.730 125.810 -1.550 ;
        RECT 126.190 -1.730 126.320 -1.550 ;
        RECT 127.680 -1.730 127.810 -1.550 ;
        RECT 128.190 -1.730 128.320 -1.550 ;
        RECT 129.680 -1.730 129.810 -1.550 ;
        RECT 130.190 -1.730 130.320 -1.550 ;
        RECT -0.320 -2.100 -0.190 -2.030 ;
        RECT -0.490 -2.400 -0.190 -2.100 ;
        RECT 0.190 -2.100 0.320 -2.030 ;
        RECT 1.680 -2.100 1.810 -2.030 ;
        RECT 0.190 -2.400 0.490 -2.100 ;
        RECT 1.510 -2.400 1.810 -2.100 ;
        RECT 2.190 -2.100 2.320 -2.030 ;
        RECT 3.680 -2.100 3.810 -2.030 ;
        RECT 2.190 -2.400 2.490 -2.100 ;
        RECT 3.510 -2.400 3.810 -2.100 ;
        RECT 4.190 -2.100 4.320 -2.030 ;
        RECT 5.680 -2.100 5.810 -2.030 ;
        RECT 4.190 -2.400 4.490 -2.100 ;
        RECT 5.510 -2.400 5.810 -2.100 ;
        RECT 6.190 -2.100 6.320 -2.030 ;
        RECT 7.680 -2.100 7.810 -2.030 ;
        RECT 6.190 -2.400 6.490 -2.100 ;
        RECT 7.510 -2.400 7.810 -2.100 ;
        RECT 8.190 -2.100 8.320 -2.030 ;
        RECT 9.680 -2.100 9.810 -2.030 ;
        RECT 8.190 -2.400 8.490 -2.100 ;
        RECT 9.510 -2.400 9.810 -2.100 ;
        RECT 10.190 -2.100 10.320 -2.030 ;
        RECT 11.680 -2.100 11.810 -2.030 ;
        RECT 10.190 -2.400 10.490 -2.100 ;
        RECT 11.510 -2.400 11.810 -2.100 ;
        RECT 12.190 -2.100 12.320 -2.030 ;
        RECT 13.680 -2.100 13.810 -2.030 ;
        RECT 12.190 -2.400 12.490 -2.100 ;
        RECT 13.510 -2.400 13.810 -2.100 ;
        RECT 14.190 -2.100 14.320 -2.030 ;
        RECT 15.680 -2.100 15.810 -2.030 ;
        RECT 14.190 -2.400 14.490 -2.100 ;
        RECT 15.510 -2.400 15.810 -2.100 ;
        RECT 16.190 -2.100 16.320 -2.030 ;
        RECT 17.680 -2.100 17.810 -2.030 ;
        RECT 16.190 -2.400 16.490 -2.100 ;
        RECT 17.510 -2.400 17.810 -2.100 ;
        RECT 18.190 -2.100 18.320 -2.030 ;
        RECT 19.680 -2.100 19.810 -2.030 ;
        RECT 18.190 -2.400 18.490 -2.100 ;
        RECT 19.510 -2.400 19.810 -2.100 ;
        RECT 20.190 -2.100 20.320 -2.030 ;
        RECT 21.680 -2.100 21.810 -2.030 ;
        RECT 20.190 -2.400 20.490 -2.100 ;
        RECT 21.510 -2.400 21.810 -2.100 ;
        RECT 22.190 -2.100 22.320 -2.030 ;
        RECT 23.680 -2.100 23.810 -2.030 ;
        RECT 22.190 -2.400 22.490 -2.100 ;
        RECT 23.510 -2.400 23.810 -2.100 ;
        RECT 24.190 -2.100 24.320 -2.030 ;
        RECT 25.680 -2.100 25.810 -2.030 ;
        RECT 24.190 -2.400 24.490 -2.100 ;
        RECT 25.510 -2.400 25.810 -2.100 ;
        RECT 26.190 -2.100 26.320 -2.030 ;
        RECT 27.680 -2.100 27.810 -2.030 ;
        RECT 26.190 -2.400 26.490 -2.100 ;
        RECT 27.510 -2.400 27.810 -2.100 ;
        RECT 28.190 -2.100 28.320 -2.030 ;
        RECT 29.680 -2.100 29.810 -2.030 ;
        RECT 28.190 -2.400 28.490 -2.100 ;
        RECT 29.510 -2.400 29.810 -2.100 ;
        RECT 30.190 -2.100 30.320 -2.030 ;
        RECT 31.680 -2.100 31.810 -2.030 ;
        RECT 30.190 -2.400 30.490 -2.100 ;
        RECT 31.510 -2.400 31.810 -2.100 ;
        RECT 32.190 -2.100 32.320 -2.030 ;
        RECT 33.680 -2.100 33.810 -2.030 ;
        RECT 32.190 -2.400 32.490 -2.100 ;
        RECT 33.510 -2.400 33.810 -2.100 ;
        RECT 34.190 -2.100 34.320 -2.030 ;
        RECT 35.680 -2.100 35.810 -2.030 ;
        RECT 34.190 -2.400 34.490 -2.100 ;
        RECT 35.510 -2.400 35.810 -2.100 ;
        RECT 36.190 -2.100 36.320 -2.030 ;
        RECT 37.680 -2.100 37.810 -2.030 ;
        RECT 36.190 -2.400 36.490 -2.100 ;
        RECT 37.510 -2.400 37.810 -2.100 ;
        RECT 38.190 -2.100 38.320 -2.030 ;
        RECT 39.680 -2.100 39.810 -2.030 ;
        RECT 38.190 -2.400 38.490 -2.100 ;
        RECT 39.510 -2.400 39.810 -2.100 ;
        RECT 40.190 -2.100 40.320 -2.030 ;
        RECT 41.680 -2.100 41.810 -2.030 ;
        RECT 40.190 -2.400 40.490 -2.100 ;
        RECT 41.510 -2.400 41.810 -2.100 ;
        RECT 42.190 -2.100 42.320 -2.030 ;
        RECT 43.680 -2.100 43.810 -2.030 ;
        RECT 42.190 -2.400 42.490 -2.100 ;
        RECT 43.510 -2.400 43.810 -2.100 ;
        RECT 44.190 -2.100 44.320 -2.030 ;
        RECT 45.680 -2.100 45.810 -2.030 ;
        RECT 44.190 -2.400 44.490 -2.100 ;
        RECT 45.510 -2.400 45.810 -2.100 ;
        RECT 46.190 -2.100 46.320 -2.030 ;
        RECT 47.680 -2.100 47.810 -2.030 ;
        RECT 46.190 -2.400 46.490 -2.100 ;
        RECT 47.510 -2.400 47.810 -2.100 ;
        RECT 48.190 -2.100 48.320 -2.030 ;
        RECT 49.680 -2.100 49.810 -2.030 ;
        RECT 48.190 -2.400 48.490 -2.100 ;
        RECT 49.510 -2.400 49.810 -2.100 ;
        RECT 50.190 -2.100 50.320 -2.030 ;
        RECT 51.680 -2.100 51.810 -2.030 ;
        RECT 50.190 -2.400 50.490 -2.100 ;
        RECT 51.510 -2.400 51.810 -2.100 ;
        RECT 52.190 -2.100 52.320 -2.030 ;
        RECT 53.680 -2.100 53.810 -2.030 ;
        RECT 52.190 -2.400 52.490 -2.100 ;
        RECT 53.510 -2.400 53.810 -2.100 ;
        RECT 54.190 -2.100 54.320 -2.030 ;
        RECT 55.680 -2.100 55.810 -2.030 ;
        RECT 54.190 -2.400 54.490 -2.100 ;
        RECT 55.510 -2.400 55.810 -2.100 ;
        RECT 56.190 -2.100 56.320 -2.030 ;
        RECT 57.680 -2.100 57.810 -2.030 ;
        RECT 56.190 -2.400 56.490 -2.100 ;
        RECT 57.510 -2.400 57.810 -2.100 ;
        RECT 58.190 -2.100 58.320 -2.030 ;
        RECT 59.680 -2.100 59.810 -2.030 ;
        RECT 58.190 -2.400 58.490 -2.100 ;
        RECT 59.510 -2.400 59.810 -2.100 ;
        RECT 60.190 -2.100 60.320 -2.030 ;
        RECT 61.680 -2.100 61.810 -2.030 ;
        RECT 60.190 -2.400 60.490 -2.100 ;
        RECT 61.510 -2.400 61.810 -2.100 ;
        RECT 62.190 -2.100 62.320 -2.030 ;
        RECT 63.680 -2.100 63.810 -2.030 ;
        RECT 62.190 -2.400 62.490 -2.100 ;
        RECT 63.510 -2.400 63.810 -2.100 ;
        RECT 64.190 -2.100 64.320 -2.030 ;
        RECT 65.680 -2.100 65.810 -2.030 ;
        RECT 64.190 -2.400 64.490 -2.100 ;
        RECT 65.510 -2.400 65.810 -2.100 ;
        RECT 66.190 -2.100 66.320 -2.030 ;
        RECT 67.680 -2.100 67.810 -2.030 ;
        RECT 66.190 -2.400 66.490 -2.100 ;
        RECT 67.510 -2.400 67.810 -2.100 ;
        RECT 68.190 -2.100 68.320 -2.030 ;
        RECT 69.680 -2.100 69.810 -2.030 ;
        RECT 68.190 -2.400 68.490 -2.100 ;
        RECT 69.510 -2.400 69.810 -2.100 ;
        RECT 70.190 -2.100 70.320 -2.030 ;
        RECT 71.680 -2.100 71.810 -2.030 ;
        RECT 70.190 -2.400 70.490 -2.100 ;
        RECT 71.510 -2.400 71.810 -2.100 ;
        RECT 72.190 -2.100 72.320 -2.030 ;
        RECT 73.680 -2.100 73.810 -2.030 ;
        RECT 72.190 -2.400 72.490 -2.100 ;
        RECT 73.510 -2.400 73.810 -2.100 ;
        RECT 74.190 -2.100 74.320 -2.030 ;
        RECT 75.680 -2.100 75.810 -2.030 ;
        RECT 74.190 -2.400 74.490 -2.100 ;
        RECT 75.510 -2.400 75.810 -2.100 ;
        RECT 76.190 -2.100 76.320 -2.030 ;
        RECT 77.680 -2.100 77.810 -2.030 ;
        RECT 76.190 -2.400 76.490 -2.100 ;
        RECT 77.510 -2.400 77.810 -2.100 ;
        RECT 78.190 -2.100 78.320 -2.030 ;
        RECT 79.680 -2.100 79.810 -2.030 ;
        RECT 78.190 -2.400 78.490 -2.100 ;
        RECT 79.510 -2.400 79.810 -2.100 ;
        RECT 80.190 -2.100 80.320 -2.030 ;
        RECT 81.680 -2.100 81.810 -2.030 ;
        RECT 80.190 -2.400 80.490 -2.100 ;
        RECT 81.510 -2.400 81.810 -2.100 ;
        RECT 82.190 -2.100 82.320 -2.030 ;
        RECT 83.680 -2.100 83.810 -2.030 ;
        RECT 82.190 -2.400 82.490 -2.100 ;
        RECT 83.510 -2.400 83.810 -2.100 ;
        RECT 84.190 -2.100 84.320 -2.030 ;
        RECT 85.680 -2.100 85.810 -2.030 ;
        RECT 84.190 -2.400 84.490 -2.100 ;
        RECT 85.510 -2.400 85.810 -2.100 ;
        RECT 86.190 -2.100 86.320 -2.030 ;
        RECT 87.680 -2.100 87.810 -2.030 ;
        RECT 86.190 -2.400 86.490 -2.100 ;
        RECT 87.510 -2.400 87.810 -2.100 ;
        RECT 88.190 -2.100 88.320 -2.030 ;
        RECT 89.680 -2.100 89.810 -2.030 ;
        RECT 88.190 -2.400 88.490 -2.100 ;
        RECT 89.510 -2.400 89.810 -2.100 ;
        RECT 90.190 -2.100 90.320 -2.030 ;
        RECT 91.680 -2.100 91.810 -2.030 ;
        RECT 90.190 -2.400 90.490 -2.100 ;
        RECT 91.510 -2.400 91.810 -2.100 ;
        RECT 92.190 -2.100 92.320 -2.030 ;
        RECT 93.680 -2.100 93.810 -2.030 ;
        RECT 92.190 -2.400 92.490 -2.100 ;
        RECT 93.510 -2.400 93.810 -2.100 ;
        RECT 94.190 -2.100 94.320 -2.030 ;
        RECT 95.680 -2.100 95.810 -2.030 ;
        RECT 94.190 -2.400 94.490 -2.100 ;
        RECT 95.510 -2.400 95.810 -2.100 ;
        RECT 96.190 -2.100 96.320 -2.030 ;
        RECT 97.680 -2.100 97.810 -2.030 ;
        RECT 96.190 -2.400 96.490 -2.100 ;
        RECT 97.510 -2.400 97.810 -2.100 ;
        RECT 98.190 -2.100 98.320 -2.030 ;
        RECT 99.680 -2.100 99.810 -2.030 ;
        RECT 98.190 -2.400 98.490 -2.100 ;
        RECT 99.510 -2.400 99.810 -2.100 ;
        RECT 100.190 -2.100 100.320 -2.030 ;
        RECT 101.680 -2.100 101.810 -2.030 ;
        RECT 100.190 -2.400 100.490 -2.100 ;
        RECT 101.510 -2.400 101.810 -2.100 ;
        RECT 102.190 -2.100 102.320 -2.030 ;
        RECT 103.680 -2.100 103.810 -2.030 ;
        RECT 102.190 -2.400 102.490 -2.100 ;
        RECT 103.510 -2.400 103.810 -2.100 ;
        RECT 104.190 -2.100 104.320 -2.030 ;
        RECT 105.680 -2.100 105.810 -2.030 ;
        RECT 104.190 -2.400 104.490 -2.100 ;
        RECT 105.510 -2.400 105.810 -2.100 ;
        RECT 106.190 -2.100 106.320 -2.030 ;
        RECT 107.680 -2.100 107.810 -2.030 ;
        RECT 106.190 -2.400 106.490 -2.100 ;
        RECT 107.510 -2.400 107.810 -2.100 ;
        RECT 108.190 -2.100 108.320 -2.030 ;
        RECT 109.680 -2.100 109.810 -2.030 ;
        RECT 108.190 -2.400 108.490 -2.100 ;
        RECT 109.510 -2.400 109.810 -2.100 ;
        RECT 110.190 -2.100 110.320 -2.030 ;
        RECT 111.680 -2.100 111.810 -2.030 ;
        RECT 110.190 -2.400 110.490 -2.100 ;
        RECT 111.510 -2.400 111.810 -2.100 ;
        RECT 112.190 -2.100 112.320 -2.030 ;
        RECT 113.680 -2.100 113.810 -2.030 ;
        RECT 112.190 -2.400 112.490 -2.100 ;
        RECT 113.510 -2.400 113.810 -2.100 ;
        RECT 114.190 -2.100 114.320 -2.030 ;
        RECT 115.680 -2.100 115.810 -2.030 ;
        RECT 114.190 -2.400 114.490 -2.100 ;
        RECT 115.510 -2.400 115.810 -2.100 ;
        RECT 116.190 -2.100 116.320 -2.030 ;
        RECT 117.680 -2.100 117.810 -2.030 ;
        RECT 116.190 -2.400 116.490 -2.100 ;
        RECT 117.510 -2.400 117.810 -2.100 ;
        RECT 118.190 -2.100 118.320 -2.030 ;
        RECT 119.680 -2.100 119.810 -2.030 ;
        RECT 118.190 -2.400 118.490 -2.100 ;
        RECT 119.510 -2.400 119.810 -2.100 ;
        RECT 120.190 -2.100 120.320 -2.030 ;
        RECT 121.680 -2.100 121.810 -2.030 ;
        RECT 120.190 -2.400 120.490 -2.100 ;
        RECT 121.510 -2.400 121.810 -2.100 ;
        RECT 122.190 -2.100 122.320 -2.030 ;
        RECT 123.680 -2.100 123.810 -2.030 ;
        RECT 122.190 -2.400 122.490 -2.100 ;
        RECT 123.510 -2.400 123.810 -2.100 ;
        RECT 124.190 -2.100 124.320 -2.030 ;
        RECT 125.680 -2.100 125.810 -2.030 ;
        RECT 124.190 -2.400 124.490 -2.100 ;
        RECT 125.510 -2.400 125.810 -2.100 ;
        RECT 126.190 -2.100 126.320 -2.030 ;
        RECT 127.680 -2.100 127.810 -2.030 ;
        RECT 126.190 -2.400 126.490 -2.100 ;
        RECT 127.510 -2.400 127.810 -2.100 ;
        RECT 128.190 -2.100 128.320 -2.030 ;
        RECT 129.680 -2.100 129.810 -2.030 ;
        RECT 128.190 -2.400 128.490 -2.100 ;
        RECT 129.510 -2.400 129.810 -2.100 ;
        RECT 130.190 -2.100 130.320 -2.030 ;
        RECT 130.190 -2.400 130.490 -2.100 ;
        RECT -0.445 -2.880 0.895 -2.580 ;
        RECT 1.555 -2.880 2.895 -2.580 ;
        RECT 3.555 -2.880 4.895 -2.580 ;
        RECT 5.555 -2.880 6.895 -2.580 ;
        RECT 7.555 -2.880 8.895 -2.580 ;
        RECT 9.555 -2.880 10.895 -2.580 ;
        RECT 11.555 -2.880 12.895 -2.580 ;
        RECT 13.555 -2.880 14.895 -2.580 ;
        RECT 15.555 -2.880 16.895 -2.580 ;
        RECT 17.555 -2.880 18.895 -2.580 ;
        RECT 19.555 -2.880 20.895 -2.580 ;
        RECT 21.555 -2.880 22.895 -2.580 ;
        RECT 23.555 -2.880 24.895 -2.580 ;
        RECT 25.555 -2.880 26.895 -2.580 ;
        RECT 27.555 -2.880 28.895 -2.580 ;
        RECT 29.555 -2.880 30.895 -2.580 ;
        RECT 31.555 -2.880 32.895 -2.580 ;
        RECT 33.555 -2.880 34.895 -2.580 ;
        RECT 35.555 -2.880 36.895 -2.580 ;
        RECT 37.555 -2.880 38.895 -2.580 ;
        RECT 39.555 -2.880 40.895 -2.580 ;
        RECT 41.555 -2.880 42.895 -2.580 ;
        RECT 43.555 -2.880 44.895 -2.580 ;
        RECT 45.555 -2.880 46.895 -2.580 ;
        RECT 47.555 -2.880 48.895 -2.580 ;
        RECT 49.555 -2.880 50.895 -2.580 ;
        RECT 51.555 -2.880 52.895 -2.580 ;
        RECT 53.555 -2.880 54.895 -2.580 ;
        RECT 55.555 -2.880 56.895 -2.580 ;
        RECT 57.555 -2.880 58.895 -2.580 ;
        RECT 59.555 -2.880 60.895 -2.580 ;
        RECT 61.555 -2.880 62.895 -2.580 ;
        RECT 63.555 -2.880 64.895 -2.580 ;
        RECT 65.555 -2.880 66.895 -2.580 ;
        RECT 67.555 -2.880 68.895 -2.580 ;
        RECT 69.555 -2.880 70.895 -2.580 ;
        RECT 71.555 -2.880 72.895 -2.580 ;
        RECT 73.555 -2.880 74.895 -2.580 ;
        RECT 75.555 -2.880 76.895 -2.580 ;
        RECT 77.555 -2.880 78.895 -2.580 ;
        RECT 79.555 -2.880 80.895 -2.580 ;
        RECT 81.555 -2.880 82.895 -2.580 ;
        RECT 83.555 -2.880 84.895 -2.580 ;
        RECT 85.555 -2.880 86.895 -2.580 ;
        RECT 87.555 -2.880 88.895 -2.580 ;
        RECT 89.555 -2.880 90.895 -2.580 ;
        RECT 91.555 -2.880 92.895 -2.580 ;
        RECT 93.555 -2.880 94.895 -2.580 ;
        RECT 95.555 -2.880 96.895 -2.580 ;
        RECT 97.555 -2.880 98.895 -2.580 ;
        RECT 99.555 -2.880 100.895 -2.580 ;
        RECT 101.555 -2.880 102.895 -2.580 ;
        RECT 103.555 -2.880 104.895 -2.580 ;
        RECT 105.555 -2.880 106.895 -2.580 ;
        RECT 107.555 -2.880 108.895 -2.580 ;
        RECT 109.555 -2.880 110.895 -2.580 ;
        RECT 111.555 -2.880 112.895 -2.580 ;
        RECT 113.555 -2.880 114.895 -2.580 ;
        RECT 115.555 -2.880 116.895 -2.580 ;
        RECT 117.555 -2.880 118.895 -2.580 ;
        RECT 119.555 -2.880 120.895 -2.580 ;
        RECT 121.555 -2.880 122.895 -2.580 ;
        RECT 123.555 -2.880 124.895 -2.580 ;
        RECT 125.555 -2.880 126.895 -2.580 ;
        RECT 127.555 -2.880 128.895 -2.580 ;
        RECT 129.555 -2.880 130.895 -2.580 ;
        RECT -0.445 -3.250 -0.145 -2.880 ;
        RECT -0.665 -3.430 -0.145 -3.250 ;
        RECT 0.145 -3.250 0.445 -3.060 ;
        RECT 1.555 -3.250 1.855 -2.880 ;
        RECT 0.145 -3.430 0.665 -3.250 ;
        RECT 1.335 -3.430 1.855 -3.250 ;
        RECT 2.145 -3.250 2.445 -3.060 ;
        RECT 3.555 -3.250 3.855 -2.880 ;
        RECT 2.145 -3.430 2.665 -3.250 ;
        RECT 3.335 -3.430 3.855 -3.250 ;
        RECT 4.145 -3.250 4.445 -3.060 ;
        RECT 5.555 -3.250 5.855 -2.880 ;
        RECT 4.145 -3.430 4.665 -3.250 ;
        RECT 5.335 -3.430 5.855 -3.250 ;
        RECT 6.145 -3.250 6.445 -3.060 ;
        RECT 7.555 -3.250 7.855 -2.880 ;
        RECT 6.145 -3.430 6.665 -3.250 ;
        RECT 7.335 -3.430 7.855 -3.250 ;
        RECT 8.145 -3.250 8.445 -3.060 ;
        RECT 9.555 -3.250 9.855 -2.880 ;
        RECT 8.145 -3.430 8.665 -3.250 ;
        RECT 9.335 -3.430 9.855 -3.250 ;
        RECT 10.145 -3.250 10.445 -3.060 ;
        RECT 11.555 -3.250 11.855 -2.880 ;
        RECT 10.145 -3.430 10.665 -3.250 ;
        RECT 11.335 -3.430 11.855 -3.250 ;
        RECT 12.145 -3.250 12.445 -3.060 ;
        RECT 13.555 -3.250 13.855 -2.880 ;
        RECT 12.145 -3.430 12.665 -3.250 ;
        RECT 13.335 -3.430 13.855 -3.250 ;
        RECT 14.145 -3.250 14.445 -3.060 ;
        RECT 15.555 -3.250 15.855 -2.880 ;
        RECT 14.145 -3.430 14.665 -3.250 ;
        RECT 15.335 -3.430 15.855 -3.250 ;
        RECT 16.145 -3.250 16.445 -3.060 ;
        RECT 17.555 -3.250 17.855 -2.880 ;
        RECT 16.145 -3.430 16.665 -3.250 ;
        RECT 17.335 -3.430 17.855 -3.250 ;
        RECT 18.145 -3.250 18.445 -3.060 ;
        RECT 19.555 -3.250 19.855 -2.880 ;
        RECT 18.145 -3.430 18.665 -3.250 ;
        RECT 19.335 -3.430 19.855 -3.250 ;
        RECT 20.145 -3.250 20.445 -3.060 ;
        RECT 21.555 -3.250 21.855 -2.880 ;
        RECT 20.145 -3.430 20.665 -3.250 ;
        RECT 21.335 -3.430 21.855 -3.250 ;
        RECT 22.145 -3.250 22.445 -3.060 ;
        RECT 23.555 -3.250 23.855 -2.880 ;
        RECT 22.145 -3.430 22.665 -3.250 ;
        RECT 23.335 -3.430 23.855 -3.250 ;
        RECT 24.145 -3.250 24.445 -3.060 ;
        RECT 25.555 -3.250 25.855 -2.880 ;
        RECT 24.145 -3.430 24.665 -3.250 ;
        RECT 25.335 -3.430 25.855 -3.250 ;
        RECT 26.145 -3.250 26.445 -3.060 ;
        RECT 27.555 -3.250 27.855 -2.880 ;
        RECT 26.145 -3.430 26.665 -3.250 ;
        RECT 27.335 -3.430 27.855 -3.250 ;
        RECT 28.145 -3.250 28.445 -3.060 ;
        RECT 29.555 -3.250 29.855 -2.880 ;
        RECT 28.145 -3.430 28.665 -3.250 ;
        RECT 29.335 -3.430 29.855 -3.250 ;
        RECT 30.145 -3.250 30.445 -3.060 ;
        RECT 31.555 -3.250 31.855 -2.880 ;
        RECT 30.145 -3.430 30.665 -3.250 ;
        RECT 31.335 -3.430 31.855 -3.250 ;
        RECT 32.145 -3.250 32.445 -3.060 ;
        RECT 33.555 -3.250 33.855 -2.880 ;
        RECT 32.145 -3.430 32.665 -3.250 ;
        RECT 33.335 -3.430 33.855 -3.250 ;
        RECT 34.145 -3.250 34.445 -3.060 ;
        RECT 35.555 -3.250 35.855 -2.880 ;
        RECT 34.145 -3.430 34.665 -3.250 ;
        RECT 35.335 -3.430 35.855 -3.250 ;
        RECT 36.145 -3.250 36.445 -3.060 ;
        RECT 37.555 -3.250 37.855 -2.880 ;
        RECT 36.145 -3.430 36.665 -3.250 ;
        RECT 37.335 -3.430 37.855 -3.250 ;
        RECT 38.145 -3.250 38.445 -3.060 ;
        RECT 39.555 -3.250 39.855 -2.880 ;
        RECT 38.145 -3.430 38.665 -3.250 ;
        RECT 39.335 -3.430 39.855 -3.250 ;
        RECT 40.145 -3.250 40.445 -3.060 ;
        RECT 41.555 -3.250 41.855 -2.880 ;
        RECT 40.145 -3.430 40.665 -3.250 ;
        RECT 41.335 -3.430 41.855 -3.250 ;
        RECT 42.145 -3.250 42.445 -3.060 ;
        RECT 43.555 -3.250 43.855 -2.880 ;
        RECT 42.145 -3.430 42.665 -3.250 ;
        RECT 43.335 -3.430 43.855 -3.250 ;
        RECT 44.145 -3.250 44.445 -3.060 ;
        RECT 45.555 -3.250 45.855 -2.880 ;
        RECT 44.145 -3.430 44.665 -3.250 ;
        RECT 45.335 -3.430 45.855 -3.250 ;
        RECT 46.145 -3.250 46.445 -3.060 ;
        RECT 47.555 -3.250 47.855 -2.880 ;
        RECT 46.145 -3.430 46.665 -3.250 ;
        RECT 47.335 -3.430 47.855 -3.250 ;
        RECT 48.145 -3.250 48.445 -3.060 ;
        RECT 49.555 -3.250 49.855 -2.880 ;
        RECT 48.145 -3.430 48.665 -3.250 ;
        RECT 49.335 -3.430 49.855 -3.250 ;
        RECT 50.145 -3.250 50.445 -3.060 ;
        RECT 51.555 -3.250 51.855 -2.880 ;
        RECT 50.145 -3.430 50.665 -3.250 ;
        RECT 51.335 -3.430 51.855 -3.250 ;
        RECT 52.145 -3.250 52.445 -3.060 ;
        RECT 53.555 -3.250 53.855 -2.880 ;
        RECT 52.145 -3.430 52.665 -3.250 ;
        RECT 53.335 -3.430 53.855 -3.250 ;
        RECT 54.145 -3.250 54.445 -3.060 ;
        RECT 55.555 -3.250 55.855 -2.880 ;
        RECT 54.145 -3.430 54.665 -3.250 ;
        RECT 55.335 -3.430 55.855 -3.250 ;
        RECT 56.145 -3.250 56.445 -3.060 ;
        RECT 57.555 -3.250 57.855 -2.880 ;
        RECT 56.145 -3.430 56.665 -3.250 ;
        RECT 57.335 -3.430 57.855 -3.250 ;
        RECT 58.145 -3.250 58.445 -3.060 ;
        RECT 59.555 -3.250 59.855 -2.880 ;
        RECT 58.145 -3.430 58.665 -3.250 ;
        RECT 59.335 -3.430 59.855 -3.250 ;
        RECT 60.145 -3.250 60.445 -3.060 ;
        RECT 61.555 -3.250 61.855 -2.880 ;
        RECT 60.145 -3.430 60.665 -3.250 ;
        RECT 61.335 -3.430 61.855 -3.250 ;
        RECT 62.145 -3.250 62.445 -3.060 ;
        RECT 63.555 -3.250 63.855 -2.880 ;
        RECT 62.145 -3.430 62.665 -3.250 ;
        RECT 63.335 -3.430 63.855 -3.250 ;
        RECT 64.145 -3.250 64.445 -3.060 ;
        RECT 65.555 -3.250 65.855 -2.880 ;
        RECT 64.145 -3.430 64.665 -3.250 ;
        RECT 65.335 -3.430 65.855 -3.250 ;
        RECT 66.145 -3.250 66.445 -3.060 ;
        RECT 67.555 -3.250 67.855 -2.880 ;
        RECT 66.145 -3.430 66.665 -3.250 ;
        RECT 67.335 -3.430 67.855 -3.250 ;
        RECT 68.145 -3.250 68.445 -3.060 ;
        RECT 69.555 -3.250 69.855 -2.880 ;
        RECT 68.145 -3.430 68.665 -3.250 ;
        RECT 69.335 -3.430 69.855 -3.250 ;
        RECT 70.145 -3.250 70.445 -3.060 ;
        RECT 71.555 -3.250 71.855 -2.880 ;
        RECT 70.145 -3.430 70.665 -3.250 ;
        RECT 71.335 -3.430 71.855 -3.250 ;
        RECT 72.145 -3.250 72.445 -3.060 ;
        RECT 73.555 -3.250 73.855 -2.880 ;
        RECT 72.145 -3.430 72.665 -3.250 ;
        RECT 73.335 -3.430 73.855 -3.250 ;
        RECT 74.145 -3.250 74.445 -3.060 ;
        RECT 75.555 -3.250 75.855 -2.880 ;
        RECT 74.145 -3.430 74.665 -3.250 ;
        RECT 75.335 -3.430 75.855 -3.250 ;
        RECT 76.145 -3.250 76.445 -3.060 ;
        RECT 77.555 -3.250 77.855 -2.880 ;
        RECT 76.145 -3.430 76.665 -3.250 ;
        RECT 77.335 -3.430 77.855 -3.250 ;
        RECT 78.145 -3.250 78.445 -3.060 ;
        RECT 79.555 -3.250 79.855 -2.880 ;
        RECT 78.145 -3.430 78.665 -3.250 ;
        RECT 79.335 -3.430 79.855 -3.250 ;
        RECT 80.145 -3.250 80.445 -3.060 ;
        RECT 81.555 -3.250 81.855 -2.880 ;
        RECT 80.145 -3.430 80.665 -3.250 ;
        RECT 81.335 -3.430 81.855 -3.250 ;
        RECT 82.145 -3.250 82.445 -3.060 ;
        RECT 83.555 -3.250 83.855 -2.880 ;
        RECT 82.145 -3.430 82.665 -3.250 ;
        RECT 83.335 -3.430 83.855 -3.250 ;
        RECT 84.145 -3.250 84.445 -3.060 ;
        RECT 85.555 -3.250 85.855 -2.880 ;
        RECT 84.145 -3.430 84.665 -3.250 ;
        RECT 85.335 -3.430 85.855 -3.250 ;
        RECT 86.145 -3.250 86.445 -3.060 ;
        RECT 87.555 -3.250 87.855 -2.880 ;
        RECT 86.145 -3.430 86.665 -3.250 ;
        RECT 87.335 -3.430 87.855 -3.250 ;
        RECT 88.145 -3.250 88.445 -3.060 ;
        RECT 89.555 -3.250 89.855 -2.880 ;
        RECT 88.145 -3.430 88.665 -3.250 ;
        RECT 89.335 -3.430 89.855 -3.250 ;
        RECT 90.145 -3.250 90.445 -3.060 ;
        RECT 91.555 -3.250 91.855 -2.880 ;
        RECT 90.145 -3.430 90.665 -3.250 ;
        RECT 91.335 -3.430 91.855 -3.250 ;
        RECT 92.145 -3.250 92.445 -3.060 ;
        RECT 93.555 -3.250 93.855 -2.880 ;
        RECT 92.145 -3.430 92.665 -3.250 ;
        RECT 93.335 -3.430 93.855 -3.250 ;
        RECT 94.145 -3.250 94.445 -3.060 ;
        RECT 95.555 -3.250 95.855 -2.880 ;
        RECT 94.145 -3.430 94.665 -3.250 ;
        RECT 95.335 -3.430 95.855 -3.250 ;
        RECT 96.145 -3.250 96.445 -3.060 ;
        RECT 97.555 -3.250 97.855 -2.880 ;
        RECT 96.145 -3.430 96.665 -3.250 ;
        RECT 97.335 -3.430 97.855 -3.250 ;
        RECT 98.145 -3.250 98.445 -3.060 ;
        RECT 99.555 -3.250 99.855 -2.880 ;
        RECT 98.145 -3.430 98.665 -3.250 ;
        RECT 99.335 -3.430 99.855 -3.250 ;
        RECT 100.145 -3.250 100.445 -3.060 ;
        RECT 101.555 -3.250 101.855 -2.880 ;
        RECT 100.145 -3.430 100.665 -3.250 ;
        RECT 101.335 -3.430 101.855 -3.250 ;
        RECT 102.145 -3.250 102.445 -3.060 ;
        RECT 103.555 -3.250 103.855 -2.880 ;
        RECT 102.145 -3.430 102.665 -3.250 ;
        RECT 103.335 -3.430 103.855 -3.250 ;
        RECT 104.145 -3.250 104.445 -3.060 ;
        RECT 105.555 -3.250 105.855 -2.880 ;
        RECT 104.145 -3.430 104.665 -3.250 ;
        RECT 105.335 -3.430 105.855 -3.250 ;
        RECT 106.145 -3.250 106.445 -3.060 ;
        RECT 107.555 -3.250 107.855 -2.880 ;
        RECT 106.145 -3.430 106.665 -3.250 ;
        RECT 107.335 -3.430 107.855 -3.250 ;
        RECT 108.145 -3.250 108.445 -3.060 ;
        RECT 109.555 -3.250 109.855 -2.880 ;
        RECT 108.145 -3.430 108.665 -3.250 ;
        RECT 109.335 -3.430 109.855 -3.250 ;
        RECT 110.145 -3.250 110.445 -3.060 ;
        RECT 111.555 -3.250 111.855 -2.880 ;
        RECT 110.145 -3.430 110.665 -3.250 ;
        RECT 111.335 -3.430 111.855 -3.250 ;
        RECT 112.145 -3.250 112.445 -3.060 ;
        RECT 113.555 -3.250 113.855 -2.880 ;
        RECT 112.145 -3.430 112.665 -3.250 ;
        RECT 113.335 -3.430 113.855 -3.250 ;
        RECT 114.145 -3.250 114.445 -3.060 ;
        RECT 115.555 -3.250 115.855 -2.880 ;
        RECT 114.145 -3.430 114.665 -3.250 ;
        RECT 115.335 -3.430 115.855 -3.250 ;
        RECT 116.145 -3.250 116.445 -3.060 ;
        RECT 117.555 -3.250 117.855 -2.880 ;
        RECT 116.145 -3.430 116.665 -3.250 ;
        RECT 117.335 -3.430 117.855 -3.250 ;
        RECT 118.145 -3.250 118.445 -3.060 ;
        RECT 119.555 -3.250 119.855 -2.880 ;
        RECT 118.145 -3.430 118.665 -3.250 ;
        RECT 119.335 -3.430 119.855 -3.250 ;
        RECT 120.145 -3.250 120.445 -3.060 ;
        RECT 121.555 -3.250 121.855 -2.880 ;
        RECT 120.145 -3.430 120.665 -3.250 ;
        RECT 121.335 -3.430 121.855 -3.250 ;
        RECT 122.145 -3.250 122.445 -3.060 ;
        RECT 123.555 -3.250 123.855 -2.880 ;
        RECT 122.145 -3.430 122.665 -3.250 ;
        RECT 123.335 -3.430 123.855 -3.250 ;
        RECT 124.145 -3.250 124.445 -3.060 ;
        RECT 125.555 -3.250 125.855 -2.880 ;
        RECT 124.145 -3.430 124.665 -3.250 ;
        RECT 125.335 -3.430 125.855 -3.250 ;
        RECT 126.145 -3.250 126.445 -3.060 ;
        RECT 127.555 -3.250 127.855 -2.880 ;
        RECT 126.145 -3.430 126.665 -3.250 ;
        RECT 127.335 -3.430 127.855 -3.250 ;
        RECT 128.145 -3.250 128.445 -3.060 ;
        RECT 129.555 -3.250 129.855 -2.880 ;
        RECT 128.145 -3.430 128.665 -3.250 ;
        RECT 129.335 -3.430 129.855 -3.250 ;
        RECT 130.145 -3.250 130.445 -3.060 ;
        RECT 130.145 -3.430 130.665 -3.250 ;
        RECT -0.665 -3.760 -0.145 -3.580 ;
        RECT 0.145 -3.760 0.665 -3.580 ;
        RECT 1.335 -3.760 1.855 -3.580 ;
        RECT 2.145 -3.760 2.665 -3.580 ;
        RECT 3.335 -3.760 3.855 -3.580 ;
        RECT 4.145 -3.760 4.665 -3.580 ;
        RECT 5.335 -3.760 5.855 -3.580 ;
        RECT 6.145 -3.760 6.665 -3.580 ;
        RECT 7.335 -3.760 7.855 -3.580 ;
        RECT 8.145 -3.760 8.665 -3.580 ;
        RECT 9.335 -3.760 9.855 -3.580 ;
        RECT 10.145 -3.760 10.665 -3.580 ;
        RECT 11.335 -3.760 11.855 -3.580 ;
        RECT 12.145 -3.760 12.665 -3.580 ;
        RECT 13.335 -3.760 13.855 -3.580 ;
        RECT 14.145 -3.760 14.665 -3.580 ;
        RECT 15.335 -3.760 15.855 -3.580 ;
        RECT 16.145 -3.760 16.665 -3.580 ;
        RECT 17.335 -3.760 17.855 -3.580 ;
        RECT 18.145 -3.760 18.665 -3.580 ;
        RECT 19.335 -3.760 19.855 -3.580 ;
        RECT 20.145 -3.760 20.665 -3.580 ;
        RECT 21.335 -3.760 21.855 -3.580 ;
        RECT 22.145 -3.760 22.665 -3.580 ;
        RECT 23.335 -3.760 23.855 -3.580 ;
        RECT 24.145 -3.760 24.665 -3.580 ;
        RECT 25.335 -3.760 25.855 -3.580 ;
        RECT 26.145 -3.760 26.665 -3.580 ;
        RECT 27.335 -3.760 27.855 -3.580 ;
        RECT 28.145 -3.760 28.665 -3.580 ;
        RECT 29.335 -3.760 29.855 -3.580 ;
        RECT 30.145 -3.760 30.665 -3.580 ;
        RECT 31.335 -3.760 31.855 -3.580 ;
        RECT 32.145 -3.760 32.665 -3.580 ;
        RECT 33.335 -3.760 33.855 -3.580 ;
        RECT 34.145 -3.760 34.665 -3.580 ;
        RECT 35.335 -3.760 35.855 -3.580 ;
        RECT 36.145 -3.760 36.665 -3.580 ;
        RECT 37.335 -3.760 37.855 -3.580 ;
        RECT 38.145 -3.760 38.665 -3.580 ;
        RECT 39.335 -3.760 39.855 -3.580 ;
        RECT 40.145 -3.760 40.665 -3.580 ;
        RECT 41.335 -3.760 41.855 -3.580 ;
        RECT 42.145 -3.760 42.665 -3.580 ;
        RECT 43.335 -3.760 43.855 -3.580 ;
        RECT 44.145 -3.760 44.665 -3.580 ;
        RECT 45.335 -3.760 45.855 -3.580 ;
        RECT 46.145 -3.760 46.665 -3.580 ;
        RECT 47.335 -3.760 47.855 -3.580 ;
        RECT 48.145 -3.760 48.665 -3.580 ;
        RECT 49.335 -3.760 49.855 -3.580 ;
        RECT 50.145 -3.760 50.665 -3.580 ;
        RECT 51.335 -3.760 51.855 -3.580 ;
        RECT 52.145 -3.760 52.665 -3.580 ;
        RECT 53.335 -3.760 53.855 -3.580 ;
        RECT 54.145 -3.760 54.665 -3.580 ;
        RECT 55.335 -3.760 55.855 -3.580 ;
        RECT 56.145 -3.760 56.665 -3.580 ;
        RECT 57.335 -3.760 57.855 -3.580 ;
        RECT 58.145 -3.760 58.665 -3.580 ;
        RECT 59.335 -3.760 59.855 -3.580 ;
        RECT 60.145 -3.760 60.665 -3.580 ;
        RECT 61.335 -3.760 61.855 -3.580 ;
        RECT 62.145 -3.760 62.665 -3.580 ;
        RECT 63.335 -3.760 63.855 -3.580 ;
        RECT 64.145 -3.760 64.665 -3.580 ;
        RECT 65.335 -3.760 65.855 -3.580 ;
        RECT 66.145 -3.760 66.665 -3.580 ;
        RECT 67.335 -3.760 67.855 -3.580 ;
        RECT 68.145 -3.760 68.665 -3.580 ;
        RECT 69.335 -3.760 69.855 -3.580 ;
        RECT 70.145 -3.760 70.665 -3.580 ;
        RECT 71.335 -3.760 71.855 -3.580 ;
        RECT 72.145 -3.760 72.665 -3.580 ;
        RECT 73.335 -3.760 73.855 -3.580 ;
        RECT 74.145 -3.760 74.665 -3.580 ;
        RECT 75.335 -3.760 75.855 -3.580 ;
        RECT 76.145 -3.760 76.665 -3.580 ;
        RECT 77.335 -3.760 77.855 -3.580 ;
        RECT 78.145 -3.760 78.665 -3.580 ;
        RECT 79.335 -3.760 79.855 -3.580 ;
        RECT 80.145 -3.760 80.665 -3.580 ;
        RECT 81.335 -3.760 81.855 -3.580 ;
        RECT 82.145 -3.760 82.665 -3.580 ;
        RECT 83.335 -3.760 83.855 -3.580 ;
        RECT 84.145 -3.760 84.665 -3.580 ;
        RECT 85.335 -3.760 85.855 -3.580 ;
        RECT 86.145 -3.760 86.665 -3.580 ;
        RECT 87.335 -3.760 87.855 -3.580 ;
        RECT 88.145 -3.760 88.665 -3.580 ;
        RECT 89.335 -3.760 89.855 -3.580 ;
        RECT 90.145 -3.760 90.665 -3.580 ;
        RECT 91.335 -3.760 91.855 -3.580 ;
        RECT 92.145 -3.760 92.665 -3.580 ;
        RECT 93.335 -3.760 93.855 -3.580 ;
        RECT 94.145 -3.760 94.665 -3.580 ;
        RECT 95.335 -3.760 95.855 -3.580 ;
        RECT 96.145 -3.760 96.665 -3.580 ;
        RECT 97.335 -3.760 97.855 -3.580 ;
        RECT 98.145 -3.760 98.665 -3.580 ;
        RECT 99.335 -3.760 99.855 -3.580 ;
        RECT 100.145 -3.760 100.665 -3.580 ;
        RECT 101.335 -3.760 101.855 -3.580 ;
        RECT 102.145 -3.760 102.665 -3.580 ;
        RECT 103.335 -3.760 103.855 -3.580 ;
        RECT 104.145 -3.760 104.665 -3.580 ;
        RECT 105.335 -3.760 105.855 -3.580 ;
        RECT 106.145 -3.760 106.665 -3.580 ;
        RECT 107.335 -3.760 107.855 -3.580 ;
        RECT 108.145 -3.760 108.665 -3.580 ;
        RECT 109.335 -3.760 109.855 -3.580 ;
        RECT 110.145 -3.760 110.665 -3.580 ;
        RECT 111.335 -3.760 111.855 -3.580 ;
        RECT 112.145 -3.760 112.665 -3.580 ;
        RECT 113.335 -3.760 113.855 -3.580 ;
        RECT 114.145 -3.760 114.665 -3.580 ;
        RECT 115.335 -3.760 115.855 -3.580 ;
        RECT 116.145 -3.760 116.665 -3.580 ;
        RECT 117.335 -3.760 117.855 -3.580 ;
        RECT 118.145 -3.760 118.665 -3.580 ;
        RECT 119.335 -3.760 119.855 -3.580 ;
        RECT 120.145 -3.760 120.665 -3.580 ;
        RECT 121.335 -3.760 121.855 -3.580 ;
        RECT 122.145 -3.760 122.665 -3.580 ;
        RECT 123.335 -3.760 123.855 -3.580 ;
        RECT 124.145 -3.760 124.665 -3.580 ;
        RECT 125.335 -3.760 125.855 -3.580 ;
        RECT 126.145 -3.760 126.665 -3.580 ;
        RECT 127.335 -3.760 127.855 -3.580 ;
        RECT 128.145 -3.760 128.665 -3.580 ;
        RECT 129.335 -3.760 129.855 -3.580 ;
        RECT 130.145 -3.760 130.665 -3.580 ;
      LAYER Metal1 ;
        RECT -0.825 18.370 -0.665 20.480 ;
        RECT -0.080 20.220 0.080 20.780 ;
        RECT 0.665 19.660 0.825 20.480 ;
        RECT -0.425 19.500 0.825 19.660 ;
        RECT -0.420 18.560 -0.130 18.850 ;
        RECT 0.130 18.560 0.420 18.850 ;
        RECT -0.420 18.490 -0.260 18.560 ;
        RECT 0.260 18.490 0.420 18.560 ;
        RECT -0.890 18.080 -0.600 18.370 ;
        RECT -0.080 17.700 0.080 18.380 ;
        RECT 0.665 18.370 0.825 19.500 ;
        RECT 1.175 18.370 1.335 20.480 ;
        RECT 1.920 20.220 2.080 20.780 ;
        RECT 2.665 19.660 2.825 20.480 ;
        RECT 1.575 19.500 2.825 19.660 ;
        RECT 1.580 18.560 1.870 18.850 ;
        RECT 2.130 18.560 2.420 18.850 ;
        RECT 1.580 18.490 1.740 18.560 ;
        RECT 2.260 18.490 2.420 18.560 ;
        RECT 0.600 18.080 0.890 18.370 ;
        RECT 1.110 18.080 1.400 18.370 ;
        RECT 1.920 17.700 2.080 18.380 ;
        RECT 2.665 18.370 2.825 19.500 ;
        RECT 3.175 18.370 3.335 20.480 ;
        RECT 3.920 20.220 4.080 20.780 ;
        RECT 4.665 19.660 4.825 20.480 ;
        RECT 3.575 19.500 4.825 19.660 ;
        RECT 3.580 18.560 3.870 18.850 ;
        RECT 4.130 18.560 4.420 18.850 ;
        RECT 3.580 18.490 3.740 18.560 ;
        RECT 4.260 18.490 4.420 18.560 ;
        RECT 2.600 18.080 2.890 18.370 ;
        RECT 3.110 18.080 3.400 18.370 ;
        RECT 3.920 17.700 4.080 18.380 ;
        RECT 4.665 18.370 4.825 19.500 ;
        RECT 5.175 18.370 5.335 20.480 ;
        RECT 5.920 20.220 6.080 20.780 ;
        RECT 6.665 19.660 6.825 20.480 ;
        RECT 5.575 19.500 6.825 19.660 ;
        RECT 5.580 18.560 5.870 18.850 ;
        RECT 6.130 18.560 6.420 18.850 ;
        RECT 5.580 18.490 5.740 18.560 ;
        RECT 6.260 18.490 6.420 18.560 ;
        RECT 4.600 18.080 4.890 18.370 ;
        RECT 5.110 18.080 5.400 18.370 ;
        RECT 5.920 17.700 6.080 18.380 ;
        RECT 6.665 18.370 6.825 19.500 ;
        RECT 7.175 18.370 7.335 20.480 ;
        RECT 7.920 20.220 8.080 20.780 ;
        RECT 8.665 19.660 8.825 20.480 ;
        RECT 7.575 19.500 8.825 19.660 ;
        RECT 7.580 18.560 7.870 18.850 ;
        RECT 8.130 18.560 8.420 18.850 ;
        RECT 7.580 18.490 7.740 18.560 ;
        RECT 8.260 18.490 8.420 18.560 ;
        RECT 6.600 18.080 6.890 18.370 ;
        RECT 7.110 18.080 7.400 18.370 ;
        RECT 7.920 17.700 8.080 18.380 ;
        RECT 8.665 18.370 8.825 19.500 ;
        RECT 9.175 18.370 9.335 20.480 ;
        RECT 9.920 20.220 10.080 20.780 ;
        RECT 10.665 19.660 10.825 20.480 ;
        RECT 9.575 19.500 10.825 19.660 ;
        RECT 9.580 18.560 9.870 18.850 ;
        RECT 10.130 18.560 10.420 18.850 ;
        RECT 9.580 18.490 9.740 18.560 ;
        RECT 10.260 18.490 10.420 18.560 ;
        RECT 8.600 18.080 8.890 18.370 ;
        RECT 9.110 18.080 9.400 18.370 ;
        RECT 9.920 17.700 10.080 18.380 ;
        RECT 10.665 18.370 10.825 19.500 ;
        RECT 11.175 18.370 11.335 20.480 ;
        RECT 11.920 20.220 12.080 20.780 ;
        RECT 12.665 19.660 12.825 20.480 ;
        RECT 11.575 19.500 12.825 19.660 ;
        RECT 11.580 18.560 11.870 18.850 ;
        RECT 12.130 18.560 12.420 18.850 ;
        RECT 11.580 18.490 11.740 18.560 ;
        RECT 12.260 18.490 12.420 18.560 ;
        RECT 10.600 18.080 10.890 18.370 ;
        RECT 11.110 18.080 11.400 18.370 ;
        RECT 11.920 17.700 12.080 18.380 ;
        RECT 12.665 18.370 12.825 19.500 ;
        RECT 13.175 18.370 13.335 20.480 ;
        RECT 13.920 20.220 14.080 20.780 ;
        RECT 14.665 19.660 14.825 20.480 ;
        RECT 13.575 19.500 14.825 19.660 ;
        RECT 13.580 18.560 13.870 18.850 ;
        RECT 14.130 18.560 14.420 18.850 ;
        RECT 13.580 18.490 13.740 18.560 ;
        RECT 14.260 18.490 14.420 18.560 ;
        RECT 12.600 18.080 12.890 18.370 ;
        RECT 13.110 18.080 13.400 18.370 ;
        RECT 13.920 17.700 14.080 18.380 ;
        RECT 14.665 18.370 14.825 19.500 ;
        RECT 15.175 18.370 15.335 20.480 ;
        RECT 15.920 20.220 16.080 20.780 ;
        RECT 16.665 19.660 16.825 20.480 ;
        RECT 15.575 19.500 16.825 19.660 ;
        RECT 15.580 18.560 15.870 18.850 ;
        RECT 16.130 18.560 16.420 18.850 ;
        RECT 15.580 18.490 15.740 18.560 ;
        RECT 16.260 18.490 16.420 18.560 ;
        RECT 14.600 18.080 14.890 18.370 ;
        RECT 15.110 18.080 15.400 18.370 ;
        RECT 15.920 17.700 16.080 18.380 ;
        RECT 16.665 18.370 16.825 19.500 ;
        RECT 17.175 18.370 17.335 20.480 ;
        RECT 17.920 20.220 18.080 20.780 ;
        RECT 18.665 19.660 18.825 20.480 ;
        RECT 17.575 19.500 18.825 19.660 ;
        RECT 17.580 18.560 17.870 18.850 ;
        RECT 18.130 18.560 18.420 18.850 ;
        RECT 17.580 18.490 17.740 18.560 ;
        RECT 18.260 18.490 18.420 18.560 ;
        RECT 16.600 18.080 16.890 18.370 ;
        RECT 17.110 18.080 17.400 18.370 ;
        RECT 17.920 17.700 18.080 18.380 ;
        RECT 18.665 18.370 18.825 19.500 ;
        RECT 19.175 18.370 19.335 20.480 ;
        RECT 19.920 20.220 20.080 20.780 ;
        RECT 20.665 19.660 20.825 20.480 ;
        RECT 19.575 19.500 20.825 19.660 ;
        RECT 19.580 18.560 19.870 18.850 ;
        RECT 20.130 18.560 20.420 18.850 ;
        RECT 19.580 18.490 19.740 18.560 ;
        RECT 20.260 18.490 20.420 18.560 ;
        RECT 18.600 18.080 18.890 18.370 ;
        RECT 19.110 18.080 19.400 18.370 ;
        RECT 19.920 17.700 20.080 18.380 ;
        RECT 20.665 18.370 20.825 19.500 ;
        RECT 21.175 18.370 21.335 20.480 ;
        RECT 21.920 20.220 22.080 20.780 ;
        RECT 22.665 19.660 22.825 20.480 ;
        RECT 21.575 19.500 22.825 19.660 ;
        RECT 21.580 18.560 21.870 18.850 ;
        RECT 22.130 18.560 22.420 18.850 ;
        RECT 21.580 18.490 21.740 18.560 ;
        RECT 22.260 18.490 22.420 18.560 ;
        RECT 20.600 18.080 20.890 18.370 ;
        RECT 21.110 18.080 21.400 18.370 ;
        RECT 21.920 17.700 22.080 18.380 ;
        RECT 22.665 18.370 22.825 19.500 ;
        RECT 23.175 18.370 23.335 20.480 ;
        RECT 23.920 20.220 24.080 20.780 ;
        RECT 24.665 19.660 24.825 20.480 ;
        RECT 23.575 19.500 24.825 19.660 ;
        RECT 23.580 18.560 23.870 18.850 ;
        RECT 24.130 18.560 24.420 18.850 ;
        RECT 23.580 18.490 23.740 18.560 ;
        RECT 24.260 18.490 24.420 18.560 ;
        RECT 22.600 18.080 22.890 18.370 ;
        RECT 23.110 18.080 23.400 18.370 ;
        RECT 23.920 17.700 24.080 18.380 ;
        RECT 24.665 18.370 24.825 19.500 ;
        RECT 25.175 18.370 25.335 20.480 ;
        RECT 25.920 20.220 26.080 20.780 ;
        RECT 26.665 19.660 26.825 20.480 ;
        RECT 25.575 19.500 26.825 19.660 ;
        RECT 25.580 18.560 25.870 18.850 ;
        RECT 26.130 18.560 26.420 18.850 ;
        RECT 25.580 18.490 25.740 18.560 ;
        RECT 26.260 18.490 26.420 18.560 ;
        RECT 24.600 18.080 24.890 18.370 ;
        RECT 25.110 18.080 25.400 18.370 ;
        RECT 25.920 17.700 26.080 18.380 ;
        RECT 26.665 18.370 26.825 19.500 ;
        RECT 27.175 18.370 27.335 20.480 ;
        RECT 27.920 20.220 28.080 20.780 ;
        RECT 28.665 19.660 28.825 20.480 ;
        RECT 27.575 19.500 28.825 19.660 ;
        RECT 27.580 18.560 27.870 18.850 ;
        RECT 28.130 18.560 28.420 18.850 ;
        RECT 27.580 18.490 27.740 18.560 ;
        RECT 28.260 18.490 28.420 18.560 ;
        RECT 26.600 18.080 26.890 18.370 ;
        RECT 27.110 18.080 27.400 18.370 ;
        RECT 27.920 17.700 28.080 18.380 ;
        RECT 28.665 18.370 28.825 19.500 ;
        RECT 29.175 18.370 29.335 20.480 ;
        RECT 29.920 20.220 30.080 20.780 ;
        RECT 30.665 19.660 30.825 20.480 ;
        RECT 29.575 19.500 30.825 19.660 ;
        RECT 29.580 18.560 29.870 18.850 ;
        RECT 30.130 18.560 30.420 18.850 ;
        RECT 29.580 18.490 29.740 18.560 ;
        RECT 30.260 18.490 30.420 18.560 ;
        RECT 28.600 18.080 28.890 18.370 ;
        RECT 29.110 18.080 29.400 18.370 ;
        RECT 29.920 17.700 30.080 18.380 ;
        RECT 30.665 18.370 30.825 19.500 ;
        RECT 31.175 18.370 31.335 20.480 ;
        RECT 31.920 20.220 32.080 20.780 ;
        RECT 32.665 19.660 32.825 20.480 ;
        RECT 31.575 19.500 32.825 19.660 ;
        RECT 31.580 18.560 31.870 18.850 ;
        RECT 32.130 18.560 32.420 18.850 ;
        RECT 31.580 18.490 31.740 18.560 ;
        RECT 32.260 18.490 32.420 18.560 ;
        RECT 30.600 18.080 30.890 18.370 ;
        RECT 31.110 18.080 31.400 18.370 ;
        RECT 31.920 17.700 32.080 18.380 ;
        RECT 32.665 18.370 32.825 19.500 ;
        RECT 33.175 18.370 33.335 20.480 ;
        RECT 33.920 20.220 34.080 20.780 ;
        RECT 34.665 19.660 34.825 20.480 ;
        RECT 33.575 19.500 34.825 19.660 ;
        RECT 33.580 18.560 33.870 18.850 ;
        RECT 34.130 18.560 34.420 18.850 ;
        RECT 33.580 18.490 33.740 18.560 ;
        RECT 34.260 18.490 34.420 18.560 ;
        RECT 32.600 18.080 32.890 18.370 ;
        RECT 33.110 18.080 33.400 18.370 ;
        RECT 33.920 17.700 34.080 18.380 ;
        RECT 34.665 18.370 34.825 19.500 ;
        RECT 35.175 18.370 35.335 20.480 ;
        RECT 35.920 20.220 36.080 20.780 ;
        RECT 36.665 19.660 36.825 20.480 ;
        RECT 35.575 19.500 36.825 19.660 ;
        RECT 35.580 18.560 35.870 18.850 ;
        RECT 36.130 18.560 36.420 18.850 ;
        RECT 35.580 18.490 35.740 18.560 ;
        RECT 36.260 18.490 36.420 18.560 ;
        RECT 34.600 18.080 34.890 18.370 ;
        RECT 35.110 18.080 35.400 18.370 ;
        RECT 35.920 17.700 36.080 18.380 ;
        RECT 36.665 18.370 36.825 19.500 ;
        RECT 37.175 18.370 37.335 20.480 ;
        RECT 37.920 20.220 38.080 20.780 ;
        RECT 38.665 19.660 38.825 20.480 ;
        RECT 37.575 19.500 38.825 19.660 ;
        RECT 37.580 18.560 37.870 18.850 ;
        RECT 38.130 18.560 38.420 18.850 ;
        RECT 37.580 18.490 37.740 18.560 ;
        RECT 38.260 18.490 38.420 18.560 ;
        RECT 36.600 18.080 36.890 18.370 ;
        RECT 37.110 18.080 37.400 18.370 ;
        RECT 37.920 17.700 38.080 18.380 ;
        RECT 38.665 18.370 38.825 19.500 ;
        RECT 39.175 18.370 39.335 20.480 ;
        RECT 39.920 20.220 40.080 20.780 ;
        RECT 40.665 19.660 40.825 20.480 ;
        RECT 39.575 19.500 40.825 19.660 ;
        RECT 39.580 18.560 39.870 18.850 ;
        RECT 40.130 18.560 40.420 18.850 ;
        RECT 39.580 18.490 39.740 18.560 ;
        RECT 40.260 18.490 40.420 18.560 ;
        RECT 38.600 18.080 38.890 18.370 ;
        RECT 39.110 18.080 39.400 18.370 ;
        RECT 39.920 17.700 40.080 18.380 ;
        RECT 40.665 18.370 40.825 19.500 ;
        RECT 41.175 18.370 41.335 20.480 ;
        RECT 41.920 20.220 42.080 20.780 ;
        RECT 42.665 19.660 42.825 20.480 ;
        RECT 41.575 19.500 42.825 19.660 ;
        RECT 41.580 18.560 41.870 18.850 ;
        RECT 42.130 18.560 42.420 18.850 ;
        RECT 41.580 18.490 41.740 18.560 ;
        RECT 42.260 18.490 42.420 18.560 ;
        RECT 40.600 18.080 40.890 18.370 ;
        RECT 41.110 18.080 41.400 18.370 ;
        RECT 41.920 17.700 42.080 18.380 ;
        RECT 42.665 18.370 42.825 19.500 ;
        RECT 43.175 18.370 43.335 20.480 ;
        RECT 43.920 20.220 44.080 20.780 ;
        RECT 44.665 19.660 44.825 20.480 ;
        RECT 43.575 19.500 44.825 19.660 ;
        RECT 43.580 18.560 43.870 18.850 ;
        RECT 44.130 18.560 44.420 18.850 ;
        RECT 43.580 18.490 43.740 18.560 ;
        RECT 44.260 18.490 44.420 18.560 ;
        RECT 42.600 18.080 42.890 18.370 ;
        RECT 43.110 18.080 43.400 18.370 ;
        RECT 43.920 17.700 44.080 18.380 ;
        RECT 44.665 18.370 44.825 19.500 ;
        RECT 45.175 18.370 45.335 20.480 ;
        RECT 45.920 20.220 46.080 20.780 ;
        RECT 46.665 19.660 46.825 20.480 ;
        RECT 45.575 19.500 46.825 19.660 ;
        RECT 45.580 18.560 45.870 18.850 ;
        RECT 46.130 18.560 46.420 18.850 ;
        RECT 45.580 18.490 45.740 18.560 ;
        RECT 46.260 18.490 46.420 18.560 ;
        RECT 44.600 18.080 44.890 18.370 ;
        RECT 45.110 18.080 45.400 18.370 ;
        RECT 45.920 17.700 46.080 18.380 ;
        RECT 46.665 18.370 46.825 19.500 ;
        RECT 47.175 18.370 47.335 20.480 ;
        RECT 47.920 20.220 48.080 20.780 ;
        RECT 48.665 19.660 48.825 20.480 ;
        RECT 47.575 19.500 48.825 19.660 ;
        RECT 47.580 18.560 47.870 18.850 ;
        RECT 48.130 18.560 48.420 18.850 ;
        RECT 47.580 18.490 47.740 18.560 ;
        RECT 48.260 18.490 48.420 18.560 ;
        RECT 46.600 18.080 46.890 18.370 ;
        RECT 47.110 18.080 47.400 18.370 ;
        RECT 47.920 17.700 48.080 18.380 ;
        RECT 48.665 18.370 48.825 19.500 ;
        RECT 49.175 18.370 49.335 20.480 ;
        RECT 49.920 20.220 50.080 20.780 ;
        RECT 50.665 19.660 50.825 20.480 ;
        RECT 49.575 19.500 50.825 19.660 ;
        RECT 49.580 18.560 49.870 18.850 ;
        RECT 50.130 18.560 50.420 18.850 ;
        RECT 49.580 18.490 49.740 18.560 ;
        RECT 50.260 18.490 50.420 18.560 ;
        RECT 48.600 18.080 48.890 18.370 ;
        RECT 49.110 18.080 49.400 18.370 ;
        RECT 49.920 17.700 50.080 18.380 ;
        RECT 50.665 18.370 50.825 19.500 ;
        RECT 51.175 18.370 51.335 20.480 ;
        RECT 51.920 20.220 52.080 20.780 ;
        RECT 52.665 19.660 52.825 20.480 ;
        RECT 51.575 19.500 52.825 19.660 ;
        RECT 51.580 18.560 51.870 18.850 ;
        RECT 52.130 18.560 52.420 18.850 ;
        RECT 51.580 18.490 51.740 18.560 ;
        RECT 52.260 18.490 52.420 18.560 ;
        RECT 50.600 18.080 50.890 18.370 ;
        RECT 51.110 18.080 51.400 18.370 ;
        RECT 51.920 17.700 52.080 18.380 ;
        RECT 52.665 18.370 52.825 19.500 ;
        RECT 53.175 18.370 53.335 20.480 ;
        RECT 53.920 20.220 54.080 20.780 ;
        RECT 54.665 19.660 54.825 20.480 ;
        RECT 53.575 19.500 54.825 19.660 ;
        RECT 53.580 18.560 53.870 18.850 ;
        RECT 54.130 18.560 54.420 18.850 ;
        RECT 53.580 18.490 53.740 18.560 ;
        RECT 54.260 18.490 54.420 18.560 ;
        RECT 52.600 18.080 52.890 18.370 ;
        RECT 53.110 18.080 53.400 18.370 ;
        RECT 53.920 17.700 54.080 18.380 ;
        RECT 54.665 18.370 54.825 19.500 ;
        RECT 55.175 18.370 55.335 20.480 ;
        RECT 55.920 20.220 56.080 20.780 ;
        RECT 56.665 19.660 56.825 20.480 ;
        RECT 55.575 19.500 56.825 19.660 ;
        RECT 55.580 18.560 55.870 18.850 ;
        RECT 56.130 18.560 56.420 18.850 ;
        RECT 55.580 18.490 55.740 18.560 ;
        RECT 56.260 18.490 56.420 18.560 ;
        RECT 54.600 18.080 54.890 18.370 ;
        RECT 55.110 18.080 55.400 18.370 ;
        RECT 55.920 17.700 56.080 18.380 ;
        RECT 56.665 18.370 56.825 19.500 ;
        RECT 57.175 18.370 57.335 20.480 ;
        RECT 57.920 20.220 58.080 20.780 ;
        RECT 58.665 19.660 58.825 20.480 ;
        RECT 57.575 19.500 58.825 19.660 ;
        RECT 57.580 18.560 57.870 18.850 ;
        RECT 58.130 18.560 58.420 18.850 ;
        RECT 57.580 18.490 57.740 18.560 ;
        RECT 58.260 18.490 58.420 18.560 ;
        RECT 56.600 18.080 56.890 18.370 ;
        RECT 57.110 18.080 57.400 18.370 ;
        RECT 57.920 17.700 58.080 18.380 ;
        RECT 58.665 18.370 58.825 19.500 ;
        RECT 59.175 18.370 59.335 20.480 ;
        RECT 59.920 20.220 60.080 20.780 ;
        RECT 60.665 19.660 60.825 20.480 ;
        RECT 59.575 19.500 60.825 19.660 ;
        RECT 59.580 18.560 59.870 18.850 ;
        RECT 60.130 18.560 60.420 18.850 ;
        RECT 59.580 18.490 59.740 18.560 ;
        RECT 60.260 18.490 60.420 18.560 ;
        RECT 58.600 18.080 58.890 18.370 ;
        RECT 59.110 18.080 59.400 18.370 ;
        RECT 59.920 17.700 60.080 18.380 ;
        RECT 60.665 18.370 60.825 19.500 ;
        RECT 61.175 18.370 61.335 20.480 ;
        RECT 61.920 20.220 62.080 20.780 ;
        RECT 62.665 19.660 62.825 20.480 ;
        RECT 61.575 19.500 62.825 19.660 ;
        RECT 61.580 18.560 61.870 18.850 ;
        RECT 62.130 18.560 62.420 18.850 ;
        RECT 61.580 18.490 61.740 18.560 ;
        RECT 62.260 18.490 62.420 18.560 ;
        RECT 60.600 18.080 60.890 18.370 ;
        RECT 61.110 18.080 61.400 18.370 ;
        RECT 61.920 17.700 62.080 18.380 ;
        RECT 62.665 18.370 62.825 19.500 ;
        RECT 63.175 18.370 63.335 20.480 ;
        RECT 63.920 20.220 64.080 20.780 ;
        RECT 64.665 19.660 64.825 20.480 ;
        RECT 63.575 19.500 64.825 19.660 ;
        RECT 63.580 18.560 63.870 18.850 ;
        RECT 64.130 18.560 64.420 18.850 ;
        RECT 63.580 18.490 63.740 18.560 ;
        RECT 64.260 18.490 64.420 18.560 ;
        RECT 62.600 18.080 62.890 18.370 ;
        RECT 63.110 18.080 63.400 18.370 ;
        RECT 63.920 17.700 64.080 18.380 ;
        RECT 64.665 18.370 64.825 19.500 ;
        RECT 65.175 18.370 65.335 20.480 ;
        RECT 65.920 20.220 66.080 20.780 ;
        RECT 66.665 19.660 66.825 20.480 ;
        RECT 65.575 19.500 66.825 19.660 ;
        RECT 65.580 18.560 65.870 18.850 ;
        RECT 66.130 18.560 66.420 18.850 ;
        RECT 65.580 18.490 65.740 18.560 ;
        RECT 66.260 18.490 66.420 18.560 ;
        RECT 64.600 18.080 64.890 18.370 ;
        RECT 65.110 18.080 65.400 18.370 ;
        RECT 65.920 17.700 66.080 18.380 ;
        RECT 66.665 18.370 66.825 19.500 ;
        RECT 67.175 18.370 67.335 20.480 ;
        RECT 67.920 20.220 68.080 20.780 ;
        RECT 68.665 19.660 68.825 20.480 ;
        RECT 67.575 19.500 68.825 19.660 ;
        RECT 67.580 18.560 67.870 18.850 ;
        RECT 68.130 18.560 68.420 18.850 ;
        RECT 67.580 18.490 67.740 18.560 ;
        RECT 68.260 18.490 68.420 18.560 ;
        RECT 66.600 18.080 66.890 18.370 ;
        RECT 67.110 18.080 67.400 18.370 ;
        RECT 67.920 17.700 68.080 18.380 ;
        RECT 68.665 18.370 68.825 19.500 ;
        RECT 69.175 18.370 69.335 20.480 ;
        RECT 69.920 20.220 70.080 20.780 ;
        RECT 70.665 19.660 70.825 20.480 ;
        RECT 69.575 19.500 70.825 19.660 ;
        RECT 69.580 18.560 69.870 18.850 ;
        RECT 70.130 18.560 70.420 18.850 ;
        RECT 69.580 18.490 69.740 18.560 ;
        RECT 70.260 18.490 70.420 18.560 ;
        RECT 68.600 18.080 68.890 18.370 ;
        RECT 69.110 18.080 69.400 18.370 ;
        RECT 69.920 17.700 70.080 18.380 ;
        RECT 70.665 18.370 70.825 19.500 ;
        RECT 71.175 18.370 71.335 20.480 ;
        RECT 71.920 20.220 72.080 20.780 ;
        RECT 72.665 19.660 72.825 20.480 ;
        RECT 71.575 19.500 72.825 19.660 ;
        RECT 71.580 18.560 71.870 18.850 ;
        RECT 72.130 18.560 72.420 18.850 ;
        RECT 71.580 18.490 71.740 18.560 ;
        RECT 72.260 18.490 72.420 18.560 ;
        RECT 70.600 18.080 70.890 18.370 ;
        RECT 71.110 18.080 71.400 18.370 ;
        RECT 71.920 17.700 72.080 18.380 ;
        RECT 72.665 18.370 72.825 19.500 ;
        RECT 73.175 18.370 73.335 20.480 ;
        RECT 73.920 20.220 74.080 20.780 ;
        RECT 74.665 19.660 74.825 20.480 ;
        RECT 73.575 19.500 74.825 19.660 ;
        RECT 73.580 18.560 73.870 18.850 ;
        RECT 74.130 18.560 74.420 18.850 ;
        RECT 73.580 18.490 73.740 18.560 ;
        RECT 74.260 18.490 74.420 18.560 ;
        RECT 72.600 18.080 72.890 18.370 ;
        RECT 73.110 18.080 73.400 18.370 ;
        RECT 73.920 17.700 74.080 18.380 ;
        RECT 74.665 18.370 74.825 19.500 ;
        RECT 75.175 18.370 75.335 20.480 ;
        RECT 75.920 20.220 76.080 20.780 ;
        RECT 76.665 19.660 76.825 20.480 ;
        RECT 75.575 19.500 76.825 19.660 ;
        RECT 75.580 18.560 75.870 18.850 ;
        RECT 76.130 18.560 76.420 18.850 ;
        RECT 75.580 18.490 75.740 18.560 ;
        RECT 76.260 18.490 76.420 18.560 ;
        RECT 74.600 18.080 74.890 18.370 ;
        RECT 75.110 18.080 75.400 18.370 ;
        RECT 75.920 17.700 76.080 18.380 ;
        RECT 76.665 18.370 76.825 19.500 ;
        RECT 77.175 18.370 77.335 20.480 ;
        RECT 77.920 20.220 78.080 20.780 ;
        RECT 78.665 19.660 78.825 20.480 ;
        RECT 77.575 19.500 78.825 19.660 ;
        RECT 77.580 18.560 77.870 18.850 ;
        RECT 78.130 18.560 78.420 18.850 ;
        RECT 77.580 18.490 77.740 18.560 ;
        RECT 78.260 18.490 78.420 18.560 ;
        RECT 76.600 18.080 76.890 18.370 ;
        RECT 77.110 18.080 77.400 18.370 ;
        RECT 77.920 17.700 78.080 18.380 ;
        RECT 78.665 18.370 78.825 19.500 ;
        RECT 79.175 18.370 79.335 20.480 ;
        RECT 79.920 20.220 80.080 20.780 ;
        RECT 80.665 19.660 80.825 20.480 ;
        RECT 79.575 19.500 80.825 19.660 ;
        RECT 79.580 18.560 79.870 18.850 ;
        RECT 80.130 18.560 80.420 18.850 ;
        RECT 79.580 18.490 79.740 18.560 ;
        RECT 80.260 18.490 80.420 18.560 ;
        RECT 78.600 18.080 78.890 18.370 ;
        RECT 79.110 18.080 79.400 18.370 ;
        RECT 79.920 17.700 80.080 18.380 ;
        RECT 80.665 18.370 80.825 19.500 ;
        RECT 81.175 18.370 81.335 20.480 ;
        RECT 81.920 20.220 82.080 20.780 ;
        RECT 82.665 19.660 82.825 20.480 ;
        RECT 81.575 19.500 82.825 19.660 ;
        RECT 81.580 18.560 81.870 18.850 ;
        RECT 82.130 18.560 82.420 18.850 ;
        RECT 81.580 18.490 81.740 18.560 ;
        RECT 82.260 18.490 82.420 18.560 ;
        RECT 80.600 18.080 80.890 18.370 ;
        RECT 81.110 18.080 81.400 18.370 ;
        RECT 81.920 17.700 82.080 18.380 ;
        RECT 82.665 18.370 82.825 19.500 ;
        RECT 83.175 18.370 83.335 20.480 ;
        RECT 83.920 20.220 84.080 20.780 ;
        RECT 84.665 19.660 84.825 20.480 ;
        RECT 83.575 19.500 84.825 19.660 ;
        RECT 83.580 18.560 83.870 18.850 ;
        RECT 84.130 18.560 84.420 18.850 ;
        RECT 83.580 18.490 83.740 18.560 ;
        RECT 84.260 18.490 84.420 18.560 ;
        RECT 82.600 18.080 82.890 18.370 ;
        RECT 83.110 18.080 83.400 18.370 ;
        RECT 83.920 17.700 84.080 18.380 ;
        RECT 84.665 18.370 84.825 19.500 ;
        RECT 85.175 18.370 85.335 20.480 ;
        RECT 85.920 20.220 86.080 20.780 ;
        RECT 86.665 19.660 86.825 20.480 ;
        RECT 85.575 19.500 86.825 19.660 ;
        RECT 85.580 18.560 85.870 18.850 ;
        RECT 86.130 18.560 86.420 18.850 ;
        RECT 85.580 18.490 85.740 18.560 ;
        RECT 86.260 18.490 86.420 18.560 ;
        RECT 84.600 18.080 84.890 18.370 ;
        RECT 85.110 18.080 85.400 18.370 ;
        RECT 85.920 17.700 86.080 18.380 ;
        RECT 86.665 18.370 86.825 19.500 ;
        RECT 87.175 18.370 87.335 20.480 ;
        RECT 87.920 20.220 88.080 20.780 ;
        RECT 88.665 19.660 88.825 20.480 ;
        RECT 87.575 19.500 88.825 19.660 ;
        RECT 87.580 18.560 87.870 18.850 ;
        RECT 88.130 18.560 88.420 18.850 ;
        RECT 87.580 18.490 87.740 18.560 ;
        RECT 88.260 18.490 88.420 18.560 ;
        RECT 86.600 18.080 86.890 18.370 ;
        RECT 87.110 18.080 87.400 18.370 ;
        RECT 87.920 17.700 88.080 18.380 ;
        RECT 88.665 18.370 88.825 19.500 ;
        RECT 89.175 18.370 89.335 20.480 ;
        RECT 89.920 20.220 90.080 20.780 ;
        RECT 90.665 19.660 90.825 20.480 ;
        RECT 89.575 19.500 90.825 19.660 ;
        RECT 89.580 18.560 89.870 18.850 ;
        RECT 90.130 18.560 90.420 18.850 ;
        RECT 89.580 18.490 89.740 18.560 ;
        RECT 90.260 18.490 90.420 18.560 ;
        RECT 88.600 18.080 88.890 18.370 ;
        RECT 89.110 18.080 89.400 18.370 ;
        RECT 89.920 17.700 90.080 18.380 ;
        RECT 90.665 18.370 90.825 19.500 ;
        RECT 91.175 18.370 91.335 20.480 ;
        RECT 91.920 20.220 92.080 20.780 ;
        RECT 92.665 19.660 92.825 20.480 ;
        RECT 91.575 19.500 92.825 19.660 ;
        RECT 91.580 18.560 91.870 18.850 ;
        RECT 92.130 18.560 92.420 18.850 ;
        RECT 91.580 18.490 91.740 18.560 ;
        RECT 92.260 18.490 92.420 18.560 ;
        RECT 90.600 18.080 90.890 18.370 ;
        RECT 91.110 18.080 91.400 18.370 ;
        RECT 91.920 17.700 92.080 18.380 ;
        RECT 92.665 18.370 92.825 19.500 ;
        RECT 93.175 18.370 93.335 20.480 ;
        RECT 93.920 20.220 94.080 20.780 ;
        RECT 94.665 19.660 94.825 20.480 ;
        RECT 93.575 19.500 94.825 19.660 ;
        RECT 93.580 18.560 93.870 18.850 ;
        RECT 94.130 18.560 94.420 18.850 ;
        RECT 93.580 18.490 93.740 18.560 ;
        RECT 94.260 18.490 94.420 18.560 ;
        RECT 92.600 18.080 92.890 18.370 ;
        RECT 93.110 18.080 93.400 18.370 ;
        RECT 93.920 17.700 94.080 18.380 ;
        RECT 94.665 18.370 94.825 19.500 ;
        RECT 95.175 18.370 95.335 20.480 ;
        RECT 95.920 20.220 96.080 20.780 ;
        RECT 96.665 19.660 96.825 20.480 ;
        RECT 95.575 19.500 96.825 19.660 ;
        RECT 95.580 18.560 95.870 18.850 ;
        RECT 96.130 18.560 96.420 18.850 ;
        RECT 95.580 18.490 95.740 18.560 ;
        RECT 96.260 18.490 96.420 18.560 ;
        RECT 94.600 18.080 94.890 18.370 ;
        RECT 95.110 18.080 95.400 18.370 ;
        RECT 95.920 17.700 96.080 18.380 ;
        RECT 96.665 18.370 96.825 19.500 ;
        RECT 97.175 18.370 97.335 20.480 ;
        RECT 97.920 20.220 98.080 20.780 ;
        RECT 98.665 19.660 98.825 20.480 ;
        RECT 97.575 19.500 98.825 19.660 ;
        RECT 97.580 18.560 97.870 18.850 ;
        RECT 98.130 18.560 98.420 18.850 ;
        RECT 97.580 18.490 97.740 18.560 ;
        RECT 98.260 18.490 98.420 18.560 ;
        RECT 96.600 18.080 96.890 18.370 ;
        RECT 97.110 18.080 97.400 18.370 ;
        RECT 97.920 17.700 98.080 18.380 ;
        RECT 98.665 18.370 98.825 19.500 ;
        RECT 99.175 18.370 99.335 20.480 ;
        RECT 99.920 20.220 100.080 20.780 ;
        RECT 100.665 19.660 100.825 20.480 ;
        RECT 99.575 19.500 100.825 19.660 ;
        RECT 99.580 18.560 99.870 18.850 ;
        RECT 100.130 18.560 100.420 18.850 ;
        RECT 99.580 18.490 99.740 18.560 ;
        RECT 100.260 18.490 100.420 18.560 ;
        RECT 98.600 18.080 98.890 18.370 ;
        RECT 99.110 18.080 99.400 18.370 ;
        RECT 99.920 17.700 100.080 18.380 ;
        RECT 100.665 18.370 100.825 19.500 ;
        RECT 101.175 18.370 101.335 20.480 ;
        RECT 101.920 20.220 102.080 20.780 ;
        RECT 102.665 19.660 102.825 20.480 ;
        RECT 101.575 19.500 102.825 19.660 ;
        RECT 101.580 18.560 101.870 18.850 ;
        RECT 102.130 18.560 102.420 18.850 ;
        RECT 101.580 18.490 101.740 18.560 ;
        RECT 102.260 18.490 102.420 18.560 ;
        RECT 100.600 18.080 100.890 18.370 ;
        RECT 101.110 18.080 101.400 18.370 ;
        RECT 101.920 17.700 102.080 18.380 ;
        RECT 102.665 18.370 102.825 19.500 ;
        RECT 103.175 18.370 103.335 20.480 ;
        RECT 103.920 20.220 104.080 20.780 ;
        RECT 104.665 19.660 104.825 20.480 ;
        RECT 103.575 19.500 104.825 19.660 ;
        RECT 103.580 18.560 103.870 18.850 ;
        RECT 104.130 18.560 104.420 18.850 ;
        RECT 103.580 18.490 103.740 18.560 ;
        RECT 104.260 18.490 104.420 18.560 ;
        RECT 102.600 18.080 102.890 18.370 ;
        RECT 103.110 18.080 103.400 18.370 ;
        RECT 103.920 17.700 104.080 18.380 ;
        RECT 104.665 18.370 104.825 19.500 ;
        RECT 105.175 18.370 105.335 20.480 ;
        RECT 105.920 20.220 106.080 20.780 ;
        RECT 106.665 19.660 106.825 20.480 ;
        RECT 105.575 19.500 106.825 19.660 ;
        RECT 105.580 18.560 105.870 18.850 ;
        RECT 106.130 18.560 106.420 18.850 ;
        RECT 105.580 18.490 105.740 18.560 ;
        RECT 106.260 18.490 106.420 18.560 ;
        RECT 104.600 18.080 104.890 18.370 ;
        RECT 105.110 18.080 105.400 18.370 ;
        RECT 105.920 17.700 106.080 18.380 ;
        RECT 106.665 18.370 106.825 19.500 ;
        RECT 107.175 18.370 107.335 20.480 ;
        RECT 107.920 20.220 108.080 20.780 ;
        RECT 108.665 19.660 108.825 20.480 ;
        RECT 107.575 19.500 108.825 19.660 ;
        RECT 107.580 18.560 107.870 18.850 ;
        RECT 108.130 18.560 108.420 18.850 ;
        RECT 107.580 18.490 107.740 18.560 ;
        RECT 108.260 18.490 108.420 18.560 ;
        RECT 106.600 18.080 106.890 18.370 ;
        RECT 107.110 18.080 107.400 18.370 ;
        RECT 107.920 17.700 108.080 18.380 ;
        RECT 108.665 18.370 108.825 19.500 ;
        RECT 109.175 18.370 109.335 20.480 ;
        RECT 109.920 20.220 110.080 20.780 ;
        RECT 110.665 19.660 110.825 20.480 ;
        RECT 109.575 19.500 110.825 19.660 ;
        RECT 109.580 18.560 109.870 18.850 ;
        RECT 110.130 18.560 110.420 18.850 ;
        RECT 109.580 18.490 109.740 18.560 ;
        RECT 110.260 18.490 110.420 18.560 ;
        RECT 108.600 18.080 108.890 18.370 ;
        RECT 109.110 18.080 109.400 18.370 ;
        RECT 109.920 17.700 110.080 18.380 ;
        RECT 110.665 18.370 110.825 19.500 ;
        RECT 111.175 18.370 111.335 20.480 ;
        RECT 111.920 20.220 112.080 20.780 ;
        RECT 112.665 19.660 112.825 20.480 ;
        RECT 111.575 19.500 112.825 19.660 ;
        RECT 111.580 18.560 111.870 18.850 ;
        RECT 112.130 18.560 112.420 18.850 ;
        RECT 111.580 18.490 111.740 18.560 ;
        RECT 112.260 18.490 112.420 18.560 ;
        RECT 110.600 18.080 110.890 18.370 ;
        RECT 111.110 18.080 111.400 18.370 ;
        RECT 111.920 17.700 112.080 18.380 ;
        RECT 112.665 18.370 112.825 19.500 ;
        RECT 113.175 18.370 113.335 20.480 ;
        RECT 113.920 20.220 114.080 20.780 ;
        RECT 114.665 19.660 114.825 20.480 ;
        RECT 113.575 19.500 114.825 19.660 ;
        RECT 113.580 18.560 113.870 18.850 ;
        RECT 114.130 18.560 114.420 18.850 ;
        RECT 113.580 18.490 113.740 18.560 ;
        RECT 114.260 18.490 114.420 18.560 ;
        RECT 112.600 18.080 112.890 18.370 ;
        RECT 113.110 18.080 113.400 18.370 ;
        RECT 113.920 17.700 114.080 18.380 ;
        RECT 114.665 18.370 114.825 19.500 ;
        RECT 115.175 18.370 115.335 20.480 ;
        RECT 115.920 20.220 116.080 20.780 ;
        RECT 116.665 19.660 116.825 20.480 ;
        RECT 115.575 19.500 116.825 19.660 ;
        RECT 115.580 18.560 115.870 18.850 ;
        RECT 116.130 18.560 116.420 18.850 ;
        RECT 115.580 18.490 115.740 18.560 ;
        RECT 116.260 18.490 116.420 18.560 ;
        RECT 114.600 18.080 114.890 18.370 ;
        RECT 115.110 18.080 115.400 18.370 ;
        RECT 115.920 17.700 116.080 18.380 ;
        RECT 116.665 18.370 116.825 19.500 ;
        RECT 117.175 18.370 117.335 20.480 ;
        RECT 117.920 20.220 118.080 20.780 ;
        RECT 118.665 19.660 118.825 20.480 ;
        RECT 117.575 19.500 118.825 19.660 ;
        RECT 117.580 18.560 117.870 18.850 ;
        RECT 118.130 18.560 118.420 18.850 ;
        RECT 117.580 18.490 117.740 18.560 ;
        RECT 118.260 18.490 118.420 18.560 ;
        RECT 116.600 18.080 116.890 18.370 ;
        RECT 117.110 18.080 117.400 18.370 ;
        RECT 117.920 17.700 118.080 18.380 ;
        RECT 118.665 18.370 118.825 19.500 ;
        RECT 119.175 18.370 119.335 20.480 ;
        RECT 119.920 20.220 120.080 20.780 ;
        RECT 120.665 19.660 120.825 20.480 ;
        RECT 119.575 19.500 120.825 19.660 ;
        RECT 119.580 18.560 119.870 18.850 ;
        RECT 120.130 18.560 120.420 18.850 ;
        RECT 119.580 18.490 119.740 18.560 ;
        RECT 120.260 18.490 120.420 18.560 ;
        RECT 118.600 18.080 118.890 18.370 ;
        RECT 119.110 18.080 119.400 18.370 ;
        RECT 119.920 17.700 120.080 18.380 ;
        RECT 120.665 18.370 120.825 19.500 ;
        RECT 121.175 18.370 121.335 20.480 ;
        RECT 121.920 20.220 122.080 20.780 ;
        RECT 122.665 19.660 122.825 20.480 ;
        RECT 121.575 19.500 122.825 19.660 ;
        RECT 121.580 18.560 121.870 18.850 ;
        RECT 122.130 18.560 122.420 18.850 ;
        RECT 121.580 18.490 121.740 18.560 ;
        RECT 122.260 18.490 122.420 18.560 ;
        RECT 120.600 18.080 120.890 18.370 ;
        RECT 121.110 18.080 121.400 18.370 ;
        RECT 121.920 17.700 122.080 18.380 ;
        RECT 122.665 18.370 122.825 19.500 ;
        RECT 123.175 18.370 123.335 20.480 ;
        RECT 123.920 20.220 124.080 20.780 ;
        RECT 124.665 19.660 124.825 20.480 ;
        RECT 123.575 19.500 124.825 19.660 ;
        RECT 123.580 18.560 123.870 18.850 ;
        RECT 124.130 18.560 124.420 18.850 ;
        RECT 123.580 18.490 123.740 18.560 ;
        RECT 124.260 18.490 124.420 18.560 ;
        RECT 122.600 18.080 122.890 18.370 ;
        RECT 123.110 18.080 123.400 18.370 ;
        RECT 123.920 17.700 124.080 18.380 ;
        RECT 124.665 18.370 124.825 19.500 ;
        RECT 125.175 18.370 125.335 20.480 ;
        RECT 125.920 20.220 126.080 20.780 ;
        RECT 126.665 19.660 126.825 20.480 ;
        RECT 125.575 19.500 126.825 19.660 ;
        RECT 125.580 18.560 125.870 18.850 ;
        RECT 126.130 18.560 126.420 18.850 ;
        RECT 125.580 18.490 125.740 18.560 ;
        RECT 126.260 18.490 126.420 18.560 ;
        RECT 124.600 18.080 124.890 18.370 ;
        RECT 125.110 18.080 125.400 18.370 ;
        RECT 125.920 17.700 126.080 18.380 ;
        RECT 126.665 18.370 126.825 19.500 ;
        RECT 127.175 18.370 127.335 20.480 ;
        RECT 127.920 20.220 128.080 20.780 ;
        RECT 128.665 19.660 128.825 20.480 ;
        RECT 127.575 19.500 128.825 19.660 ;
        RECT 127.580 18.560 127.870 18.850 ;
        RECT 128.130 18.560 128.420 18.850 ;
        RECT 127.580 18.490 127.740 18.560 ;
        RECT 128.260 18.490 128.420 18.560 ;
        RECT 126.600 18.080 126.890 18.370 ;
        RECT 127.110 18.080 127.400 18.370 ;
        RECT 127.920 17.700 128.080 18.380 ;
        RECT 128.665 18.370 128.825 19.500 ;
        RECT 129.175 18.370 129.335 20.480 ;
        RECT 129.920 20.220 130.080 20.780 ;
        RECT 130.665 19.660 130.825 20.480 ;
        RECT 129.575 19.500 130.825 19.660 ;
        RECT 129.580 18.560 129.870 18.850 ;
        RECT 130.130 18.560 130.420 18.850 ;
        RECT 129.580 18.490 129.740 18.560 ;
        RECT 130.260 18.490 130.420 18.560 ;
        RECT 128.600 18.080 128.890 18.370 ;
        RECT 129.110 18.080 129.400 18.370 ;
        RECT 129.920 17.700 130.080 18.380 ;
        RECT 130.665 18.370 130.825 19.500 ;
        RECT 130.600 18.080 130.890 18.370 ;
        RECT -0.930 16.500 -0.670 17.200 ;
        RECT -0.490 16.720 -0.190 17.020 ;
        RECT 0.190 16.720 0.490 17.020 ;
        RECT -0.930 16.240 -0.430 16.500 ;
        RECT -0.150 16.220 0.150 16.520 ;
        RECT 0.360 16.220 0.660 16.520 ;
        RECT 1.070 16.500 1.330 17.200 ;
        RECT 1.510 16.720 1.810 17.020 ;
        RECT 2.190 16.720 2.490 17.020 ;
        RECT 1.070 16.240 1.570 16.500 ;
        RECT 1.850 16.220 2.150 16.520 ;
        RECT 2.360 16.220 2.660 16.520 ;
        RECT 3.070 16.500 3.330 17.200 ;
        RECT 3.510 16.720 3.810 17.020 ;
        RECT 4.190 16.720 4.490 17.020 ;
        RECT 3.070 16.240 3.570 16.500 ;
        RECT 3.850 16.220 4.150 16.520 ;
        RECT 4.360 16.220 4.660 16.520 ;
        RECT 5.070 16.500 5.330 17.200 ;
        RECT 5.510 16.720 5.810 17.020 ;
        RECT 6.190 16.720 6.490 17.020 ;
        RECT 5.070 16.240 5.570 16.500 ;
        RECT 5.850 16.220 6.150 16.520 ;
        RECT 6.360 16.220 6.660 16.520 ;
        RECT 7.070 16.500 7.330 17.200 ;
        RECT 7.510 16.720 7.810 17.020 ;
        RECT 8.190 16.720 8.490 17.020 ;
        RECT 7.070 16.240 7.570 16.500 ;
        RECT 7.850 16.220 8.150 16.520 ;
        RECT 8.360 16.220 8.660 16.520 ;
        RECT 9.070 16.500 9.330 17.200 ;
        RECT 9.510 16.720 9.810 17.020 ;
        RECT 10.190 16.720 10.490 17.020 ;
        RECT 9.070 16.240 9.570 16.500 ;
        RECT 9.850 16.220 10.150 16.520 ;
        RECT 10.360 16.220 10.660 16.520 ;
        RECT 11.070 16.500 11.330 17.200 ;
        RECT 11.510 16.720 11.810 17.020 ;
        RECT 12.190 16.720 12.490 17.020 ;
        RECT 11.070 16.240 11.570 16.500 ;
        RECT 11.850 16.220 12.150 16.520 ;
        RECT 12.360 16.220 12.660 16.520 ;
        RECT 13.070 16.500 13.330 17.200 ;
        RECT 13.510 16.720 13.810 17.020 ;
        RECT 14.190 16.720 14.490 17.020 ;
        RECT 13.070 16.240 13.570 16.500 ;
        RECT 13.850 16.220 14.150 16.520 ;
        RECT 14.360 16.220 14.660 16.520 ;
        RECT 15.070 16.500 15.330 17.200 ;
        RECT 15.510 16.720 15.810 17.020 ;
        RECT 16.190 16.720 16.490 17.020 ;
        RECT 15.070 16.240 15.570 16.500 ;
        RECT 15.850 16.220 16.150 16.520 ;
        RECT 16.360 16.220 16.660 16.520 ;
        RECT 17.070 16.500 17.330 17.200 ;
        RECT 17.510 16.720 17.810 17.020 ;
        RECT 18.190 16.720 18.490 17.020 ;
        RECT 17.070 16.240 17.570 16.500 ;
        RECT 17.850 16.220 18.150 16.520 ;
        RECT 18.360 16.220 18.660 16.520 ;
        RECT 19.070 16.500 19.330 17.200 ;
        RECT 19.510 16.720 19.810 17.020 ;
        RECT 20.190 16.720 20.490 17.020 ;
        RECT 19.070 16.240 19.570 16.500 ;
        RECT 19.850 16.220 20.150 16.520 ;
        RECT 20.360 16.220 20.660 16.520 ;
        RECT 21.070 16.500 21.330 17.200 ;
        RECT 21.510 16.720 21.810 17.020 ;
        RECT 22.190 16.720 22.490 17.020 ;
        RECT 21.070 16.240 21.570 16.500 ;
        RECT 21.850 16.220 22.150 16.520 ;
        RECT 22.360 16.220 22.660 16.520 ;
        RECT 23.070 16.500 23.330 17.200 ;
        RECT 23.510 16.720 23.810 17.020 ;
        RECT 24.190 16.720 24.490 17.020 ;
        RECT 23.070 16.240 23.570 16.500 ;
        RECT 23.850 16.220 24.150 16.520 ;
        RECT 24.360 16.220 24.660 16.520 ;
        RECT 25.070 16.500 25.330 17.200 ;
        RECT 25.510 16.720 25.810 17.020 ;
        RECT 26.190 16.720 26.490 17.020 ;
        RECT 25.070 16.240 25.570 16.500 ;
        RECT 25.850 16.220 26.150 16.520 ;
        RECT 26.360 16.220 26.660 16.520 ;
        RECT 27.070 16.500 27.330 17.200 ;
        RECT 27.510 16.720 27.810 17.020 ;
        RECT 28.190 16.720 28.490 17.020 ;
        RECT 27.070 16.240 27.570 16.500 ;
        RECT 27.850 16.220 28.150 16.520 ;
        RECT 28.360 16.220 28.660 16.520 ;
        RECT 29.070 16.500 29.330 17.200 ;
        RECT 29.510 16.720 29.810 17.020 ;
        RECT 30.190 16.720 30.490 17.020 ;
        RECT 29.070 16.240 29.570 16.500 ;
        RECT 29.850 16.220 30.150 16.520 ;
        RECT 30.360 16.220 30.660 16.520 ;
        RECT 31.070 16.500 31.330 17.200 ;
        RECT 31.510 16.720 31.810 17.020 ;
        RECT 32.190 16.720 32.490 17.020 ;
        RECT 31.070 16.240 31.570 16.500 ;
        RECT 31.850 16.220 32.150 16.520 ;
        RECT 32.360 16.220 32.660 16.520 ;
        RECT 33.070 16.500 33.330 17.200 ;
        RECT 33.510 16.720 33.810 17.020 ;
        RECT 34.190 16.720 34.490 17.020 ;
        RECT 33.070 16.240 33.570 16.500 ;
        RECT 33.850 16.220 34.150 16.520 ;
        RECT 34.360 16.220 34.660 16.520 ;
        RECT 35.070 16.500 35.330 17.200 ;
        RECT 35.510 16.720 35.810 17.020 ;
        RECT 36.190 16.720 36.490 17.020 ;
        RECT 35.070 16.240 35.570 16.500 ;
        RECT 35.850 16.220 36.150 16.520 ;
        RECT 36.360 16.220 36.660 16.520 ;
        RECT 37.070 16.500 37.330 17.200 ;
        RECT 37.510 16.720 37.810 17.020 ;
        RECT 38.190 16.720 38.490 17.020 ;
        RECT 37.070 16.240 37.570 16.500 ;
        RECT 37.850 16.220 38.150 16.520 ;
        RECT 38.360 16.220 38.660 16.520 ;
        RECT 39.070 16.500 39.330 17.200 ;
        RECT 39.510 16.720 39.810 17.020 ;
        RECT 40.190 16.720 40.490 17.020 ;
        RECT 39.070 16.240 39.570 16.500 ;
        RECT 39.850 16.220 40.150 16.520 ;
        RECT 40.360 16.220 40.660 16.520 ;
        RECT 41.070 16.500 41.330 17.200 ;
        RECT 41.510 16.720 41.810 17.020 ;
        RECT 42.190 16.720 42.490 17.020 ;
        RECT 41.070 16.240 41.570 16.500 ;
        RECT 41.850 16.220 42.150 16.520 ;
        RECT 42.360 16.220 42.660 16.520 ;
        RECT 43.070 16.500 43.330 17.200 ;
        RECT 43.510 16.720 43.810 17.020 ;
        RECT 44.190 16.720 44.490 17.020 ;
        RECT 43.070 16.240 43.570 16.500 ;
        RECT 43.850 16.220 44.150 16.520 ;
        RECT 44.360 16.220 44.660 16.520 ;
        RECT 45.070 16.500 45.330 17.200 ;
        RECT 45.510 16.720 45.810 17.020 ;
        RECT 46.190 16.720 46.490 17.020 ;
        RECT 45.070 16.240 45.570 16.500 ;
        RECT 45.850 16.220 46.150 16.520 ;
        RECT 46.360 16.220 46.660 16.520 ;
        RECT 47.070 16.500 47.330 17.200 ;
        RECT 47.510 16.720 47.810 17.020 ;
        RECT 48.190 16.720 48.490 17.020 ;
        RECT 47.070 16.240 47.570 16.500 ;
        RECT 47.850 16.220 48.150 16.520 ;
        RECT 48.360 16.220 48.660 16.520 ;
        RECT 49.070 16.500 49.330 17.200 ;
        RECT 49.510 16.720 49.810 17.020 ;
        RECT 50.190 16.720 50.490 17.020 ;
        RECT 49.070 16.240 49.570 16.500 ;
        RECT 49.850 16.220 50.150 16.520 ;
        RECT 50.360 16.220 50.660 16.520 ;
        RECT 51.070 16.500 51.330 17.200 ;
        RECT 51.510 16.720 51.810 17.020 ;
        RECT 52.190 16.720 52.490 17.020 ;
        RECT 51.070 16.240 51.570 16.500 ;
        RECT 51.850 16.220 52.150 16.520 ;
        RECT 52.360 16.220 52.660 16.520 ;
        RECT 53.070 16.500 53.330 17.200 ;
        RECT 53.510 16.720 53.810 17.020 ;
        RECT 54.190 16.720 54.490 17.020 ;
        RECT 53.070 16.240 53.570 16.500 ;
        RECT 53.850 16.220 54.150 16.520 ;
        RECT 54.360 16.220 54.660 16.520 ;
        RECT 55.070 16.500 55.330 17.200 ;
        RECT 55.510 16.720 55.810 17.020 ;
        RECT 56.190 16.720 56.490 17.020 ;
        RECT 55.070 16.240 55.570 16.500 ;
        RECT 55.850 16.220 56.150 16.520 ;
        RECT 56.360 16.220 56.660 16.520 ;
        RECT 57.070 16.500 57.330 17.200 ;
        RECT 57.510 16.720 57.810 17.020 ;
        RECT 58.190 16.720 58.490 17.020 ;
        RECT 57.070 16.240 57.570 16.500 ;
        RECT 57.850 16.220 58.150 16.520 ;
        RECT 58.360 16.220 58.660 16.520 ;
        RECT 59.070 16.500 59.330 17.200 ;
        RECT 59.510 16.720 59.810 17.020 ;
        RECT 60.190 16.720 60.490 17.020 ;
        RECT 59.070 16.240 59.570 16.500 ;
        RECT 59.850 16.220 60.150 16.520 ;
        RECT 60.360 16.220 60.660 16.520 ;
        RECT 61.070 16.500 61.330 17.200 ;
        RECT 61.510 16.720 61.810 17.020 ;
        RECT 62.190 16.720 62.490 17.020 ;
        RECT 61.070 16.240 61.570 16.500 ;
        RECT 61.850 16.220 62.150 16.520 ;
        RECT 62.360 16.220 62.660 16.520 ;
        RECT 63.070 16.500 63.330 17.200 ;
        RECT 63.510 16.720 63.810 17.020 ;
        RECT 64.190 16.720 64.490 17.020 ;
        RECT 63.070 16.240 63.570 16.500 ;
        RECT 63.850 16.220 64.150 16.520 ;
        RECT 64.360 16.220 64.660 16.520 ;
        RECT 65.070 16.500 65.330 17.200 ;
        RECT 65.510 16.720 65.810 17.020 ;
        RECT 66.190 16.720 66.490 17.020 ;
        RECT 65.070 16.240 65.570 16.500 ;
        RECT 65.850 16.220 66.150 16.520 ;
        RECT 66.360 16.220 66.660 16.520 ;
        RECT 67.070 16.500 67.330 17.200 ;
        RECT 67.510 16.720 67.810 17.020 ;
        RECT 68.190 16.720 68.490 17.020 ;
        RECT 67.070 16.240 67.570 16.500 ;
        RECT 67.850 16.220 68.150 16.520 ;
        RECT 68.360 16.220 68.660 16.520 ;
        RECT 69.070 16.500 69.330 17.200 ;
        RECT 69.510 16.720 69.810 17.020 ;
        RECT 70.190 16.720 70.490 17.020 ;
        RECT 69.070 16.240 69.570 16.500 ;
        RECT 69.850 16.220 70.150 16.520 ;
        RECT 70.360 16.220 70.660 16.520 ;
        RECT 71.070 16.500 71.330 17.200 ;
        RECT 71.510 16.720 71.810 17.020 ;
        RECT 72.190 16.720 72.490 17.020 ;
        RECT 71.070 16.240 71.570 16.500 ;
        RECT 71.850 16.220 72.150 16.520 ;
        RECT 72.360 16.220 72.660 16.520 ;
        RECT 73.070 16.500 73.330 17.200 ;
        RECT 73.510 16.720 73.810 17.020 ;
        RECT 74.190 16.720 74.490 17.020 ;
        RECT 73.070 16.240 73.570 16.500 ;
        RECT 73.850 16.220 74.150 16.520 ;
        RECT 74.360 16.220 74.660 16.520 ;
        RECT 75.070 16.500 75.330 17.200 ;
        RECT 75.510 16.720 75.810 17.020 ;
        RECT 76.190 16.720 76.490 17.020 ;
        RECT 75.070 16.240 75.570 16.500 ;
        RECT 75.850 16.220 76.150 16.520 ;
        RECT 76.360 16.220 76.660 16.520 ;
        RECT 77.070 16.500 77.330 17.200 ;
        RECT 77.510 16.720 77.810 17.020 ;
        RECT 78.190 16.720 78.490 17.020 ;
        RECT 77.070 16.240 77.570 16.500 ;
        RECT 77.850 16.220 78.150 16.520 ;
        RECT 78.360 16.220 78.660 16.520 ;
        RECT 79.070 16.500 79.330 17.200 ;
        RECT 79.510 16.720 79.810 17.020 ;
        RECT 80.190 16.720 80.490 17.020 ;
        RECT 79.070 16.240 79.570 16.500 ;
        RECT 79.850 16.220 80.150 16.520 ;
        RECT 80.360 16.220 80.660 16.520 ;
        RECT 81.070 16.500 81.330 17.200 ;
        RECT 81.510 16.720 81.810 17.020 ;
        RECT 82.190 16.720 82.490 17.020 ;
        RECT 81.070 16.240 81.570 16.500 ;
        RECT 81.850 16.220 82.150 16.520 ;
        RECT 82.360 16.220 82.660 16.520 ;
        RECT 83.070 16.500 83.330 17.200 ;
        RECT 83.510 16.720 83.810 17.020 ;
        RECT 84.190 16.720 84.490 17.020 ;
        RECT 83.070 16.240 83.570 16.500 ;
        RECT 83.850 16.220 84.150 16.520 ;
        RECT 84.360 16.220 84.660 16.520 ;
        RECT 85.070 16.500 85.330 17.200 ;
        RECT 85.510 16.720 85.810 17.020 ;
        RECT 86.190 16.720 86.490 17.020 ;
        RECT 85.070 16.240 85.570 16.500 ;
        RECT 85.850 16.220 86.150 16.520 ;
        RECT 86.360 16.220 86.660 16.520 ;
        RECT 87.070 16.500 87.330 17.200 ;
        RECT 87.510 16.720 87.810 17.020 ;
        RECT 88.190 16.720 88.490 17.020 ;
        RECT 87.070 16.240 87.570 16.500 ;
        RECT 87.850 16.220 88.150 16.520 ;
        RECT 88.360 16.220 88.660 16.520 ;
        RECT 89.070 16.500 89.330 17.200 ;
        RECT 89.510 16.720 89.810 17.020 ;
        RECT 90.190 16.720 90.490 17.020 ;
        RECT 89.070 16.240 89.570 16.500 ;
        RECT 89.850 16.220 90.150 16.520 ;
        RECT 90.360 16.220 90.660 16.520 ;
        RECT 91.070 16.500 91.330 17.200 ;
        RECT 91.510 16.720 91.810 17.020 ;
        RECT 92.190 16.720 92.490 17.020 ;
        RECT 91.070 16.240 91.570 16.500 ;
        RECT 91.850 16.220 92.150 16.520 ;
        RECT 92.360 16.220 92.660 16.520 ;
        RECT 93.070 16.500 93.330 17.200 ;
        RECT 93.510 16.720 93.810 17.020 ;
        RECT 94.190 16.720 94.490 17.020 ;
        RECT 93.070 16.240 93.570 16.500 ;
        RECT 93.850 16.220 94.150 16.520 ;
        RECT 94.360 16.220 94.660 16.520 ;
        RECT 95.070 16.500 95.330 17.200 ;
        RECT 95.510 16.720 95.810 17.020 ;
        RECT 96.190 16.720 96.490 17.020 ;
        RECT 95.070 16.240 95.570 16.500 ;
        RECT 95.850 16.220 96.150 16.520 ;
        RECT 96.360 16.220 96.660 16.520 ;
        RECT 97.070 16.500 97.330 17.200 ;
        RECT 97.510 16.720 97.810 17.020 ;
        RECT 98.190 16.720 98.490 17.020 ;
        RECT 97.070 16.240 97.570 16.500 ;
        RECT 97.850 16.220 98.150 16.520 ;
        RECT 98.360 16.220 98.660 16.520 ;
        RECT 99.070 16.500 99.330 17.200 ;
        RECT 99.510 16.720 99.810 17.020 ;
        RECT 100.190 16.720 100.490 17.020 ;
        RECT 99.070 16.240 99.570 16.500 ;
        RECT 99.850 16.220 100.150 16.520 ;
        RECT 100.360 16.220 100.660 16.520 ;
        RECT 101.070 16.500 101.330 17.200 ;
        RECT 101.510 16.720 101.810 17.020 ;
        RECT 102.190 16.720 102.490 17.020 ;
        RECT 101.070 16.240 101.570 16.500 ;
        RECT 101.850 16.220 102.150 16.520 ;
        RECT 102.360 16.220 102.660 16.520 ;
        RECT 103.070 16.500 103.330 17.200 ;
        RECT 103.510 16.720 103.810 17.020 ;
        RECT 104.190 16.720 104.490 17.020 ;
        RECT 103.070 16.240 103.570 16.500 ;
        RECT 103.850 16.220 104.150 16.520 ;
        RECT 104.360 16.220 104.660 16.520 ;
        RECT 105.070 16.500 105.330 17.200 ;
        RECT 105.510 16.720 105.810 17.020 ;
        RECT 106.190 16.720 106.490 17.020 ;
        RECT 105.070 16.240 105.570 16.500 ;
        RECT 105.850 16.220 106.150 16.520 ;
        RECT 106.360 16.220 106.660 16.520 ;
        RECT 107.070 16.500 107.330 17.200 ;
        RECT 107.510 16.720 107.810 17.020 ;
        RECT 108.190 16.720 108.490 17.020 ;
        RECT 107.070 16.240 107.570 16.500 ;
        RECT 107.850 16.220 108.150 16.520 ;
        RECT 108.360 16.220 108.660 16.520 ;
        RECT 109.070 16.500 109.330 17.200 ;
        RECT 109.510 16.720 109.810 17.020 ;
        RECT 110.190 16.720 110.490 17.020 ;
        RECT 109.070 16.240 109.570 16.500 ;
        RECT 109.850 16.220 110.150 16.520 ;
        RECT 110.360 16.220 110.660 16.520 ;
        RECT 111.070 16.500 111.330 17.200 ;
        RECT 111.510 16.720 111.810 17.020 ;
        RECT 112.190 16.720 112.490 17.020 ;
        RECT 111.070 16.240 111.570 16.500 ;
        RECT 111.850 16.220 112.150 16.520 ;
        RECT 112.360 16.220 112.660 16.520 ;
        RECT 113.070 16.500 113.330 17.200 ;
        RECT 113.510 16.720 113.810 17.020 ;
        RECT 114.190 16.720 114.490 17.020 ;
        RECT 113.070 16.240 113.570 16.500 ;
        RECT 113.850 16.220 114.150 16.520 ;
        RECT 114.360 16.220 114.660 16.520 ;
        RECT 115.070 16.500 115.330 17.200 ;
        RECT 115.510 16.720 115.810 17.020 ;
        RECT 116.190 16.720 116.490 17.020 ;
        RECT 115.070 16.240 115.570 16.500 ;
        RECT 115.850 16.220 116.150 16.520 ;
        RECT 116.360 16.220 116.660 16.520 ;
        RECT 117.070 16.500 117.330 17.200 ;
        RECT 117.510 16.720 117.810 17.020 ;
        RECT 118.190 16.720 118.490 17.020 ;
        RECT 117.070 16.240 117.570 16.500 ;
        RECT 117.850 16.220 118.150 16.520 ;
        RECT 118.360 16.220 118.660 16.520 ;
        RECT 119.070 16.500 119.330 17.200 ;
        RECT 119.510 16.720 119.810 17.020 ;
        RECT 120.190 16.720 120.490 17.020 ;
        RECT 119.070 16.240 119.570 16.500 ;
        RECT 119.850 16.220 120.150 16.520 ;
        RECT 120.360 16.220 120.660 16.520 ;
        RECT 121.070 16.500 121.330 17.200 ;
        RECT 121.510 16.720 121.810 17.020 ;
        RECT 122.190 16.720 122.490 17.020 ;
        RECT 121.070 16.240 121.570 16.500 ;
        RECT 121.850 16.220 122.150 16.520 ;
        RECT 122.360 16.220 122.660 16.520 ;
        RECT 123.070 16.500 123.330 17.200 ;
        RECT 123.510 16.720 123.810 17.020 ;
        RECT 124.190 16.720 124.490 17.020 ;
        RECT 123.070 16.240 123.570 16.500 ;
        RECT 123.850 16.220 124.150 16.520 ;
        RECT 124.360 16.220 124.660 16.520 ;
        RECT 125.070 16.500 125.330 17.200 ;
        RECT 125.510 16.720 125.810 17.020 ;
        RECT 126.190 16.720 126.490 17.020 ;
        RECT 125.070 16.240 125.570 16.500 ;
        RECT 125.850 16.220 126.150 16.520 ;
        RECT 126.360 16.220 126.660 16.520 ;
        RECT 127.070 16.500 127.330 17.200 ;
        RECT 127.510 16.720 127.810 17.020 ;
        RECT 128.190 16.720 128.490 17.020 ;
        RECT 127.070 16.240 127.570 16.500 ;
        RECT 127.850 16.220 128.150 16.520 ;
        RECT 128.360 16.220 128.660 16.520 ;
        RECT 129.070 16.500 129.330 17.200 ;
        RECT 129.510 16.720 129.810 17.020 ;
        RECT 130.190 16.720 130.490 17.020 ;
        RECT 129.070 16.240 129.570 16.500 ;
        RECT 129.850 16.220 130.150 16.520 ;
        RECT 130.360 16.220 130.660 16.520 ;
        RECT -1.895 8.760 -1.605 14.970 ;
        RECT -1.300 10.040 -1.000 14.610 ;
        RECT 131.000 10.040 131.300 14.610 ;
        RECT -1.300 8.760 -1.140 10.040 ;
        RECT -0.815 8.755 0.375 10.040 ;
        RECT 0.560 9.145 0.780 9.855 ;
        RECT 2.560 9.145 2.780 9.855 ;
        RECT 4.560 9.145 4.780 9.855 ;
        RECT 6.560 9.145 6.780 9.855 ;
        RECT 8.560 9.145 8.780 9.855 ;
        RECT 10.560 9.145 10.780 9.855 ;
        RECT 12.560 9.145 12.780 9.855 ;
        RECT 14.560 9.145 14.780 9.855 ;
        RECT 16.560 9.145 16.780 9.855 ;
        RECT 18.560 9.145 18.780 9.855 ;
        RECT 20.560 9.145 20.780 9.855 ;
        RECT 22.560 9.145 22.780 9.855 ;
        RECT 24.560 9.145 24.780 9.855 ;
        RECT 26.560 9.145 26.780 9.855 ;
        RECT 28.560 9.145 28.780 9.855 ;
        RECT 30.560 9.145 30.780 9.855 ;
        RECT 32.560 9.145 32.780 9.855 ;
        RECT 34.560 9.145 34.780 9.855 ;
        RECT 36.560 9.145 36.780 9.855 ;
        RECT 38.560 9.145 38.780 9.855 ;
        RECT 40.560 9.145 40.780 9.855 ;
        RECT 42.560 9.145 42.780 9.855 ;
        RECT 44.560 9.145 44.780 9.855 ;
        RECT 46.560 9.145 46.780 9.855 ;
        RECT 48.560 9.145 48.780 9.855 ;
        RECT 50.560 9.145 50.780 9.855 ;
        RECT 52.560 9.145 52.780 9.855 ;
        RECT 54.560 9.145 54.780 9.855 ;
        RECT 56.560 9.145 56.780 9.855 ;
        RECT 58.560 9.145 58.780 9.855 ;
        RECT 60.560 9.145 60.780 9.855 ;
        RECT 62.560 9.145 62.780 9.855 ;
        RECT 64.560 9.145 64.780 9.855 ;
        RECT 66.560 9.145 66.780 9.855 ;
        RECT 68.560 9.145 68.780 9.855 ;
        RECT 70.560 9.145 70.780 9.855 ;
        RECT 72.560 9.145 72.780 9.855 ;
        RECT 74.560 9.145 74.780 9.855 ;
        RECT 76.560 9.145 76.780 9.855 ;
        RECT 78.560 9.145 78.780 9.855 ;
        RECT 80.560 9.145 80.780 9.855 ;
        RECT 82.560 9.145 82.780 9.855 ;
        RECT 84.560 9.145 84.780 9.855 ;
        RECT 86.560 9.145 86.780 9.855 ;
        RECT 88.560 9.145 88.780 9.855 ;
        RECT 90.560 9.145 90.780 9.855 ;
        RECT 92.560 9.145 92.780 9.855 ;
        RECT 94.560 9.145 94.780 9.855 ;
        RECT 96.560 9.145 96.780 9.855 ;
        RECT 98.560 9.145 98.780 9.855 ;
        RECT 100.560 9.145 100.780 9.855 ;
        RECT 102.560 9.145 102.780 9.855 ;
        RECT 104.560 9.145 104.780 9.855 ;
        RECT 106.560 9.145 106.780 9.855 ;
        RECT 108.560 9.145 108.780 9.855 ;
        RECT 110.560 9.145 110.780 9.855 ;
        RECT 112.560 9.145 112.780 9.855 ;
        RECT 114.560 9.145 114.780 9.855 ;
        RECT 116.560 9.145 116.780 9.855 ;
        RECT 118.560 9.145 118.780 9.855 ;
        RECT 120.560 9.145 120.780 9.855 ;
        RECT 122.560 9.145 122.780 9.855 ;
        RECT 124.560 9.145 124.780 9.855 ;
        RECT 126.560 9.145 126.780 9.855 ;
        RECT 128.560 9.145 128.780 9.855 ;
        RECT 1.185 8.535 128.375 8.965 ;
        RECT 129.185 8.755 130.375 10.040 ;
        RECT 130.560 9.145 130.780 9.855 ;
        RECT 131.140 8.760 131.300 10.040 ;
        RECT 131.605 8.760 131.895 14.970 ;
        RECT -1.895 1.400 -1.605 7.610 ;
        RECT -1.300 6.330 -1.140 7.610 ;
        RECT -0.780 6.515 -0.560 7.225 ;
        RECT -0.375 6.330 0.815 7.615 ;
        RECT 1.625 7.405 128.815 7.835 ;
        RECT 1.220 6.515 1.440 7.225 ;
        RECT 3.220 6.515 3.440 7.225 ;
        RECT 5.220 6.515 5.440 7.225 ;
        RECT 7.220 6.515 7.440 7.225 ;
        RECT 9.220 6.515 9.440 7.225 ;
        RECT 11.220 6.515 11.440 7.225 ;
        RECT 13.220 6.515 13.440 7.225 ;
        RECT 15.220 6.515 15.440 7.225 ;
        RECT 17.220 6.515 17.440 7.225 ;
        RECT 19.220 6.515 19.440 7.225 ;
        RECT 21.220 6.515 21.440 7.225 ;
        RECT 23.220 6.515 23.440 7.225 ;
        RECT 25.220 6.515 25.440 7.225 ;
        RECT 27.220 6.515 27.440 7.225 ;
        RECT 29.220 6.515 29.440 7.225 ;
        RECT 31.220 6.515 31.440 7.225 ;
        RECT 33.220 6.515 33.440 7.225 ;
        RECT 35.220 6.515 35.440 7.225 ;
        RECT 37.220 6.515 37.440 7.225 ;
        RECT 39.220 6.515 39.440 7.225 ;
        RECT 41.220 6.515 41.440 7.225 ;
        RECT 43.220 6.515 43.440 7.225 ;
        RECT 45.220 6.515 45.440 7.225 ;
        RECT 47.220 6.515 47.440 7.225 ;
        RECT 49.220 6.515 49.440 7.225 ;
        RECT 51.220 6.515 51.440 7.225 ;
        RECT 53.220 6.515 53.440 7.225 ;
        RECT 55.220 6.515 55.440 7.225 ;
        RECT 57.220 6.515 57.440 7.225 ;
        RECT 59.220 6.515 59.440 7.225 ;
        RECT 61.220 6.515 61.440 7.225 ;
        RECT 63.220 6.515 63.440 7.225 ;
        RECT 65.220 6.515 65.440 7.225 ;
        RECT 67.220 6.515 67.440 7.225 ;
        RECT 69.220 6.515 69.440 7.225 ;
        RECT 71.220 6.515 71.440 7.225 ;
        RECT 73.220 6.515 73.440 7.225 ;
        RECT 75.220 6.515 75.440 7.225 ;
        RECT 77.220 6.515 77.440 7.225 ;
        RECT 79.220 6.515 79.440 7.225 ;
        RECT 81.220 6.515 81.440 7.225 ;
        RECT 83.220 6.515 83.440 7.225 ;
        RECT 85.220 6.515 85.440 7.225 ;
        RECT 87.220 6.515 87.440 7.225 ;
        RECT 89.220 6.515 89.440 7.225 ;
        RECT 91.220 6.515 91.440 7.225 ;
        RECT 93.220 6.515 93.440 7.225 ;
        RECT 95.220 6.515 95.440 7.225 ;
        RECT 97.220 6.515 97.440 7.225 ;
        RECT 99.220 6.515 99.440 7.225 ;
        RECT 101.220 6.515 101.440 7.225 ;
        RECT 103.220 6.515 103.440 7.225 ;
        RECT 105.220 6.515 105.440 7.225 ;
        RECT 107.220 6.515 107.440 7.225 ;
        RECT 109.220 6.515 109.440 7.225 ;
        RECT 111.220 6.515 111.440 7.225 ;
        RECT 113.220 6.515 113.440 7.225 ;
        RECT 115.220 6.515 115.440 7.225 ;
        RECT 117.220 6.515 117.440 7.225 ;
        RECT 119.220 6.515 119.440 7.225 ;
        RECT 121.220 6.515 121.440 7.225 ;
        RECT 123.220 6.515 123.440 7.225 ;
        RECT 125.220 6.515 125.440 7.225 ;
        RECT 127.220 6.515 127.440 7.225 ;
        RECT 129.220 6.515 129.440 7.225 ;
        RECT 129.625 6.330 130.815 7.615 ;
        RECT 131.140 6.330 131.300 7.610 ;
        RECT -1.300 1.760 -1.000 6.330 ;
        RECT 131.000 1.760 131.300 6.330 ;
        RECT 131.605 1.400 131.895 7.610 ;
        RECT -0.660 -0.150 -0.360 0.150 ;
        RECT -0.150 -0.150 0.150 0.150 ;
        RECT 0.430 -0.130 0.930 0.130 ;
        RECT -0.490 -0.650 -0.190 -0.350 ;
        RECT 0.190 -0.650 0.490 -0.350 ;
        RECT 0.670 -0.830 0.930 -0.130 ;
        RECT 1.340 -0.150 1.640 0.150 ;
        RECT 1.850 -0.150 2.150 0.150 ;
        RECT 2.430 -0.130 2.930 0.130 ;
        RECT 1.510 -0.650 1.810 -0.350 ;
        RECT 2.190 -0.650 2.490 -0.350 ;
        RECT 2.670 -0.830 2.930 -0.130 ;
        RECT 3.340 -0.150 3.640 0.150 ;
        RECT 3.850 -0.150 4.150 0.150 ;
        RECT 4.430 -0.130 4.930 0.130 ;
        RECT 3.510 -0.650 3.810 -0.350 ;
        RECT 4.190 -0.650 4.490 -0.350 ;
        RECT 4.670 -0.830 4.930 -0.130 ;
        RECT 5.340 -0.150 5.640 0.150 ;
        RECT 5.850 -0.150 6.150 0.150 ;
        RECT 6.430 -0.130 6.930 0.130 ;
        RECT 5.510 -0.650 5.810 -0.350 ;
        RECT 6.190 -0.650 6.490 -0.350 ;
        RECT 6.670 -0.830 6.930 -0.130 ;
        RECT 7.340 -0.150 7.640 0.150 ;
        RECT 7.850 -0.150 8.150 0.150 ;
        RECT 8.430 -0.130 8.930 0.130 ;
        RECT 7.510 -0.650 7.810 -0.350 ;
        RECT 8.190 -0.650 8.490 -0.350 ;
        RECT 8.670 -0.830 8.930 -0.130 ;
        RECT 9.340 -0.150 9.640 0.150 ;
        RECT 9.850 -0.150 10.150 0.150 ;
        RECT 10.430 -0.130 10.930 0.130 ;
        RECT 9.510 -0.650 9.810 -0.350 ;
        RECT 10.190 -0.650 10.490 -0.350 ;
        RECT 10.670 -0.830 10.930 -0.130 ;
        RECT 11.340 -0.150 11.640 0.150 ;
        RECT 11.850 -0.150 12.150 0.150 ;
        RECT 12.430 -0.130 12.930 0.130 ;
        RECT 11.510 -0.650 11.810 -0.350 ;
        RECT 12.190 -0.650 12.490 -0.350 ;
        RECT 12.670 -0.830 12.930 -0.130 ;
        RECT 13.340 -0.150 13.640 0.150 ;
        RECT 13.850 -0.150 14.150 0.150 ;
        RECT 14.430 -0.130 14.930 0.130 ;
        RECT 13.510 -0.650 13.810 -0.350 ;
        RECT 14.190 -0.650 14.490 -0.350 ;
        RECT 14.670 -0.830 14.930 -0.130 ;
        RECT 15.340 -0.150 15.640 0.150 ;
        RECT 15.850 -0.150 16.150 0.150 ;
        RECT 16.430 -0.130 16.930 0.130 ;
        RECT 15.510 -0.650 15.810 -0.350 ;
        RECT 16.190 -0.650 16.490 -0.350 ;
        RECT 16.670 -0.830 16.930 -0.130 ;
        RECT 17.340 -0.150 17.640 0.150 ;
        RECT 17.850 -0.150 18.150 0.150 ;
        RECT 18.430 -0.130 18.930 0.130 ;
        RECT 17.510 -0.650 17.810 -0.350 ;
        RECT 18.190 -0.650 18.490 -0.350 ;
        RECT 18.670 -0.830 18.930 -0.130 ;
        RECT 19.340 -0.150 19.640 0.150 ;
        RECT 19.850 -0.150 20.150 0.150 ;
        RECT 20.430 -0.130 20.930 0.130 ;
        RECT 19.510 -0.650 19.810 -0.350 ;
        RECT 20.190 -0.650 20.490 -0.350 ;
        RECT 20.670 -0.830 20.930 -0.130 ;
        RECT 21.340 -0.150 21.640 0.150 ;
        RECT 21.850 -0.150 22.150 0.150 ;
        RECT 22.430 -0.130 22.930 0.130 ;
        RECT 21.510 -0.650 21.810 -0.350 ;
        RECT 22.190 -0.650 22.490 -0.350 ;
        RECT 22.670 -0.830 22.930 -0.130 ;
        RECT 23.340 -0.150 23.640 0.150 ;
        RECT 23.850 -0.150 24.150 0.150 ;
        RECT 24.430 -0.130 24.930 0.130 ;
        RECT 23.510 -0.650 23.810 -0.350 ;
        RECT 24.190 -0.650 24.490 -0.350 ;
        RECT 24.670 -0.830 24.930 -0.130 ;
        RECT 25.340 -0.150 25.640 0.150 ;
        RECT 25.850 -0.150 26.150 0.150 ;
        RECT 26.430 -0.130 26.930 0.130 ;
        RECT 25.510 -0.650 25.810 -0.350 ;
        RECT 26.190 -0.650 26.490 -0.350 ;
        RECT 26.670 -0.830 26.930 -0.130 ;
        RECT 27.340 -0.150 27.640 0.150 ;
        RECT 27.850 -0.150 28.150 0.150 ;
        RECT 28.430 -0.130 28.930 0.130 ;
        RECT 27.510 -0.650 27.810 -0.350 ;
        RECT 28.190 -0.650 28.490 -0.350 ;
        RECT 28.670 -0.830 28.930 -0.130 ;
        RECT 29.340 -0.150 29.640 0.150 ;
        RECT 29.850 -0.150 30.150 0.150 ;
        RECT 30.430 -0.130 30.930 0.130 ;
        RECT 29.510 -0.650 29.810 -0.350 ;
        RECT 30.190 -0.650 30.490 -0.350 ;
        RECT 30.670 -0.830 30.930 -0.130 ;
        RECT 31.340 -0.150 31.640 0.150 ;
        RECT 31.850 -0.150 32.150 0.150 ;
        RECT 32.430 -0.130 32.930 0.130 ;
        RECT 31.510 -0.650 31.810 -0.350 ;
        RECT 32.190 -0.650 32.490 -0.350 ;
        RECT 32.670 -0.830 32.930 -0.130 ;
        RECT 33.340 -0.150 33.640 0.150 ;
        RECT 33.850 -0.150 34.150 0.150 ;
        RECT 34.430 -0.130 34.930 0.130 ;
        RECT 33.510 -0.650 33.810 -0.350 ;
        RECT 34.190 -0.650 34.490 -0.350 ;
        RECT 34.670 -0.830 34.930 -0.130 ;
        RECT 35.340 -0.150 35.640 0.150 ;
        RECT 35.850 -0.150 36.150 0.150 ;
        RECT 36.430 -0.130 36.930 0.130 ;
        RECT 35.510 -0.650 35.810 -0.350 ;
        RECT 36.190 -0.650 36.490 -0.350 ;
        RECT 36.670 -0.830 36.930 -0.130 ;
        RECT 37.340 -0.150 37.640 0.150 ;
        RECT 37.850 -0.150 38.150 0.150 ;
        RECT 38.430 -0.130 38.930 0.130 ;
        RECT 37.510 -0.650 37.810 -0.350 ;
        RECT 38.190 -0.650 38.490 -0.350 ;
        RECT 38.670 -0.830 38.930 -0.130 ;
        RECT 39.340 -0.150 39.640 0.150 ;
        RECT 39.850 -0.150 40.150 0.150 ;
        RECT 40.430 -0.130 40.930 0.130 ;
        RECT 39.510 -0.650 39.810 -0.350 ;
        RECT 40.190 -0.650 40.490 -0.350 ;
        RECT 40.670 -0.830 40.930 -0.130 ;
        RECT 41.340 -0.150 41.640 0.150 ;
        RECT 41.850 -0.150 42.150 0.150 ;
        RECT 42.430 -0.130 42.930 0.130 ;
        RECT 41.510 -0.650 41.810 -0.350 ;
        RECT 42.190 -0.650 42.490 -0.350 ;
        RECT 42.670 -0.830 42.930 -0.130 ;
        RECT 43.340 -0.150 43.640 0.150 ;
        RECT 43.850 -0.150 44.150 0.150 ;
        RECT 44.430 -0.130 44.930 0.130 ;
        RECT 43.510 -0.650 43.810 -0.350 ;
        RECT 44.190 -0.650 44.490 -0.350 ;
        RECT 44.670 -0.830 44.930 -0.130 ;
        RECT 45.340 -0.150 45.640 0.150 ;
        RECT 45.850 -0.150 46.150 0.150 ;
        RECT 46.430 -0.130 46.930 0.130 ;
        RECT 45.510 -0.650 45.810 -0.350 ;
        RECT 46.190 -0.650 46.490 -0.350 ;
        RECT 46.670 -0.830 46.930 -0.130 ;
        RECT 47.340 -0.150 47.640 0.150 ;
        RECT 47.850 -0.150 48.150 0.150 ;
        RECT 48.430 -0.130 48.930 0.130 ;
        RECT 47.510 -0.650 47.810 -0.350 ;
        RECT 48.190 -0.650 48.490 -0.350 ;
        RECT 48.670 -0.830 48.930 -0.130 ;
        RECT 49.340 -0.150 49.640 0.150 ;
        RECT 49.850 -0.150 50.150 0.150 ;
        RECT 50.430 -0.130 50.930 0.130 ;
        RECT 49.510 -0.650 49.810 -0.350 ;
        RECT 50.190 -0.650 50.490 -0.350 ;
        RECT 50.670 -0.830 50.930 -0.130 ;
        RECT 51.340 -0.150 51.640 0.150 ;
        RECT 51.850 -0.150 52.150 0.150 ;
        RECT 52.430 -0.130 52.930 0.130 ;
        RECT 51.510 -0.650 51.810 -0.350 ;
        RECT 52.190 -0.650 52.490 -0.350 ;
        RECT 52.670 -0.830 52.930 -0.130 ;
        RECT 53.340 -0.150 53.640 0.150 ;
        RECT 53.850 -0.150 54.150 0.150 ;
        RECT 54.430 -0.130 54.930 0.130 ;
        RECT 53.510 -0.650 53.810 -0.350 ;
        RECT 54.190 -0.650 54.490 -0.350 ;
        RECT 54.670 -0.830 54.930 -0.130 ;
        RECT 55.340 -0.150 55.640 0.150 ;
        RECT 55.850 -0.150 56.150 0.150 ;
        RECT 56.430 -0.130 56.930 0.130 ;
        RECT 55.510 -0.650 55.810 -0.350 ;
        RECT 56.190 -0.650 56.490 -0.350 ;
        RECT 56.670 -0.830 56.930 -0.130 ;
        RECT 57.340 -0.150 57.640 0.150 ;
        RECT 57.850 -0.150 58.150 0.150 ;
        RECT 58.430 -0.130 58.930 0.130 ;
        RECT 57.510 -0.650 57.810 -0.350 ;
        RECT 58.190 -0.650 58.490 -0.350 ;
        RECT 58.670 -0.830 58.930 -0.130 ;
        RECT 59.340 -0.150 59.640 0.150 ;
        RECT 59.850 -0.150 60.150 0.150 ;
        RECT 60.430 -0.130 60.930 0.130 ;
        RECT 59.510 -0.650 59.810 -0.350 ;
        RECT 60.190 -0.650 60.490 -0.350 ;
        RECT 60.670 -0.830 60.930 -0.130 ;
        RECT 61.340 -0.150 61.640 0.150 ;
        RECT 61.850 -0.150 62.150 0.150 ;
        RECT 62.430 -0.130 62.930 0.130 ;
        RECT 61.510 -0.650 61.810 -0.350 ;
        RECT 62.190 -0.650 62.490 -0.350 ;
        RECT 62.670 -0.830 62.930 -0.130 ;
        RECT 63.340 -0.150 63.640 0.150 ;
        RECT 63.850 -0.150 64.150 0.150 ;
        RECT 64.430 -0.130 64.930 0.130 ;
        RECT 63.510 -0.650 63.810 -0.350 ;
        RECT 64.190 -0.650 64.490 -0.350 ;
        RECT 64.670 -0.830 64.930 -0.130 ;
        RECT 65.340 -0.150 65.640 0.150 ;
        RECT 65.850 -0.150 66.150 0.150 ;
        RECT 66.430 -0.130 66.930 0.130 ;
        RECT 65.510 -0.650 65.810 -0.350 ;
        RECT 66.190 -0.650 66.490 -0.350 ;
        RECT 66.670 -0.830 66.930 -0.130 ;
        RECT 67.340 -0.150 67.640 0.150 ;
        RECT 67.850 -0.150 68.150 0.150 ;
        RECT 68.430 -0.130 68.930 0.130 ;
        RECT 67.510 -0.650 67.810 -0.350 ;
        RECT 68.190 -0.650 68.490 -0.350 ;
        RECT 68.670 -0.830 68.930 -0.130 ;
        RECT 69.340 -0.150 69.640 0.150 ;
        RECT 69.850 -0.150 70.150 0.150 ;
        RECT 70.430 -0.130 70.930 0.130 ;
        RECT 69.510 -0.650 69.810 -0.350 ;
        RECT 70.190 -0.650 70.490 -0.350 ;
        RECT 70.670 -0.830 70.930 -0.130 ;
        RECT 71.340 -0.150 71.640 0.150 ;
        RECT 71.850 -0.150 72.150 0.150 ;
        RECT 72.430 -0.130 72.930 0.130 ;
        RECT 71.510 -0.650 71.810 -0.350 ;
        RECT 72.190 -0.650 72.490 -0.350 ;
        RECT 72.670 -0.830 72.930 -0.130 ;
        RECT 73.340 -0.150 73.640 0.150 ;
        RECT 73.850 -0.150 74.150 0.150 ;
        RECT 74.430 -0.130 74.930 0.130 ;
        RECT 73.510 -0.650 73.810 -0.350 ;
        RECT 74.190 -0.650 74.490 -0.350 ;
        RECT 74.670 -0.830 74.930 -0.130 ;
        RECT 75.340 -0.150 75.640 0.150 ;
        RECT 75.850 -0.150 76.150 0.150 ;
        RECT 76.430 -0.130 76.930 0.130 ;
        RECT 75.510 -0.650 75.810 -0.350 ;
        RECT 76.190 -0.650 76.490 -0.350 ;
        RECT 76.670 -0.830 76.930 -0.130 ;
        RECT 77.340 -0.150 77.640 0.150 ;
        RECT 77.850 -0.150 78.150 0.150 ;
        RECT 78.430 -0.130 78.930 0.130 ;
        RECT 77.510 -0.650 77.810 -0.350 ;
        RECT 78.190 -0.650 78.490 -0.350 ;
        RECT 78.670 -0.830 78.930 -0.130 ;
        RECT 79.340 -0.150 79.640 0.150 ;
        RECT 79.850 -0.150 80.150 0.150 ;
        RECT 80.430 -0.130 80.930 0.130 ;
        RECT 79.510 -0.650 79.810 -0.350 ;
        RECT 80.190 -0.650 80.490 -0.350 ;
        RECT 80.670 -0.830 80.930 -0.130 ;
        RECT 81.340 -0.150 81.640 0.150 ;
        RECT 81.850 -0.150 82.150 0.150 ;
        RECT 82.430 -0.130 82.930 0.130 ;
        RECT 81.510 -0.650 81.810 -0.350 ;
        RECT 82.190 -0.650 82.490 -0.350 ;
        RECT 82.670 -0.830 82.930 -0.130 ;
        RECT 83.340 -0.150 83.640 0.150 ;
        RECT 83.850 -0.150 84.150 0.150 ;
        RECT 84.430 -0.130 84.930 0.130 ;
        RECT 83.510 -0.650 83.810 -0.350 ;
        RECT 84.190 -0.650 84.490 -0.350 ;
        RECT 84.670 -0.830 84.930 -0.130 ;
        RECT 85.340 -0.150 85.640 0.150 ;
        RECT 85.850 -0.150 86.150 0.150 ;
        RECT 86.430 -0.130 86.930 0.130 ;
        RECT 85.510 -0.650 85.810 -0.350 ;
        RECT 86.190 -0.650 86.490 -0.350 ;
        RECT 86.670 -0.830 86.930 -0.130 ;
        RECT 87.340 -0.150 87.640 0.150 ;
        RECT 87.850 -0.150 88.150 0.150 ;
        RECT 88.430 -0.130 88.930 0.130 ;
        RECT 87.510 -0.650 87.810 -0.350 ;
        RECT 88.190 -0.650 88.490 -0.350 ;
        RECT 88.670 -0.830 88.930 -0.130 ;
        RECT 89.340 -0.150 89.640 0.150 ;
        RECT 89.850 -0.150 90.150 0.150 ;
        RECT 90.430 -0.130 90.930 0.130 ;
        RECT 89.510 -0.650 89.810 -0.350 ;
        RECT 90.190 -0.650 90.490 -0.350 ;
        RECT 90.670 -0.830 90.930 -0.130 ;
        RECT 91.340 -0.150 91.640 0.150 ;
        RECT 91.850 -0.150 92.150 0.150 ;
        RECT 92.430 -0.130 92.930 0.130 ;
        RECT 91.510 -0.650 91.810 -0.350 ;
        RECT 92.190 -0.650 92.490 -0.350 ;
        RECT 92.670 -0.830 92.930 -0.130 ;
        RECT 93.340 -0.150 93.640 0.150 ;
        RECT 93.850 -0.150 94.150 0.150 ;
        RECT 94.430 -0.130 94.930 0.130 ;
        RECT 93.510 -0.650 93.810 -0.350 ;
        RECT 94.190 -0.650 94.490 -0.350 ;
        RECT 94.670 -0.830 94.930 -0.130 ;
        RECT 95.340 -0.150 95.640 0.150 ;
        RECT 95.850 -0.150 96.150 0.150 ;
        RECT 96.430 -0.130 96.930 0.130 ;
        RECT 95.510 -0.650 95.810 -0.350 ;
        RECT 96.190 -0.650 96.490 -0.350 ;
        RECT 96.670 -0.830 96.930 -0.130 ;
        RECT 97.340 -0.150 97.640 0.150 ;
        RECT 97.850 -0.150 98.150 0.150 ;
        RECT 98.430 -0.130 98.930 0.130 ;
        RECT 97.510 -0.650 97.810 -0.350 ;
        RECT 98.190 -0.650 98.490 -0.350 ;
        RECT 98.670 -0.830 98.930 -0.130 ;
        RECT 99.340 -0.150 99.640 0.150 ;
        RECT 99.850 -0.150 100.150 0.150 ;
        RECT 100.430 -0.130 100.930 0.130 ;
        RECT 99.510 -0.650 99.810 -0.350 ;
        RECT 100.190 -0.650 100.490 -0.350 ;
        RECT 100.670 -0.830 100.930 -0.130 ;
        RECT 101.340 -0.150 101.640 0.150 ;
        RECT 101.850 -0.150 102.150 0.150 ;
        RECT 102.430 -0.130 102.930 0.130 ;
        RECT 101.510 -0.650 101.810 -0.350 ;
        RECT 102.190 -0.650 102.490 -0.350 ;
        RECT 102.670 -0.830 102.930 -0.130 ;
        RECT 103.340 -0.150 103.640 0.150 ;
        RECT 103.850 -0.150 104.150 0.150 ;
        RECT 104.430 -0.130 104.930 0.130 ;
        RECT 103.510 -0.650 103.810 -0.350 ;
        RECT 104.190 -0.650 104.490 -0.350 ;
        RECT 104.670 -0.830 104.930 -0.130 ;
        RECT 105.340 -0.150 105.640 0.150 ;
        RECT 105.850 -0.150 106.150 0.150 ;
        RECT 106.430 -0.130 106.930 0.130 ;
        RECT 105.510 -0.650 105.810 -0.350 ;
        RECT 106.190 -0.650 106.490 -0.350 ;
        RECT 106.670 -0.830 106.930 -0.130 ;
        RECT 107.340 -0.150 107.640 0.150 ;
        RECT 107.850 -0.150 108.150 0.150 ;
        RECT 108.430 -0.130 108.930 0.130 ;
        RECT 107.510 -0.650 107.810 -0.350 ;
        RECT 108.190 -0.650 108.490 -0.350 ;
        RECT 108.670 -0.830 108.930 -0.130 ;
        RECT 109.340 -0.150 109.640 0.150 ;
        RECT 109.850 -0.150 110.150 0.150 ;
        RECT 110.430 -0.130 110.930 0.130 ;
        RECT 109.510 -0.650 109.810 -0.350 ;
        RECT 110.190 -0.650 110.490 -0.350 ;
        RECT 110.670 -0.830 110.930 -0.130 ;
        RECT 111.340 -0.150 111.640 0.150 ;
        RECT 111.850 -0.150 112.150 0.150 ;
        RECT 112.430 -0.130 112.930 0.130 ;
        RECT 111.510 -0.650 111.810 -0.350 ;
        RECT 112.190 -0.650 112.490 -0.350 ;
        RECT 112.670 -0.830 112.930 -0.130 ;
        RECT 113.340 -0.150 113.640 0.150 ;
        RECT 113.850 -0.150 114.150 0.150 ;
        RECT 114.430 -0.130 114.930 0.130 ;
        RECT 113.510 -0.650 113.810 -0.350 ;
        RECT 114.190 -0.650 114.490 -0.350 ;
        RECT 114.670 -0.830 114.930 -0.130 ;
        RECT 115.340 -0.150 115.640 0.150 ;
        RECT 115.850 -0.150 116.150 0.150 ;
        RECT 116.430 -0.130 116.930 0.130 ;
        RECT 115.510 -0.650 115.810 -0.350 ;
        RECT 116.190 -0.650 116.490 -0.350 ;
        RECT 116.670 -0.830 116.930 -0.130 ;
        RECT 117.340 -0.150 117.640 0.150 ;
        RECT 117.850 -0.150 118.150 0.150 ;
        RECT 118.430 -0.130 118.930 0.130 ;
        RECT 117.510 -0.650 117.810 -0.350 ;
        RECT 118.190 -0.650 118.490 -0.350 ;
        RECT 118.670 -0.830 118.930 -0.130 ;
        RECT 119.340 -0.150 119.640 0.150 ;
        RECT 119.850 -0.150 120.150 0.150 ;
        RECT 120.430 -0.130 120.930 0.130 ;
        RECT 119.510 -0.650 119.810 -0.350 ;
        RECT 120.190 -0.650 120.490 -0.350 ;
        RECT 120.670 -0.830 120.930 -0.130 ;
        RECT 121.340 -0.150 121.640 0.150 ;
        RECT 121.850 -0.150 122.150 0.150 ;
        RECT 122.430 -0.130 122.930 0.130 ;
        RECT 121.510 -0.650 121.810 -0.350 ;
        RECT 122.190 -0.650 122.490 -0.350 ;
        RECT 122.670 -0.830 122.930 -0.130 ;
        RECT 123.340 -0.150 123.640 0.150 ;
        RECT 123.850 -0.150 124.150 0.150 ;
        RECT 124.430 -0.130 124.930 0.130 ;
        RECT 123.510 -0.650 123.810 -0.350 ;
        RECT 124.190 -0.650 124.490 -0.350 ;
        RECT 124.670 -0.830 124.930 -0.130 ;
        RECT 125.340 -0.150 125.640 0.150 ;
        RECT 125.850 -0.150 126.150 0.150 ;
        RECT 126.430 -0.130 126.930 0.130 ;
        RECT 125.510 -0.650 125.810 -0.350 ;
        RECT 126.190 -0.650 126.490 -0.350 ;
        RECT 126.670 -0.830 126.930 -0.130 ;
        RECT 127.340 -0.150 127.640 0.150 ;
        RECT 127.850 -0.150 128.150 0.150 ;
        RECT 128.430 -0.130 128.930 0.130 ;
        RECT 127.510 -0.650 127.810 -0.350 ;
        RECT 128.190 -0.650 128.490 -0.350 ;
        RECT 128.670 -0.830 128.930 -0.130 ;
        RECT 129.340 -0.150 129.640 0.150 ;
        RECT 129.850 -0.150 130.150 0.150 ;
        RECT 130.430 -0.130 130.930 0.130 ;
        RECT 129.510 -0.650 129.810 -0.350 ;
        RECT 130.190 -0.650 130.490 -0.350 ;
        RECT 130.670 -0.830 130.930 -0.130 ;
        RECT -0.890 -2.000 -0.600 -1.710 ;
        RECT -0.825 -3.130 -0.665 -2.000 ;
        RECT -0.080 -2.010 0.080 -1.330 ;
        RECT 0.600 -2.000 0.890 -1.710 ;
        RECT 1.110 -2.000 1.400 -1.710 ;
        RECT -0.420 -2.190 -0.260 -2.120 ;
        RECT 0.260 -2.190 0.420 -2.120 ;
        RECT -0.420 -2.480 -0.130 -2.190 ;
        RECT 0.130 -2.480 0.420 -2.190 ;
        RECT -0.825 -3.290 0.425 -3.130 ;
        RECT -0.825 -4.110 -0.665 -3.290 ;
        RECT -0.080 -4.410 0.080 -3.850 ;
        RECT 0.665 -4.110 0.825 -2.000 ;
        RECT 1.175 -3.130 1.335 -2.000 ;
        RECT 1.920 -2.010 2.080 -1.330 ;
        RECT 2.600 -2.000 2.890 -1.710 ;
        RECT 3.110 -2.000 3.400 -1.710 ;
        RECT 1.580 -2.190 1.740 -2.120 ;
        RECT 2.260 -2.190 2.420 -2.120 ;
        RECT 1.580 -2.480 1.870 -2.190 ;
        RECT 2.130 -2.480 2.420 -2.190 ;
        RECT 1.175 -3.290 2.425 -3.130 ;
        RECT 1.175 -4.110 1.335 -3.290 ;
        RECT 1.920 -4.410 2.080 -3.850 ;
        RECT 2.665 -4.110 2.825 -2.000 ;
        RECT 3.175 -3.130 3.335 -2.000 ;
        RECT 3.920 -2.010 4.080 -1.330 ;
        RECT 4.600 -2.000 4.890 -1.710 ;
        RECT 5.110 -2.000 5.400 -1.710 ;
        RECT 3.580 -2.190 3.740 -2.120 ;
        RECT 4.260 -2.190 4.420 -2.120 ;
        RECT 3.580 -2.480 3.870 -2.190 ;
        RECT 4.130 -2.480 4.420 -2.190 ;
        RECT 3.175 -3.290 4.425 -3.130 ;
        RECT 3.175 -4.110 3.335 -3.290 ;
        RECT 3.920 -4.410 4.080 -3.850 ;
        RECT 4.665 -4.110 4.825 -2.000 ;
        RECT 5.175 -3.130 5.335 -2.000 ;
        RECT 5.920 -2.010 6.080 -1.330 ;
        RECT 6.600 -2.000 6.890 -1.710 ;
        RECT 7.110 -2.000 7.400 -1.710 ;
        RECT 5.580 -2.190 5.740 -2.120 ;
        RECT 6.260 -2.190 6.420 -2.120 ;
        RECT 5.580 -2.480 5.870 -2.190 ;
        RECT 6.130 -2.480 6.420 -2.190 ;
        RECT 5.175 -3.290 6.425 -3.130 ;
        RECT 5.175 -4.110 5.335 -3.290 ;
        RECT 5.920 -4.410 6.080 -3.850 ;
        RECT 6.665 -4.110 6.825 -2.000 ;
        RECT 7.175 -3.130 7.335 -2.000 ;
        RECT 7.920 -2.010 8.080 -1.330 ;
        RECT 8.600 -2.000 8.890 -1.710 ;
        RECT 9.110 -2.000 9.400 -1.710 ;
        RECT 7.580 -2.190 7.740 -2.120 ;
        RECT 8.260 -2.190 8.420 -2.120 ;
        RECT 7.580 -2.480 7.870 -2.190 ;
        RECT 8.130 -2.480 8.420 -2.190 ;
        RECT 7.175 -3.290 8.425 -3.130 ;
        RECT 7.175 -4.110 7.335 -3.290 ;
        RECT 7.920 -4.410 8.080 -3.850 ;
        RECT 8.665 -4.110 8.825 -2.000 ;
        RECT 9.175 -3.130 9.335 -2.000 ;
        RECT 9.920 -2.010 10.080 -1.330 ;
        RECT 10.600 -2.000 10.890 -1.710 ;
        RECT 11.110 -2.000 11.400 -1.710 ;
        RECT 9.580 -2.190 9.740 -2.120 ;
        RECT 10.260 -2.190 10.420 -2.120 ;
        RECT 9.580 -2.480 9.870 -2.190 ;
        RECT 10.130 -2.480 10.420 -2.190 ;
        RECT 9.175 -3.290 10.425 -3.130 ;
        RECT 9.175 -4.110 9.335 -3.290 ;
        RECT 9.920 -4.410 10.080 -3.850 ;
        RECT 10.665 -4.110 10.825 -2.000 ;
        RECT 11.175 -3.130 11.335 -2.000 ;
        RECT 11.920 -2.010 12.080 -1.330 ;
        RECT 12.600 -2.000 12.890 -1.710 ;
        RECT 13.110 -2.000 13.400 -1.710 ;
        RECT 11.580 -2.190 11.740 -2.120 ;
        RECT 12.260 -2.190 12.420 -2.120 ;
        RECT 11.580 -2.480 11.870 -2.190 ;
        RECT 12.130 -2.480 12.420 -2.190 ;
        RECT 11.175 -3.290 12.425 -3.130 ;
        RECT 11.175 -4.110 11.335 -3.290 ;
        RECT 11.920 -4.410 12.080 -3.850 ;
        RECT 12.665 -4.110 12.825 -2.000 ;
        RECT 13.175 -3.130 13.335 -2.000 ;
        RECT 13.920 -2.010 14.080 -1.330 ;
        RECT 14.600 -2.000 14.890 -1.710 ;
        RECT 15.110 -2.000 15.400 -1.710 ;
        RECT 13.580 -2.190 13.740 -2.120 ;
        RECT 14.260 -2.190 14.420 -2.120 ;
        RECT 13.580 -2.480 13.870 -2.190 ;
        RECT 14.130 -2.480 14.420 -2.190 ;
        RECT 13.175 -3.290 14.425 -3.130 ;
        RECT 13.175 -4.110 13.335 -3.290 ;
        RECT 13.920 -4.410 14.080 -3.850 ;
        RECT 14.665 -4.110 14.825 -2.000 ;
        RECT 15.175 -3.130 15.335 -2.000 ;
        RECT 15.920 -2.010 16.080 -1.330 ;
        RECT 16.600 -2.000 16.890 -1.710 ;
        RECT 17.110 -2.000 17.400 -1.710 ;
        RECT 15.580 -2.190 15.740 -2.120 ;
        RECT 16.260 -2.190 16.420 -2.120 ;
        RECT 15.580 -2.480 15.870 -2.190 ;
        RECT 16.130 -2.480 16.420 -2.190 ;
        RECT 15.175 -3.290 16.425 -3.130 ;
        RECT 15.175 -4.110 15.335 -3.290 ;
        RECT 15.920 -4.410 16.080 -3.850 ;
        RECT 16.665 -4.110 16.825 -2.000 ;
        RECT 17.175 -3.130 17.335 -2.000 ;
        RECT 17.920 -2.010 18.080 -1.330 ;
        RECT 18.600 -2.000 18.890 -1.710 ;
        RECT 19.110 -2.000 19.400 -1.710 ;
        RECT 17.580 -2.190 17.740 -2.120 ;
        RECT 18.260 -2.190 18.420 -2.120 ;
        RECT 17.580 -2.480 17.870 -2.190 ;
        RECT 18.130 -2.480 18.420 -2.190 ;
        RECT 17.175 -3.290 18.425 -3.130 ;
        RECT 17.175 -4.110 17.335 -3.290 ;
        RECT 17.920 -4.410 18.080 -3.850 ;
        RECT 18.665 -4.110 18.825 -2.000 ;
        RECT 19.175 -3.130 19.335 -2.000 ;
        RECT 19.920 -2.010 20.080 -1.330 ;
        RECT 20.600 -2.000 20.890 -1.710 ;
        RECT 21.110 -2.000 21.400 -1.710 ;
        RECT 19.580 -2.190 19.740 -2.120 ;
        RECT 20.260 -2.190 20.420 -2.120 ;
        RECT 19.580 -2.480 19.870 -2.190 ;
        RECT 20.130 -2.480 20.420 -2.190 ;
        RECT 19.175 -3.290 20.425 -3.130 ;
        RECT 19.175 -4.110 19.335 -3.290 ;
        RECT 19.920 -4.410 20.080 -3.850 ;
        RECT 20.665 -4.110 20.825 -2.000 ;
        RECT 21.175 -3.130 21.335 -2.000 ;
        RECT 21.920 -2.010 22.080 -1.330 ;
        RECT 22.600 -2.000 22.890 -1.710 ;
        RECT 23.110 -2.000 23.400 -1.710 ;
        RECT 21.580 -2.190 21.740 -2.120 ;
        RECT 22.260 -2.190 22.420 -2.120 ;
        RECT 21.580 -2.480 21.870 -2.190 ;
        RECT 22.130 -2.480 22.420 -2.190 ;
        RECT 21.175 -3.290 22.425 -3.130 ;
        RECT 21.175 -4.110 21.335 -3.290 ;
        RECT 21.920 -4.410 22.080 -3.850 ;
        RECT 22.665 -4.110 22.825 -2.000 ;
        RECT 23.175 -3.130 23.335 -2.000 ;
        RECT 23.920 -2.010 24.080 -1.330 ;
        RECT 24.600 -2.000 24.890 -1.710 ;
        RECT 25.110 -2.000 25.400 -1.710 ;
        RECT 23.580 -2.190 23.740 -2.120 ;
        RECT 24.260 -2.190 24.420 -2.120 ;
        RECT 23.580 -2.480 23.870 -2.190 ;
        RECT 24.130 -2.480 24.420 -2.190 ;
        RECT 23.175 -3.290 24.425 -3.130 ;
        RECT 23.175 -4.110 23.335 -3.290 ;
        RECT 23.920 -4.410 24.080 -3.850 ;
        RECT 24.665 -4.110 24.825 -2.000 ;
        RECT 25.175 -3.130 25.335 -2.000 ;
        RECT 25.920 -2.010 26.080 -1.330 ;
        RECT 26.600 -2.000 26.890 -1.710 ;
        RECT 27.110 -2.000 27.400 -1.710 ;
        RECT 25.580 -2.190 25.740 -2.120 ;
        RECT 26.260 -2.190 26.420 -2.120 ;
        RECT 25.580 -2.480 25.870 -2.190 ;
        RECT 26.130 -2.480 26.420 -2.190 ;
        RECT 25.175 -3.290 26.425 -3.130 ;
        RECT 25.175 -4.110 25.335 -3.290 ;
        RECT 25.920 -4.410 26.080 -3.850 ;
        RECT 26.665 -4.110 26.825 -2.000 ;
        RECT 27.175 -3.130 27.335 -2.000 ;
        RECT 27.920 -2.010 28.080 -1.330 ;
        RECT 28.600 -2.000 28.890 -1.710 ;
        RECT 29.110 -2.000 29.400 -1.710 ;
        RECT 27.580 -2.190 27.740 -2.120 ;
        RECT 28.260 -2.190 28.420 -2.120 ;
        RECT 27.580 -2.480 27.870 -2.190 ;
        RECT 28.130 -2.480 28.420 -2.190 ;
        RECT 27.175 -3.290 28.425 -3.130 ;
        RECT 27.175 -4.110 27.335 -3.290 ;
        RECT 27.920 -4.410 28.080 -3.850 ;
        RECT 28.665 -4.110 28.825 -2.000 ;
        RECT 29.175 -3.130 29.335 -2.000 ;
        RECT 29.920 -2.010 30.080 -1.330 ;
        RECT 30.600 -2.000 30.890 -1.710 ;
        RECT 31.110 -2.000 31.400 -1.710 ;
        RECT 29.580 -2.190 29.740 -2.120 ;
        RECT 30.260 -2.190 30.420 -2.120 ;
        RECT 29.580 -2.480 29.870 -2.190 ;
        RECT 30.130 -2.480 30.420 -2.190 ;
        RECT 29.175 -3.290 30.425 -3.130 ;
        RECT 29.175 -4.110 29.335 -3.290 ;
        RECT 29.920 -4.410 30.080 -3.850 ;
        RECT 30.665 -4.110 30.825 -2.000 ;
        RECT 31.175 -3.130 31.335 -2.000 ;
        RECT 31.920 -2.010 32.080 -1.330 ;
        RECT 32.600 -2.000 32.890 -1.710 ;
        RECT 33.110 -2.000 33.400 -1.710 ;
        RECT 31.580 -2.190 31.740 -2.120 ;
        RECT 32.260 -2.190 32.420 -2.120 ;
        RECT 31.580 -2.480 31.870 -2.190 ;
        RECT 32.130 -2.480 32.420 -2.190 ;
        RECT 31.175 -3.290 32.425 -3.130 ;
        RECT 31.175 -4.110 31.335 -3.290 ;
        RECT 31.920 -4.410 32.080 -3.850 ;
        RECT 32.665 -4.110 32.825 -2.000 ;
        RECT 33.175 -3.130 33.335 -2.000 ;
        RECT 33.920 -2.010 34.080 -1.330 ;
        RECT 34.600 -2.000 34.890 -1.710 ;
        RECT 35.110 -2.000 35.400 -1.710 ;
        RECT 33.580 -2.190 33.740 -2.120 ;
        RECT 34.260 -2.190 34.420 -2.120 ;
        RECT 33.580 -2.480 33.870 -2.190 ;
        RECT 34.130 -2.480 34.420 -2.190 ;
        RECT 33.175 -3.290 34.425 -3.130 ;
        RECT 33.175 -4.110 33.335 -3.290 ;
        RECT 33.920 -4.410 34.080 -3.850 ;
        RECT 34.665 -4.110 34.825 -2.000 ;
        RECT 35.175 -3.130 35.335 -2.000 ;
        RECT 35.920 -2.010 36.080 -1.330 ;
        RECT 36.600 -2.000 36.890 -1.710 ;
        RECT 37.110 -2.000 37.400 -1.710 ;
        RECT 35.580 -2.190 35.740 -2.120 ;
        RECT 36.260 -2.190 36.420 -2.120 ;
        RECT 35.580 -2.480 35.870 -2.190 ;
        RECT 36.130 -2.480 36.420 -2.190 ;
        RECT 35.175 -3.290 36.425 -3.130 ;
        RECT 35.175 -4.110 35.335 -3.290 ;
        RECT 35.920 -4.410 36.080 -3.850 ;
        RECT 36.665 -4.110 36.825 -2.000 ;
        RECT 37.175 -3.130 37.335 -2.000 ;
        RECT 37.920 -2.010 38.080 -1.330 ;
        RECT 38.600 -2.000 38.890 -1.710 ;
        RECT 39.110 -2.000 39.400 -1.710 ;
        RECT 37.580 -2.190 37.740 -2.120 ;
        RECT 38.260 -2.190 38.420 -2.120 ;
        RECT 37.580 -2.480 37.870 -2.190 ;
        RECT 38.130 -2.480 38.420 -2.190 ;
        RECT 37.175 -3.290 38.425 -3.130 ;
        RECT 37.175 -4.110 37.335 -3.290 ;
        RECT 37.920 -4.410 38.080 -3.850 ;
        RECT 38.665 -4.110 38.825 -2.000 ;
        RECT 39.175 -3.130 39.335 -2.000 ;
        RECT 39.920 -2.010 40.080 -1.330 ;
        RECT 40.600 -2.000 40.890 -1.710 ;
        RECT 41.110 -2.000 41.400 -1.710 ;
        RECT 39.580 -2.190 39.740 -2.120 ;
        RECT 40.260 -2.190 40.420 -2.120 ;
        RECT 39.580 -2.480 39.870 -2.190 ;
        RECT 40.130 -2.480 40.420 -2.190 ;
        RECT 39.175 -3.290 40.425 -3.130 ;
        RECT 39.175 -4.110 39.335 -3.290 ;
        RECT 39.920 -4.410 40.080 -3.850 ;
        RECT 40.665 -4.110 40.825 -2.000 ;
        RECT 41.175 -3.130 41.335 -2.000 ;
        RECT 41.920 -2.010 42.080 -1.330 ;
        RECT 42.600 -2.000 42.890 -1.710 ;
        RECT 43.110 -2.000 43.400 -1.710 ;
        RECT 41.580 -2.190 41.740 -2.120 ;
        RECT 42.260 -2.190 42.420 -2.120 ;
        RECT 41.580 -2.480 41.870 -2.190 ;
        RECT 42.130 -2.480 42.420 -2.190 ;
        RECT 41.175 -3.290 42.425 -3.130 ;
        RECT 41.175 -4.110 41.335 -3.290 ;
        RECT 41.920 -4.410 42.080 -3.850 ;
        RECT 42.665 -4.110 42.825 -2.000 ;
        RECT 43.175 -3.130 43.335 -2.000 ;
        RECT 43.920 -2.010 44.080 -1.330 ;
        RECT 44.600 -2.000 44.890 -1.710 ;
        RECT 45.110 -2.000 45.400 -1.710 ;
        RECT 43.580 -2.190 43.740 -2.120 ;
        RECT 44.260 -2.190 44.420 -2.120 ;
        RECT 43.580 -2.480 43.870 -2.190 ;
        RECT 44.130 -2.480 44.420 -2.190 ;
        RECT 43.175 -3.290 44.425 -3.130 ;
        RECT 43.175 -4.110 43.335 -3.290 ;
        RECT 43.920 -4.410 44.080 -3.850 ;
        RECT 44.665 -4.110 44.825 -2.000 ;
        RECT 45.175 -3.130 45.335 -2.000 ;
        RECT 45.920 -2.010 46.080 -1.330 ;
        RECT 46.600 -2.000 46.890 -1.710 ;
        RECT 47.110 -2.000 47.400 -1.710 ;
        RECT 45.580 -2.190 45.740 -2.120 ;
        RECT 46.260 -2.190 46.420 -2.120 ;
        RECT 45.580 -2.480 45.870 -2.190 ;
        RECT 46.130 -2.480 46.420 -2.190 ;
        RECT 45.175 -3.290 46.425 -3.130 ;
        RECT 45.175 -4.110 45.335 -3.290 ;
        RECT 45.920 -4.410 46.080 -3.850 ;
        RECT 46.665 -4.110 46.825 -2.000 ;
        RECT 47.175 -3.130 47.335 -2.000 ;
        RECT 47.920 -2.010 48.080 -1.330 ;
        RECT 48.600 -2.000 48.890 -1.710 ;
        RECT 49.110 -2.000 49.400 -1.710 ;
        RECT 47.580 -2.190 47.740 -2.120 ;
        RECT 48.260 -2.190 48.420 -2.120 ;
        RECT 47.580 -2.480 47.870 -2.190 ;
        RECT 48.130 -2.480 48.420 -2.190 ;
        RECT 47.175 -3.290 48.425 -3.130 ;
        RECT 47.175 -4.110 47.335 -3.290 ;
        RECT 47.920 -4.410 48.080 -3.850 ;
        RECT 48.665 -4.110 48.825 -2.000 ;
        RECT 49.175 -3.130 49.335 -2.000 ;
        RECT 49.920 -2.010 50.080 -1.330 ;
        RECT 50.600 -2.000 50.890 -1.710 ;
        RECT 51.110 -2.000 51.400 -1.710 ;
        RECT 49.580 -2.190 49.740 -2.120 ;
        RECT 50.260 -2.190 50.420 -2.120 ;
        RECT 49.580 -2.480 49.870 -2.190 ;
        RECT 50.130 -2.480 50.420 -2.190 ;
        RECT 49.175 -3.290 50.425 -3.130 ;
        RECT 49.175 -4.110 49.335 -3.290 ;
        RECT 49.920 -4.410 50.080 -3.850 ;
        RECT 50.665 -4.110 50.825 -2.000 ;
        RECT 51.175 -3.130 51.335 -2.000 ;
        RECT 51.920 -2.010 52.080 -1.330 ;
        RECT 52.600 -2.000 52.890 -1.710 ;
        RECT 53.110 -2.000 53.400 -1.710 ;
        RECT 51.580 -2.190 51.740 -2.120 ;
        RECT 52.260 -2.190 52.420 -2.120 ;
        RECT 51.580 -2.480 51.870 -2.190 ;
        RECT 52.130 -2.480 52.420 -2.190 ;
        RECT 51.175 -3.290 52.425 -3.130 ;
        RECT 51.175 -4.110 51.335 -3.290 ;
        RECT 51.920 -4.410 52.080 -3.850 ;
        RECT 52.665 -4.110 52.825 -2.000 ;
        RECT 53.175 -3.130 53.335 -2.000 ;
        RECT 53.920 -2.010 54.080 -1.330 ;
        RECT 54.600 -2.000 54.890 -1.710 ;
        RECT 55.110 -2.000 55.400 -1.710 ;
        RECT 53.580 -2.190 53.740 -2.120 ;
        RECT 54.260 -2.190 54.420 -2.120 ;
        RECT 53.580 -2.480 53.870 -2.190 ;
        RECT 54.130 -2.480 54.420 -2.190 ;
        RECT 53.175 -3.290 54.425 -3.130 ;
        RECT 53.175 -4.110 53.335 -3.290 ;
        RECT 53.920 -4.410 54.080 -3.850 ;
        RECT 54.665 -4.110 54.825 -2.000 ;
        RECT 55.175 -3.130 55.335 -2.000 ;
        RECT 55.920 -2.010 56.080 -1.330 ;
        RECT 56.600 -2.000 56.890 -1.710 ;
        RECT 57.110 -2.000 57.400 -1.710 ;
        RECT 55.580 -2.190 55.740 -2.120 ;
        RECT 56.260 -2.190 56.420 -2.120 ;
        RECT 55.580 -2.480 55.870 -2.190 ;
        RECT 56.130 -2.480 56.420 -2.190 ;
        RECT 55.175 -3.290 56.425 -3.130 ;
        RECT 55.175 -4.110 55.335 -3.290 ;
        RECT 55.920 -4.410 56.080 -3.850 ;
        RECT 56.665 -4.110 56.825 -2.000 ;
        RECT 57.175 -3.130 57.335 -2.000 ;
        RECT 57.920 -2.010 58.080 -1.330 ;
        RECT 58.600 -2.000 58.890 -1.710 ;
        RECT 59.110 -2.000 59.400 -1.710 ;
        RECT 57.580 -2.190 57.740 -2.120 ;
        RECT 58.260 -2.190 58.420 -2.120 ;
        RECT 57.580 -2.480 57.870 -2.190 ;
        RECT 58.130 -2.480 58.420 -2.190 ;
        RECT 57.175 -3.290 58.425 -3.130 ;
        RECT 57.175 -4.110 57.335 -3.290 ;
        RECT 57.920 -4.410 58.080 -3.850 ;
        RECT 58.665 -4.110 58.825 -2.000 ;
        RECT 59.175 -3.130 59.335 -2.000 ;
        RECT 59.920 -2.010 60.080 -1.330 ;
        RECT 60.600 -2.000 60.890 -1.710 ;
        RECT 61.110 -2.000 61.400 -1.710 ;
        RECT 59.580 -2.190 59.740 -2.120 ;
        RECT 60.260 -2.190 60.420 -2.120 ;
        RECT 59.580 -2.480 59.870 -2.190 ;
        RECT 60.130 -2.480 60.420 -2.190 ;
        RECT 59.175 -3.290 60.425 -3.130 ;
        RECT 59.175 -4.110 59.335 -3.290 ;
        RECT 59.920 -4.410 60.080 -3.850 ;
        RECT 60.665 -4.110 60.825 -2.000 ;
        RECT 61.175 -3.130 61.335 -2.000 ;
        RECT 61.920 -2.010 62.080 -1.330 ;
        RECT 62.600 -2.000 62.890 -1.710 ;
        RECT 63.110 -2.000 63.400 -1.710 ;
        RECT 61.580 -2.190 61.740 -2.120 ;
        RECT 62.260 -2.190 62.420 -2.120 ;
        RECT 61.580 -2.480 61.870 -2.190 ;
        RECT 62.130 -2.480 62.420 -2.190 ;
        RECT 61.175 -3.290 62.425 -3.130 ;
        RECT 61.175 -4.110 61.335 -3.290 ;
        RECT 61.920 -4.410 62.080 -3.850 ;
        RECT 62.665 -4.110 62.825 -2.000 ;
        RECT 63.175 -3.130 63.335 -2.000 ;
        RECT 63.920 -2.010 64.080 -1.330 ;
        RECT 64.600 -2.000 64.890 -1.710 ;
        RECT 65.110 -2.000 65.400 -1.710 ;
        RECT 63.580 -2.190 63.740 -2.120 ;
        RECT 64.260 -2.190 64.420 -2.120 ;
        RECT 63.580 -2.480 63.870 -2.190 ;
        RECT 64.130 -2.480 64.420 -2.190 ;
        RECT 63.175 -3.290 64.425 -3.130 ;
        RECT 63.175 -4.110 63.335 -3.290 ;
        RECT 63.920 -4.410 64.080 -3.850 ;
        RECT 64.665 -4.110 64.825 -2.000 ;
        RECT 65.175 -3.130 65.335 -2.000 ;
        RECT 65.920 -2.010 66.080 -1.330 ;
        RECT 66.600 -2.000 66.890 -1.710 ;
        RECT 67.110 -2.000 67.400 -1.710 ;
        RECT 65.580 -2.190 65.740 -2.120 ;
        RECT 66.260 -2.190 66.420 -2.120 ;
        RECT 65.580 -2.480 65.870 -2.190 ;
        RECT 66.130 -2.480 66.420 -2.190 ;
        RECT 65.175 -3.290 66.425 -3.130 ;
        RECT 65.175 -4.110 65.335 -3.290 ;
        RECT 65.920 -4.410 66.080 -3.850 ;
        RECT 66.665 -4.110 66.825 -2.000 ;
        RECT 67.175 -3.130 67.335 -2.000 ;
        RECT 67.920 -2.010 68.080 -1.330 ;
        RECT 68.600 -2.000 68.890 -1.710 ;
        RECT 69.110 -2.000 69.400 -1.710 ;
        RECT 67.580 -2.190 67.740 -2.120 ;
        RECT 68.260 -2.190 68.420 -2.120 ;
        RECT 67.580 -2.480 67.870 -2.190 ;
        RECT 68.130 -2.480 68.420 -2.190 ;
        RECT 67.175 -3.290 68.425 -3.130 ;
        RECT 67.175 -4.110 67.335 -3.290 ;
        RECT 67.920 -4.410 68.080 -3.850 ;
        RECT 68.665 -4.110 68.825 -2.000 ;
        RECT 69.175 -3.130 69.335 -2.000 ;
        RECT 69.920 -2.010 70.080 -1.330 ;
        RECT 70.600 -2.000 70.890 -1.710 ;
        RECT 71.110 -2.000 71.400 -1.710 ;
        RECT 69.580 -2.190 69.740 -2.120 ;
        RECT 70.260 -2.190 70.420 -2.120 ;
        RECT 69.580 -2.480 69.870 -2.190 ;
        RECT 70.130 -2.480 70.420 -2.190 ;
        RECT 69.175 -3.290 70.425 -3.130 ;
        RECT 69.175 -4.110 69.335 -3.290 ;
        RECT 69.920 -4.410 70.080 -3.850 ;
        RECT 70.665 -4.110 70.825 -2.000 ;
        RECT 71.175 -3.130 71.335 -2.000 ;
        RECT 71.920 -2.010 72.080 -1.330 ;
        RECT 72.600 -2.000 72.890 -1.710 ;
        RECT 73.110 -2.000 73.400 -1.710 ;
        RECT 71.580 -2.190 71.740 -2.120 ;
        RECT 72.260 -2.190 72.420 -2.120 ;
        RECT 71.580 -2.480 71.870 -2.190 ;
        RECT 72.130 -2.480 72.420 -2.190 ;
        RECT 71.175 -3.290 72.425 -3.130 ;
        RECT 71.175 -4.110 71.335 -3.290 ;
        RECT 71.920 -4.410 72.080 -3.850 ;
        RECT 72.665 -4.110 72.825 -2.000 ;
        RECT 73.175 -3.130 73.335 -2.000 ;
        RECT 73.920 -2.010 74.080 -1.330 ;
        RECT 74.600 -2.000 74.890 -1.710 ;
        RECT 75.110 -2.000 75.400 -1.710 ;
        RECT 73.580 -2.190 73.740 -2.120 ;
        RECT 74.260 -2.190 74.420 -2.120 ;
        RECT 73.580 -2.480 73.870 -2.190 ;
        RECT 74.130 -2.480 74.420 -2.190 ;
        RECT 73.175 -3.290 74.425 -3.130 ;
        RECT 73.175 -4.110 73.335 -3.290 ;
        RECT 73.920 -4.410 74.080 -3.850 ;
        RECT 74.665 -4.110 74.825 -2.000 ;
        RECT 75.175 -3.130 75.335 -2.000 ;
        RECT 75.920 -2.010 76.080 -1.330 ;
        RECT 76.600 -2.000 76.890 -1.710 ;
        RECT 77.110 -2.000 77.400 -1.710 ;
        RECT 75.580 -2.190 75.740 -2.120 ;
        RECT 76.260 -2.190 76.420 -2.120 ;
        RECT 75.580 -2.480 75.870 -2.190 ;
        RECT 76.130 -2.480 76.420 -2.190 ;
        RECT 75.175 -3.290 76.425 -3.130 ;
        RECT 75.175 -4.110 75.335 -3.290 ;
        RECT 75.920 -4.410 76.080 -3.850 ;
        RECT 76.665 -4.110 76.825 -2.000 ;
        RECT 77.175 -3.130 77.335 -2.000 ;
        RECT 77.920 -2.010 78.080 -1.330 ;
        RECT 78.600 -2.000 78.890 -1.710 ;
        RECT 79.110 -2.000 79.400 -1.710 ;
        RECT 77.580 -2.190 77.740 -2.120 ;
        RECT 78.260 -2.190 78.420 -2.120 ;
        RECT 77.580 -2.480 77.870 -2.190 ;
        RECT 78.130 -2.480 78.420 -2.190 ;
        RECT 77.175 -3.290 78.425 -3.130 ;
        RECT 77.175 -4.110 77.335 -3.290 ;
        RECT 77.920 -4.410 78.080 -3.850 ;
        RECT 78.665 -4.110 78.825 -2.000 ;
        RECT 79.175 -3.130 79.335 -2.000 ;
        RECT 79.920 -2.010 80.080 -1.330 ;
        RECT 80.600 -2.000 80.890 -1.710 ;
        RECT 81.110 -2.000 81.400 -1.710 ;
        RECT 79.580 -2.190 79.740 -2.120 ;
        RECT 80.260 -2.190 80.420 -2.120 ;
        RECT 79.580 -2.480 79.870 -2.190 ;
        RECT 80.130 -2.480 80.420 -2.190 ;
        RECT 79.175 -3.290 80.425 -3.130 ;
        RECT 79.175 -4.110 79.335 -3.290 ;
        RECT 79.920 -4.410 80.080 -3.850 ;
        RECT 80.665 -4.110 80.825 -2.000 ;
        RECT 81.175 -3.130 81.335 -2.000 ;
        RECT 81.920 -2.010 82.080 -1.330 ;
        RECT 82.600 -2.000 82.890 -1.710 ;
        RECT 83.110 -2.000 83.400 -1.710 ;
        RECT 81.580 -2.190 81.740 -2.120 ;
        RECT 82.260 -2.190 82.420 -2.120 ;
        RECT 81.580 -2.480 81.870 -2.190 ;
        RECT 82.130 -2.480 82.420 -2.190 ;
        RECT 81.175 -3.290 82.425 -3.130 ;
        RECT 81.175 -4.110 81.335 -3.290 ;
        RECT 81.920 -4.410 82.080 -3.850 ;
        RECT 82.665 -4.110 82.825 -2.000 ;
        RECT 83.175 -3.130 83.335 -2.000 ;
        RECT 83.920 -2.010 84.080 -1.330 ;
        RECT 84.600 -2.000 84.890 -1.710 ;
        RECT 85.110 -2.000 85.400 -1.710 ;
        RECT 83.580 -2.190 83.740 -2.120 ;
        RECT 84.260 -2.190 84.420 -2.120 ;
        RECT 83.580 -2.480 83.870 -2.190 ;
        RECT 84.130 -2.480 84.420 -2.190 ;
        RECT 83.175 -3.290 84.425 -3.130 ;
        RECT 83.175 -4.110 83.335 -3.290 ;
        RECT 83.920 -4.410 84.080 -3.850 ;
        RECT 84.665 -4.110 84.825 -2.000 ;
        RECT 85.175 -3.130 85.335 -2.000 ;
        RECT 85.920 -2.010 86.080 -1.330 ;
        RECT 86.600 -2.000 86.890 -1.710 ;
        RECT 87.110 -2.000 87.400 -1.710 ;
        RECT 85.580 -2.190 85.740 -2.120 ;
        RECT 86.260 -2.190 86.420 -2.120 ;
        RECT 85.580 -2.480 85.870 -2.190 ;
        RECT 86.130 -2.480 86.420 -2.190 ;
        RECT 85.175 -3.290 86.425 -3.130 ;
        RECT 85.175 -4.110 85.335 -3.290 ;
        RECT 85.920 -4.410 86.080 -3.850 ;
        RECT 86.665 -4.110 86.825 -2.000 ;
        RECT 87.175 -3.130 87.335 -2.000 ;
        RECT 87.920 -2.010 88.080 -1.330 ;
        RECT 88.600 -2.000 88.890 -1.710 ;
        RECT 89.110 -2.000 89.400 -1.710 ;
        RECT 87.580 -2.190 87.740 -2.120 ;
        RECT 88.260 -2.190 88.420 -2.120 ;
        RECT 87.580 -2.480 87.870 -2.190 ;
        RECT 88.130 -2.480 88.420 -2.190 ;
        RECT 87.175 -3.290 88.425 -3.130 ;
        RECT 87.175 -4.110 87.335 -3.290 ;
        RECT 87.920 -4.410 88.080 -3.850 ;
        RECT 88.665 -4.110 88.825 -2.000 ;
        RECT 89.175 -3.130 89.335 -2.000 ;
        RECT 89.920 -2.010 90.080 -1.330 ;
        RECT 90.600 -2.000 90.890 -1.710 ;
        RECT 91.110 -2.000 91.400 -1.710 ;
        RECT 89.580 -2.190 89.740 -2.120 ;
        RECT 90.260 -2.190 90.420 -2.120 ;
        RECT 89.580 -2.480 89.870 -2.190 ;
        RECT 90.130 -2.480 90.420 -2.190 ;
        RECT 89.175 -3.290 90.425 -3.130 ;
        RECT 89.175 -4.110 89.335 -3.290 ;
        RECT 89.920 -4.410 90.080 -3.850 ;
        RECT 90.665 -4.110 90.825 -2.000 ;
        RECT 91.175 -3.130 91.335 -2.000 ;
        RECT 91.920 -2.010 92.080 -1.330 ;
        RECT 92.600 -2.000 92.890 -1.710 ;
        RECT 93.110 -2.000 93.400 -1.710 ;
        RECT 91.580 -2.190 91.740 -2.120 ;
        RECT 92.260 -2.190 92.420 -2.120 ;
        RECT 91.580 -2.480 91.870 -2.190 ;
        RECT 92.130 -2.480 92.420 -2.190 ;
        RECT 91.175 -3.290 92.425 -3.130 ;
        RECT 91.175 -4.110 91.335 -3.290 ;
        RECT 91.920 -4.410 92.080 -3.850 ;
        RECT 92.665 -4.110 92.825 -2.000 ;
        RECT 93.175 -3.130 93.335 -2.000 ;
        RECT 93.920 -2.010 94.080 -1.330 ;
        RECT 94.600 -2.000 94.890 -1.710 ;
        RECT 95.110 -2.000 95.400 -1.710 ;
        RECT 93.580 -2.190 93.740 -2.120 ;
        RECT 94.260 -2.190 94.420 -2.120 ;
        RECT 93.580 -2.480 93.870 -2.190 ;
        RECT 94.130 -2.480 94.420 -2.190 ;
        RECT 93.175 -3.290 94.425 -3.130 ;
        RECT 93.175 -4.110 93.335 -3.290 ;
        RECT 93.920 -4.410 94.080 -3.850 ;
        RECT 94.665 -4.110 94.825 -2.000 ;
        RECT 95.175 -3.130 95.335 -2.000 ;
        RECT 95.920 -2.010 96.080 -1.330 ;
        RECT 96.600 -2.000 96.890 -1.710 ;
        RECT 97.110 -2.000 97.400 -1.710 ;
        RECT 95.580 -2.190 95.740 -2.120 ;
        RECT 96.260 -2.190 96.420 -2.120 ;
        RECT 95.580 -2.480 95.870 -2.190 ;
        RECT 96.130 -2.480 96.420 -2.190 ;
        RECT 95.175 -3.290 96.425 -3.130 ;
        RECT 95.175 -4.110 95.335 -3.290 ;
        RECT 95.920 -4.410 96.080 -3.850 ;
        RECT 96.665 -4.110 96.825 -2.000 ;
        RECT 97.175 -3.130 97.335 -2.000 ;
        RECT 97.920 -2.010 98.080 -1.330 ;
        RECT 98.600 -2.000 98.890 -1.710 ;
        RECT 99.110 -2.000 99.400 -1.710 ;
        RECT 97.580 -2.190 97.740 -2.120 ;
        RECT 98.260 -2.190 98.420 -2.120 ;
        RECT 97.580 -2.480 97.870 -2.190 ;
        RECT 98.130 -2.480 98.420 -2.190 ;
        RECT 97.175 -3.290 98.425 -3.130 ;
        RECT 97.175 -4.110 97.335 -3.290 ;
        RECT 97.920 -4.410 98.080 -3.850 ;
        RECT 98.665 -4.110 98.825 -2.000 ;
        RECT 99.175 -3.130 99.335 -2.000 ;
        RECT 99.920 -2.010 100.080 -1.330 ;
        RECT 100.600 -2.000 100.890 -1.710 ;
        RECT 101.110 -2.000 101.400 -1.710 ;
        RECT 99.580 -2.190 99.740 -2.120 ;
        RECT 100.260 -2.190 100.420 -2.120 ;
        RECT 99.580 -2.480 99.870 -2.190 ;
        RECT 100.130 -2.480 100.420 -2.190 ;
        RECT 99.175 -3.290 100.425 -3.130 ;
        RECT 99.175 -4.110 99.335 -3.290 ;
        RECT 99.920 -4.410 100.080 -3.850 ;
        RECT 100.665 -4.110 100.825 -2.000 ;
        RECT 101.175 -3.130 101.335 -2.000 ;
        RECT 101.920 -2.010 102.080 -1.330 ;
        RECT 102.600 -2.000 102.890 -1.710 ;
        RECT 103.110 -2.000 103.400 -1.710 ;
        RECT 101.580 -2.190 101.740 -2.120 ;
        RECT 102.260 -2.190 102.420 -2.120 ;
        RECT 101.580 -2.480 101.870 -2.190 ;
        RECT 102.130 -2.480 102.420 -2.190 ;
        RECT 101.175 -3.290 102.425 -3.130 ;
        RECT 101.175 -4.110 101.335 -3.290 ;
        RECT 101.920 -4.410 102.080 -3.850 ;
        RECT 102.665 -4.110 102.825 -2.000 ;
        RECT 103.175 -3.130 103.335 -2.000 ;
        RECT 103.920 -2.010 104.080 -1.330 ;
        RECT 104.600 -2.000 104.890 -1.710 ;
        RECT 105.110 -2.000 105.400 -1.710 ;
        RECT 103.580 -2.190 103.740 -2.120 ;
        RECT 104.260 -2.190 104.420 -2.120 ;
        RECT 103.580 -2.480 103.870 -2.190 ;
        RECT 104.130 -2.480 104.420 -2.190 ;
        RECT 103.175 -3.290 104.425 -3.130 ;
        RECT 103.175 -4.110 103.335 -3.290 ;
        RECT 103.920 -4.410 104.080 -3.850 ;
        RECT 104.665 -4.110 104.825 -2.000 ;
        RECT 105.175 -3.130 105.335 -2.000 ;
        RECT 105.920 -2.010 106.080 -1.330 ;
        RECT 106.600 -2.000 106.890 -1.710 ;
        RECT 107.110 -2.000 107.400 -1.710 ;
        RECT 105.580 -2.190 105.740 -2.120 ;
        RECT 106.260 -2.190 106.420 -2.120 ;
        RECT 105.580 -2.480 105.870 -2.190 ;
        RECT 106.130 -2.480 106.420 -2.190 ;
        RECT 105.175 -3.290 106.425 -3.130 ;
        RECT 105.175 -4.110 105.335 -3.290 ;
        RECT 105.920 -4.410 106.080 -3.850 ;
        RECT 106.665 -4.110 106.825 -2.000 ;
        RECT 107.175 -3.130 107.335 -2.000 ;
        RECT 107.920 -2.010 108.080 -1.330 ;
        RECT 108.600 -2.000 108.890 -1.710 ;
        RECT 109.110 -2.000 109.400 -1.710 ;
        RECT 107.580 -2.190 107.740 -2.120 ;
        RECT 108.260 -2.190 108.420 -2.120 ;
        RECT 107.580 -2.480 107.870 -2.190 ;
        RECT 108.130 -2.480 108.420 -2.190 ;
        RECT 107.175 -3.290 108.425 -3.130 ;
        RECT 107.175 -4.110 107.335 -3.290 ;
        RECT 107.920 -4.410 108.080 -3.850 ;
        RECT 108.665 -4.110 108.825 -2.000 ;
        RECT 109.175 -3.130 109.335 -2.000 ;
        RECT 109.920 -2.010 110.080 -1.330 ;
        RECT 110.600 -2.000 110.890 -1.710 ;
        RECT 111.110 -2.000 111.400 -1.710 ;
        RECT 109.580 -2.190 109.740 -2.120 ;
        RECT 110.260 -2.190 110.420 -2.120 ;
        RECT 109.580 -2.480 109.870 -2.190 ;
        RECT 110.130 -2.480 110.420 -2.190 ;
        RECT 109.175 -3.290 110.425 -3.130 ;
        RECT 109.175 -4.110 109.335 -3.290 ;
        RECT 109.920 -4.410 110.080 -3.850 ;
        RECT 110.665 -4.110 110.825 -2.000 ;
        RECT 111.175 -3.130 111.335 -2.000 ;
        RECT 111.920 -2.010 112.080 -1.330 ;
        RECT 112.600 -2.000 112.890 -1.710 ;
        RECT 113.110 -2.000 113.400 -1.710 ;
        RECT 111.580 -2.190 111.740 -2.120 ;
        RECT 112.260 -2.190 112.420 -2.120 ;
        RECT 111.580 -2.480 111.870 -2.190 ;
        RECT 112.130 -2.480 112.420 -2.190 ;
        RECT 111.175 -3.290 112.425 -3.130 ;
        RECT 111.175 -4.110 111.335 -3.290 ;
        RECT 111.920 -4.410 112.080 -3.850 ;
        RECT 112.665 -4.110 112.825 -2.000 ;
        RECT 113.175 -3.130 113.335 -2.000 ;
        RECT 113.920 -2.010 114.080 -1.330 ;
        RECT 114.600 -2.000 114.890 -1.710 ;
        RECT 115.110 -2.000 115.400 -1.710 ;
        RECT 113.580 -2.190 113.740 -2.120 ;
        RECT 114.260 -2.190 114.420 -2.120 ;
        RECT 113.580 -2.480 113.870 -2.190 ;
        RECT 114.130 -2.480 114.420 -2.190 ;
        RECT 113.175 -3.290 114.425 -3.130 ;
        RECT 113.175 -4.110 113.335 -3.290 ;
        RECT 113.920 -4.410 114.080 -3.850 ;
        RECT 114.665 -4.110 114.825 -2.000 ;
        RECT 115.175 -3.130 115.335 -2.000 ;
        RECT 115.920 -2.010 116.080 -1.330 ;
        RECT 116.600 -2.000 116.890 -1.710 ;
        RECT 117.110 -2.000 117.400 -1.710 ;
        RECT 115.580 -2.190 115.740 -2.120 ;
        RECT 116.260 -2.190 116.420 -2.120 ;
        RECT 115.580 -2.480 115.870 -2.190 ;
        RECT 116.130 -2.480 116.420 -2.190 ;
        RECT 115.175 -3.290 116.425 -3.130 ;
        RECT 115.175 -4.110 115.335 -3.290 ;
        RECT 115.920 -4.410 116.080 -3.850 ;
        RECT 116.665 -4.110 116.825 -2.000 ;
        RECT 117.175 -3.130 117.335 -2.000 ;
        RECT 117.920 -2.010 118.080 -1.330 ;
        RECT 118.600 -2.000 118.890 -1.710 ;
        RECT 119.110 -2.000 119.400 -1.710 ;
        RECT 117.580 -2.190 117.740 -2.120 ;
        RECT 118.260 -2.190 118.420 -2.120 ;
        RECT 117.580 -2.480 117.870 -2.190 ;
        RECT 118.130 -2.480 118.420 -2.190 ;
        RECT 117.175 -3.290 118.425 -3.130 ;
        RECT 117.175 -4.110 117.335 -3.290 ;
        RECT 117.920 -4.410 118.080 -3.850 ;
        RECT 118.665 -4.110 118.825 -2.000 ;
        RECT 119.175 -3.130 119.335 -2.000 ;
        RECT 119.920 -2.010 120.080 -1.330 ;
        RECT 120.600 -2.000 120.890 -1.710 ;
        RECT 121.110 -2.000 121.400 -1.710 ;
        RECT 119.580 -2.190 119.740 -2.120 ;
        RECT 120.260 -2.190 120.420 -2.120 ;
        RECT 119.580 -2.480 119.870 -2.190 ;
        RECT 120.130 -2.480 120.420 -2.190 ;
        RECT 119.175 -3.290 120.425 -3.130 ;
        RECT 119.175 -4.110 119.335 -3.290 ;
        RECT 119.920 -4.410 120.080 -3.850 ;
        RECT 120.665 -4.110 120.825 -2.000 ;
        RECT 121.175 -3.130 121.335 -2.000 ;
        RECT 121.920 -2.010 122.080 -1.330 ;
        RECT 122.600 -2.000 122.890 -1.710 ;
        RECT 123.110 -2.000 123.400 -1.710 ;
        RECT 121.580 -2.190 121.740 -2.120 ;
        RECT 122.260 -2.190 122.420 -2.120 ;
        RECT 121.580 -2.480 121.870 -2.190 ;
        RECT 122.130 -2.480 122.420 -2.190 ;
        RECT 121.175 -3.290 122.425 -3.130 ;
        RECT 121.175 -4.110 121.335 -3.290 ;
        RECT 121.920 -4.410 122.080 -3.850 ;
        RECT 122.665 -4.110 122.825 -2.000 ;
        RECT 123.175 -3.130 123.335 -2.000 ;
        RECT 123.920 -2.010 124.080 -1.330 ;
        RECT 124.600 -2.000 124.890 -1.710 ;
        RECT 125.110 -2.000 125.400 -1.710 ;
        RECT 123.580 -2.190 123.740 -2.120 ;
        RECT 124.260 -2.190 124.420 -2.120 ;
        RECT 123.580 -2.480 123.870 -2.190 ;
        RECT 124.130 -2.480 124.420 -2.190 ;
        RECT 123.175 -3.290 124.425 -3.130 ;
        RECT 123.175 -4.110 123.335 -3.290 ;
        RECT 123.920 -4.410 124.080 -3.850 ;
        RECT 124.665 -4.110 124.825 -2.000 ;
        RECT 125.175 -3.130 125.335 -2.000 ;
        RECT 125.920 -2.010 126.080 -1.330 ;
        RECT 126.600 -2.000 126.890 -1.710 ;
        RECT 127.110 -2.000 127.400 -1.710 ;
        RECT 125.580 -2.190 125.740 -2.120 ;
        RECT 126.260 -2.190 126.420 -2.120 ;
        RECT 125.580 -2.480 125.870 -2.190 ;
        RECT 126.130 -2.480 126.420 -2.190 ;
        RECT 125.175 -3.290 126.425 -3.130 ;
        RECT 125.175 -4.110 125.335 -3.290 ;
        RECT 125.920 -4.410 126.080 -3.850 ;
        RECT 126.665 -4.110 126.825 -2.000 ;
        RECT 127.175 -3.130 127.335 -2.000 ;
        RECT 127.920 -2.010 128.080 -1.330 ;
        RECT 128.600 -2.000 128.890 -1.710 ;
        RECT 129.110 -2.000 129.400 -1.710 ;
        RECT 127.580 -2.190 127.740 -2.120 ;
        RECT 128.260 -2.190 128.420 -2.120 ;
        RECT 127.580 -2.480 127.870 -2.190 ;
        RECT 128.130 -2.480 128.420 -2.190 ;
        RECT 127.175 -3.290 128.425 -3.130 ;
        RECT 127.175 -4.110 127.335 -3.290 ;
        RECT 127.920 -4.410 128.080 -3.850 ;
        RECT 128.665 -4.110 128.825 -2.000 ;
        RECT 129.175 -3.130 129.335 -2.000 ;
        RECT 129.920 -2.010 130.080 -1.330 ;
        RECT 130.600 -2.000 130.890 -1.710 ;
        RECT 129.580 -2.190 129.740 -2.120 ;
        RECT 130.260 -2.190 130.420 -2.120 ;
        RECT 129.580 -2.480 129.870 -2.190 ;
        RECT 130.130 -2.480 130.420 -2.190 ;
        RECT 129.175 -3.290 130.425 -3.130 ;
        RECT 129.175 -4.110 129.335 -3.290 ;
        RECT 129.920 -4.410 130.080 -3.850 ;
        RECT 130.665 -4.110 130.825 -2.000 ;
      LAYER Metal2 ;
        RECT -0.420 18.560 -0.130 20.990 ;
        RECT 0.130 18.560 0.420 20.990 ;
        RECT 1.580 18.560 1.870 20.990 ;
        RECT 2.130 18.560 2.420 20.990 ;
        RECT 3.580 18.560 3.870 20.990 ;
        RECT 4.130 18.560 4.420 20.990 ;
        RECT 5.580 18.560 5.870 20.990 ;
        RECT 6.130 18.560 6.420 20.990 ;
        RECT 7.580 18.560 7.870 20.990 ;
        RECT 8.130 18.560 8.420 20.990 ;
        RECT 9.580 18.560 9.870 20.990 ;
        RECT 10.130 18.560 10.420 20.990 ;
        RECT 11.580 18.560 11.870 20.990 ;
        RECT 12.130 18.560 12.420 20.990 ;
        RECT 13.580 18.560 13.870 20.990 ;
        RECT 14.130 18.560 14.420 20.990 ;
        RECT 15.580 18.560 15.870 20.990 ;
        RECT 16.130 18.560 16.420 20.990 ;
        RECT 17.580 18.560 17.870 20.990 ;
        RECT 18.130 18.560 18.420 20.990 ;
        RECT 19.580 18.560 19.870 20.990 ;
        RECT 20.130 18.560 20.420 20.990 ;
        RECT 21.580 18.560 21.870 20.990 ;
        RECT 22.130 18.560 22.420 20.990 ;
        RECT 23.580 18.560 23.870 20.990 ;
        RECT 24.130 18.560 24.420 20.990 ;
        RECT 25.580 18.560 25.870 20.990 ;
        RECT 26.130 18.560 26.420 20.990 ;
        RECT 27.580 18.560 27.870 20.990 ;
        RECT 28.130 18.560 28.420 20.990 ;
        RECT 29.580 18.560 29.870 20.990 ;
        RECT 30.130 18.560 30.420 20.990 ;
        RECT 31.580 18.560 31.870 20.990 ;
        RECT 32.130 18.560 32.420 20.990 ;
        RECT 33.580 18.560 33.870 20.990 ;
        RECT 34.130 18.560 34.420 20.990 ;
        RECT 35.580 18.560 35.870 20.990 ;
        RECT 36.130 18.560 36.420 20.990 ;
        RECT 37.580 18.560 37.870 20.990 ;
        RECT 38.130 18.560 38.420 20.990 ;
        RECT 39.580 18.560 39.870 20.990 ;
        RECT 40.130 18.560 40.420 20.990 ;
        RECT 41.580 18.560 41.870 20.990 ;
        RECT 42.130 18.560 42.420 20.990 ;
        RECT 43.580 18.560 43.870 20.990 ;
        RECT 44.130 18.560 44.420 20.990 ;
        RECT 45.580 18.560 45.870 20.990 ;
        RECT 46.130 18.560 46.420 20.990 ;
        RECT 47.580 18.560 47.870 20.990 ;
        RECT 48.130 18.560 48.420 20.990 ;
        RECT 49.580 18.560 49.870 20.990 ;
        RECT 50.130 18.560 50.420 20.990 ;
        RECT 51.580 18.560 51.870 20.990 ;
        RECT 52.130 18.560 52.420 20.990 ;
        RECT 53.580 18.560 53.870 20.990 ;
        RECT 54.130 18.560 54.420 20.990 ;
        RECT 55.580 18.560 55.870 20.990 ;
        RECT 56.130 18.560 56.420 20.990 ;
        RECT 57.580 18.560 57.870 20.990 ;
        RECT 58.130 18.560 58.420 20.990 ;
        RECT 59.580 18.560 59.870 20.990 ;
        RECT 60.130 18.560 60.420 20.990 ;
        RECT 61.580 18.560 61.870 20.990 ;
        RECT 62.130 18.560 62.420 20.990 ;
        RECT 63.580 18.560 63.870 20.990 ;
        RECT 64.130 18.560 64.420 20.990 ;
        RECT 65.580 18.560 65.870 20.990 ;
        RECT 66.130 18.560 66.420 20.990 ;
        RECT 67.580 18.560 67.870 20.990 ;
        RECT 68.130 18.560 68.420 20.990 ;
        RECT 69.580 18.560 69.870 20.990 ;
        RECT 70.130 18.560 70.420 20.990 ;
        RECT 71.580 18.560 71.870 20.990 ;
        RECT 72.130 18.560 72.420 20.990 ;
        RECT 73.580 18.560 73.870 20.990 ;
        RECT 74.130 18.560 74.420 20.990 ;
        RECT 75.580 18.560 75.870 20.990 ;
        RECT 76.130 18.560 76.420 20.990 ;
        RECT 77.580 18.560 77.870 20.990 ;
        RECT 78.130 18.560 78.420 20.990 ;
        RECT 79.580 18.560 79.870 20.990 ;
        RECT 80.130 18.560 80.420 20.990 ;
        RECT 81.580 18.560 81.870 20.990 ;
        RECT 82.130 18.560 82.420 20.990 ;
        RECT 83.580 18.560 83.870 20.990 ;
        RECT 84.130 18.560 84.420 20.990 ;
        RECT 85.580 18.560 85.870 20.990 ;
        RECT 86.130 18.560 86.420 20.990 ;
        RECT 87.580 18.560 87.870 20.990 ;
        RECT 88.130 18.560 88.420 20.990 ;
        RECT 89.580 18.560 89.870 20.990 ;
        RECT 90.130 18.560 90.420 20.990 ;
        RECT 91.580 18.560 91.870 20.990 ;
        RECT 92.130 18.560 92.420 20.990 ;
        RECT 93.580 18.560 93.870 20.990 ;
        RECT 94.130 18.560 94.420 20.990 ;
        RECT 95.580 18.560 95.870 20.990 ;
        RECT 96.130 18.560 96.420 20.990 ;
        RECT 97.580 18.560 97.870 20.990 ;
        RECT 98.130 18.560 98.420 20.990 ;
        RECT 99.580 18.560 99.870 20.990 ;
        RECT 100.130 18.560 100.420 20.990 ;
        RECT 101.580 18.560 101.870 20.990 ;
        RECT 102.130 18.560 102.420 20.990 ;
        RECT 103.580 18.560 103.870 20.990 ;
        RECT 104.130 18.560 104.420 20.990 ;
        RECT 105.580 18.560 105.870 20.990 ;
        RECT 106.130 18.560 106.420 20.990 ;
        RECT 107.580 18.560 107.870 20.990 ;
        RECT 108.130 18.560 108.420 20.990 ;
        RECT 109.580 18.560 109.870 20.990 ;
        RECT 110.130 18.560 110.420 20.990 ;
        RECT 111.580 18.560 111.870 20.990 ;
        RECT 112.130 18.560 112.420 20.990 ;
        RECT 113.580 18.560 113.870 20.990 ;
        RECT 114.130 18.560 114.420 20.990 ;
        RECT 115.580 18.560 115.870 20.990 ;
        RECT 116.130 18.560 116.420 20.990 ;
        RECT 117.580 18.560 117.870 20.990 ;
        RECT 118.130 18.560 118.420 20.990 ;
        RECT 119.580 18.560 119.870 20.990 ;
        RECT 120.130 18.560 120.420 20.990 ;
        RECT 121.580 18.560 121.870 20.990 ;
        RECT 122.130 18.560 122.420 20.990 ;
        RECT 123.580 18.560 123.870 20.990 ;
        RECT 124.130 18.560 124.420 20.990 ;
        RECT 125.580 18.560 125.870 20.990 ;
        RECT 126.130 18.560 126.420 20.990 ;
        RECT 127.580 18.560 127.870 20.990 ;
        RECT 128.130 18.560 128.420 20.990 ;
        RECT 129.580 18.560 129.870 20.990 ;
        RECT 130.130 18.560 130.420 20.990 ;
        RECT -0.890 18.080 -0.600 18.370 ;
        RECT 0.600 18.080 0.890 18.370 ;
        RECT 1.110 18.080 1.400 18.370 ;
        RECT 2.600 18.080 2.890 18.370 ;
        RECT 3.110 18.080 3.400 18.370 ;
        RECT 4.600 18.080 4.890 18.370 ;
        RECT 5.110 18.080 5.400 18.370 ;
        RECT 6.600 18.080 6.890 18.370 ;
        RECT 7.110 18.080 7.400 18.370 ;
        RECT 8.600 18.080 8.890 18.370 ;
        RECT 9.110 18.080 9.400 18.370 ;
        RECT 10.600 18.080 10.890 18.370 ;
        RECT 11.110 18.080 11.400 18.370 ;
        RECT 12.600 18.080 12.890 18.370 ;
        RECT 13.110 18.080 13.400 18.370 ;
        RECT 14.600 18.080 14.890 18.370 ;
        RECT 15.110 18.080 15.400 18.370 ;
        RECT 16.600 18.080 16.890 18.370 ;
        RECT 17.110 18.080 17.400 18.370 ;
        RECT 18.600 18.080 18.890 18.370 ;
        RECT 19.110 18.080 19.400 18.370 ;
        RECT 20.600 18.080 20.890 18.370 ;
        RECT 21.110 18.080 21.400 18.370 ;
        RECT 22.600 18.080 22.890 18.370 ;
        RECT 23.110 18.080 23.400 18.370 ;
        RECT 24.600 18.080 24.890 18.370 ;
        RECT 25.110 18.080 25.400 18.370 ;
        RECT 26.600 18.080 26.890 18.370 ;
        RECT 27.110 18.080 27.400 18.370 ;
        RECT 28.600 18.080 28.890 18.370 ;
        RECT 29.110 18.080 29.400 18.370 ;
        RECT 30.600 18.080 30.890 18.370 ;
        RECT 31.110 18.080 31.400 18.370 ;
        RECT 32.600 18.080 32.890 18.370 ;
        RECT 33.110 18.080 33.400 18.370 ;
        RECT 34.600 18.080 34.890 18.370 ;
        RECT 35.110 18.080 35.400 18.370 ;
        RECT 36.600 18.080 36.890 18.370 ;
        RECT 37.110 18.080 37.400 18.370 ;
        RECT 38.600 18.080 38.890 18.370 ;
        RECT 39.110 18.080 39.400 18.370 ;
        RECT 40.600 18.080 40.890 18.370 ;
        RECT 41.110 18.080 41.400 18.370 ;
        RECT 42.600 18.080 42.890 18.370 ;
        RECT 43.110 18.080 43.400 18.370 ;
        RECT 44.600 18.080 44.890 18.370 ;
        RECT 45.110 18.080 45.400 18.370 ;
        RECT 46.600 18.080 46.890 18.370 ;
        RECT 47.110 18.080 47.400 18.370 ;
        RECT 48.600 18.080 48.890 18.370 ;
        RECT 49.110 18.080 49.400 18.370 ;
        RECT 50.600 18.080 50.890 18.370 ;
        RECT 51.110 18.080 51.400 18.370 ;
        RECT 52.600 18.080 52.890 18.370 ;
        RECT 53.110 18.080 53.400 18.370 ;
        RECT 54.600 18.080 54.890 18.370 ;
        RECT 55.110 18.080 55.400 18.370 ;
        RECT 56.600 18.080 56.890 18.370 ;
        RECT 57.110 18.080 57.400 18.370 ;
        RECT 58.600 18.080 58.890 18.370 ;
        RECT 59.110 18.080 59.400 18.370 ;
        RECT 60.600 18.080 60.890 18.370 ;
        RECT 61.110 18.080 61.400 18.370 ;
        RECT 62.600 18.080 62.890 18.370 ;
        RECT 63.110 18.080 63.400 18.370 ;
        RECT 64.600 18.080 64.890 18.370 ;
        RECT 65.110 18.080 65.400 18.370 ;
        RECT 66.600 18.080 66.890 18.370 ;
        RECT 67.110 18.080 67.400 18.370 ;
        RECT 68.600 18.080 68.890 18.370 ;
        RECT 69.110 18.080 69.400 18.370 ;
        RECT 70.600 18.080 70.890 18.370 ;
        RECT 71.110 18.080 71.400 18.370 ;
        RECT 72.600 18.080 72.890 18.370 ;
        RECT 73.110 18.080 73.400 18.370 ;
        RECT 74.600 18.080 74.890 18.370 ;
        RECT 75.110 18.080 75.400 18.370 ;
        RECT 76.600 18.080 76.890 18.370 ;
        RECT 77.110 18.080 77.400 18.370 ;
        RECT 78.600 18.080 78.890 18.370 ;
        RECT 79.110 18.080 79.400 18.370 ;
        RECT 80.600 18.080 80.890 18.370 ;
        RECT 81.110 18.080 81.400 18.370 ;
        RECT 82.600 18.080 82.890 18.370 ;
        RECT 83.110 18.080 83.400 18.370 ;
        RECT 84.600 18.080 84.890 18.370 ;
        RECT 85.110 18.080 85.400 18.370 ;
        RECT 86.600 18.080 86.890 18.370 ;
        RECT 87.110 18.080 87.400 18.370 ;
        RECT 88.600 18.080 88.890 18.370 ;
        RECT 89.110 18.080 89.400 18.370 ;
        RECT 90.600 18.080 90.890 18.370 ;
        RECT 91.110 18.080 91.400 18.370 ;
        RECT 92.600 18.080 92.890 18.370 ;
        RECT 93.110 18.080 93.400 18.370 ;
        RECT 94.600 18.080 94.890 18.370 ;
        RECT 95.110 18.080 95.400 18.370 ;
        RECT 96.600 18.080 96.890 18.370 ;
        RECT 97.110 18.080 97.400 18.370 ;
        RECT 98.600 18.080 98.890 18.370 ;
        RECT 99.110 18.080 99.400 18.370 ;
        RECT 100.600 18.080 100.890 18.370 ;
        RECT 101.110 18.080 101.400 18.370 ;
        RECT 102.600 18.080 102.890 18.370 ;
        RECT 103.110 18.080 103.400 18.370 ;
        RECT 104.600 18.080 104.890 18.370 ;
        RECT 105.110 18.080 105.400 18.370 ;
        RECT 106.600 18.080 106.890 18.370 ;
        RECT 107.110 18.080 107.400 18.370 ;
        RECT 108.600 18.080 108.890 18.370 ;
        RECT 109.110 18.080 109.400 18.370 ;
        RECT 110.600 18.080 110.890 18.370 ;
        RECT 111.110 18.080 111.400 18.370 ;
        RECT 112.600 18.080 112.890 18.370 ;
        RECT 113.110 18.080 113.400 18.370 ;
        RECT 114.600 18.080 114.890 18.370 ;
        RECT 115.110 18.080 115.400 18.370 ;
        RECT 116.600 18.080 116.890 18.370 ;
        RECT 117.110 18.080 117.400 18.370 ;
        RECT 118.600 18.080 118.890 18.370 ;
        RECT 119.110 18.080 119.400 18.370 ;
        RECT 120.600 18.080 120.890 18.370 ;
        RECT 121.110 18.080 121.400 18.370 ;
        RECT 122.600 18.080 122.890 18.370 ;
        RECT 123.110 18.080 123.400 18.370 ;
        RECT 124.600 18.080 124.890 18.370 ;
        RECT 125.110 18.080 125.400 18.370 ;
        RECT 126.600 18.080 126.890 18.370 ;
        RECT 127.110 18.080 127.400 18.370 ;
        RECT 128.600 18.080 128.890 18.370 ;
        RECT 129.110 18.080 129.400 18.370 ;
        RECT 130.600 18.080 130.890 18.370 ;
        RECT -0.840 17.015 -0.640 18.080 ;
        RECT 0.645 17.015 0.845 18.080 ;
        RECT -0.840 16.815 -0.195 17.015 ;
        RECT -0.485 16.725 -0.195 16.815 ;
        RECT 0.195 16.815 0.845 17.015 ;
        RECT 1.160 17.015 1.360 18.080 ;
        RECT 2.645 17.015 2.845 18.080 ;
        RECT 1.160 16.815 1.805 17.015 ;
        RECT 0.195 16.725 0.485 16.815 ;
        RECT 1.515 16.725 1.805 16.815 ;
        RECT 2.195 16.815 2.845 17.015 ;
        RECT 3.160 17.015 3.360 18.080 ;
        RECT 4.645 17.015 4.845 18.080 ;
        RECT 3.160 16.815 3.805 17.015 ;
        RECT 2.195 16.725 2.485 16.815 ;
        RECT 3.515 16.725 3.805 16.815 ;
        RECT 4.195 16.815 4.845 17.015 ;
        RECT 5.160 17.015 5.360 18.080 ;
        RECT 6.645 17.015 6.845 18.080 ;
        RECT 5.160 16.815 5.805 17.015 ;
        RECT 4.195 16.725 4.485 16.815 ;
        RECT 5.515 16.725 5.805 16.815 ;
        RECT 6.195 16.815 6.845 17.015 ;
        RECT 7.160 17.015 7.360 18.080 ;
        RECT 8.645 17.015 8.845 18.080 ;
        RECT 7.160 16.815 7.805 17.015 ;
        RECT 6.195 16.725 6.485 16.815 ;
        RECT 7.515 16.725 7.805 16.815 ;
        RECT 8.195 16.815 8.845 17.015 ;
        RECT 9.160 17.015 9.360 18.080 ;
        RECT 10.645 17.015 10.845 18.080 ;
        RECT 9.160 16.815 9.805 17.015 ;
        RECT 8.195 16.725 8.485 16.815 ;
        RECT 9.515 16.725 9.805 16.815 ;
        RECT 10.195 16.815 10.845 17.015 ;
        RECT 11.160 17.015 11.360 18.080 ;
        RECT 12.645 17.015 12.845 18.080 ;
        RECT 11.160 16.815 11.805 17.015 ;
        RECT 10.195 16.725 10.485 16.815 ;
        RECT 11.515 16.725 11.805 16.815 ;
        RECT 12.195 16.815 12.845 17.015 ;
        RECT 13.160 17.015 13.360 18.080 ;
        RECT 14.645 17.015 14.845 18.080 ;
        RECT 13.160 16.815 13.805 17.015 ;
        RECT 12.195 16.725 12.485 16.815 ;
        RECT 13.515 16.725 13.805 16.815 ;
        RECT 14.195 16.815 14.845 17.015 ;
        RECT 15.160 17.015 15.360 18.080 ;
        RECT 16.645 17.015 16.845 18.080 ;
        RECT 15.160 16.815 15.805 17.015 ;
        RECT 14.195 16.725 14.485 16.815 ;
        RECT 15.515 16.725 15.805 16.815 ;
        RECT 16.195 16.815 16.845 17.015 ;
        RECT 17.160 17.015 17.360 18.080 ;
        RECT 18.645 17.015 18.845 18.080 ;
        RECT 17.160 16.815 17.805 17.015 ;
        RECT 16.195 16.725 16.485 16.815 ;
        RECT 17.515 16.725 17.805 16.815 ;
        RECT 18.195 16.815 18.845 17.015 ;
        RECT 19.160 17.015 19.360 18.080 ;
        RECT 20.645 17.015 20.845 18.080 ;
        RECT 19.160 16.815 19.805 17.015 ;
        RECT 18.195 16.725 18.485 16.815 ;
        RECT 19.515 16.725 19.805 16.815 ;
        RECT 20.195 16.815 20.845 17.015 ;
        RECT 21.160 17.015 21.360 18.080 ;
        RECT 22.645 17.015 22.845 18.080 ;
        RECT 21.160 16.815 21.805 17.015 ;
        RECT 20.195 16.725 20.485 16.815 ;
        RECT 21.515 16.725 21.805 16.815 ;
        RECT 22.195 16.815 22.845 17.015 ;
        RECT 23.160 17.015 23.360 18.080 ;
        RECT 24.645 17.015 24.845 18.080 ;
        RECT 23.160 16.815 23.805 17.015 ;
        RECT 22.195 16.725 22.485 16.815 ;
        RECT 23.515 16.725 23.805 16.815 ;
        RECT 24.195 16.815 24.845 17.015 ;
        RECT 25.160 17.015 25.360 18.080 ;
        RECT 26.645 17.015 26.845 18.080 ;
        RECT 25.160 16.815 25.805 17.015 ;
        RECT 24.195 16.725 24.485 16.815 ;
        RECT 25.515 16.725 25.805 16.815 ;
        RECT 26.195 16.815 26.845 17.015 ;
        RECT 27.160 17.015 27.360 18.080 ;
        RECT 28.645 17.015 28.845 18.080 ;
        RECT 27.160 16.815 27.805 17.015 ;
        RECT 26.195 16.725 26.485 16.815 ;
        RECT 27.515 16.725 27.805 16.815 ;
        RECT 28.195 16.815 28.845 17.015 ;
        RECT 29.160 17.015 29.360 18.080 ;
        RECT 30.645 17.015 30.845 18.080 ;
        RECT 29.160 16.815 29.805 17.015 ;
        RECT 28.195 16.725 28.485 16.815 ;
        RECT 29.515 16.725 29.805 16.815 ;
        RECT 30.195 16.815 30.845 17.015 ;
        RECT 31.160 17.015 31.360 18.080 ;
        RECT 32.645 17.015 32.845 18.080 ;
        RECT 31.160 16.815 31.805 17.015 ;
        RECT 30.195 16.725 30.485 16.815 ;
        RECT 31.515 16.725 31.805 16.815 ;
        RECT 32.195 16.815 32.845 17.015 ;
        RECT 33.160 17.015 33.360 18.080 ;
        RECT 34.645 17.015 34.845 18.080 ;
        RECT 33.160 16.815 33.805 17.015 ;
        RECT 32.195 16.725 32.485 16.815 ;
        RECT 33.515 16.725 33.805 16.815 ;
        RECT 34.195 16.815 34.845 17.015 ;
        RECT 35.160 17.015 35.360 18.080 ;
        RECT 36.645 17.015 36.845 18.080 ;
        RECT 35.160 16.815 35.805 17.015 ;
        RECT 34.195 16.725 34.485 16.815 ;
        RECT 35.515 16.725 35.805 16.815 ;
        RECT 36.195 16.815 36.845 17.015 ;
        RECT 37.160 17.015 37.360 18.080 ;
        RECT 38.645 17.015 38.845 18.080 ;
        RECT 37.160 16.815 37.805 17.015 ;
        RECT 36.195 16.725 36.485 16.815 ;
        RECT 37.515 16.725 37.805 16.815 ;
        RECT 38.195 16.815 38.845 17.015 ;
        RECT 39.160 17.015 39.360 18.080 ;
        RECT 40.645 17.015 40.845 18.080 ;
        RECT 39.160 16.815 39.805 17.015 ;
        RECT 38.195 16.725 38.485 16.815 ;
        RECT 39.515 16.725 39.805 16.815 ;
        RECT 40.195 16.815 40.845 17.015 ;
        RECT 41.160 17.015 41.360 18.080 ;
        RECT 42.645 17.015 42.845 18.080 ;
        RECT 41.160 16.815 41.805 17.015 ;
        RECT 40.195 16.725 40.485 16.815 ;
        RECT 41.515 16.725 41.805 16.815 ;
        RECT 42.195 16.815 42.845 17.015 ;
        RECT 43.160 17.015 43.360 18.080 ;
        RECT 44.645 17.015 44.845 18.080 ;
        RECT 43.160 16.815 43.805 17.015 ;
        RECT 42.195 16.725 42.485 16.815 ;
        RECT 43.515 16.725 43.805 16.815 ;
        RECT 44.195 16.815 44.845 17.015 ;
        RECT 45.160 17.015 45.360 18.080 ;
        RECT 46.645 17.015 46.845 18.080 ;
        RECT 45.160 16.815 45.805 17.015 ;
        RECT 44.195 16.725 44.485 16.815 ;
        RECT 45.515 16.725 45.805 16.815 ;
        RECT 46.195 16.815 46.845 17.015 ;
        RECT 47.160 17.015 47.360 18.080 ;
        RECT 48.645 17.015 48.845 18.080 ;
        RECT 47.160 16.815 47.805 17.015 ;
        RECT 46.195 16.725 46.485 16.815 ;
        RECT 47.515 16.725 47.805 16.815 ;
        RECT 48.195 16.815 48.845 17.015 ;
        RECT 49.160 17.015 49.360 18.080 ;
        RECT 50.645 17.015 50.845 18.080 ;
        RECT 49.160 16.815 49.805 17.015 ;
        RECT 48.195 16.725 48.485 16.815 ;
        RECT 49.515 16.725 49.805 16.815 ;
        RECT 50.195 16.815 50.845 17.015 ;
        RECT 51.160 17.015 51.360 18.080 ;
        RECT 52.645 17.015 52.845 18.080 ;
        RECT 51.160 16.815 51.805 17.015 ;
        RECT 50.195 16.725 50.485 16.815 ;
        RECT 51.515 16.725 51.805 16.815 ;
        RECT 52.195 16.815 52.845 17.015 ;
        RECT 53.160 17.015 53.360 18.080 ;
        RECT 54.645 17.015 54.845 18.080 ;
        RECT 53.160 16.815 53.805 17.015 ;
        RECT 52.195 16.725 52.485 16.815 ;
        RECT 53.515 16.725 53.805 16.815 ;
        RECT 54.195 16.815 54.845 17.015 ;
        RECT 55.160 17.015 55.360 18.080 ;
        RECT 56.645 17.015 56.845 18.080 ;
        RECT 55.160 16.815 55.805 17.015 ;
        RECT 54.195 16.725 54.485 16.815 ;
        RECT 55.515 16.725 55.805 16.815 ;
        RECT 56.195 16.815 56.845 17.015 ;
        RECT 57.160 17.015 57.360 18.080 ;
        RECT 58.645 17.015 58.845 18.080 ;
        RECT 57.160 16.815 57.805 17.015 ;
        RECT 56.195 16.725 56.485 16.815 ;
        RECT 57.515 16.725 57.805 16.815 ;
        RECT 58.195 16.815 58.845 17.015 ;
        RECT 59.160 17.015 59.360 18.080 ;
        RECT 60.645 17.015 60.845 18.080 ;
        RECT 59.160 16.815 59.805 17.015 ;
        RECT 58.195 16.725 58.485 16.815 ;
        RECT 59.515 16.725 59.805 16.815 ;
        RECT 60.195 16.815 60.845 17.015 ;
        RECT 61.160 17.015 61.360 18.080 ;
        RECT 62.645 17.015 62.845 18.080 ;
        RECT 61.160 16.815 61.805 17.015 ;
        RECT 60.195 16.725 60.485 16.815 ;
        RECT 61.515 16.725 61.805 16.815 ;
        RECT 62.195 16.815 62.845 17.015 ;
        RECT 63.160 17.015 63.360 18.080 ;
        RECT 64.645 17.015 64.845 18.080 ;
        RECT 63.160 16.815 63.805 17.015 ;
        RECT 62.195 16.725 62.485 16.815 ;
        RECT 63.515 16.725 63.805 16.815 ;
        RECT 64.195 16.815 64.845 17.015 ;
        RECT 65.160 17.015 65.360 18.080 ;
        RECT 66.645 17.015 66.845 18.080 ;
        RECT 65.160 16.815 65.805 17.015 ;
        RECT 64.195 16.725 64.485 16.815 ;
        RECT 65.515 16.725 65.805 16.815 ;
        RECT 66.195 16.815 66.845 17.015 ;
        RECT 67.160 17.015 67.360 18.080 ;
        RECT 68.645 17.015 68.845 18.080 ;
        RECT 67.160 16.815 67.805 17.015 ;
        RECT 66.195 16.725 66.485 16.815 ;
        RECT 67.515 16.725 67.805 16.815 ;
        RECT 68.195 16.815 68.845 17.015 ;
        RECT 69.160 17.015 69.360 18.080 ;
        RECT 70.645 17.015 70.845 18.080 ;
        RECT 69.160 16.815 69.805 17.015 ;
        RECT 68.195 16.725 68.485 16.815 ;
        RECT 69.515 16.725 69.805 16.815 ;
        RECT 70.195 16.815 70.845 17.015 ;
        RECT 71.160 17.015 71.360 18.080 ;
        RECT 72.645 17.015 72.845 18.080 ;
        RECT 71.160 16.815 71.805 17.015 ;
        RECT 70.195 16.725 70.485 16.815 ;
        RECT 71.515 16.725 71.805 16.815 ;
        RECT 72.195 16.815 72.845 17.015 ;
        RECT 73.160 17.015 73.360 18.080 ;
        RECT 74.645 17.015 74.845 18.080 ;
        RECT 73.160 16.815 73.805 17.015 ;
        RECT 72.195 16.725 72.485 16.815 ;
        RECT 73.515 16.725 73.805 16.815 ;
        RECT 74.195 16.815 74.845 17.015 ;
        RECT 75.160 17.015 75.360 18.080 ;
        RECT 76.645 17.015 76.845 18.080 ;
        RECT 75.160 16.815 75.805 17.015 ;
        RECT 74.195 16.725 74.485 16.815 ;
        RECT 75.515 16.725 75.805 16.815 ;
        RECT 76.195 16.815 76.845 17.015 ;
        RECT 77.160 17.015 77.360 18.080 ;
        RECT 78.645 17.015 78.845 18.080 ;
        RECT 77.160 16.815 77.805 17.015 ;
        RECT 76.195 16.725 76.485 16.815 ;
        RECT 77.515 16.725 77.805 16.815 ;
        RECT 78.195 16.815 78.845 17.015 ;
        RECT 79.160 17.015 79.360 18.080 ;
        RECT 80.645 17.015 80.845 18.080 ;
        RECT 79.160 16.815 79.805 17.015 ;
        RECT 78.195 16.725 78.485 16.815 ;
        RECT 79.515 16.725 79.805 16.815 ;
        RECT 80.195 16.815 80.845 17.015 ;
        RECT 81.160 17.015 81.360 18.080 ;
        RECT 82.645 17.015 82.845 18.080 ;
        RECT 81.160 16.815 81.805 17.015 ;
        RECT 80.195 16.725 80.485 16.815 ;
        RECT 81.515 16.725 81.805 16.815 ;
        RECT 82.195 16.815 82.845 17.015 ;
        RECT 83.160 17.015 83.360 18.080 ;
        RECT 84.645 17.015 84.845 18.080 ;
        RECT 83.160 16.815 83.805 17.015 ;
        RECT 82.195 16.725 82.485 16.815 ;
        RECT 83.515 16.725 83.805 16.815 ;
        RECT 84.195 16.815 84.845 17.015 ;
        RECT 85.160 17.015 85.360 18.080 ;
        RECT 86.645 17.015 86.845 18.080 ;
        RECT 85.160 16.815 85.805 17.015 ;
        RECT 84.195 16.725 84.485 16.815 ;
        RECT 85.515 16.725 85.805 16.815 ;
        RECT 86.195 16.815 86.845 17.015 ;
        RECT 87.160 17.015 87.360 18.080 ;
        RECT 88.645 17.015 88.845 18.080 ;
        RECT 87.160 16.815 87.805 17.015 ;
        RECT 86.195 16.725 86.485 16.815 ;
        RECT 87.515 16.725 87.805 16.815 ;
        RECT 88.195 16.815 88.845 17.015 ;
        RECT 89.160 17.015 89.360 18.080 ;
        RECT 90.645 17.015 90.845 18.080 ;
        RECT 89.160 16.815 89.805 17.015 ;
        RECT 88.195 16.725 88.485 16.815 ;
        RECT 89.515 16.725 89.805 16.815 ;
        RECT 90.195 16.815 90.845 17.015 ;
        RECT 91.160 17.015 91.360 18.080 ;
        RECT 92.645 17.015 92.845 18.080 ;
        RECT 91.160 16.815 91.805 17.015 ;
        RECT 90.195 16.725 90.485 16.815 ;
        RECT 91.515 16.725 91.805 16.815 ;
        RECT 92.195 16.815 92.845 17.015 ;
        RECT 93.160 17.015 93.360 18.080 ;
        RECT 94.645 17.015 94.845 18.080 ;
        RECT 93.160 16.815 93.805 17.015 ;
        RECT 92.195 16.725 92.485 16.815 ;
        RECT 93.515 16.725 93.805 16.815 ;
        RECT 94.195 16.815 94.845 17.015 ;
        RECT 95.160 17.015 95.360 18.080 ;
        RECT 96.645 17.015 96.845 18.080 ;
        RECT 95.160 16.815 95.805 17.015 ;
        RECT 94.195 16.725 94.485 16.815 ;
        RECT 95.515 16.725 95.805 16.815 ;
        RECT 96.195 16.815 96.845 17.015 ;
        RECT 97.160 17.015 97.360 18.080 ;
        RECT 98.645 17.015 98.845 18.080 ;
        RECT 97.160 16.815 97.805 17.015 ;
        RECT 96.195 16.725 96.485 16.815 ;
        RECT 97.515 16.725 97.805 16.815 ;
        RECT 98.195 16.815 98.845 17.015 ;
        RECT 99.160 17.015 99.360 18.080 ;
        RECT 100.645 17.015 100.845 18.080 ;
        RECT 99.160 16.815 99.805 17.015 ;
        RECT 98.195 16.725 98.485 16.815 ;
        RECT 99.515 16.725 99.805 16.815 ;
        RECT 100.195 16.815 100.845 17.015 ;
        RECT 101.160 17.015 101.360 18.080 ;
        RECT 102.645 17.015 102.845 18.080 ;
        RECT 101.160 16.815 101.805 17.015 ;
        RECT 100.195 16.725 100.485 16.815 ;
        RECT 101.515 16.725 101.805 16.815 ;
        RECT 102.195 16.815 102.845 17.015 ;
        RECT 103.160 17.015 103.360 18.080 ;
        RECT 104.645 17.015 104.845 18.080 ;
        RECT 103.160 16.815 103.805 17.015 ;
        RECT 102.195 16.725 102.485 16.815 ;
        RECT 103.515 16.725 103.805 16.815 ;
        RECT 104.195 16.815 104.845 17.015 ;
        RECT 105.160 17.015 105.360 18.080 ;
        RECT 106.645 17.015 106.845 18.080 ;
        RECT 105.160 16.815 105.805 17.015 ;
        RECT 104.195 16.725 104.485 16.815 ;
        RECT 105.515 16.725 105.805 16.815 ;
        RECT 106.195 16.815 106.845 17.015 ;
        RECT 107.160 17.015 107.360 18.080 ;
        RECT 108.645 17.015 108.845 18.080 ;
        RECT 107.160 16.815 107.805 17.015 ;
        RECT 106.195 16.725 106.485 16.815 ;
        RECT 107.515 16.725 107.805 16.815 ;
        RECT 108.195 16.815 108.845 17.015 ;
        RECT 109.160 17.015 109.360 18.080 ;
        RECT 110.645 17.015 110.845 18.080 ;
        RECT 109.160 16.815 109.805 17.015 ;
        RECT 108.195 16.725 108.485 16.815 ;
        RECT 109.515 16.725 109.805 16.815 ;
        RECT 110.195 16.815 110.845 17.015 ;
        RECT 111.160 17.015 111.360 18.080 ;
        RECT 112.645 17.015 112.845 18.080 ;
        RECT 111.160 16.815 111.805 17.015 ;
        RECT 110.195 16.725 110.485 16.815 ;
        RECT 111.515 16.725 111.805 16.815 ;
        RECT 112.195 16.815 112.845 17.015 ;
        RECT 113.160 17.015 113.360 18.080 ;
        RECT 114.645 17.015 114.845 18.080 ;
        RECT 113.160 16.815 113.805 17.015 ;
        RECT 112.195 16.725 112.485 16.815 ;
        RECT 113.515 16.725 113.805 16.815 ;
        RECT 114.195 16.815 114.845 17.015 ;
        RECT 115.160 17.015 115.360 18.080 ;
        RECT 116.645 17.015 116.845 18.080 ;
        RECT 115.160 16.815 115.805 17.015 ;
        RECT 114.195 16.725 114.485 16.815 ;
        RECT 115.515 16.725 115.805 16.815 ;
        RECT 116.195 16.815 116.845 17.015 ;
        RECT 117.160 17.015 117.360 18.080 ;
        RECT 118.645 17.015 118.845 18.080 ;
        RECT 117.160 16.815 117.805 17.015 ;
        RECT 116.195 16.725 116.485 16.815 ;
        RECT 117.515 16.725 117.805 16.815 ;
        RECT 118.195 16.815 118.845 17.015 ;
        RECT 119.160 17.015 119.360 18.080 ;
        RECT 120.645 17.015 120.845 18.080 ;
        RECT 119.160 16.815 119.805 17.015 ;
        RECT 118.195 16.725 118.485 16.815 ;
        RECT 119.515 16.725 119.805 16.815 ;
        RECT 120.195 16.815 120.845 17.015 ;
        RECT 121.160 17.015 121.360 18.080 ;
        RECT 122.645 17.015 122.845 18.080 ;
        RECT 121.160 16.815 121.805 17.015 ;
        RECT 120.195 16.725 120.485 16.815 ;
        RECT 121.515 16.725 121.805 16.815 ;
        RECT 122.195 16.815 122.845 17.015 ;
        RECT 123.160 17.015 123.360 18.080 ;
        RECT 124.645 17.015 124.845 18.080 ;
        RECT 123.160 16.815 123.805 17.015 ;
        RECT 122.195 16.725 122.485 16.815 ;
        RECT 123.515 16.725 123.805 16.815 ;
        RECT 124.195 16.815 124.845 17.015 ;
        RECT 125.160 17.015 125.360 18.080 ;
        RECT 126.645 17.015 126.845 18.080 ;
        RECT 125.160 16.815 125.805 17.015 ;
        RECT 124.195 16.725 124.485 16.815 ;
        RECT 125.515 16.725 125.805 16.815 ;
        RECT 126.195 16.815 126.845 17.015 ;
        RECT 127.160 17.015 127.360 18.080 ;
        RECT 128.645 17.015 128.845 18.080 ;
        RECT 127.160 16.815 127.805 17.015 ;
        RECT 126.195 16.725 126.485 16.815 ;
        RECT 127.515 16.725 127.805 16.815 ;
        RECT 128.195 16.815 128.845 17.015 ;
        RECT 129.160 17.015 129.360 18.080 ;
        RECT 130.645 17.015 130.845 18.080 ;
        RECT 129.160 16.815 129.805 17.015 ;
        RECT 128.195 16.725 128.485 16.815 ;
        RECT 129.515 16.725 129.805 16.815 ;
        RECT 130.195 16.815 130.845 17.015 ;
        RECT 130.195 16.725 130.485 16.815 ;
        RECT -1.895 8.920 -1.605 16.720 ;
        RECT -0.145 16.225 0.145 16.515 ;
        RECT -0.100 15.585 0.100 16.225 ;
        RECT 0.365 16.165 0.845 16.515 ;
        RECT 1.855 16.225 2.145 16.515 ;
        RECT 1.900 15.585 2.100 16.225 ;
        RECT 2.365 16.165 2.845 16.515 ;
        RECT 3.855 16.225 4.145 16.515 ;
        RECT 3.900 15.585 4.100 16.225 ;
        RECT 4.365 16.165 4.845 16.515 ;
        RECT 5.855 16.225 6.145 16.515 ;
        RECT 5.900 15.585 6.100 16.225 ;
        RECT 6.365 16.165 6.845 16.515 ;
        RECT 7.855 16.225 8.145 16.515 ;
        RECT 7.900 15.585 8.100 16.225 ;
        RECT 8.365 16.165 8.845 16.515 ;
        RECT 9.855 16.225 10.145 16.515 ;
        RECT 9.900 15.585 10.100 16.225 ;
        RECT 10.365 16.165 10.845 16.515 ;
        RECT 11.855 16.225 12.145 16.515 ;
        RECT 11.900 15.585 12.100 16.225 ;
        RECT 12.365 16.165 12.845 16.515 ;
        RECT 13.855 16.225 14.145 16.515 ;
        RECT 13.900 15.585 14.100 16.225 ;
        RECT 14.365 16.165 14.845 16.515 ;
        RECT 15.855 16.225 16.145 16.515 ;
        RECT 15.900 15.585 16.100 16.225 ;
        RECT 16.365 16.165 16.845 16.515 ;
        RECT 17.855 16.225 18.145 16.515 ;
        RECT 17.900 15.585 18.100 16.225 ;
        RECT 18.365 16.165 18.845 16.515 ;
        RECT 19.855 16.225 20.145 16.515 ;
        RECT 19.900 15.585 20.100 16.225 ;
        RECT 20.365 16.165 20.845 16.515 ;
        RECT 21.855 16.225 22.145 16.515 ;
        RECT 21.900 15.585 22.100 16.225 ;
        RECT 22.365 16.165 22.845 16.515 ;
        RECT 23.855 16.225 24.145 16.515 ;
        RECT 23.900 15.585 24.100 16.225 ;
        RECT 24.365 16.165 24.845 16.515 ;
        RECT 25.855 16.225 26.145 16.515 ;
        RECT 25.900 15.585 26.100 16.225 ;
        RECT 26.365 16.165 26.845 16.515 ;
        RECT 27.855 16.225 28.145 16.515 ;
        RECT 27.900 15.585 28.100 16.225 ;
        RECT 28.365 16.165 28.845 16.515 ;
        RECT 29.855 16.225 30.145 16.515 ;
        RECT 29.900 15.585 30.100 16.225 ;
        RECT 30.365 16.165 30.845 16.515 ;
        RECT 31.855 16.225 32.145 16.515 ;
        RECT 31.900 15.585 32.100 16.225 ;
        RECT 32.365 16.165 32.845 16.515 ;
        RECT 33.855 16.225 34.145 16.515 ;
        RECT 33.900 15.585 34.100 16.225 ;
        RECT 34.365 16.165 34.845 16.515 ;
        RECT 35.855 16.225 36.145 16.515 ;
        RECT 35.900 15.585 36.100 16.225 ;
        RECT 36.365 16.165 36.845 16.515 ;
        RECT 37.855 16.225 38.145 16.515 ;
        RECT 37.900 15.585 38.100 16.225 ;
        RECT 38.365 16.165 38.845 16.515 ;
        RECT 39.855 16.225 40.145 16.515 ;
        RECT 39.900 15.585 40.100 16.225 ;
        RECT 40.365 16.165 40.845 16.515 ;
        RECT 41.855 16.225 42.145 16.515 ;
        RECT 41.900 15.585 42.100 16.225 ;
        RECT 42.365 16.165 42.845 16.515 ;
        RECT 43.855 16.225 44.145 16.515 ;
        RECT 43.900 15.585 44.100 16.225 ;
        RECT 44.365 16.165 44.845 16.515 ;
        RECT 45.855 16.225 46.145 16.515 ;
        RECT 45.900 15.585 46.100 16.225 ;
        RECT 46.365 16.165 46.845 16.515 ;
        RECT 47.855 16.225 48.145 16.515 ;
        RECT 47.900 15.585 48.100 16.225 ;
        RECT 48.365 16.165 48.845 16.515 ;
        RECT 49.855 16.225 50.145 16.515 ;
        RECT 49.900 15.585 50.100 16.225 ;
        RECT 50.365 16.165 50.845 16.515 ;
        RECT 51.855 16.225 52.145 16.515 ;
        RECT 51.900 15.585 52.100 16.225 ;
        RECT 52.365 16.165 52.845 16.515 ;
        RECT 53.855 16.225 54.145 16.515 ;
        RECT 53.900 15.585 54.100 16.225 ;
        RECT 54.365 16.165 54.845 16.515 ;
        RECT 55.855 16.225 56.145 16.515 ;
        RECT 55.900 15.585 56.100 16.225 ;
        RECT 56.365 16.165 56.845 16.515 ;
        RECT 57.855 16.225 58.145 16.515 ;
        RECT 57.900 15.585 58.100 16.225 ;
        RECT 58.365 16.165 58.845 16.515 ;
        RECT 59.855 16.225 60.145 16.515 ;
        RECT 59.900 15.585 60.100 16.225 ;
        RECT 60.365 16.165 60.845 16.515 ;
        RECT 61.855 16.225 62.145 16.515 ;
        RECT 61.900 15.585 62.100 16.225 ;
        RECT 62.365 16.165 62.845 16.515 ;
        RECT 63.855 16.225 64.145 16.515 ;
        RECT 63.900 15.585 64.100 16.225 ;
        RECT 64.365 16.165 64.845 16.515 ;
        RECT 65.855 16.225 66.145 16.515 ;
        RECT 65.900 15.585 66.100 16.225 ;
        RECT 66.365 16.165 66.845 16.515 ;
        RECT 67.855 16.225 68.145 16.515 ;
        RECT 67.900 15.585 68.100 16.225 ;
        RECT 68.365 16.165 68.845 16.515 ;
        RECT 69.855 16.225 70.145 16.515 ;
        RECT 69.900 15.585 70.100 16.225 ;
        RECT 70.365 16.165 70.845 16.515 ;
        RECT 71.855 16.225 72.145 16.515 ;
        RECT 71.900 15.585 72.100 16.225 ;
        RECT 72.365 16.165 72.845 16.515 ;
        RECT 73.855 16.225 74.145 16.515 ;
        RECT 73.900 15.585 74.100 16.225 ;
        RECT 74.365 16.165 74.845 16.515 ;
        RECT 75.855 16.225 76.145 16.515 ;
        RECT 75.900 15.585 76.100 16.225 ;
        RECT 76.365 16.165 76.845 16.515 ;
        RECT 77.855 16.225 78.145 16.515 ;
        RECT 77.900 15.585 78.100 16.225 ;
        RECT 78.365 16.165 78.845 16.515 ;
        RECT 79.855 16.225 80.145 16.515 ;
        RECT 79.900 15.585 80.100 16.225 ;
        RECT 80.365 16.165 80.845 16.515 ;
        RECT 81.855 16.225 82.145 16.515 ;
        RECT 81.900 15.585 82.100 16.225 ;
        RECT 82.365 16.165 82.845 16.515 ;
        RECT 83.855 16.225 84.145 16.515 ;
        RECT 83.900 15.585 84.100 16.225 ;
        RECT 84.365 16.165 84.845 16.515 ;
        RECT 85.855 16.225 86.145 16.515 ;
        RECT 85.900 15.585 86.100 16.225 ;
        RECT 86.365 16.165 86.845 16.515 ;
        RECT 87.855 16.225 88.145 16.515 ;
        RECT 87.900 15.585 88.100 16.225 ;
        RECT 88.365 16.165 88.845 16.515 ;
        RECT 89.855 16.225 90.145 16.515 ;
        RECT 89.900 15.585 90.100 16.225 ;
        RECT 90.365 16.165 90.845 16.515 ;
        RECT 91.855 16.225 92.145 16.515 ;
        RECT 91.900 15.585 92.100 16.225 ;
        RECT 92.365 16.165 92.845 16.515 ;
        RECT 93.855 16.225 94.145 16.515 ;
        RECT 93.900 15.585 94.100 16.225 ;
        RECT 94.365 16.165 94.845 16.515 ;
        RECT 95.855 16.225 96.145 16.515 ;
        RECT 95.900 15.585 96.100 16.225 ;
        RECT 96.365 16.165 96.845 16.515 ;
        RECT 97.855 16.225 98.145 16.515 ;
        RECT 97.900 15.585 98.100 16.225 ;
        RECT 98.365 16.165 98.845 16.515 ;
        RECT 99.855 16.225 100.145 16.515 ;
        RECT 99.900 15.585 100.100 16.225 ;
        RECT 100.365 16.165 100.845 16.515 ;
        RECT 101.855 16.225 102.145 16.515 ;
        RECT 101.900 15.585 102.100 16.225 ;
        RECT 102.365 16.165 102.845 16.515 ;
        RECT 103.855 16.225 104.145 16.515 ;
        RECT 103.900 15.585 104.100 16.225 ;
        RECT 104.365 16.165 104.845 16.515 ;
        RECT 105.855 16.225 106.145 16.515 ;
        RECT 105.900 15.585 106.100 16.225 ;
        RECT 106.365 16.165 106.845 16.515 ;
        RECT 107.855 16.225 108.145 16.515 ;
        RECT 107.900 15.585 108.100 16.225 ;
        RECT 108.365 16.165 108.845 16.515 ;
        RECT 109.855 16.225 110.145 16.515 ;
        RECT 109.900 15.585 110.100 16.225 ;
        RECT 110.365 16.165 110.845 16.515 ;
        RECT 111.855 16.225 112.145 16.515 ;
        RECT 111.900 15.585 112.100 16.225 ;
        RECT 112.365 16.165 112.845 16.515 ;
        RECT 113.855 16.225 114.145 16.515 ;
        RECT 113.900 15.585 114.100 16.225 ;
        RECT 114.365 16.165 114.845 16.515 ;
        RECT 115.855 16.225 116.145 16.515 ;
        RECT 115.900 15.585 116.100 16.225 ;
        RECT 116.365 16.165 116.845 16.515 ;
        RECT 117.855 16.225 118.145 16.515 ;
        RECT 117.900 15.585 118.100 16.225 ;
        RECT 118.365 16.165 118.845 16.515 ;
        RECT 119.855 16.225 120.145 16.515 ;
        RECT 119.900 15.585 120.100 16.225 ;
        RECT 120.365 16.165 120.845 16.515 ;
        RECT 121.855 16.225 122.145 16.515 ;
        RECT 121.900 15.585 122.100 16.225 ;
        RECT 122.365 16.165 122.845 16.515 ;
        RECT 123.855 16.225 124.145 16.515 ;
        RECT 123.900 15.585 124.100 16.225 ;
        RECT 124.365 16.165 124.845 16.515 ;
        RECT 125.855 16.225 126.145 16.515 ;
        RECT 125.900 15.585 126.100 16.225 ;
        RECT 126.365 16.165 126.845 16.515 ;
        RECT 127.855 16.225 128.145 16.515 ;
        RECT 127.900 15.585 128.100 16.225 ;
        RECT 128.365 16.165 128.845 16.515 ;
        RECT 129.855 16.225 130.145 16.515 ;
        RECT 129.900 15.585 130.100 16.225 ;
        RECT 130.365 16.165 130.845 16.515 ;
        RECT -0.100 15.385 0.770 15.585 ;
        RECT 1.900 15.385 2.770 15.585 ;
        RECT 3.900 15.385 4.770 15.585 ;
        RECT 5.900 15.385 6.770 15.585 ;
        RECT 7.900 15.385 8.770 15.585 ;
        RECT 9.900 15.385 10.770 15.585 ;
        RECT 11.900 15.385 12.770 15.585 ;
        RECT 13.900 15.385 14.770 15.585 ;
        RECT 15.900 15.385 16.770 15.585 ;
        RECT 17.900 15.385 18.770 15.585 ;
        RECT 19.900 15.385 20.770 15.585 ;
        RECT 21.900 15.385 22.770 15.585 ;
        RECT 23.900 15.385 24.770 15.585 ;
        RECT 25.900 15.385 26.770 15.585 ;
        RECT 27.900 15.385 28.770 15.585 ;
        RECT 29.900 15.385 30.770 15.585 ;
        RECT 31.900 15.385 32.770 15.585 ;
        RECT 33.900 15.385 34.770 15.585 ;
        RECT 35.900 15.385 36.770 15.585 ;
        RECT 37.900 15.385 38.770 15.585 ;
        RECT 39.900 15.385 40.770 15.585 ;
        RECT 41.900 15.385 42.770 15.585 ;
        RECT 43.900 15.385 44.770 15.585 ;
        RECT 45.900 15.385 46.770 15.585 ;
        RECT 47.900 15.385 48.770 15.585 ;
        RECT 49.900 15.385 50.770 15.585 ;
        RECT 51.900 15.385 52.770 15.585 ;
        RECT 53.900 15.385 54.770 15.585 ;
        RECT 55.900 15.385 56.770 15.585 ;
        RECT 57.900 15.385 58.770 15.585 ;
        RECT 59.900 15.385 60.770 15.585 ;
        RECT 61.900 15.385 62.770 15.585 ;
        RECT 63.900 15.385 64.770 15.585 ;
        RECT 65.900 15.385 66.770 15.585 ;
        RECT 67.900 15.385 68.770 15.585 ;
        RECT 69.900 15.385 70.770 15.585 ;
        RECT 71.900 15.385 72.770 15.585 ;
        RECT 73.900 15.385 74.770 15.585 ;
        RECT 75.900 15.385 76.770 15.585 ;
        RECT 77.900 15.385 78.770 15.585 ;
        RECT 79.900 15.385 80.770 15.585 ;
        RECT 81.900 15.385 82.770 15.585 ;
        RECT 83.900 15.385 84.770 15.585 ;
        RECT 85.900 15.385 86.770 15.585 ;
        RECT 87.900 15.385 88.770 15.585 ;
        RECT 89.900 15.385 90.770 15.585 ;
        RECT 91.900 15.385 92.770 15.585 ;
        RECT 93.900 15.385 94.770 15.585 ;
        RECT 95.900 15.385 96.770 15.585 ;
        RECT 97.900 15.385 98.770 15.585 ;
        RECT 99.900 15.385 100.770 15.585 ;
        RECT 101.900 15.385 102.770 15.585 ;
        RECT 103.900 15.385 104.770 15.585 ;
        RECT 105.900 15.385 106.770 15.585 ;
        RECT 107.900 15.385 108.770 15.585 ;
        RECT 109.900 15.385 110.770 15.585 ;
        RECT 111.900 15.385 112.770 15.585 ;
        RECT 113.900 15.385 114.770 15.585 ;
        RECT 115.900 15.385 116.770 15.585 ;
        RECT 117.900 15.385 118.770 15.585 ;
        RECT 119.900 15.385 120.770 15.585 ;
        RECT 121.900 15.385 122.770 15.585 ;
        RECT 123.900 15.385 124.770 15.585 ;
        RECT 125.900 15.385 126.770 15.585 ;
        RECT 127.900 15.385 128.770 15.585 ;
        RECT 129.900 15.385 130.770 15.585 ;
        RECT 0.570 9.735 0.770 15.385 ;
        RECT 2.570 9.735 2.770 15.385 ;
        RECT 4.570 9.735 4.770 15.385 ;
        RECT 6.570 9.735 6.770 15.385 ;
        RECT 8.570 9.735 8.770 15.385 ;
        RECT 10.570 9.735 10.770 15.385 ;
        RECT 12.570 9.735 12.770 15.385 ;
        RECT 14.570 9.735 14.770 15.385 ;
        RECT 16.570 9.735 16.770 15.385 ;
        RECT 18.570 9.735 18.770 15.385 ;
        RECT 20.570 9.735 20.770 15.385 ;
        RECT 22.570 9.735 22.770 15.385 ;
        RECT 24.570 9.735 24.770 15.385 ;
        RECT 26.570 9.735 26.770 15.385 ;
        RECT 28.570 9.735 28.770 15.385 ;
        RECT 30.570 9.735 30.770 15.385 ;
        RECT 32.570 9.735 32.770 15.385 ;
        RECT 34.570 9.735 34.770 15.385 ;
        RECT 36.570 9.735 36.770 15.385 ;
        RECT 38.570 9.735 38.770 15.385 ;
        RECT 40.570 9.735 40.770 15.385 ;
        RECT 42.570 9.735 42.770 15.385 ;
        RECT 44.570 9.735 44.770 15.385 ;
        RECT 46.570 9.735 46.770 15.385 ;
        RECT 48.570 9.735 48.770 15.385 ;
        RECT 50.570 9.735 50.770 15.385 ;
        RECT 52.570 9.735 52.770 15.385 ;
        RECT 54.570 9.735 54.770 15.385 ;
        RECT 56.570 9.735 56.770 15.385 ;
        RECT 58.570 9.735 58.770 15.385 ;
        RECT 60.570 9.735 60.770 15.385 ;
        RECT 62.570 9.735 62.770 15.385 ;
        RECT 64.570 9.735 64.770 15.385 ;
        RECT 66.570 9.735 66.770 15.385 ;
        RECT 68.570 9.735 68.770 15.385 ;
        RECT 70.570 9.735 70.770 15.385 ;
        RECT 72.570 9.735 72.770 15.385 ;
        RECT 74.570 9.735 74.770 15.385 ;
        RECT 76.570 9.735 76.770 15.385 ;
        RECT 78.570 9.735 78.770 15.385 ;
        RECT 80.570 9.735 80.770 15.385 ;
        RECT 82.570 9.735 82.770 15.385 ;
        RECT 84.570 9.735 84.770 15.385 ;
        RECT 86.570 9.735 86.770 15.385 ;
        RECT 88.570 9.735 88.770 15.385 ;
        RECT 90.570 9.735 90.770 15.385 ;
        RECT 92.570 9.735 92.770 15.385 ;
        RECT 94.570 9.735 94.770 15.385 ;
        RECT 96.570 9.735 96.770 15.385 ;
        RECT 98.570 9.735 98.770 15.385 ;
        RECT 100.570 9.735 100.770 15.385 ;
        RECT 102.570 9.735 102.770 15.385 ;
        RECT 104.570 9.735 104.770 15.385 ;
        RECT 106.570 9.735 106.770 15.385 ;
        RECT 108.570 9.735 108.770 15.385 ;
        RECT 110.570 9.735 110.770 15.385 ;
        RECT 112.570 9.735 112.770 15.385 ;
        RECT 114.570 9.735 114.770 15.385 ;
        RECT 116.570 9.735 116.770 15.385 ;
        RECT 118.570 9.735 118.770 15.385 ;
        RECT 120.570 9.735 120.770 15.385 ;
        RECT 122.570 9.735 122.770 15.385 ;
        RECT 124.570 9.735 124.770 15.385 ;
        RECT 126.570 9.735 126.770 15.385 ;
        RECT 128.570 9.735 128.770 15.385 ;
        RECT 130.570 9.735 130.770 15.385 ;
        RECT 0.560 9.145 0.780 9.735 ;
        RECT 2.560 9.145 2.780 9.735 ;
        RECT 4.560 9.145 4.780 9.735 ;
        RECT 6.560 9.145 6.780 9.735 ;
        RECT 8.560 9.145 8.780 9.735 ;
        RECT 10.560 9.145 10.780 9.735 ;
        RECT 12.560 9.145 12.780 9.735 ;
        RECT 14.560 9.145 14.780 9.735 ;
        RECT 16.560 9.145 16.780 9.735 ;
        RECT 18.560 9.145 18.780 9.735 ;
        RECT 20.560 9.145 20.780 9.735 ;
        RECT 22.560 9.145 22.780 9.735 ;
        RECT 24.560 9.145 24.780 9.735 ;
        RECT 26.560 9.145 26.780 9.735 ;
        RECT 28.560 9.145 28.780 9.735 ;
        RECT 30.560 9.145 30.780 9.735 ;
        RECT 32.560 9.145 32.780 9.735 ;
        RECT 34.560 9.145 34.780 9.735 ;
        RECT 36.560 9.145 36.780 9.735 ;
        RECT 38.560 9.145 38.780 9.735 ;
        RECT 40.560 9.145 40.780 9.735 ;
        RECT 42.560 9.145 42.780 9.735 ;
        RECT 44.560 9.145 44.780 9.735 ;
        RECT 46.560 9.145 46.780 9.735 ;
        RECT 48.560 9.145 48.780 9.735 ;
        RECT 50.560 9.145 50.780 9.735 ;
        RECT 52.560 9.145 52.780 9.735 ;
        RECT 54.560 9.145 54.780 9.735 ;
        RECT 56.560 9.145 56.780 9.735 ;
        RECT 58.560 9.145 58.780 9.735 ;
        RECT 60.560 9.145 60.780 9.735 ;
        RECT 62.560 9.145 62.780 9.735 ;
        RECT 64.560 9.145 64.780 9.735 ;
        RECT 66.560 9.145 66.780 9.735 ;
        RECT 68.560 9.145 68.780 9.735 ;
        RECT 70.560 9.145 70.780 9.735 ;
        RECT 72.560 9.145 72.780 9.735 ;
        RECT 74.560 9.145 74.780 9.735 ;
        RECT 76.560 9.145 76.780 9.735 ;
        RECT 78.560 9.145 78.780 9.735 ;
        RECT 80.560 9.145 80.780 9.735 ;
        RECT 82.560 9.145 82.780 9.735 ;
        RECT 84.560 9.145 84.780 9.735 ;
        RECT 86.560 9.145 86.780 9.735 ;
        RECT 88.560 9.145 88.780 9.735 ;
        RECT 90.560 9.145 90.780 9.735 ;
        RECT 92.560 9.145 92.780 9.735 ;
        RECT 94.560 9.145 94.780 9.735 ;
        RECT 96.560 9.145 96.780 9.735 ;
        RECT 98.560 9.145 98.780 9.735 ;
        RECT 100.560 9.145 100.780 9.735 ;
        RECT 102.560 9.145 102.780 9.735 ;
        RECT 104.560 9.145 104.780 9.735 ;
        RECT 106.560 9.145 106.780 9.735 ;
        RECT 108.560 9.145 108.780 9.735 ;
        RECT 110.560 9.145 110.780 9.735 ;
        RECT 112.560 9.145 112.780 9.735 ;
        RECT 114.560 9.145 114.780 9.735 ;
        RECT 116.560 9.145 116.780 9.735 ;
        RECT 118.560 9.145 118.780 9.735 ;
        RECT 120.560 9.145 120.780 9.735 ;
        RECT 122.560 9.145 122.780 9.735 ;
        RECT 124.560 9.145 124.780 9.735 ;
        RECT 126.560 9.145 126.780 9.735 ;
        RECT 128.560 9.145 128.780 9.735 ;
        RECT 130.560 9.145 130.780 9.735 ;
        RECT 131.605 8.920 131.895 16.720 ;
        RECT -1.895 -0.350 -1.605 7.450 ;
        RECT -0.780 6.635 -0.560 7.225 ;
        RECT 1.220 6.635 1.440 7.225 ;
        RECT 3.220 6.635 3.440 7.225 ;
        RECT 5.220 6.635 5.440 7.225 ;
        RECT 7.220 6.635 7.440 7.225 ;
        RECT 9.220 6.635 9.440 7.225 ;
        RECT 11.220 6.635 11.440 7.225 ;
        RECT 13.220 6.635 13.440 7.225 ;
        RECT 15.220 6.635 15.440 7.225 ;
        RECT 17.220 6.635 17.440 7.225 ;
        RECT 19.220 6.635 19.440 7.225 ;
        RECT 21.220 6.635 21.440 7.225 ;
        RECT 23.220 6.635 23.440 7.225 ;
        RECT 25.220 6.635 25.440 7.225 ;
        RECT 27.220 6.635 27.440 7.225 ;
        RECT 29.220 6.635 29.440 7.225 ;
        RECT 31.220 6.635 31.440 7.225 ;
        RECT 33.220 6.635 33.440 7.225 ;
        RECT 35.220 6.635 35.440 7.225 ;
        RECT 37.220 6.635 37.440 7.225 ;
        RECT 39.220 6.635 39.440 7.225 ;
        RECT 41.220 6.635 41.440 7.225 ;
        RECT 43.220 6.635 43.440 7.225 ;
        RECT 45.220 6.635 45.440 7.225 ;
        RECT 47.220 6.635 47.440 7.225 ;
        RECT 49.220 6.635 49.440 7.225 ;
        RECT 51.220 6.635 51.440 7.225 ;
        RECT 53.220 6.635 53.440 7.225 ;
        RECT 55.220 6.635 55.440 7.225 ;
        RECT 57.220 6.635 57.440 7.225 ;
        RECT 59.220 6.635 59.440 7.225 ;
        RECT 61.220 6.635 61.440 7.225 ;
        RECT 63.220 6.635 63.440 7.225 ;
        RECT 65.220 6.635 65.440 7.225 ;
        RECT 67.220 6.635 67.440 7.225 ;
        RECT 69.220 6.635 69.440 7.225 ;
        RECT 71.220 6.635 71.440 7.225 ;
        RECT 73.220 6.635 73.440 7.225 ;
        RECT 75.220 6.635 75.440 7.225 ;
        RECT 77.220 6.635 77.440 7.225 ;
        RECT 79.220 6.635 79.440 7.225 ;
        RECT 81.220 6.635 81.440 7.225 ;
        RECT 83.220 6.635 83.440 7.225 ;
        RECT 85.220 6.635 85.440 7.225 ;
        RECT 87.220 6.635 87.440 7.225 ;
        RECT 89.220 6.635 89.440 7.225 ;
        RECT 91.220 6.635 91.440 7.225 ;
        RECT 93.220 6.635 93.440 7.225 ;
        RECT 95.220 6.635 95.440 7.225 ;
        RECT 97.220 6.635 97.440 7.225 ;
        RECT 99.220 6.635 99.440 7.225 ;
        RECT 101.220 6.635 101.440 7.225 ;
        RECT 103.220 6.635 103.440 7.225 ;
        RECT 105.220 6.635 105.440 7.225 ;
        RECT 107.220 6.635 107.440 7.225 ;
        RECT 109.220 6.635 109.440 7.225 ;
        RECT 111.220 6.635 111.440 7.225 ;
        RECT 113.220 6.635 113.440 7.225 ;
        RECT 115.220 6.635 115.440 7.225 ;
        RECT 117.220 6.635 117.440 7.225 ;
        RECT 119.220 6.635 119.440 7.225 ;
        RECT 121.220 6.635 121.440 7.225 ;
        RECT 123.220 6.635 123.440 7.225 ;
        RECT 125.220 6.635 125.440 7.225 ;
        RECT 127.220 6.635 127.440 7.225 ;
        RECT 129.220 6.635 129.440 7.225 ;
        RECT -0.770 0.985 -0.570 6.635 ;
        RECT 1.230 0.985 1.430 6.635 ;
        RECT 3.230 0.985 3.430 6.635 ;
        RECT 5.230 0.985 5.430 6.635 ;
        RECT 7.230 0.985 7.430 6.635 ;
        RECT 9.230 0.985 9.430 6.635 ;
        RECT 11.230 0.985 11.430 6.635 ;
        RECT 13.230 0.985 13.430 6.635 ;
        RECT 15.230 0.985 15.430 6.635 ;
        RECT 17.230 0.985 17.430 6.635 ;
        RECT 19.230 0.985 19.430 6.635 ;
        RECT 21.230 0.985 21.430 6.635 ;
        RECT 23.230 0.985 23.430 6.635 ;
        RECT 25.230 0.985 25.430 6.635 ;
        RECT 27.230 0.985 27.430 6.635 ;
        RECT 29.230 0.985 29.430 6.635 ;
        RECT 31.230 0.985 31.430 6.635 ;
        RECT 33.230 0.985 33.430 6.635 ;
        RECT 35.230 0.985 35.430 6.635 ;
        RECT 37.230 0.985 37.430 6.635 ;
        RECT 39.230 0.985 39.430 6.635 ;
        RECT 41.230 0.985 41.430 6.635 ;
        RECT 43.230 0.985 43.430 6.635 ;
        RECT 45.230 0.985 45.430 6.635 ;
        RECT 47.230 0.985 47.430 6.635 ;
        RECT 49.230 0.985 49.430 6.635 ;
        RECT 51.230 0.985 51.430 6.635 ;
        RECT 53.230 0.985 53.430 6.635 ;
        RECT 55.230 0.985 55.430 6.635 ;
        RECT 57.230 0.985 57.430 6.635 ;
        RECT 59.230 0.985 59.430 6.635 ;
        RECT 61.230 0.985 61.430 6.635 ;
        RECT 63.230 0.985 63.430 6.635 ;
        RECT 65.230 0.985 65.430 6.635 ;
        RECT 67.230 0.985 67.430 6.635 ;
        RECT 69.230 0.985 69.430 6.635 ;
        RECT 71.230 0.985 71.430 6.635 ;
        RECT 73.230 0.985 73.430 6.635 ;
        RECT 75.230 0.985 75.430 6.635 ;
        RECT 77.230 0.985 77.430 6.635 ;
        RECT 79.230 0.985 79.430 6.635 ;
        RECT 81.230 0.985 81.430 6.635 ;
        RECT 83.230 0.985 83.430 6.635 ;
        RECT 85.230 0.985 85.430 6.635 ;
        RECT 87.230 0.985 87.430 6.635 ;
        RECT 89.230 0.985 89.430 6.635 ;
        RECT 91.230 0.985 91.430 6.635 ;
        RECT 93.230 0.985 93.430 6.635 ;
        RECT 95.230 0.985 95.430 6.635 ;
        RECT 97.230 0.985 97.430 6.635 ;
        RECT 99.230 0.985 99.430 6.635 ;
        RECT 101.230 0.985 101.430 6.635 ;
        RECT 103.230 0.985 103.430 6.635 ;
        RECT 105.230 0.985 105.430 6.635 ;
        RECT 107.230 0.985 107.430 6.635 ;
        RECT 109.230 0.985 109.430 6.635 ;
        RECT 111.230 0.985 111.430 6.635 ;
        RECT 113.230 0.985 113.430 6.635 ;
        RECT 115.230 0.985 115.430 6.635 ;
        RECT 117.230 0.985 117.430 6.635 ;
        RECT 119.230 0.985 119.430 6.635 ;
        RECT 121.230 0.985 121.430 6.635 ;
        RECT 123.230 0.985 123.430 6.635 ;
        RECT 125.230 0.985 125.430 6.635 ;
        RECT 127.230 0.985 127.430 6.635 ;
        RECT 129.230 0.985 129.430 6.635 ;
        RECT -0.770 0.785 0.100 0.985 ;
        RECT 1.230 0.785 2.100 0.985 ;
        RECT 3.230 0.785 4.100 0.985 ;
        RECT 5.230 0.785 6.100 0.985 ;
        RECT 7.230 0.785 8.100 0.985 ;
        RECT 9.230 0.785 10.100 0.985 ;
        RECT 11.230 0.785 12.100 0.985 ;
        RECT 13.230 0.785 14.100 0.985 ;
        RECT 15.230 0.785 16.100 0.985 ;
        RECT 17.230 0.785 18.100 0.985 ;
        RECT 19.230 0.785 20.100 0.985 ;
        RECT 21.230 0.785 22.100 0.985 ;
        RECT 23.230 0.785 24.100 0.985 ;
        RECT 25.230 0.785 26.100 0.985 ;
        RECT 27.230 0.785 28.100 0.985 ;
        RECT 29.230 0.785 30.100 0.985 ;
        RECT 31.230 0.785 32.100 0.985 ;
        RECT 33.230 0.785 34.100 0.985 ;
        RECT 35.230 0.785 36.100 0.985 ;
        RECT 37.230 0.785 38.100 0.985 ;
        RECT 39.230 0.785 40.100 0.985 ;
        RECT 41.230 0.785 42.100 0.985 ;
        RECT 43.230 0.785 44.100 0.985 ;
        RECT 45.230 0.785 46.100 0.985 ;
        RECT 47.230 0.785 48.100 0.985 ;
        RECT 49.230 0.785 50.100 0.985 ;
        RECT 51.230 0.785 52.100 0.985 ;
        RECT 53.230 0.785 54.100 0.985 ;
        RECT 55.230 0.785 56.100 0.985 ;
        RECT 57.230 0.785 58.100 0.985 ;
        RECT 59.230 0.785 60.100 0.985 ;
        RECT 61.230 0.785 62.100 0.985 ;
        RECT 63.230 0.785 64.100 0.985 ;
        RECT 65.230 0.785 66.100 0.985 ;
        RECT 67.230 0.785 68.100 0.985 ;
        RECT 69.230 0.785 70.100 0.985 ;
        RECT 71.230 0.785 72.100 0.985 ;
        RECT 73.230 0.785 74.100 0.985 ;
        RECT 75.230 0.785 76.100 0.985 ;
        RECT 77.230 0.785 78.100 0.985 ;
        RECT 79.230 0.785 80.100 0.985 ;
        RECT 81.230 0.785 82.100 0.985 ;
        RECT 83.230 0.785 84.100 0.985 ;
        RECT 85.230 0.785 86.100 0.985 ;
        RECT 87.230 0.785 88.100 0.985 ;
        RECT 89.230 0.785 90.100 0.985 ;
        RECT 91.230 0.785 92.100 0.985 ;
        RECT 93.230 0.785 94.100 0.985 ;
        RECT 95.230 0.785 96.100 0.985 ;
        RECT 97.230 0.785 98.100 0.985 ;
        RECT 99.230 0.785 100.100 0.985 ;
        RECT 101.230 0.785 102.100 0.985 ;
        RECT 103.230 0.785 104.100 0.985 ;
        RECT 105.230 0.785 106.100 0.985 ;
        RECT 107.230 0.785 108.100 0.985 ;
        RECT 109.230 0.785 110.100 0.985 ;
        RECT 111.230 0.785 112.100 0.985 ;
        RECT 113.230 0.785 114.100 0.985 ;
        RECT 115.230 0.785 116.100 0.985 ;
        RECT 117.230 0.785 118.100 0.985 ;
        RECT 119.230 0.785 120.100 0.985 ;
        RECT 121.230 0.785 122.100 0.985 ;
        RECT 123.230 0.785 124.100 0.985 ;
        RECT 125.230 0.785 126.100 0.985 ;
        RECT 127.230 0.785 128.100 0.985 ;
        RECT 129.230 0.785 130.100 0.985 ;
        RECT -0.845 -0.145 -0.365 0.205 ;
        RECT -0.100 0.145 0.100 0.785 ;
        RECT -0.145 -0.145 0.145 0.145 ;
        RECT 1.155 -0.145 1.635 0.205 ;
        RECT 1.900 0.145 2.100 0.785 ;
        RECT 1.855 -0.145 2.145 0.145 ;
        RECT 3.155 -0.145 3.635 0.205 ;
        RECT 3.900 0.145 4.100 0.785 ;
        RECT 3.855 -0.145 4.145 0.145 ;
        RECT 5.155 -0.145 5.635 0.205 ;
        RECT 5.900 0.145 6.100 0.785 ;
        RECT 5.855 -0.145 6.145 0.145 ;
        RECT 7.155 -0.145 7.635 0.205 ;
        RECT 7.900 0.145 8.100 0.785 ;
        RECT 7.855 -0.145 8.145 0.145 ;
        RECT 9.155 -0.145 9.635 0.205 ;
        RECT 9.900 0.145 10.100 0.785 ;
        RECT 9.855 -0.145 10.145 0.145 ;
        RECT 11.155 -0.145 11.635 0.205 ;
        RECT 11.900 0.145 12.100 0.785 ;
        RECT 11.855 -0.145 12.145 0.145 ;
        RECT 13.155 -0.145 13.635 0.205 ;
        RECT 13.900 0.145 14.100 0.785 ;
        RECT 13.855 -0.145 14.145 0.145 ;
        RECT 15.155 -0.145 15.635 0.205 ;
        RECT 15.900 0.145 16.100 0.785 ;
        RECT 15.855 -0.145 16.145 0.145 ;
        RECT 17.155 -0.145 17.635 0.205 ;
        RECT 17.900 0.145 18.100 0.785 ;
        RECT 17.855 -0.145 18.145 0.145 ;
        RECT 19.155 -0.145 19.635 0.205 ;
        RECT 19.900 0.145 20.100 0.785 ;
        RECT 19.855 -0.145 20.145 0.145 ;
        RECT 21.155 -0.145 21.635 0.205 ;
        RECT 21.900 0.145 22.100 0.785 ;
        RECT 21.855 -0.145 22.145 0.145 ;
        RECT 23.155 -0.145 23.635 0.205 ;
        RECT 23.900 0.145 24.100 0.785 ;
        RECT 23.855 -0.145 24.145 0.145 ;
        RECT 25.155 -0.145 25.635 0.205 ;
        RECT 25.900 0.145 26.100 0.785 ;
        RECT 25.855 -0.145 26.145 0.145 ;
        RECT 27.155 -0.145 27.635 0.205 ;
        RECT 27.900 0.145 28.100 0.785 ;
        RECT 27.855 -0.145 28.145 0.145 ;
        RECT 29.155 -0.145 29.635 0.205 ;
        RECT 29.900 0.145 30.100 0.785 ;
        RECT 29.855 -0.145 30.145 0.145 ;
        RECT 31.155 -0.145 31.635 0.205 ;
        RECT 31.900 0.145 32.100 0.785 ;
        RECT 31.855 -0.145 32.145 0.145 ;
        RECT 33.155 -0.145 33.635 0.205 ;
        RECT 33.900 0.145 34.100 0.785 ;
        RECT 33.855 -0.145 34.145 0.145 ;
        RECT 35.155 -0.145 35.635 0.205 ;
        RECT 35.900 0.145 36.100 0.785 ;
        RECT 35.855 -0.145 36.145 0.145 ;
        RECT 37.155 -0.145 37.635 0.205 ;
        RECT 37.900 0.145 38.100 0.785 ;
        RECT 37.855 -0.145 38.145 0.145 ;
        RECT 39.155 -0.145 39.635 0.205 ;
        RECT 39.900 0.145 40.100 0.785 ;
        RECT 39.855 -0.145 40.145 0.145 ;
        RECT 41.155 -0.145 41.635 0.205 ;
        RECT 41.900 0.145 42.100 0.785 ;
        RECT 41.855 -0.145 42.145 0.145 ;
        RECT 43.155 -0.145 43.635 0.205 ;
        RECT 43.900 0.145 44.100 0.785 ;
        RECT 43.855 -0.145 44.145 0.145 ;
        RECT 45.155 -0.145 45.635 0.205 ;
        RECT 45.900 0.145 46.100 0.785 ;
        RECT 45.855 -0.145 46.145 0.145 ;
        RECT 47.155 -0.145 47.635 0.205 ;
        RECT 47.900 0.145 48.100 0.785 ;
        RECT 47.855 -0.145 48.145 0.145 ;
        RECT 49.155 -0.145 49.635 0.205 ;
        RECT 49.900 0.145 50.100 0.785 ;
        RECT 49.855 -0.145 50.145 0.145 ;
        RECT 51.155 -0.145 51.635 0.205 ;
        RECT 51.900 0.145 52.100 0.785 ;
        RECT 51.855 -0.145 52.145 0.145 ;
        RECT 53.155 -0.145 53.635 0.205 ;
        RECT 53.900 0.145 54.100 0.785 ;
        RECT 53.855 -0.145 54.145 0.145 ;
        RECT 55.155 -0.145 55.635 0.205 ;
        RECT 55.900 0.145 56.100 0.785 ;
        RECT 55.855 -0.145 56.145 0.145 ;
        RECT 57.155 -0.145 57.635 0.205 ;
        RECT 57.900 0.145 58.100 0.785 ;
        RECT 57.855 -0.145 58.145 0.145 ;
        RECT 59.155 -0.145 59.635 0.205 ;
        RECT 59.900 0.145 60.100 0.785 ;
        RECT 59.855 -0.145 60.145 0.145 ;
        RECT 61.155 -0.145 61.635 0.205 ;
        RECT 61.900 0.145 62.100 0.785 ;
        RECT 61.855 -0.145 62.145 0.145 ;
        RECT 63.155 -0.145 63.635 0.205 ;
        RECT 63.900 0.145 64.100 0.785 ;
        RECT 63.855 -0.145 64.145 0.145 ;
        RECT 65.155 -0.145 65.635 0.205 ;
        RECT 65.900 0.145 66.100 0.785 ;
        RECT 65.855 -0.145 66.145 0.145 ;
        RECT 67.155 -0.145 67.635 0.205 ;
        RECT 67.900 0.145 68.100 0.785 ;
        RECT 67.855 -0.145 68.145 0.145 ;
        RECT 69.155 -0.145 69.635 0.205 ;
        RECT 69.900 0.145 70.100 0.785 ;
        RECT 69.855 -0.145 70.145 0.145 ;
        RECT 71.155 -0.145 71.635 0.205 ;
        RECT 71.900 0.145 72.100 0.785 ;
        RECT 71.855 -0.145 72.145 0.145 ;
        RECT 73.155 -0.145 73.635 0.205 ;
        RECT 73.900 0.145 74.100 0.785 ;
        RECT 73.855 -0.145 74.145 0.145 ;
        RECT 75.155 -0.145 75.635 0.205 ;
        RECT 75.900 0.145 76.100 0.785 ;
        RECT 75.855 -0.145 76.145 0.145 ;
        RECT 77.155 -0.145 77.635 0.205 ;
        RECT 77.900 0.145 78.100 0.785 ;
        RECT 77.855 -0.145 78.145 0.145 ;
        RECT 79.155 -0.145 79.635 0.205 ;
        RECT 79.900 0.145 80.100 0.785 ;
        RECT 79.855 -0.145 80.145 0.145 ;
        RECT 81.155 -0.145 81.635 0.205 ;
        RECT 81.900 0.145 82.100 0.785 ;
        RECT 81.855 -0.145 82.145 0.145 ;
        RECT 83.155 -0.145 83.635 0.205 ;
        RECT 83.900 0.145 84.100 0.785 ;
        RECT 83.855 -0.145 84.145 0.145 ;
        RECT 85.155 -0.145 85.635 0.205 ;
        RECT 85.900 0.145 86.100 0.785 ;
        RECT 85.855 -0.145 86.145 0.145 ;
        RECT 87.155 -0.145 87.635 0.205 ;
        RECT 87.900 0.145 88.100 0.785 ;
        RECT 87.855 -0.145 88.145 0.145 ;
        RECT 89.155 -0.145 89.635 0.205 ;
        RECT 89.900 0.145 90.100 0.785 ;
        RECT 89.855 -0.145 90.145 0.145 ;
        RECT 91.155 -0.145 91.635 0.205 ;
        RECT 91.900 0.145 92.100 0.785 ;
        RECT 91.855 -0.145 92.145 0.145 ;
        RECT 93.155 -0.145 93.635 0.205 ;
        RECT 93.900 0.145 94.100 0.785 ;
        RECT 93.855 -0.145 94.145 0.145 ;
        RECT 95.155 -0.145 95.635 0.205 ;
        RECT 95.900 0.145 96.100 0.785 ;
        RECT 95.855 -0.145 96.145 0.145 ;
        RECT 97.155 -0.145 97.635 0.205 ;
        RECT 97.900 0.145 98.100 0.785 ;
        RECT 97.855 -0.145 98.145 0.145 ;
        RECT 99.155 -0.145 99.635 0.205 ;
        RECT 99.900 0.145 100.100 0.785 ;
        RECT 99.855 -0.145 100.145 0.145 ;
        RECT 101.155 -0.145 101.635 0.205 ;
        RECT 101.900 0.145 102.100 0.785 ;
        RECT 101.855 -0.145 102.145 0.145 ;
        RECT 103.155 -0.145 103.635 0.205 ;
        RECT 103.900 0.145 104.100 0.785 ;
        RECT 103.855 -0.145 104.145 0.145 ;
        RECT 105.155 -0.145 105.635 0.205 ;
        RECT 105.900 0.145 106.100 0.785 ;
        RECT 105.855 -0.145 106.145 0.145 ;
        RECT 107.155 -0.145 107.635 0.205 ;
        RECT 107.900 0.145 108.100 0.785 ;
        RECT 107.855 -0.145 108.145 0.145 ;
        RECT 109.155 -0.145 109.635 0.205 ;
        RECT 109.900 0.145 110.100 0.785 ;
        RECT 109.855 -0.145 110.145 0.145 ;
        RECT 111.155 -0.145 111.635 0.205 ;
        RECT 111.900 0.145 112.100 0.785 ;
        RECT 111.855 -0.145 112.145 0.145 ;
        RECT 113.155 -0.145 113.635 0.205 ;
        RECT 113.900 0.145 114.100 0.785 ;
        RECT 113.855 -0.145 114.145 0.145 ;
        RECT 115.155 -0.145 115.635 0.205 ;
        RECT 115.900 0.145 116.100 0.785 ;
        RECT 115.855 -0.145 116.145 0.145 ;
        RECT 117.155 -0.145 117.635 0.205 ;
        RECT 117.900 0.145 118.100 0.785 ;
        RECT 117.855 -0.145 118.145 0.145 ;
        RECT 119.155 -0.145 119.635 0.205 ;
        RECT 119.900 0.145 120.100 0.785 ;
        RECT 119.855 -0.145 120.145 0.145 ;
        RECT 121.155 -0.145 121.635 0.205 ;
        RECT 121.900 0.145 122.100 0.785 ;
        RECT 121.855 -0.145 122.145 0.145 ;
        RECT 123.155 -0.145 123.635 0.205 ;
        RECT 123.900 0.145 124.100 0.785 ;
        RECT 123.855 -0.145 124.145 0.145 ;
        RECT 125.155 -0.145 125.635 0.205 ;
        RECT 125.900 0.145 126.100 0.785 ;
        RECT 125.855 -0.145 126.145 0.145 ;
        RECT 127.155 -0.145 127.635 0.205 ;
        RECT 127.900 0.145 128.100 0.785 ;
        RECT 127.855 -0.145 128.145 0.145 ;
        RECT 129.155 -0.145 129.635 0.205 ;
        RECT 129.900 0.145 130.100 0.785 ;
        RECT 129.855 -0.145 130.145 0.145 ;
        RECT 131.605 -0.350 131.895 7.450 ;
        RECT -0.485 -0.445 -0.195 -0.355 ;
        RECT -0.845 -0.645 -0.195 -0.445 ;
        RECT 0.195 -0.445 0.485 -0.355 ;
        RECT 1.515 -0.445 1.805 -0.355 ;
        RECT 0.195 -0.645 0.840 -0.445 ;
        RECT -0.845 -1.710 -0.645 -0.645 ;
        RECT 0.640 -1.710 0.840 -0.645 ;
        RECT 1.155 -0.645 1.805 -0.445 ;
        RECT 2.195 -0.445 2.485 -0.355 ;
        RECT 3.515 -0.445 3.805 -0.355 ;
        RECT 2.195 -0.645 2.840 -0.445 ;
        RECT 1.155 -1.710 1.355 -0.645 ;
        RECT 2.640 -1.710 2.840 -0.645 ;
        RECT 3.155 -0.645 3.805 -0.445 ;
        RECT 4.195 -0.445 4.485 -0.355 ;
        RECT 5.515 -0.445 5.805 -0.355 ;
        RECT 4.195 -0.645 4.840 -0.445 ;
        RECT 3.155 -1.710 3.355 -0.645 ;
        RECT 4.640 -1.710 4.840 -0.645 ;
        RECT 5.155 -0.645 5.805 -0.445 ;
        RECT 6.195 -0.445 6.485 -0.355 ;
        RECT 7.515 -0.445 7.805 -0.355 ;
        RECT 6.195 -0.645 6.840 -0.445 ;
        RECT 5.155 -1.710 5.355 -0.645 ;
        RECT 6.640 -1.710 6.840 -0.645 ;
        RECT 7.155 -0.645 7.805 -0.445 ;
        RECT 8.195 -0.445 8.485 -0.355 ;
        RECT 9.515 -0.445 9.805 -0.355 ;
        RECT 8.195 -0.645 8.840 -0.445 ;
        RECT 7.155 -1.710 7.355 -0.645 ;
        RECT 8.640 -1.710 8.840 -0.645 ;
        RECT 9.155 -0.645 9.805 -0.445 ;
        RECT 10.195 -0.445 10.485 -0.355 ;
        RECT 11.515 -0.445 11.805 -0.355 ;
        RECT 10.195 -0.645 10.840 -0.445 ;
        RECT 9.155 -1.710 9.355 -0.645 ;
        RECT 10.640 -1.710 10.840 -0.645 ;
        RECT 11.155 -0.645 11.805 -0.445 ;
        RECT 12.195 -0.445 12.485 -0.355 ;
        RECT 13.515 -0.445 13.805 -0.355 ;
        RECT 12.195 -0.645 12.840 -0.445 ;
        RECT 11.155 -1.710 11.355 -0.645 ;
        RECT 12.640 -1.710 12.840 -0.645 ;
        RECT 13.155 -0.645 13.805 -0.445 ;
        RECT 14.195 -0.445 14.485 -0.355 ;
        RECT 15.515 -0.445 15.805 -0.355 ;
        RECT 14.195 -0.645 14.840 -0.445 ;
        RECT 13.155 -1.710 13.355 -0.645 ;
        RECT 14.640 -1.710 14.840 -0.645 ;
        RECT 15.155 -0.645 15.805 -0.445 ;
        RECT 16.195 -0.445 16.485 -0.355 ;
        RECT 17.515 -0.445 17.805 -0.355 ;
        RECT 16.195 -0.645 16.840 -0.445 ;
        RECT 15.155 -1.710 15.355 -0.645 ;
        RECT 16.640 -1.710 16.840 -0.645 ;
        RECT 17.155 -0.645 17.805 -0.445 ;
        RECT 18.195 -0.445 18.485 -0.355 ;
        RECT 19.515 -0.445 19.805 -0.355 ;
        RECT 18.195 -0.645 18.840 -0.445 ;
        RECT 17.155 -1.710 17.355 -0.645 ;
        RECT 18.640 -1.710 18.840 -0.645 ;
        RECT 19.155 -0.645 19.805 -0.445 ;
        RECT 20.195 -0.445 20.485 -0.355 ;
        RECT 21.515 -0.445 21.805 -0.355 ;
        RECT 20.195 -0.645 20.840 -0.445 ;
        RECT 19.155 -1.710 19.355 -0.645 ;
        RECT 20.640 -1.710 20.840 -0.645 ;
        RECT 21.155 -0.645 21.805 -0.445 ;
        RECT 22.195 -0.445 22.485 -0.355 ;
        RECT 23.515 -0.445 23.805 -0.355 ;
        RECT 22.195 -0.645 22.840 -0.445 ;
        RECT 21.155 -1.710 21.355 -0.645 ;
        RECT 22.640 -1.710 22.840 -0.645 ;
        RECT 23.155 -0.645 23.805 -0.445 ;
        RECT 24.195 -0.445 24.485 -0.355 ;
        RECT 25.515 -0.445 25.805 -0.355 ;
        RECT 24.195 -0.645 24.840 -0.445 ;
        RECT 23.155 -1.710 23.355 -0.645 ;
        RECT 24.640 -1.710 24.840 -0.645 ;
        RECT 25.155 -0.645 25.805 -0.445 ;
        RECT 26.195 -0.445 26.485 -0.355 ;
        RECT 27.515 -0.445 27.805 -0.355 ;
        RECT 26.195 -0.645 26.840 -0.445 ;
        RECT 25.155 -1.710 25.355 -0.645 ;
        RECT 26.640 -1.710 26.840 -0.645 ;
        RECT 27.155 -0.645 27.805 -0.445 ;
        RECT 28.195 -0.445 28.485 -0.355 ;
        RECT 29.515 -0.445 29.805 -0.355 ;
        RECT 28.195 -0.645 28.840 -0.445 ;
        RECT 27.155 -1.710 27.355 -0.645 ;
        RECT 28.640 -1.710 28.840 -0.645 ;
        RECT 29.155 -0.645 29.805 -0.445 ;
        RECT 30.195 -0.445 30.485 -0.355 ;
        RECT 31.515 -0.445 31.805 -0.355 ;
        RECT 30.195 -0.645 30.840 -0.445 ;
        RECT 29.155 -1.710 29.355 -0.645 ;
        RECT 30.640 -1.710 30.840 -0.645 ;
        RECT 31.155 -0.645 31.805 -0.445 ;
        RECT 32.195 -0.445 32.485 -0.355 ;
        RECT 33.515 -0.445 33.805 -0.355 ;
        RECT 32.195 -0.645 32.840 -0.445 ;
        RECT 31.155 -1.710 31.355 -0.645 ;
        RECT 32.640 -1.710 32.840 -0.645 ;
        RECT 33.155 -0.645 33.805 -0.445 ;
        RECT 34.195 -0.445 34.485 -0.355 ;
        RECT 35.515 -0.445 35.805 -0.355 ;
        RECT 34.195 -0.645 34.840 -0.445 ;
        RECT 33.155 -1.710 33.355 -0.645 ;
        RECT 34.640 -1.710 34.840 -0.645 ;
        RECT 35.155 -0.645 35.805 -0.445 ;
        RECT 36.195 -0.445 36.485 -0.355 ;
        RECT 37.515 -0.445 37.805 -0.355 ;
        RECT 36.195 -0.645 36.840 -0.445 ;
        RECT 35.155 -1.710 35.355 -0.645 ;
        RECT 36.640 -1.710 36.840 -0.645 ;
        RECT 37.155 -0.645 37.805 -0.445 ;
        RECT 38.195 -0.445 38.485 -0.355 ;
        RECT 39.515 -0.445 39.805 -0.355 ;
        RECT 38.195 -0.645 38.840 -0.445 ;
        RECT 37.155 -1.710 37.355 -0.645 ;
        RECT 38.640 -1.710 38.840 -0.645 ;
        RECT 39.155 -0.645 39.805 -0.445 ;
        RECT 40.195 -0.445 40.485 -0.355 ;
        RECT 41.515 -0.445 41.805 -0.355 ;
        RECT 40.195 -0.645 40.840 -0.445 ;
        RECT 39.155 -1.710 39.355 -0.645 ;
        RECT 40.640 -1.710 40.840 -0.645 ;
        RECT 41.155 -0.645 41.805 -0.445 ;
        RECT 42.195 -0.445 42.485 -0.355 ;
        RECT 43.515 -0.445 43.805 -0.355 ;
        RECT 42.195 -0.645 42.840 -0.445 ;
        RECT 41.155 -1.710 41.355 -0.645 ;
        RECT 42.640 -1.710 42.840 -0.645 ;
        RECT 43.155 -0.645 43.805 -0.445 ;
        RECT 44.195 -0.445 44.485 -0.355 ;
        RECT 45.515 -0.445 45.805 -0.355 ;
        RECT 44.195 -0.645 44.840 -0.445 ;
        RECT 43.155 -1.710 43.355 -0.645 ;
        RECT 44.640 -1.710 44.840 -0.645 ;
        RECT 45.155 -0.645 45.805 -0.445 ;
        RECT 46.195 -0.445 46.485 -0.355 ;
        RECT 47.515 -0.445 47.805 -0.355 ;
        RECT 46.195 -0.645 46.840 -0.445 ;
        RECT 45.155 -1.710 45.355 -0.645 ;
        RECT 46.640 -1.710 46.840 -0.645 ;
        RECT 47.155 -0.645 47.805 -0.445 ;
        RECT 48.195 -0.445 48.485 -0.355 ;
        RECT 49.515 -0.445 49.805 -0.355 ;
        RECT 48.195 -0.645 48.840 -0.445 ;
        RECT 47.155 -1.710 47.355 -0.645 ;
        RECT 48.640 -1.710 48.840 -0.645 ;
        RECT 49.155 -0.645 49.805 -0.445 ;
        RECT 50.195 -0.445 50.485 -0.355 ;
        RECT 51.515 -0.445 51.805 -0.355 ;
        RECT 50.195 -0.645 50.840 -0.445 ;
        RECT 49.155 -1.710 49.355 -0.645 ;
        RECT 50.640 -1.710 50.840 -0.645 ;
        RECT 51.155 -0.645 51.805 -0.445 ;
        RECT 52.195 -0.445 52.485 -0.355 ;
        RECT 53.515 -0.445 53.805 -0.355 ;
        RECT 52.195 -0.645 52.840 -0.445 ;
        RECT 51.155 -1.710 51.355 -0.645 ;
        RECT 52.640 -1.710 52.840 -0.645 ;
        RECT 53.155 -0.645 53.805 -0.445 ;
        RECT 54.195 -0.445 54.485 -0.355 ;
        RECT 55.515 -0.445 55.805 -0.355 ;
        RECT 54.195 -0.645 54.840 -0.445 ;
        RECT 53.155 -1.710 53.355 -0.645 ;
        RECT 54.640 -1.710 54.840 -0.645 ;
        RECT 55.155 -0.645 55.805 -0.445 ;
        RECT 56.195 -0.445 56.485 -0.355 ;
        RECT 57.515 -0.445 57.805 -0.355 ;
        RECT 56.195 -0.645 56.840 -0.445 ;
        RECT 55.155 -1.710 55.355 -0.645 ;
        RECT 56.640 -1.710 56.840 -0.645 ;
        RECT 57.155 -0.645 57.805 -0.445 ;
        RECT 58.195 -0.445 58.485 -0.355 ;
        RECT 59.515 -0.445 59.805 -0.355 ;
        RECT 58.195 -0.645 58.840 -0.445 ;
        RECT 57.155 -1.710 57.355 -0.645 ;
        RECT 58.640 -1.710 58.840 -0.645 ;
        RECT 59.155 -0.645 59.805 -0.445 ;
        RECT 60.195 -0.445 60.485 -0.355 ;
        RECT 61.515 -0.445 61.805 -0.355 ;
        RECT 60.195 -0.645 60.840 -0.445 ;
        RECT 59.155 -1.710 59.355 -0.645 ;
        RECT 60.640 -1.710 60.840 -0.645 ;
        RECT 61.155 -0.645 61.805 -0.445 ;
        RECT 62.195 -0.445 62.485 -0.355 ;
        RECT 63.515 -0.445 63.805 -0.355 ;
        RECT 62.195 -0.645 62.840 -0.445 ;
        RECT 61.155 -1.710 61.355 -0.645 ;
        RECT 62.640 -1.710 62.840 -0.645 ;
        RECT 63.155 -0.645 63.805 -0.445 ;
        RECT 64.195 -0.445 64.485 -0.355 ;
        RECT 65.515 -0.445 65.805 -0.355 ;
        RECT 64.195 -0.645 64.840 -0.445 ;
        RECT 63.155 -1.710 63.355 -0.645 ;
        RECT 64.640 -1.710 64.840 -0.645 ;
        RECT 65.155 -0.645 65.805 -0.445 ;
        RECT 66.195 -0.445 66.485 -0.355 ;
        RECT 67.515 -0.445 67.805 -0.355 ;
        RECT 66.195 -0.645 66.840 -0.445 ;
        RECT 65.155 -1.710 65.355 -0.645 ;
        RECT 66.640 -1.710 66.840 -0.645 ;
        RECT 67.155 -0.645 67.805 -0.445 ;
        RECT 68.195 -0.445 68.485 -0.355 ;
        RECT 69.515 -0.445 69.805 -0.355 ;
        RECT 68.195 -0.645 68.840 -0.445 ;
        RECT 67.155 -1.710 67.355 -0.645 ;
        RECT 68.640 -1.710 68.840 -0.645 ;
        RECT 69.155 -0.645 69.805 -0.445 ;
        RECT 70.195 -0.445 70.485 -0.355 ;
        RECT 71.515 -0.445 71.805 -0.355 ;
        RECT 70.195 -0.645 70.840 -0.445 ;
        RECT 69.155 -1.710 69.355 -0.645 ;
        RECT 70.640 -1.710 70.840 -0.645 ;
        RECT 71.155 -0.645 71.805 -0.445 ;
        RECT 72.195 -0.445 72.485 -0.355 ;
        RECT 73.515 -0.445 73.805 -0.355 ;
        RECT 72.195 -0.645 72.840 -0.445 ;
        RECT 71.155 -1.710 71.355 -0.645 ;
        RECT 72.640 -1.710 72.840 -0.645 ;
        RECT 73.155 -0.645 73.805 -0.445 ;
        RECT 74.195 -0.445 74.485 -0.355 ;
        RECT 75.515 -0.445 75.805 -0.355 ;
        RECT 74.195 -0.645 74.840 -0.445 ;
        RECT 73.155 -1.710 73.355 -0.645 ;
        RECT 74.640 -1.710 74.840 -0.645 ;
        RECT 75.155 -0.645 75.805 -0.445 ;
        RECT 76.195 -0.445 76.485 -0.355 ;
        RECT 77.515 -0.445 77.805 -0.355 ;
        RECT 76.195 -0.645 76.840 -0.445 ;
        RECT 75.155 -1.710 75.355 -0.645 ;
        RECT 76.640 -1.710 76.840 -0.645 ;
        RECT 77.155 -0.645 77.805 -0.445 ;
        RECT 78.195 -0.445 78.485 -0.355 ;
        RECT 79.515 -0.445 79.805 -0.355 ;
        RECT 78.195 -0.645 78.840 -0.445 ;
        RECT 77.155 -1.710 77.355 -0.645 ;
        RECT 78.640 -1.710 78.840 -0.645 ;
        RECT 79.155 -0.645 79.805 -0.445 ;
        RECT 80.195 -0.445 80.485 -0.355 ;
        RECT 81.515 -0.445 81.805 -0.355 ;
        RECT 80.195 -0.645 80.840 -0.445 ;
        RECT 79.155 -1.710 79.355 -0.645 ;
        RECT 80.640 -1.710 80.840 -0.645 ;
        RECT 81.155 -0.645 81.805 -0.445 ;
        RECT 82.195 -0.445 82.485 -0.355 ;
        RECT 83.515 -0.445 83.805 -0.355 ;
        RECT 82.195 -0.645 82.840 -0.445 ;
        RECT 81.155 -1.710 81.355 -0.645 ;
        RECT 82.640 -1.710 82.840 -0.645 ;
        RECT 83.155 -0.645 83.805 -0.445 ;
        RECT 84.195 -0.445 84.485 -0.355 ;
        RECT 85.515 -0.445 85.805 -0.355 ;
        RECT 84.195 -0.645 84.840 -0.445 ;
        RECT 83.155 -1.710 83.355 -0.645 ;
        RECT 84.640 -1.710 84.840 -0.645 ;
        RECT 85.155 -0.645 85.805 -0.445 ;
        RECT 86.195 -0.445 86.485 -0.355 ;
        RECT 87.515 -0.445 87.805 -0.355 ;
        RECT 86.195 -0.645 86.840 -0.445 ;
        RECT 85.155 -1.710 85.355 -0.645 ;
        RECT 86.640 -1.710 86.840 -0.645 ;
        RECT 87.155 -0.645 87.805 -0.445 ;
        RECT 88.195 -0.445 88.485 -0.355 ;
        RECT 89.515 -0.445 89.805 -0.355 ;
        RECT 88.195 -0.645 88.840 -0.445 ;
        RECT 87.155 -1.710 87.355 -0.645 ;
        RECT 88.640 -1.710 88.840 -0.645 ;
        RECT 89.155 -0.645 89.805 -0.445 ;
        RECT 90.195 -0.445 90.485 -0.355 ;
        RECT 91.515 -0.445 91.805 -0.355 ;
        RECT 90.195 -0.645 90.840 -0.445 ;
        RECT 89.155 -1.710 89.355 -0.645 ;
        RECT 90.640 -1.710 90.840 -0.645 ;
        RECT 91.155 -0.645 91.805 -0.445 ;
        RECT 92.195 -0.445 92.485 -0.355 ;
        RECT 93.515 -0.445 93.805 -0.355 ;
        RECT 92.195 -0.645 92.840 -0.445 ;
        RECT 91.155 -1.710 91.355 -0.645 ;
        RECT 92.640 -1.710 92.840 -0.645 ;
        RECT 93.155 -0.645 93.805 -0.445 ;
        RECT 94.195 -0.445 94.485 -0.355 ;
        RECT 95.515 -0.445 95.805 -0.355 ;
        RECT 94.195 -0.645 94.840 -0.445 ;
        RECT 93.155 -1.710 93.355 -0.645 ;
        RECT 94.640 -1.710 94.840 -0.645 ;
        RECT 95.155 -0.645 95.805 -0.445 ;
        RECT 96.195 -0.445 96.485 -0.355 ;
        RECT 97.515 -0.445 97.805 -0.355 ;
        RECT 96.195 -0.645 96.840 -0.445 ;
        RECT 95.155 -1.710 95.355 -0.645 ;
        RECT 96.640 -1.710 96.840 -0.645 ;
        RECT 97.155 -0.645 97.805 -0.445 ;
        RECT 98.195 -0.445 98.485 -0.355 ;
        RECT 99.515 -0.445 99.805 -0.355 ;
        RECT 98.195 -0.645 98.840 -0.445 ;
        RECT 97.155 -1.710 97.355 -0.645 ;
        RECT 98.640 -1.710 98.840 -0.645 ;
        RECT 99.155 -0.645 99.805 -0.445 ;
        RECT 100.195 -0.445 100.485 -0.355 ;
        RECT 101.515 -0.445 101.805 -0.355 ;
        RECT 100.195 -0.645 100.840 -0.445 ;
        RECT 99.155 -1.710 99.355 -0.645 ;
        RECT 100.640 -1.710 100.840 -0.645 ;
        RECT 101.155 -0.645 101.805 -0.445 ;
        RECT 102.195 -0.445 102.485 -0.355 ;
        RECT 103.515 -0.445 103.805 -0.355 ;
        RECT 102.195 -0.645 102.840 -0.445 ;
        RECT 101.155 -1.710 101.355 -0.645 ;
        RECT 102.640 -1.710 102.840 -0.645 ;
        RECT 103.155 -0.645 103.805 -0.445 ;
        RECT 104.195 -0.445 104.485 -0.355 ;
        RECT 105.515 -0.445 105.805 -0.355 ;
        RECT 104.195 -0.645 104.840 -0.445 ;
        RECT 103.155 -1.710 103.355 -0.645 ;
        RECT 104.640 -1.710 104.840 -0.645 ;
        RECT 105.155 -0.645 105.805 -0.445 ;
        RECT 106.195 -0.445 106.485 -0.355 ;
        RECT 107.515 -0.445 107.805 -0.355 ;
        RECT 106.195 -0.645 106.840 -0.445 ;
        RECT 105.155 -1.710 105.355 -0.645 ;
        RECT 106.640 -1.710 106.840 -0.645 ;
        RECT 107.155 -0.645 107.805 -0.445 ;
        RECT 108.195 -0.445 108.485 -0.355 ;
        RECT 109.515 -0.445 109.805 -0.355 ;
        RECT 108.195 -0.645 108.840 -0.445 ;
        RECT 107.155 -1.710 107.355 -0.645 ;
        RECT 108.640 -1.710 108.840 -0.645 ;
        RECT 109.155 -0.645 109.805 -0.445 ;
        RECT 110.195 -0.445 110.485 -0.355 ;
        RECT 111.515 -0.445 111.805 -0.355 ;
        RECT 110.195 -0.645 110.840 -0.445 ;
        RECT 109.155 -1.710 109.355 -0.645 ;
        RECT 110.640 -1.710 110.840 -0.645 ;
        RECT 111.155 -0.645 111.805 -0.445 ;
        RECT 112.195 -0.445 112.485 -0.355 ;
        RECT 113.515 -0.445 113.805 -0.355 ;
        RECT 112.195 -0.645 112.840 -0.445 ;
        RECT 111.155 -1.710 111.355 -0.645 ;
        RECT 112.640 -1.710 112.840 -0.645 ;
        RECT 113.155 -0.645 113.805 -0.445 ;
        RECT 114.195 -0.445 114.485 -0.355 ;
        RECT 115.515 -0.445 115.805 -0.355 ;
        RECT 114.195 -0.645 114.840 -0.445 ;
        RECT 113.155 -1.710 113.355 -0.645 ;
        RECT 114.640 -1.710 114.840 -0.645 ;
        RECT 115.155 -0.645 115.805 -0.445 ;
        RECT 116.195 -0.445 116.485 -0.355 ;
        RECT 117.515 -0.445 117.805 -0.355 ;
        RECT 116.195 -0.645 116.840 -0.445 ;
        RECT 115.155 -1.710 115.355 -0.645 ;
        RECT 116.640 -1.710 116.840 -0.645 ;
        RECT 117.155 -0.645 117.805 -0.445 ;
        RECT 118.195 -0.445 118.485 -0.355 ;
        RECT 119.515 -0.445 119.805 -0.355 ;
        RECT 118.195 -0.645 118.840 -0.445 ;
        RECT 117.155 -1.710 117.355 -0.645 ;
        RECT 118.640 -1.710 118.840 -0.645 ;
        RECT 119.155 -0.645 119.805 -0.445 ;
        RECT 120.195 -0.445 120.485 -0.355 ;
        RECT 121.515 -0.445 121.805 -0.355 ;
        RECT 120.195 -0.645 120.840 -0.445 ;
        RECT 119.155 -1.710 119.355 -0.645 ;
        RECT 120.640 -1.710 120.840 -0.645 ;
        RECT 121.155 -0.645 121.805 -0.445 ;
        RECT 122.195 -0.445 122.485 -0.355 ;
        RECT 123.515 -0.445 123.805 -0.355 ;
        RECT 122.195 -0.645 122.840 -0.445 ;
        RECT 121.155 -1.710 121.355 -0.645 ;
        RECT 122.640 -1.710 122.840 -0.645 ;
        RECT 123.155 -0.645 123.805 -0.445 ;
        RECT 124.195 -0.445 124.485 -0.355 ;
        RECT 125.515 -0.445 125.805 -0.355 ;
        RECT 124.195 -0.645 124.840 -0.445 ;
        RECT 123.155 -1.710 123.355 -0.645 ;
        RECT 124.640 -1.710 124.840 -0.645 ;
        RECT 125.155 -0.645 125.805 -0.445 ;
        RECT 126.195 -0.445 126.485 -0.355 ;
        RECT 127.515 -0.445 127.805 -0.355 ;
        RECT 126.195 -0.645 126.840 -0.445 ;
        RECT 125.155 -1.710 125.355 -0.645 ;
        RECT 126.640 -1.710 126.840 -0.645 ;
        RECT 127.155 -0.645 127.805 -0.445 ;
        RECT 128.195 -0.445 128.485 -0.355 ;
        RECT 129.515 -0.445 129.805 -0.355 ;
        RECT 128.195 -0.645 128.840 -0.445 ;
        RECT 127.155 -1.710 127.355 -0.645 ;
        RECT 128.640 -1.710 128.840 -0.645 ;
        RECT 129.155 -0.645 129.805 -0.445 ;
        RECT 130.195 -0.445 130.485 -0.355 ;
        RECT 130.195 -0.645 130.840 -0.445 ;
        RECT 129.155 -1.710 129.355 -0.645 ;
        RECT 130.640 -1.710 130.840 -0.645 ;
        RECT -0.890 -2.000 -0.600 -1.710 ;
        RECT 0.600 -2.000 0.890 -1.710 ;
        RECT 1.110 -2.000 1.400 -1.710 ;
        RECT 2.600 -2.000 2.890 -1.710 ;
        RECT 3.110 -2.000 3.400 -1.710 ;
        RECT 4.600 -2.000 4.890 -1.710 ;
        RECT 5.110 -2.000 5.400 -1.710 ;
        RECT 6.600 -2.000 6.890 -1.710 ;
        RECT 7.110 -2.000 7.400 -1.710 ;
        RECT 8.600 -2.000 8.890 -1.710 ;
        RECT 9.110 -2.000 9.400 -1.710 ;
        RECT 10.600 -2.000 10.890 -1.710 ;
        RECT 11.110 -2.000 11.400 -1.710 ;
        RECT 12.600 -2.000 12.890 -1.710 ;
        RECT 13.110 -2.000 13.400 -1.710 ;
        RECT 14.600 -2.000 14.890 -1.710 ;
        RECT 15.110 -2.000 15.400 -1.710 ;
        RECT 16.600 -2.000 16.890 -1.710 ;
        RECT 17.110 -2.000 17.400 -1.710 ;
        RECT 18.600 -2.000 18.890 -1.710 ;
        RECT 19.110 -2.000 19.400 -1.710 ;
        RECT 20.600 -2.000 20.890 -1.710 ;
        RECT 21.110 -2.000 21.400 -1.710 ;
        RECT 22.600 -2.000 22.890 -1.710 ;
        RECT 23.110 -2.000 23.400 -1.710 ;
        RECT 24.600 -2.000 24.890 -1.710 ;
        RECT 25.110 -2.000 25.400 -1.710 ;
        RECT 26.600 -2.000 26.890 -1.710 ;
        RECT 27.110 -2.000 27.400 -1.710 ;
        RECT 28.600 -2.000 28.890 -1.710 ;
        RECT 29.110 -2.000 29.400 -1.710 ;
        RECT 30.600 -2.000 30.890 -1.710 ;
        RECT 31.110 -2.000 31.400 -1.710 ;
        RECT 32.600 -2.000 32.890 -1.710 ;
        RECT 33.110 -2.000 33.400 -1.710 ;
        RECT 34.600 -2.000 34.890 -1.710 ;
        RECT 35.110 -2.000 35.400 -1.710 ;
        RECT 36.600 -2.000 36.890 -1.710 ;
        RECT 37.110 -2.000 37.400 -1.710 ;
        RECT 38.600 -2.000 38.890 -1.710 ;
        RECT 39.110 -2.000 39.400 -1.710 ;
        RECT 40.600 -2.000 40.890 -1.710 ;
        RECT 41.110 -2.000 41.400 -1.710 ;
        RECT 42.600 -2.000 42.890 -1.710 ;
        RECT 43.110 -2.000 43.400 -1.710 ;
        RECT 44.600 -2.000 44.890 -1.710 ;
        RECT 45.110 -2.000 45.400 -1.710 ;
        RECT 46.600 -2.000 46.890 -1.710 ;
        RECT 47.110 -2.000 47.400 -1.710 ;
        RECT 48.600 -2.000 48.890 -1.710 ;
        RECT 49.110 -2.000 49.400 -1.710 ;
        RECT 50.600 -2.000 50.890 -1.710 ;
        RECT 51.110 -2.000 51.400 -1.710 ;
        RECT 52.600 -2.000 52.890 -1.710 ;
        RECT 53.110 -2.000 53.400 -1.710 ;
        RECT 54.600 -2.000 54.890 -1.710 ;
        RECT 55.110 -2.000 55.400 -1.710 ;
        RECT 56.600 -2.000 56.890 -1.710 ;
        RECT 57.110 -2.000 57.400 -1.710 ;
        RECT 58.600 -2.000 58.890 -1.710 ;
        RECT 59.110 -2.000 59.400 -1.710 ;
        RECT 60.600 -2.000 60.890 -1.710 ;
        RECT 61.110 -2.000 61.400 -1.710 ;
        RECT 62.600 -2.000 62.890 -1.710 ;
        RECT 63.110 -2.000 63.400 -1.710 ;
        RECT 64.600 -2.000 64.890 -1.710 ;
        RECT 65.110 -2.000 65.400 -1.710 ;
        RECT 66.600 -2.000 66.890 -1.710 ;
        RECT 67.110 -2.000 67.400 -1.710 ;
        RECT 68.600 -2.000 68.890 -1.710 ;
        RECT 69.110 -2.000 69.400 -1.710 ;
        RECT 70.600 -2.000 70.890 -1.710 ;
        RECT 71.110 -2.000 71.400 -1.710 ;
        RECT 72.600 -2.000 72.890 -1.710 ;
        RECT 73.110 -2.000 73.400 -1.710 ;
        RECT 74.600 -2.000 74.890 -1.710 ;
        RECT 75.110 -2.000 75.400 -1.710 ;
        RECT 76.600 -2.000 76.890 -1.710 ;
        RECT 77.110 -2.000 77.400 -1.710 ;
        RECT 78.600 -2.000 78.890 -1.710 ;
        RECT 79.110 -2.000 79.400 -1.710 ;
        RECT 80.600 -2.000 80.890 -1.710 ;
        RECT 81.110 -2.000 81.400 -1.710 ;
        RECT 82.600 -2.000 82.890 -1.710 ;
        RECT 83.110 -2.000 83.400 -1.710 ;
        RECT 84.600 -2.000 84.890 -1.710 ;
        RECT 85.110 -2.000 85.400 -1.710 ;
        RECT 86.600 -2.000 86.890 -1.710 ;
        RECT 87.110 -2.000 87.400 -1.710 ;
        RECT 88.600 -2.000 88.890 -1.710 ;
        RECT 89.110 -2.000 89.400 -1.710 ;
        RECT 90.600 -2.000 90.890 -1.710 ;
        RECT 91.110 -2.000 91.400 -1.710 ;
        RECT 92.600 -2.000 92.890 -1.710 ;
        RECT 93.110 -2.000 93.400 -1.710 ;
        RECT 94.600 -2.000 94.890 -1.710 ;
        RECT 95.110 -2.000 95.400 -1.710 ;
        RECT 96.600 -2.000 96.890 -1.710 ;
        RECT 97.110 -2.000 97.400 -1.710 ;
        RECT 98.600 -2.000 98.890 -1.710 ;
        RECT 99.110 -2.000 99.400 -1.710 ;
        RECT 100.600 -2.000 100.890 -1.710 ;
        RECT 101.110 -2.000 101.400 -1.710 ;
        RECT 102.600 -2.000 102.890 -1.710 ;
        RECT 103.110 -2.000 103.400 -1.710 ;
        RECT 104.600 -2.000 104.890 -1.710 ;
        RECT 105.110 -2.000 105.400 -1.710 ;
        RECT 106.600 -2.000 106.890 -1.710 ;
        RECT 107.110 -2.000 107.400 -1.710 ;
        RECT 108.600 -2.000 108.890 -1.710 ;
        RECT 109.110 -2.000 109.400 -1.710 ;
        RECT 110.600 -2.000 110.890 -1.710 ;
        RECT 111.110 -2.000 111.400 -1.710 ;
        RECT 112.600 -2.000 112.890 -1.710 ;
        RECT 113.110 -2.000 113.400 -1.710 ;
        RECT 114.600 -2.000 114.890 -1.710 ;
        RECT 115.110 -2.000 115.400 -1.710 ;
        RECT 116.600 -2.000 116.890 -1.710 ;
        RECT 117.110 -2.000 117.400 -1.710 ;
        RECT 118.600 -2.000 118.890 -1.710 ;
        RECT 119.110 -2.000 119.400 -1.710 ;
        RECT 120.600 -2.000 120.890 -1.710 ;
        RECT 121.110 -2.000 121.400 -1.710 ;
        RECT 122.600 -2.000 122.890 -1.710 ;
        RECT 123.110 -2.000 123.400 -1.710 ;
        RECT 124.600 -2.000 124.890 -1.710 ;
        RECT 125.110 -2.000 125.400 -1.710 ;
        RECT 126.600 -2.000 126.890 -1.710 ;
        RECT 127.110 -2.000 127.400 -1.710 ;
        RECT 128.600 -2.000 128.890 -1.710 ;
        RECT 129.110 -2.000 129.400 -1.710 ;
        RECT 130.600 -2.000 130.890 -1.710 ;
        RECT -0.420 -4.620 -0.130 -2.190 ;
        RECT 0.130 -4.620 0.420 -2.190 ;
        RECT 1.580 -4.620 1.870 -2.190 ;
        RECT 2.130 -4.620 2.420 -2.190 ;
        RECT 3.580 -4.620 3.870 -2.190 ;
        RECT 4.130 -4.620 4.420 -2.190 ;
        RECT 5.580 -4.620 5.870 -2.190 ;
        RECT 6.130 -4.620 6.420 -2.190 ;
        RECT 7.580 -4.620 7.870 -2.190 ;
        RECT 8.130 -4.620 8.420 -2.190 ;
        RECT 9.580 -4.620 9.870 -2.190 ;
        RECT 10.130 -4.620 10.420 -2.190 ;
        RECT 11.580 -4.620 11.870 -2.190 ;
        RECT 12.130 -4.620 12.420 -2.190 ;
        RECT 13.580 -4.620 13.870 -2.190 ;
        RECT 14.130 -4.620 14.420 -2.190 ;
        RECT 15.580 -4.620 15.870 -2.190 ;
        RECT 16.130 -4.620 16.420 -2.190 ;
        RECT 17.580 -4.620 17.870 -2.190 ;
        RECT 18.130 -4.620 18.420 -2.190 ;
        RECT 19.580 -4.620 19.870 -2.190 ;
        RECT 20.130 -4.620 20.420 -2.190 ;
        RECT 21.580 -4.620 21.870 -2.190 ;
        RECT 22.130 -4.620 22.420 -2.190 ;
        RECT 23.580 -4.620 23.870 -2.190 ;
        RECT 24.130 -4.620 24.420 -2.190 ;
        RECT 25.580 -4.620 25.870 -2.190 ;
        RECT 26.130 -4.620 26.420 -2.190 ;
        RECT 27.580 -4.620 27.870 -2.190 ;
        RECT 28.130 -4.620 28.420 -2.190 ;
        RECT 29.580 -4.620 29.870 -2.190 ;
        RECT 30.130 -4.620 30.420 -2.190 ;
        RECT 31.580 -4.620 31.870 -2.190 ;
        RECT 32.130 -4.620 32.420 -2.190 ;
        RECT 33.580 -4.620 33.870 -2.190 ;
        RECT 34.130 -4.620 34.420 -2.190 ;
        RECT 35.580 -4.620 35.870 -2.190 ;
        RECT 36.130 -4.620 36.420 -2.190 ;
        RECT 37.580 -4.620 37.870 -2.190 ;
        RECT 38.130 -4.620 38.420 -2.190 ;
        RECT 39.580 -4.620 39.870 -2.190 ;
        RECT 40.130 -4.620 40.420 -2.190 ;
        RECT 41.580 -4.620 41.870 -2.190 ;
        RECT 42.130 -4.620 42.420 -2.190 ;
        RECT 43.580 -4.620 43.870 -2.190 ;
        RECT 44.130 -4.620 44.420 -2.190 ;
        RECT 45.580 -4.620 45.870 -2.190 ;
        RECT 46.130 -4.620 46.420 -2.190 ;
        RECT 47.580 -4.620 47.870 -2.190 ;
        RECT 48.130 -4.620 48.420 -2.190 ;
        RECT 49.580 -4.620 49.870 -2.190 ;
        RECT 50.130 -4.620 50.420 -2.190 ;
        RECT 51.580 -4.620 51.870 -2.190 ;
        RECT 52.130 -4.620 52.420 -2.190 ;
        RECT 53.580 -4.620 53.870 -2.190 ;
        RECT 54.130 -4.620 54.420 -2.190 ;
        RECT 55.580 -4.620 55.870 -2.190 ;
        RECT 56.130 -4.620 56.420 -2.190 ;
        RECT 57.580 -4.620 57.870 -2.190 ;
        RECT 58.130 -4.620 58.420 -2.190 ;
        RECT 59.580 -4.620 59.870 -2.190 ;
        RECT 60.130 -4.620 60.420 -2.190 ;
        RECT 61.580 -4.620 61.870 -2.190 ;
        RECT 62.130 -4.620 62.420 -2.190 ;
        RECT 63.580 -4.620 63.870 -2.190 ;
        RECT 64.130 -4.620 64.420 -2.190 ;
        RECT 65.580 -4.620 65.870 -2.190 ;
        RECT 66.130 -4.620 66.420 -2.190 ;
        RECT 67.580 -4.620 67.870 -2.190 ;
        RECT 68.130 -4.620 68.420 -2.190 ;
        RECT 69.580 -4.620 69.870 -2.190 ;
        RECT 70.130 -4.620 70.420 -2.190 ;
        RECT 71.580 -4.620 71.870 -2.190 ;
        RECT 72.130 -4.620 72.420 -2.190 ;
        RECT 73.580 -4.620 73.870 -2.190 ;
        RECT 74.130 -4.620 74.420 -2.190 ;
        RECT 75.580 -4.620 75.870 -2.190 ;
        RECT 76.130 -4.620 76.420 -2.190 ;
        RECT 77.580 -4.620 77.870 -2.190 ;
        RECT 78.130 -4.620 78.420 -2.190 ;
        RECT 79.580 -4.620 79.870 -2.190 ;
        RECT 80.130 -4.620 80.420 -2.190 ;
        RECT 81.580 -4.620 81.870 -2.190 ;
        RECT 82.130 -4.620 82.420 -2.190 ;
        RECT 83.580 -4.620 83.870 -2.190 ;
        RECT 84.130 -4.620 84.420 -2.190 ;
        RECT 85.580 -4.620 85.870 -2.190 ;
        RECT 86.130 -4.620 86.420 -2.190 ;
        RECT 87.580 -4.620 87.870 -2.190 ;
        RECT 88.130 -4.620 88.420 -2.190 ;
        RECT 89.580 -4.620 89.870 -2.190 ;
        RECT 90.130 -4.620 90.420 -2.190 ;
        RECT 91.580 -4.620 91.870 -2.190 ;
        RECT 92.130 -4.620 92.420 -2.190 ;
        RECT 93.580 -4.620 93.870 -2.190 ;
        RECT 94.130 -4.620 94.420 -2.190 ;
        RECT 95.580 -4.620 95.870 -2.190 ;
        RECT 96.130 -4.620 96.420 -2.190 ;
        RECT 97.580 -4.620 97.870 -2.190 ;
        RECT 98.130 -4.620 98.420 -2.190 ;
        RECT 99.580 -4.620 99.870 -2.190 ;
        RECT 100.130 -4.620 100.420 -2.190 ;
        RECT 101.580 -4.620 101.870 -2.190 ;
        RECT 102.130 -4.620 102.420 -2.190 ;
        RECT 103.580 -4.620 103.870 -2.190 ;
        RECT 104.130 -4.620 104.420 -2.190 ;
        RECT 105.580 -4.620 105.870 -2.190 ;
        RECT 106.130 -4.620 106.420 -2.190 ;
        RECT 107.580 -4.620 107.870 -2.190 ;
        RECT 108.130 -4.620 108.420 -2.190 ;
        RECT 109.580 -4.620 109.870 -2.190 ;
        RECT 110.130 -4.620 110.420 -2.190 ;
        RECT 111.580 -4.620 111.870 -2.190 ;
        RECT 112.130 -4.620 112.420 -2.190 ;
        RECT 113.580 -4.620 113.870 -2.190 ;
        RECT 114.130 -4.620 114.420 -2.190 ;
        RECT 115.580 -4.620 115.870 -2.190 ;
        RECT 116.130 -4.620 116.420 -2.190 ;
        RECT 117.580 -4.620 117.870 -2.190 ;
        RECT 118.130 -4.620 118.420 -2.190 ;
        RECT 119.580 -4.620 119.870 -2.190 ;
        RECT 120.130 -4.620 120.420 -2.190 ;
        RECT 121.580 -4.620 121.870 -2.190 ;
        RECT 122.130 -4.620 122.420 -2.190 ;
        RECT 123.580 -4.620 123.870 -2.190 ;
        RECT 124.130 -4.620 124.420 -2.190 ;
        RECT 125.580 -4.620 125.870 -2.190 ;
        RECT 126.130 -4.620 126.420 -2.190 ;
        RECT 127.580 -4.620 127.870 -2.190 ;
        RECT 128.130 -4.620 128.420 -2.190 ;
        RECT 129.580 -4.620 129.870 -2.190 ;
        RECT 130.130 -4.620 130.420 -2.190 ;
  END
END DAC2U128OUT4IN
END LIBRARY

