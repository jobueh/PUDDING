* Extracted by KLayout with SG13G2 LVS runset on : 31/08/2025 06:12

.SUBCKT DAC2U64OUT2IN
M$1 \$2 \$3 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p PS=2.16u
+ PD=1.14u
M$2 \$1 \$2 \$3 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p PS=1.14u
+ PD=2.16u
M$3 \$4 \$5 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p PS=2.16u
+ PD=1.14u
M$4 \$1 \$4 \$5 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p PS=1.14u
+ PD=2.16u
M$5 \$6 \$7 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p PS=2.16u
+ PD=1.14u
M$6 \$1 \$6 \$7 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p PS=1.14u
+ PD=2.16u
M$7 \$8 \$9 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p PS=2.16u
+ PD=1.14u
M$8 \$1 \$8 \$9 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p PS=1.14u
+ PD=2.16u
M$9 \$10 \$11 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$10 \$1 \$10 \$11 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$11 \$12 \$13 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$12 \$1 \$12 \$13 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$13 \$14 \$15 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$14 \$1 \$14 \$15 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$15 \$16 \$17 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$16 \$1 \$16 \$17 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$17 \$18 \$19 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$18 \$1 \$18 \$19 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$19 \$20 \$21 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$20 \$1 \$20 \$21 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$21 \$22 \$23 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$22 \$1 \$22 \$23 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$23 \$24 \$25 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$24 \$1 \$24 \$25 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$25 \$26 \$27 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$26 \$1 \$26 \$27 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$27 \$28 \$29 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$28 \$1 \$28 \$29 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$29 \$30 \$31 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$30 \$1 \$30 \$31 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$31 \$32 \$33 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$32 \$1 \$32 \$33 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$33 \$34 \$35 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$34 \$1 \$34 \$35 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$35 \$36 \$37 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$36 \$1 \$36 \$37 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$37 \$38 \$39 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$38 \$1 \$38 \$39 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$39 \$40 \$41 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$40 \$1 \$40 \$41 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$41 \$42 \$43 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$42 \$1 \$42 \$43 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$43 \$44 \$45 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$44 \$1 \$44 \$45 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$45 \$46 \$47 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$46 \$1 \$46 \$47 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$47 \$48 \$49 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$48 \$1 \$48 \$49 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$49 \$50 \$51 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$50 \$1 \$50 \$51 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$51 \$52 \$53 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$52 \$1 \$52 \$53 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$53 \$54 \$55 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$54 \$1 \$54 \$55 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$55 \$56 \$57 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$56 \$1 \$56 \$57 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$57 \$58 \$59 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$58 \$1 \$58 \$59 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$59 \$60 \$61 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$60 \$1 \$60 \$61 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$61 \$62 \$63 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$62 \$1 \$62 \$63 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$63 \$64 \$65 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$64 \$1 \$64 \$65 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$65 \$66 \$67 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$66 \$1 \$66 \$67 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$67 \$68 \$69 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$68 \$1 \$68 \$69 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$69 \$70 \$71 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$70 \$1 \$70 \$71 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$71 \$72 \$73 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$72 \$1 \$72 \$73 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$73 \$74 \$75 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$74 \$1 \$74 \$75 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$75 \$76 \$77 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$76 \$1 \$76 \$77 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$77 \$78 \$79 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$78 \$1 \$78 \$79 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$79 \$80 \$81 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$80 \$1 \$80 \$81 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$81 \$82 \$83 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$82 \$1 \$82 \$83 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$83 \$84 \$85 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$84 \$1 \$84 \$85 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$85 \$86 \$87 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$86 \$1 \$86 \$87 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$87 \$88 \$89 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$88 \$1 \$88 \$89 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$89 \$90 \$91 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$90 \$1 \$90 \$91 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$91 \$92 \$93 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$92 \$1 \$92 \$93 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$93 \$94 \$95 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$94 \$1 \$94 \$95 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$95 \$96 \$97 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$96 \$1 \$96 \$97 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$97 \$98 \$99 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$98 \$1 \$98 \$99 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$99 \$100 \$101 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$100 \$1 \$100 \$101 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$101 \$102 \$103 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$102 \$1 \$102 \$103 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$103 \$104 \$105 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$104 \$1 \$104 \$105 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$105 \$106 \$107 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$106 \$1 \$106 \$107 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$107 \$108 \$109 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$108 \$1 \$108 \$109 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$109 \$110 \$111 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$110 \$1 \$110 \$111 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$111 \$112 \$113 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$112 \$1 \$112 \$113 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$113 \$114 \$115 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$114 \$1 \$114 \$115 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$115 \$116 \$117 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$116 \$1 \$116 \$117 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$117 \$118 \$119 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$118 \$1 \$118 \$119 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$119 \$120 \$121 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$120 \$1 \$120 \$121 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$121 \$122 \$123 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$122 \$1 \$122 \$123 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$123 \$124 \$125 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$124 \$1 \$124 \$125 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$125 \$126 \$127 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$126 \$1 \$126 \$127 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$127 \$128 \$129 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$128 \$1 \$128 \$129 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$129 \$130 \$131 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$130 \$1 \$130 \$131 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$131 \$132 \$133 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$132 \$1 \$132 \$133 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$133 \$2 \$134 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$134 \$266 \$135 \$3 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$135 \$4 \$136 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$136 \$266 \$137 \$5 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$137 \$6 \$138 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$138 \$266 \$139 \$7 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$139 \$8 \$140 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$140 \$266 \$141 \$9 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$141 \$10 \$142 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$142 \$266 \$143 \$11 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$143 \$12 \$144 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$144 \$266 \$145 \$13 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$145 \$14 \$146 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$146 \$266 \$147 \$15 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$147 \$16 \$148 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$148 \$266 \$149 \$17 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$149 \$18 \$150 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$150 \$266 \$151 \$19 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$151 \$20 \$152 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$152 \$266 \$153 \$21 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$153 \$22 \$154 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$154 \$266 \$155 \$23 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$155 \$24 \$156 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$156 \$266 \$157 \$25 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$157 \$26 \$158 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$158 \$266 \$159 \$27 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$159 \$28 \$160 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$160 \$266 \$161 \$29 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$161 \$30 \$162 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$162 \$266 \$163 \$31 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$163 \$32 \$164 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$164 \$266 \$165 \$33 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$165 \$34 \$166 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$166 \$266 \$167 \$35 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$167 \$36 \$168 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$168 \$266 \$169 \$37 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$169 \$38 \$170 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$170 \$266 \$171 \$39 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$171 \$40 \$172 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$172 \$266 \$173 \$41 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$173 \$42 \$174 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$174 \$266 \$175 \$43 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$175 \$44 \$176 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$176 \$266 \$177 \$45 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$177 \$46 \$178 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$178 \$266 \$179 \$47 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$179 \$48 \$180 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$180 \$266 \$181 \$49 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$181 \$50 \$182 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$182 \$266 \$183 \$51 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$183 \$52 \$184 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$184 \$266 \$185 \$53 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$185 \$54 \$186 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$186 \$266 \$187 \$55 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$187 \$56 \$188 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$188 \$266 \$189 \$57 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$189 \$58 \$190 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$190 \$266 \$191 \$59 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$191 \$60 \$192 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$192 \$266 \$193 \$61 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$193 \$62 \$194 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$194 \$266 \$195 \$63 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$195 \$64 \$196 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$196 \$266 \$197 \$65 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$197 \$66 \$198 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$198 \$266 \$199 \$67 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$199 \$68 \$200 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$200 \$266 \$201 \$69 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$201 \$70 \$202 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$202 \$266 \$203 \$71 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$203 \$72 \$204 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$204 \$266 \$205 \$73 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$205 \$74 \$206 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$206 \$266 \$207 \$75 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$207 \$76 \$208 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$208 \$266 \$209 \$77 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$209 \$78 \$210 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$210 \$266 \$211 \$79 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$211 \$80 \$212 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$212 \$266 \$213 \$81 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$213 \$82 \$214 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$214 \$266 \$215 \$83 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$215 \$84 \$216 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$216 \$266 \$217 \$85 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$217 \$86 \$218 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$218 \$266 \$219 \$87 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$219 \$88 \$220 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$220 \$266 \$221 \$89 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$221 \$90 \$222 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$222 \$266 \$223 \$91 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$223 \$92 \$224 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$224 \$266 \$225 \$93 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$225 \$94 \$226 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$226 \$266 \$227 \$95 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$227 \$96 \$228 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$228 \$266 \$229 \$97 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$229 \$98 \$230 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$230 \$266 \$231 \$99 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$231 \$100 \$232 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$232 \$266 \$233 \$101 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$233 \$102 \$234 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$234 \$266 \$235 \$103 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$235 \$104 \$236 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$236 \$266 \$237 \$105 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$237 \$106 \$238 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$238 \$266 \$239 \$107 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$239 \$108 \$240 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$240 \$266 \$241 \$109 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$241 \$110 \$242 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$242 \$266 \$243 \$111 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$243 \$112 \$244 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$244 \$266 \$245 \$113 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$245 \$114 \$246 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$246 \$266 \$247 \$115 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$247 \$116 \$248 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$248 \$266 \$249 \$117 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$249 \$118 \$250 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$250 \$266 \$251 \$119 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$251 \$120 \$252 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$252 \$266 \$253 \$121 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$253 \$122 \$254 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$254 \$266 \$255 \$123 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$255 \$124 \$256 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$256 \$266 \$257 \$125 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$257 \$126 \$258 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$258 \$266 \$259 \$127 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$259 \$128 \$260 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$260 \$266 \$261 \$129 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$261 \$130 \$262 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$262 \$266 \$263 \$131 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$263 \$132 \$264 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$264 \$266 \$265 \$133 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$265 \$267 \$2 \$268 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$266 \$268 \$3 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$267 \$267 \$4 \$269 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$268 \$269 \$5 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$269 \$267 \$6 \$270 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$270 \$270 \$7 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$271 \$267 \$8 \$271 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$272 \$271 \$9 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$273 \$267 \$10 \$272 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$274 \$272 \$11 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$275 \$267 \$12 \$273 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$276 \$273 \$13 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$277 \$267 \$14 \$274 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$278 \$274 \$15 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$279 \$267 \$16 \$275 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$280 \$275 \$17 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$281 \$267 \$18 \$276 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$282 \$276 \$19 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$283 \$267 \$20 \$277 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$284 \$277 \$21 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$285 \$267 \$22 \$278 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$286 \$278 \$23 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$287 \$267 \$24 \$279 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$288 \$279 \$25 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$289 \$267 \$26 \$280 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$290 \$280 \$27 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$291 \$267 \$28 \$281 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$292 \$281 \$29 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$293 \$267 \$30 \$282 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$294 \$282 \$31 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$295 \$267 \$32 \$283 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$296 \$283 \$33 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$297 \$267 \$34 \$284 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$298 \$284 \$35 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$299 \$267 \$36 \$285 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$300 \$285 \$37 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$301 \$267 \$38 \$286 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$302 \$286 \$39 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$303 \$267 \$40 \$287 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$304 \$287 \$41 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$305 \$267 \$42 \$288 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$306 \$288 \$43 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$307 \$267 \$44 \$289 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$308 \$289 \$45 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$309 \$267 \$46 \$290 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$310 \$290 \$47 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$311 \$267 \$48 \$291 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$312 \$291 \$49 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$313 \$267 \$50 \$292 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$314 \$292 \$51 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$315 \$267 \$52 \$293 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$316 \$293 \$53 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$317 \$267 \$54 \$294 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$318 \$294 \$55 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$319 \$267 \$56 \$295 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$320 \$295 \$57 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$321 \$267 \$58 \$296 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$322 \$296 \$59 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$323 \$267 \$60 \$297 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$324 \$297 \$61 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$325 \$267 \$62 \$298 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$326 \$298 \$63 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$327 \$267 \$64 \$299 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$328 \$299 \$65 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$329 \$267 \$66 \$300 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$330 \$300 \$67 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$331 \$267 \$68 \$301 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$332 \$301 \$69 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$333 \$267 \$70 \$302 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$334 \$302 \$71 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$335 \$267 \$72 \$303 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$336 \$303 \$73 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$337 \$267 \$74 \$304 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$338 \$304 \$75 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$339 \$267 \$76 \$305 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$340 \$305 \$77 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$341 \$267 \$78 \$306 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$342 \$306 \$79 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$343 \$267 \$80 \$307 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$344 \$307 \$81 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$345 \$267 \$82 \$308 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$346 \$308 \$83 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$347 \$267 \$84 \$309 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$348 \$309 \$85 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$349 \$267 \$86 \$310 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$350 \$310 \$87 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$351 \$267 \$88 \$311 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$352 \$311 \$89 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$353 \$267 \$90 \$312 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$354 \$312 \$91 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$355 \$267 \$92 \$313 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$356 \$313 \$93 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$357 \$267 \$94 \$314 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$358 \$314 \$95 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$359 \$267 \$96 \$315 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$360 \$315 \$97 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$361 \$267 \$98 \$316 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$362 \$316 \$99 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$363 \$267 \$100 \$317 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$364 \$317 \$101 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$365 \$267 \$102 \$318 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$366 \$318 \$103 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$367 \$267 \$104 \$319 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$368 \$319 \$105 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$369 \$267 \$106 \$320 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$370 \$320 \$107 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$371 \$267 \$108 \$321 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$372 \$321 \$109 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$373 \$267 \$110 \$322 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$374 \$322 \$111 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$375 \$267 \$112 \$323 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$376 \$323 \$113 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$377 \$267 \$114 \$324 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$378 \$324 \$115 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$379 \$267 \$116 \$325 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$380 \$325 \$117 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$381 \$267 \$118 \$326 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$382 \$326 \$119 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$383 \$267 \$120 \$327 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$384 \$327 \$121 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$385 \$267 \$122 \$328 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$386 \$328 \$123 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$387 \$267 \$124 \$329 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$388 \$329 \$125 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$389 \$267 \$126 \$330 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$390 \$330 \$127 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$391 \$267 \$128 \$331 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$392 \$331 \$129 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$393 \$267 \$130 \$332 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$394 \$332 \$131 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$395 \$267 \$132 \$333 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$396 \$333 \$133 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$397 \$267 \$267 \$334 \$266 sg13_lv_pmos L=0.15u W=11.7u AS=3.978p AD=3.978p
+ PS=24.76u PD=24.76u
M$398 \$266 \$334 \$346 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$399 \$346 \$268 \$334 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$400 \$266 \$334 \$339 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$401 \$339 \$269 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$402 \$266 \$334 \$349 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$403 \$349 \$270 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$404 \$266 \$334 \$354 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$405 \$354 \$271 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$406 \$266 \$334 \$359 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$407 \$359 \$272 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$408 \$266 \$334 \$364 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$409 \$364 \$273 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$410 \$266 \$334 \$369 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$411 \$369 \$274 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$412 \$266 \$334 \$374 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$413 \$374 \$275 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$414 \$266 \$334 \$379 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$415 \$379 \$276 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$416 \$266 \$334 \$384 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$417 \$384 \$277 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$418 \$266 \$334 \$389 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$419 \$389 \$278 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$420 \$266 \$334 \$394 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$421 \$394 \$279 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$422 \$266 \$334 \$399 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$423 \$399 \$280 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$424 \$266 \$334 \$400 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$425 \$400 \$281 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$426 \$266 \$334 \$398 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$427 \$398 \$282 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$428 \$266 \$334 \$397 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$429 \$397 \$283 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$430 \$266 \$334 \$396 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$431 \$396 \$284 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$432 \$266 \$334 \$395 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$433 \$395 \$285 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$434 \$266 \$334 \$393 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$435 \$393 \$286 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$436 \$266 \$334 \$392 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$437 \$392 \$287 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$438 \$266 \$334 \$391 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$439 \$391 \$288 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$440 \$266 \$334 \$390 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$441 \$390 \$289 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$442 \$266 \$334 \$388 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$443 \$388 \$290 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$444 \$266 \$334 \$387 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$445 \$387 \$291 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$446 \$266 \$334 \$386 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$447 \$386 \$292 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$448 \$266 \$334 \$385 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$449 \$385 \$293 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$450 \$266 \$334 \$383 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$451 \$383 \$294 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$452 \$266 \$334 \$382 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$453 \$382 \$295 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$454 \$266 \$334 \$381 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$455 \$381 \$296 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$456 \$266 \$334 \$380 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$457 \$380 \$297 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$458 \$266 \$334 \$378 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$459 \$378 \$298 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$460 \$266 \$334 \$377 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$461 \$377 \$299 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$462 \$266 \$334 \$376 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$463 \$376 \$300 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$464 \$266 \$334 \$375 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$465 \$375 \$301 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$466 \$266 \$334 \$373 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$467 \$373 \$302 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$468 \$266 \$334 \$372 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$469 \$372 \$303 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$470 \$266 \$334 \$371 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$471 \$371 \$304 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$472 \$266 \$334 \$370 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$473 \$370 \$305 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$474 \$266 \$334 \$368 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$475 \$368 \$306 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$476 \$266 \$334 \$367 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$477 \$367 \$307 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$478 \$266 \$334 \$366 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$479 \$366 \$308 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$480 \$266 \$334 \$365 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$481 \$365 \$309 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$482 \$266 \$334 \$363 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$483 \$363 \$310 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$484 \$266 \$334 \$362 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$485 \$362 \$311 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$486 \$266 \$334 \$361 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$487 \$361 \$312 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$488 \$266 \$334 \$360 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$489 \$360 \$313 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$490 \$266 \$334 \$358 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$491 \$358 \$314 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$492 \$266 \$334 \$357 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$493 \$357 \$315 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$494 \$266 \$334 \$356 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$495 \$356 \$316 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$496 \$266 \$334 \$355 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$497 \$355 \$317 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$498 \$266 \$334 \$353 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$499 \$353 \$318 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$500 \$266 \$334 \$352 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$501 \$352 \$319 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$502 \$266 \$334 \$351 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$503 \$351 \$320 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$504 \$266 \$334 \$350 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$505 \$350 \$321 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$506 \$266 \$334 \$348 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$507 \$348 \$322 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$508 \$266 \$334 \$347 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$509 \$347 \$323 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$510 \$266 \$334 \$345 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$511 \$345 \$324 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$512 \$266 \$334 \$344 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$513 \$344 \$325 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$514 \$266 \$334 \$343 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$515 \$343 \$326 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$516 \$266 \$334 \$342 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$517 \$342 \$327 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$518 \$266 \$334 \$341 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$519 \$341 \$328 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$520 \$266 \$334 \$340 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$521 \$340 \$329 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$522 \$266 \$334 \$338 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$523 \$338 \$330 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$524 \$266 \$334 \$337 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$525 \$337 \$331 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$526 \$266 \$334 \$336 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$527 \$336 \$332 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$528 \$266 \$334 \$335 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$529 \$335 \$333 \$334 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
.ENDS DAC2U64OUT2IN
