magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757286748
<< metal1 >>
rect 576 38576 99360 38600
rect 576 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 8352 38576
rect 8392 38536 8434 38576
rect 8474 38536 8516 38576
rect 8556 38536 8598 38576
rect 8638 38536 8680 38576
rect 8720 38536 12352 38576
rect 12392 38536 12434 38576
rect 12474 38536 12516 38576
rect 12556 38536 12598 38576
rect 12638 38536 12680 38576
rect 12720 38536 16352 38576
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16720 38536 20352 38576
rect 20392 38536 20434 38576
rect 20474 38536 20516 38576
rect 20556 38536 20598 38576
rect 20638 38536 20680 38576
rect 20720 38536 24352 38576
rect 24392 38536 24434 38576
rect 24474 38536 24516 38576
rect 24556 38536 24598 38576
rect 24638 38536 24680 38576
rect 24720 38536 28352 38576
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28720 38536 32352 38576
rect 32392 38536 32434 38576
rect 32474 38536 32516 38576
rect 32556 38536 32598 38576
rect 32638 38536 32680 38576
rect 32720 38536 36352 38576
rect 36392 38536 36434 38576
rect 36474 38536 36516 38576
rect 36556 38536 36598 38576
rect 36638 38536 36680 38576
rect 36720 38536 40352 38576
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40720 38536 44352 38576
rect 44392 38536 44434 38576
rect 44474 38536 44516 38576
rect 44556 38536 44598 38576
rect 44638 38536 44680 38576
rect 44720 38536 48352 38576
rect 48392 38536 48434 38576
rect 48474 38536 48516 38576
rect 48556 38536 48598 38576
rect 48638 38536 48680 38576
rect 48720 38536 52352 38576
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52720 38536 56352 38576
rect 56392 38536 56434 38576
rect 56474 38536 56516 38576
rect 56556 38536 56598 38576
rect 56638 38536 56680 38576
rect 56720 38536 60352 38576
rect 60392 38536 60434 38576
rect 60474 38536 60516 38576
rect 60556 38536 60598 38576
rect 60638 38536 60680 38576
rect 60720 38536 64352 38576
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64720 38536 68352 38576
rect 68392 38536 68434 38576
rect 68474 38536 68516 38576
rect 68556 38536 68598 38576
rect 68638 38536 68680 38576
rect 68720 38536 72352 38576
rect 72392 38536 72434 38576
rect 72474 38536 72516 38576
rect 72556 38536 72598 38576
rect 72638 38536 72680 38576
rect 72720 38536 76352 38576
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76720 38536 80352 38576
rect 80392 38536 80434 38576
rect 80474 38536 80516 38576
rect 80556 38536 80598 38576
rect 80638 38536 80680 38576
rect 80720 38536 84352 38576
rect 84392 38536 84434 38576
rect 84474 38536 84516 38576
rect 84556 38536 84598 38576
rect 84638 38536 84680 38576
rect 84720 38536 88352 38576
rect 88392 38536 88434 38576
rect 88474 38536 88516 38576
rect 88556 38536 88598 38576
rect 88638 38536 88680 38576
rect 88720 38536 92352 38576
rect 92392 38536 92434 38576
rect 92474 38536 92516 38576
rect 92556 38536 92598 38576
rect 92638 38536 92680 38576
rect 92720 38536 96352 38576
rect 96392 38536 96434 38576
rect 96474 38536 96516 38576
rect 96556 38536 96598 38576
rect 96638 38536 96680 38576
rect 96720 38536 99360 38576
rect 576 38512 99360 38536
rect 576 37820 99516 37844
rect 576 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 7112 37820
rect 7152 37780 7194 37820
rect 7234 37780 7276 37820
rect 7316 37780 7358 37820
rect 7398 37780 7440 37820
rect 7480 37780 11112 37820
rect 11152 37780 11194 37820
rect 11234 37780 11276 37820
rect 11316 37780 11358 37820
rect 11398 37780 11440 37820
rect 11480 37780 15112 37820
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15480 37780 19112 37820
rect 19152 37780 19194 37820
rect 19234 37780 19276 37820
rect 19316 37780 19358 37820
rect 19398 37780 19440 37820
rect 19480 37780 23112 37820
rect 23152 37780 23194 37820
rect 23234 37780 23276 37820
rect 23316 37780 23358 37820
rect 23398 37780 23440 37820
rect 23480 37780 27112 37820
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27480 37780 31112 37820
rect 31152 37780 31194 37820
rect 31234 37780 31276 37820
rect 31316 37780 31358 37820
rect 31398 37780 31440 37820
rect 31480 37780 35112 37820
rect 35152 37780 35194 37820
rect 35234 37780 35276 37820
rect 35316 37780 35358 37820
rect 35398 37780 35440 37820
rect 35480 37780 39112 37820
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39480 37780 43112 37820
rect 43152 37780 43194 37820
rect 43234 37780 43276 37820
rect 43316 37780 43358 37820
rect 43398 37780 43440 37820
rect 43480 37780 47112 37820
rect 47152 37780 47194 37820
rect 47234 37780 47276 37820
rect 47316 37780 47358 37820
rect 47398 37780 47440 37820
rect 47480 37780 51112 37820
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51480 37780 55112 37820
rect 55152 37780 55194 37820
rect 55234 37780 55276 37820
rect 55316 37780 55358 37820
rect 55398 37780 55440 37820
rect 55480 37780 59112 37820
rect 59152 37780 59194 37820
rect 59234 37780 59276 37820
rect 59316 37780 59358 37820
rect 59398 37780 59440 37820
rect 59480 37780 63112 37820
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63480 37780 67112 37820
rect 67152 37780 67194 37820
rect 67234 37780 67276 37820
rect 67316 37780 67358 37820
rect 67398 37780 67440 37820
rect 67480 37780 71112 37820
rect 71152 37780 71194 37820
rect 71234 37780 71276 37820
rect 71316 37780 71358 37820
rect 71398 37780 71440 37820
rect 71480 37780 75112 37820
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75480 37780 79112 37820
rect 79152 37780 79194 37820
rect 79234 37780 79276 37820
rect 79316 37780 79358 37820
rect 79398 37780 79440 37820
rect 79480 37780 83112 37820
rect 83152 37780 83194 37820
rect 83234 37780 83276 37820
rect 83316 37780 83358 37820
rect 83398 37780 83440 37820
rect 83480 37780 87112 37820
rect 87152 37780 87194 37820
rect 87234 37780 87276 37820
rect 87316 37780 87358 37820
rect 87398 37780 87440 37820
rect 87480 37780 91112 37820
rect 91152 37780 91194 37820
rect 91234 37780 91276 37820
rect 91316 37780 91358 37820
rect 91398 37780 91440 37820
rect 91480 37780 95112 37820
rect 95152 37780 95194 37820
rect 95234 37780 95276 37820
rect 95316 37780 95358 37820
rect 95398 37780 95440 37820
rect 95480 37780 99112 37820
rect 99152 37780 99194 37820
rect 99234 37780 99276 37820
rect 99316 37780 99358 37820
rect 99398 37780 99440 37820
rect 99480 37780 99516 37820
rect 576 37756 99516 37780
rect 576 37064 99360 37088
rect 576 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 8352 37064
rect 8392 37024 8434 37064
rect 8474 37024 8516 37064
rect 8556 37024 8598 37064
rect 8638 37024 8680 37064
rect 8720 37024 12352 37064
rect 12392 37024 12434 37064
rect 12474 37024 12516 37064
rect 12556 37024 12598 37064
rect 12638 37024 12680 37064
rect 12720 37024 16352 37064
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16720 37024 20352 37064
rect 20392 37024 20434 37064
rect 20474 37024 20516 37064
rect 20556 37024 20598 37064
rect 20638 37024 20680 37064
rect 20720 37024 24352 37064
rect 24392 37024 24434 37064
rect 24474 37024 24516 37064
rect 24556 37024 24598 37064
rect 24638 37024 24680 37064
rect 24720 37024 28352 37064
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28720 37024 32352 37064
rect 32392 37024 32434 37064
rect 32474 37024 32516 37064
rect 32556 37024 32598 37064
rect 32638 37024 32680 37064
rect 32720 37024 36352 37064
rect 36392 37024 36434 37064
rect 36474 37024 36516 37064
rect 36556 37024 36598 37064
rect 36638 37024 36680 37064
rect 36720 37024 40352 37064
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40720 37024 44352 37064
rect 44392 37024 44434 37064
rect 44474 37024 44516 37064
rect 44556 37024 44598 37064
rect 44638 37024 44680 37064
rect 44720 37024 48352 37064
rect 48392 37024 48434 37064
rect 48474 37024 48516 37064
rect 48556 37024 48598 37064
rect 48638 37024 48680 37064
rect 48720 37024 52352 37064
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52720 37024 56352 37064
rect 56392 37024 56434 37064
rect 56474 37024 56516 37064
rect 56556 37024 56598 37064
rect 56638 37024 56680 37064
rect 56720 37024 60352 37064
rect 60392 37024 60434 37064
rect 60474 37024 60516 37064
rect 60556 37024 60598 37064
rect 60638 37024 60680 37064
rect 60720 37024 64352 37064
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64720 37024 68352 37064
rect 68392 37024 68434 37064
rect 68474 37024 68516 37064
rect 68556 37024 68598 37064
rect 68638 37024 68680 37064
rect 68720 37024 72352 37064
rect 72392 37024 72434 37064
rect 72474 37024 72516 37064
rect 72556 37024 72598 37064
rect 72638 37024 72680 37064
rect 72720 37024 76352 37064
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76720 37024 80352 37064
rect 80392 37024 80434 37064
rect 80474 37024 80516 37064
rect 80556 37024 80598 37064
rect 80638 37024 80680 37064
rect 80720 37024 84352 37064
rect 84392 37024 84434 37064
rect 84474 37024 84516 37064
rect 84556 37024 84598 37064
rect 84638 37024 84680 37064
rect 84720 37024 88352 37064
rect 88392 37024 88434 37064
rect 88474 37024 88516 37064
rect 88556 37024 88598 37064
rect 88638 37024 88680 37064
rect 88720 37024 92352 37064
rect 92392 37024 92434 37064
rect 92474 37024 92516 37064
rect 92556 37024 92598 37064
rect 92638 37024 92680 37064
rect 92720 37024 96352 37064
rect 96392 37024 96434 37064
rect 96474 37024 96516 37064
rect 96556 37024 96598 37064
rect 96638 37024 96680 37064
rect 96720 37024 99360 37064
rect 576 37000 99360 37024
rect 576 36308 99516 36332
rect 576 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 7112 36308
rect 7152 36268 7194 36308
rect 7234 36268 7276 36308
rect 7316 36268 7358 36308
rect 7398 36268 7440 36308
rect 7480 36268 11112 36308
rect 11152 36268 11194 36308
rect 11234 36268 11276 36308
rect 11316 36268 11358 36308
rect 11398 36268 11440 36308
rect 11480 36268 15112 36308
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15480 36268 19112 36308
rect 19152 36268 19194 36308
rect 19234 36268 19276 36308
rect 19316 36268 19358 36308
rect 19398 36268 19440 36308
rect 19480 36268 23112 36308
rect 23152 36268 23194 36308
rect 23234 36268 23276 36308
rect 23316 36268 23358 36308
rect 23398 36268 23440 36308
rect 23480 36268 27112 36308
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27480 36268 31112 36308
rect 31152 36268 31194 36308
rect 31234 36268 31276 36308
rect 31316 36268 31358 36308
rect 31398 36268 31440 36308
rect 31480 36268 35112 36308
rect 35152 36268 35194 36308
rect 35234 36268 35276 36308
rect 35316 36268 35358 36308
rect 35398 36268 35440 36308
rect 35480 36268 39112 36308
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39480 36268 43112 36308
rect 43152 36268 43194 36308
rect 43234 36268 43276 36308
rect 43316 36268 43358 36308
rect 43398 36268 43440 36308
rect 43480 36268 47112 36308
rect 47152 36268 47194 36308
rect 47234 36268 47276 36308
rect 47316 36268 47358 36308
rect 47398 36268 47440 36308
rect 47480 36268 51112 36308
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51480 36268 55112 36308
rect 55152 36268 55194 36308
rect 55234 36268 55276 36308
rect 55316 36268 55358 36308
rect 55398 36268 55440 36308
rect 55480 36268 59112 36308
rect 59152 36268 59194 36308
rect 59234 36268 59276 36308
rect 59316 36268 59358 36308
rect 59398 36268 59440 36308
rect 59480 36268 63112 36308
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63480 36268 67112 36308
rect 67152 36268 67194 36308
rect 67234 36268 67276 36308
rect 67316 36268 67358 36308
rect 67398 36268 67440 36308
rect 67480 36268 71112 36308
rect 71152 36268 71194 36308
rect 71234 36268 71276 36308
rect 71316 36268 71358 36308
rect 71398 36268 71440 36308
rect 71480 36268 75112 36308
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75480 36268 79112 36308
rect 79152 36268 79194 36308
rect 79234 36268 79276 36308
rect 79316 36268 79358 36308
rect 79398 36268 79440 36308
rect 79480 36268 83112 36308
rect 83152 36268 83194 36308
rect 83234 36268 83276 36308
rect 83316 36268 83358 36308
rect 83398 36268 83440 36308
rect 83480 36268 87112 36308
rect 87152 36268 87194 36308
rect 87234 36268 87276 36308
rect 87316 36268 87358 36308
rect 87398 36268 87440 36308
rect 87480 36268 91112 36308
rect 91152 36268 91194 36308
rect 91234 36268 91276 36308
rect 91316 36268 91358 36308
rect 91398 36268 91440 36308
rect 91480 36268 95112 36308
rect 95152 36268 95194 36308
rect 95234 36268 95276 36308
rect 95316 36268 95358 36308
rect 95398 36268 95440 36308
rect 95480 36268 99112 36308
rect 99152 36268 99194 36308
rect 99234 36268 99276 36308
rect 99316 36268 99358 36308
rect 99398 36268 99440 36308
rect 99480 36268 99516 36308
rect 576 36244 99516 36268
rect 576 35552 99360 35576
rect 576 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 8352 35552
rect 8392 35512 8434 35552
rect 8474 35512 8516 35552
rect 8556 35512 8598 35552
rect 8638 35512 8680 35552
rect 8720 35512 12352 35552
rect 12392 35512 12434 35552
rect 12474 35512 12516 35552
rect 12556 35512 12598 35552
rect 12638 35512 12680 35552
rect 12720 35512 16352 35552
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16720 35512 20352 35552
rect 20392 35512 20434 35552
rect 20474 35512 20516 35552
rect 20556 35512 20598 35552
rect 20638 35512 20680 35552
rect 20720 35512 24352 35552
rect 24392 35512 24434 35552
rect 24474 35512 24516 35552
rect 24556 35512 24598 35552
rect 24638 35512 24680 35552
rect 24720 35512 28352 35552
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28720 35512 32352 35552
rect 32392 35512 32434 35552
rect 32474 35512 32516 35552
rect 32556 35512 32598 35552
rect 32638 35512 32680 35552
rect 32720 35512 36352 35552
rect 36392 35512 36434 35552
rect 36474 35512 36516 35552
rect 36556 35512 36598 35552
rect 36638 35512 36680 35552
rect 36720 35512 40352 35552
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40720 35512 44352 35552
rect 44392 35512 44434 35552
rect 44474 35512 44516 35552
rect 44556 35512 44598 35552
rect 44638 35512 44680 35552
rect 44720 35512 48352 35552
rect 48392 35512 48434 35552
rect 48474 35512 48516 35552
rect 48556 35512 48598 35552
rect 48638 35512 48680 35552
rect 48720 35512 52352 35552
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52720 35512 56352 35552
rect 56392 35512 56434 35552
rect 56474 35512 56516 35552
rect 56556 35512 56598 35552
rect 56638 35512 56680 35552
rect 56720 35512 60352 35552
rect 60392 35512 60434 35552
rect 60474 35512 60516 35552
rect 60556 35512 60598 35552
rect 60638 35512 60680 35552
rect 60720 35512 64352 35552
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64720 35512 68352 35552
rect 68392 35512 68434 35552
rect 68474 35512 68516 35552
rect 68556 35512 68598 35552
rect 68638 35512 68680 35552
rect 68720 35512 72352 35552
rect 72392 35512 72434 35552
rect 72474 35512 72516 35552
rect 72556 35512 72598 35552
rect 72638 35512 72680 35552
rect 72720 35512 76352 35552
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76720 35512 80352 35552
rect 80392 35512 80434 35552
rect 80474 35512 80516 35552
rect 80556 35512 80598 35552
rect 80638 35512 80680 35552
rect 80720 35512 84352 35552
rect 84392 35512 84434 35552
rect 84474 35512 84516 35552
rect 84556 35512 84598 35552
rect 84638 35512 84680 35552
rect 84720 35512 88352 35552
rect 88392 35512 88434 35552
rect 88474 35512 88516 35552
rect 88556 35512 88598 35552
rect 88638 35512 88680 35552
rect 88720 35512 92352 35552
rect 92392 35512 92434 35552
rect 92474 35512 92516 35552
rect 92556 35512 92598 35552
rect 92638 35512 92680 35552
rect 92720 35512 96352 35552
rect 96392 35512 96434 35552
rect 96474 35512 96516 35552
rect 96556 35512 96598 35552
rect 96638 35512 96680 35552
rect 96720 35512 99360 35552
rect 576 35488 99360 35512
rect 576 34796 99516 34820
rect 576 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 7112 34796
rect 7152 34756 7194 34796
rect 7234 34756 7276 34796
rect 7316 34756 7358 34796
rect 7398 34756 7440 34796
rect 7480 34756 11112 34796
rect 11152 34756 11194 34796
rect 11234 34756 11276 34796
rect 11316 34756 11358 34796
rect 11398 34756 11440 34796
rect 11480 34756 15112 34796
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15480 34756 19112 34796
rect 19152 34756 19194 34796
rect 19234 34756 19276 34796
rect 19316 34756 19358 34796
rect 19398 34756 19440 34796
rect 19480 34756 23112 34796
rect 23152 34756 23194 34796
rect 23234 34756 23276 34796
rect 23316 34756 23358 34796
rect 23398 34756 23440 34796
rect 23480 34756 27112 34796
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27480 34756 31112 34796
rect 31152 34756 31194 34796
rect 31234 34756 31276 34796
rect 31316 34756 31358 34796
rect 31398 34756 31440 34796
rect 31480 34756 35112 34796
rect 35152 34756 35194 34796
rect 35234 34756 35276 34796
rect 35316 34756 35358 34796
rect 35398 34756 35440 34796
rect 35480 34756 39112 34796
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39480 34756 43112 34796
rect 43152 34756 43194 34796
rect 43234 34756 43276 34796
rect 43316 34756 43358 34796
rect 43398 34756 43440 34796
rect 43480 34756 47112 34796
rect 47152 34756 47194 34796
rect 47234 34756 47276 34796
rect 47316 34756 47358 34796
rect 47398 34756 47440 34796
rect 47480 34756 51112 34796
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51480 34756 55112 34796
rect 55152 34756 55194 34796
rect 55234 34756 55276 34796
rect 55316 34756 55358 34796
rect 55398 34756 55440 34796
rect 55480 34756 59112 34796
rect 59152 34756 59194 34796
rect 59234 34756 59276 34796
rect 59316 34756 59358 34796
rect 59398 34756 59440 34796
rect 59480 34756 63112 34796
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63480 34756 67112 34796
rect 67152 34756 67194 34796
rect 67234 34756 67276 34796
rect 67316 34756 67358 34796
rect 67398 34756 67440 34796
rect 67480 34756 71112 34796
rect 71152 34756 71194 34796
rect 71234 34756 71276 34796
rect 71316 34756 71358 34796
rect 71398 34756 71440 34796
rect 71480 34756 75112 34796
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75480 34756 79112 34796
rect 79152 34756 79194 34796
rect 79234 34756 79276 34796
rect 79316 34756 79358 34796
rect 79398 34756 79440 34796
rect 79480 34756 83112 34796
rect 83152 34756 83194 34796
rect 83234 34756 83276 34796
rect 83316 34756 83358 34796
rect 83398 34756 83440 34796
rect 83480 34756 87112 34796
rect 87152 34756 87194 34796
rect 87234 34756 87276 34796
rect 87316 34756 87358 34796
rect 87398 34756 87440 34796
rect 87480 34756 91112 34796
rect 91152 34756 91194 34796
rect 91234 34756 91276 34796
rect 91316 34756 91358 34796
rect 91398 34756 91440 34796
rect 91480 34756 95112 34796
rect 95152 34756 95194 34796
rect 95234 34756 95276 34796
rect 95316 34756 95358 34796
rect 95398 34756 95440 34796
rect 95480 34756 99112 34796
rect 99152 34756 99194 34796
rect 99234 34756 99276 34796
rect 99316 34756 99358 34796
rect 99398 34756 99440 34796
rect 99480 34756 99516 34796
rect 576 34732 99516 34756
rect 91459 34460 91517 34461
rect 91459 34420 91468 34460
rect 91508 34420 91517 34460
rect 91459 34419 91517 34420
rect 93379 34460 93437 34461
rect 93379 34420 93388 34460
rect 93428 34420 93437 34460
rect 93379 34419 93437 34420
rect 91659 34208 91701 34217
rect 91659 34168 91660 34208
rect 91700 34168 91701 34208
rect 91659 34159 91701 34168
rect 93579 34208 93621 34217
rect 93579 34168 93580 34208
rect 93620 34168 93621 34208
rect 93579 34159 93621 34168
rect 576 34040 99360 34064
rect 576 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 8352 34040
rect 8392 34000 8434 34040
rect 8474 34000 8516 34040
rect 8556 34000 8598 34040
rect 8638 34000 8680 34040
rect 8720 34000 12352 34040
rect 12392 34000 12434 34040
rect 12474 34000 12516 34040
rect 12556 34000 12598 34040
rect 12638 34000 12680 34040
rect 12720 34000 16352 34040
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16720 34000 20352 34040
rect 20392 34000 20434 34040
rect 20474 34000 20516 34040
rect 20556 34000 20598 34040
rect 20638 34000 20680 34040
rect 20720 34000 24352 34040
rect 24392 34000 24434 34040
rect 24474 34000 24516 34040
rect 24556 34000 24598 34040
rect 24638 34000 24680 34040
rect 24720 34000 28352 34040
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28720 34000 32352 34040
rect 32392 34000 32434 34040
rect 32474 34000 32516 34040
rect 32556 34000 32598 34040
rect 32638 34000 32680 34040
rect 32720 34000 36352 34040
rect 36392 34000 36434 34040
rect 36474 34000 36516 34040
rect 36556 34000 36598 34040
rect 36638 34000 36680 34040
rect 36720 34000 40352 34040
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40720 34000 44352 34040
rect 44392 34000 44434 34040
rect 44474 34000 44516 34040
rect 44556 34000 44598 34040
rect 44638 34000 44680 34040
rect 44720 34000 48352 34040
rect 48392 34000 48434 34040
rect 48474 34000 48516 34040
rect 48556 34000 48598 34040
rect 48638 34000 48680 34040
rect 48720 34000 52352 34040
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52720 34000 56352 34040
rect 56392 34000 56434 34040
rect 56474 34000 56516 34040
rect 56556 34000 56598 34040
rect 56638 34000 56680 34040
rect 56720 34000 60352 34040
rect 60392 34000 60434 34040
rect 60474 34000 60516 34040
rect 60556 34000 60598 34040
rect 60638 34000 60680 34040
rect 60720 34000 64352 34040
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64720 34000 68352 34040
rect 68392 34000 68434 34040
rect 68474 34000 68516 34040
rect 68556 34000 68598 34040
rect 68638 34000 68680 34040
rect 68720 34000 99360 34040
rect 576 33976 99360 34000
rect 95499 33872 95541 33881
rect 95499 33832 95500 33872
rect 95540 33832 95541 33872
rect 95499 33823 95541 33832
rect 73219 33620 73277 33621
rect 73219 33580 73228 33620
rect 73268 33580 73277 33620
rect 73219 33579 73277 33580
rect 73603 33620 73661 33621
rect 73603 33580 73612 33620
rect 73652 33580 73661 33620
rect 73603 33579 73661 33580
rect 74083 33620 74141 33621
rect 74083 33580 74092 33620
rect 74132 33580 74141 33620
rect 74083 33579 74141 33580
rect 74467 33620 74525 33621
rect 74467 33580 74476 33620
rect 74516 33580 74525 33620
rect 74467 33579 74525 33580
rect 74851 33620 74909 33621
rect 74851 33580 74860 33620
rect 74900 33580 74909 33620
rect 74851 33579 74909 33580
rect 75331 33620 75389 33621
rect 75331 33580 75340 33620
rect 75380 33580 75389 33620
rect 75331 33579 75389 33580
rect 75811 33620 75869 33621
rect 75811 33580 75820 33620
rect 75860 33580 75869 33620
rect 75811 33579 75869 33580
rect 76195 33620 76253 33621
rect 76195 33580 76204 33620
rect 76244 33580 76253 33620
rect 76195 33579 76253 33580
rect 76579 33620 76637 33621
rect 76579 33580 76588 33620
rect 76628 33580 76637 33620
rect 76579 33579 76637 33580
rect 76963 33620 77021 33621
rect 76963 33580 76972 33620
rect 77012 33580 77021 33620
rect 76963 33579 77021 33580
rect 77443 33620 77501 33621
rect 77443 33580 77452 33620
rect 77492 33580 77501 33620
rect 77443 33579 77501 33580
rect 77827 33620 77885 33621
rect 77827 33580 77836 33620
rect 77876 33580 77885 33620
rect 77827 33579 77885 33580
rect 78211 33620 78269 33621
rect 78211 33580 78220 33620
rect 78260 33580 78269 33620
rect 78211 33579 78269 33580
rect 78595 33620 78653 33621
rect 78595 33580 78604 33620
rect 78644 33580 78653 33620
rect 78595 33579 78653 33580
rect 78979 33620 79037 33621
rect 78979 33580 78988 33620
rect 79028 33580 79037 33620
rect 78979 33579 79037 33580
rect 79363 33620 79421 33621
rect 79363 33580 79372 33620
rect 79412 33580 79421 33620
rect 79363 33579 79421 33580
rect 79747 33620 79805 33621
rect 79747 33580 79756 33620
rect 79796 33580 79805 33620
rect 79747 33579 79805 33580
rect 80323 33620 80381 33621
rect 80323 33580 80332 33620
rect 80372 33580 80381 33620
rect 80323 33579 80381 33580
rect 80899 33620 80957 33621
rect 80899 33580 80908 33620
rect 80948 33580 80957 33620
rect 80899 33579 80957 33580
rect 81091 33620 81149 33621
rect 81091 33580 81100 33620
rect 81140 33580 81149 33620
rect 81091 33579 81149 33580
rect 81667 33620 81725 33621
rect 81667 33580 81676 33620
rect 81716 33580 81725 33620
rect 81667 33579 81725 33580
rect 82051 33620 82109 33621
rect 82051 33580 82060 33620
rect 82100 33580 82109 33620
rect 82051 33579 82109 33580
rect 82435 33620 82493 33621
rect 82435 33580 82444 33620
rect 82484 33580 82493 33620
rect 82435 33579 82493 33580
rect 82819 33620 82877 33621
rect 82819 33580 82828 33620
rect 82868 33580 82877 33620
rect 82819 33579 82877 33580
rect 83203 33620 83261 33621
rect 83203 33580 83212 33620
rect 83252 33580 83261 33620
rect 83203 33579 83261 33580
rect 83587 33620 83645 33621
rect 83587 33580 83596 33620
rect 83636 33580 83645 33620
rect 83587 33579 83645 33580
rect 83971 33620 84029 33621
rect 83971 33580 83980 33620
rect 84020 33580 84029 33620
rect 83971 33579 84029 33580
rect 84355 33620 84413 33621
rect 84355 33580 84364 33620
rect 84404 33580 84413 33620
rect 84355 33579 84413 33580
rect 84739 33620 84797 33621
rect 84739 33580 84748 33620
rect 84788 33580 84797 33620
rect 84739 33579 84797 33580
rect 85123 33620 85181 33621
rect 85123 33580 85132 33620
rect 85172 33580 85181 33620
rect 85123 33579 85181 33580
rect 85507 33620 85565 33621
rect 85507 33580 85516 33620
rect 85556 33580 85565 33620
rect 85507 33579 85565 33580
rect 85891 33620 85949 33621
rect 85891 33580 85900 33620
rect 85940 33580 85949 33620
rect 85891 33579 85949 33580
rect 86275 33620 86333 33621
rect 86275 33580 86284 33620
rect 86324 33580 86333 33620
rect 86275 33579 86333 33580
rect 86659 33620 86717 33621
rect 86659 33580 86668 33620
rect 86708 33580 86717 33620
rect 86659 33579 86717 33580
rect 87043 33620 87101 33621
rect 87043 33580 87052 33620
rect 87092 33580 87101 33620
rect 87043 33579 87101 33580
rect 87427 33620 87485 33621
rect 87427 33580 87436 33620
rect 87476 33580 87485 33620
rect 87427 33579 87485 33580
rect 87811 33620 87869 33621
rect 87811 33580 87820 33620
rect 87860 33580 87869 33620
rect 87811 33579 87869 33580
rect 88195 33620 88253 33621
rect 88195 33580 88204 33620
rect 88244 33580 88253 33620
rect 88195 33579 88253 33580
rect 88579 33620 88637 33621
rect 88579 33580 88588 33620
rect 88628 33580 88637 33620
rect 88579 33579 88637 33580
rect 88963 33620 89021 33621
rect 88963 33580 88972 33620
rect 89012 33580 89021 33620
rect 88963 33579 89021 33580
rect 89347 33620 89405 33621
rect 89347 33580 89356 33620
rect 89396 33580 89405 33620
rect 89347 33579 89405 33580
rect 89731 33620 89789 33621
rect 89731 33580 89740 33620
rect 89780 33580 89789 33620
rect 89731 33579 89789 33580
rect 90115 33620 90173 33621
rect 90115 33580 90124 33620
rect 90164 33580 90173 33620
rect 90115 33579 90173 33580
rect 90499 33620 90557 33621
rect 90499 33580 90508 33620
rect 90548 33580 90557 33620
rect 90499 33579 90557 33580
rect 90883 33620 90941 33621
rect 90883 33580 90892 33620
rect 90932 33580 90941 33620
rect 90883 33579 90941 33580
rect 91267 33620 91325 33621
rect 91267 33580 91276 33620
rect 91316 33580 91325 33620
rect 91267 33579 91325 33580
rect 91651 33620 91709 33621
rect 91651 33580 91660 33620
rect 91700 33580 91709 33620
rect 91651 33579 91709 33580
rect 91843 33620 91901 33621
rect 91843 33580 91852 33620
rect 91892 33580 91901 33620
rect 91843 33579 91901 33580
rect 92227 33620 92285 33621
rect 92227 33580 92236 33620
rect 92276 33580 92285 33620
rect 92227 33579 92285 33580
rect 92611 33620 92669 33621
rect 92611 33580 92620 33620
rect 92660 33580 92669 33620
rect 92611 33579 92669 33580
rect 93187 33620 93245 33621
rect 93187 33580 93196 33620
rect 93236 33580 93245 33620
rect 93187 33579 93245 33580
rect 93571 33620 93629 33621
rect 93571 33580 93580 33620
rect 93620 33580 93629 33620
rect 93571 33579 93629 33580
rect 94051 33620 94109 33621
rect 94051 33580 94060 33620
rect 94100 33580 94109 33620
rect 94051 33579 94109 33580
rect 94243 33620 94301 33621
rect 94243 33580 94252 33620
rect 94292 33580 94301 33620
rect 94243 33579 94301 33580
rect 94627 33620 94685 33621
rect 94627 33580 94636 33620
rect 94676 33580 94685 33620
rect 94627 33579 94685 33580
rect 95299 33620 95357 33621
rect 95299 33580 95308 33620
rect 95348 33580 95357 33620
rect 95299 33579 95357 33580
rect 95683 33620 95741 33621
rect 95683 33580 95692 33620
rect 95732 33580 95741 33620
rect 95683 33579 95741 33580
rect 96067 33620 96125 33621
rect 96067 33580 96076 33620
rect 96116 33580 96125 33620
rect 96067 33579 96125 33580
rect 96451 33620 96509 33621
rect 96451 33580 96460 33620
rect 96500 33580 96509 33620
rect 96451 33579 96509 33580
rect 96835 33620 96893 33621
rect 96835 33580 96844 33620
rect 96884 33580 96893 33620
rect 96835 33579 96893 33580
rect 97219 33620 97277 33621
rect 97219 33580 97228 33620
rect 97268 33580 97277 33620
rect 97219 33579 97277 33580
rect 97603 33620 97661 33621
rect 97603 33580 97612 33620
rect 97652 33580 97661 33620
rect 97603 33579 97661 33580
rect 97987 33620 98045 33621
rect 97987 33580 97996 33620
rect 98036 33580 98045 33620
rect 97987 33579 98045 33580
rect 98371 33620 98429 33621
rect 98371 33580 98380 33620
rect 98420 33580 98429 33620
rect 98371 33579 98429 33580
rect 80523 33536 80565 33545
rect 80523 33496 80524 33536
rect 80564 33496 80565 33536
rect 80523 33487 80565 33496
rect 81291 33536 81333 33545
rect 81291 33496 81292 33536
rect 81332 33496 81333 33536
rect 81291 33487 81333 33496
rect 82251 33536 82293 33545
rect 82251 33496 82252 33536
rect 82292 33496 82293 33536
rect 82251 33487 82293 33496
rect 92811 33536 92853 33545
rect 92811 33496 92812 33536
rect 92852 33496 92853 33536
rect 92811 33487 92853 33496
rect 73419 33452 73461 33461
rect 73419 33412 73420 33452
rect 73460 33412 73461 33452
rect 73419 33403 73461 33412
rect 73803 33452 73845 33461
rect 73803 33412 73804 33452
rect 73844 33412 73845 33452
rect 73803 33403 73845 33412
rect 74283 33452 74325 33461
rect 74283 33412 74284 33452
rect 74324 33412 74325 33452
rect 74283 33403 74325 33412
rect 74667 33452 74709 33461
rect 74667 33412 74668 33452
rect 74708 33412 74709 33452
rect 74667 33403 74709 33412
rect 75051 33452 75093 33461
rect 75051 33412 75052 33452
rect 75092 33412 75093 33452
rect 75051 33403 75093 33412
rect 75531 33452 75573 33461
rect 75531 33412 75532 33452
rect 75572 33412 75573 33452
rect 75531 33403 75573 33412
rect 76011 33452 76053 33461
rect 76011 33412 76012 33452
rect 76052 33412 76053 33452
rect 76011 33403 76053 33412
rect 76395 33452 76437 33461
rect 76395 33412 76396 33452
rect 76436 33412 76437 33452
rect 76395 33403 76437 33412
rect 76779 33452 76821 33461
rect 76779 33412 76780 33452
rect 76820 33412 76821 33452
rect 76779 33403 76821 33412
rect 77163 33452 77205 33461
rect 77163 33412 77164 33452
rect 77204 33412 77205 33452
rect 77163 33403 77205 33412
rect 77643 33452 77685 33461
rect 77643 33412 77644 33452
rect 77684 33412 77685 33452
rect 77643 33403 77685 33412
rect 78027 33452 78069 33461
rect 78027 33412 78028 33452
rect 78068 33412 78069 33452
rect 78027 33403 78069 33412
rect 78411 33452 78453 33461
rect 78411 33412 78412 33452
rect 78452 33412 78453 33452
rect 78411 33403 78453 33412
rect 78795 33452 78837 33461
rect 78795 33412 78796 33452
rect 78836 33412 78837 33452
rect 78795 33403 78837 33412
rect 79179 33452 79221 33461
rect 79179 33412 79180 33452
rect 79220 33412 79221 33452
rect 79179 33403 79221 33412
rect 79563 33452 79605 33461
rect 79563 33412 79564 33452
rect 79604 33412 79605 33452
rect 79563 33403 79605 33412
rect 79947 33452 79989 33461
rect 79947 33412 79948 33452
rect 79988 33412 79989 33452
rect 79947 33403 79989 33412
rect 80715 33452 80757 33461
rect 80715 33412 80716 33452
rect 80756 33412 80757 33452
rect 80715 33403 80757 33412
rect 81483 33452 81525 33461
rect 81483 33412 81484 33452
rect 81524 33412 81525 33452
rect 81483 33403 81525 33412
rect 81867 33452 81909 33461
rect 81867 33412 81868 33452
rect 81908 33412 81909 33452
rect 81867 33403 81909 33412
rect 82635 33452 82677 33461
rect 82635 33412 82636 33452
rect 82676 33412 82677 33452
rect 82635 33403 82677 33412
rect 83019 33452 83061 33461
rect 83019 33412 83020 33452
rect 83060 33412 83061 33452
rect 83019 33403 83061 33412
rect 83403 33452 83445 33461
rect 83403 33412 83404 33452
rect 83444 33412 83445 33452
rect 83403 33403 83445 33412
rect 83787 33452 83829 33461
rect 83787 33412 83788 33452
rect 83828 33412 83829 33452
rect 83787 33403 83829 33412
rect 84171 33452 84213 33461
rect 84171 33412 84172 33452
rect 84212 33412 84213 33452
rect 84171 33403 84213 33412
rect 84555 33452 84597 33461
rect 84555 33412 84556 33452
rect 84596 33412 84597 33452
rect 84555 33403 84597 33412
rect 84939 33452 84981 33461
rect 84939 33412 84940 33452
rect 84980 33412 84981 33452
rect 84939 33403 84981 33412
rect 85323 33452 85365 33461
rect 85323 33412 85324 33452
rect 85364 33412 85365 33452
rect 85323 33403 85365 33412
rect 85707 33452 85749 33461
rect 85707 33412 85708 33452
rect 85748 33412 85749 33452
rect 85707 33403 85749 33412
rect 86091 33452 86133 33461
rect 86091 33412 86092 33452
rect 86132 33412 86133 33452
rect 86091 33403 86133 33412
rect 86475 33452 86517 33461
rect 86475 33412 86476 33452
rect 86516 33412 86517 33452
rect 86475 33403 86517 33412
rect 86859 33452 86901 33461
rect 86859 33412 86860 33452
rect 86900 33412 86901 33452
rect 86859 33403 86901 33412
rect 87243 33452 87285 33461
rect 87243 33412 87244 33452
rect 87284 33412 87285 33452
rect 87243 33403 87285 33412
rect 87627 33452 87669 33461
rect 87627 33412 87628 33452
rect 87668 33412 87669 33452
rect 87627 33403 87669 33412
rect 88011 33452 88053 33461
rect 88011 33412 88012 33452
rect 88052 33412 88053 33452
rect 88011 33403 88053 33412
rect 88395 33452 88437 33461
rect 88395 33412 88396 33452
rect 88436 33412 88437 33452
rect 88395 33403 88437 33412
rect 88779 33452 88821 33461
rect 88779 33412 88780 33452
rect 88820 33412 88821 33452
rect 88779 33403 88821 33412
rect 89163 33452 89205 33461
rect 89163 33412 89164 33452
rect 89204 33412 89205 33452
rect 89163 33403 89205 33412
rect 89547 33452 89589 33461
rect 89547 33412 89548 33452
rect 89588 33412 89589 33452
rect 89547 33403 89589 33412
rect 89931 33452 89973 33461
rect 89931 33412 89932 33452
rect 89972 33412 89973 33452
rect 89931 33403 89973 33412
rect 90315 33452 90357 33461
rect 90315 33412 90316 33452
rect 90356 33412 90357 33452
rect 90315 33403 90357 33412
rect 90699 33452 90741 33461
rect 90699 33412 90700 33452
rect 90740 33412 90741 33452
rect 90699 33403 90741 33412
rect 91083 33452 91125 33461
rect 91083 33412 91084 33452
rect 91124 33412 91125 33452
rect 91083 33403 91125 33412
rect 91467 33452 91509 33461
rect 91467 33412 91468 33452
rect 91508 33412 91509 33452
rect 91467 33403 91509 33412
rect 92043 33452 92085 33461
rect 92043 33412 92044 33452
rect 92084 33412 92085 33452
rect 92043 33403 92085 33412
rect 92427 33452 92469 33461
rect 92427 33412 92428 33452
rect 92468 33412 92469 33452
rect 92427 33403 92469 33412
rect 93003 33452 93045 33461
rect 93003 33412 93004 33452
rect 93044 33412 93045 33452
rect 93003 33403 93045 33412
rect 93387 33452 93429 33461
rect 93387 33412 93388 33452
rect 93428 33412 93429 33452
rect 93387 33403 93429 33412
rect 93867 33452 93909 33461
rect 93867 33412 93868 33452
rect 93908 33412 93909 33452
rect 93867 33403 93909 33412
rect 94443 33452 94485 33461
rect 94443 33412 94444 33452
rect 94484 33412 94485 33452
rect 94443 33403 94485 33412
rect 94827 33452 94869 33461
rect 94827 33412 94828 33452
rect 94868 33412 94869 33452
rect 94827 33403 94869 33412
rect 95115 33452 95157 33461
rect 95115 33412 95116 33452
rect 95156 33412 95157 33452
rect 95115 33403 95157 33412
rect 95883 33452 95925 33461
rect 95883 33412 95884 33452
rect 95924 33412 95925 33452
rect 95883 33403 95925 33412
rect 96267 33452 96309 33461
rect 96267 33412 96268 33452
rect 96308 33412 96309 33452
rect 96267 33403 96309 33412
rect 96651 33452 96693 33461
rect 96651 33412 96652 33452
rect 96692 33412 96693 33452
rect 96651 33403 96693 33412
rect 97035 33452 97077 33461
rect 97035 33412 97036 33452
rect 97076 33412 97077 33452
rect 97035 33403 97077 33412
rect 97419 33452 97461 33461
rect 97419 33412 97420 33452
rect 97460 33412 97461 33452
rect 97419 33403 97461 33412
rect 97803 33452 97845 33461
rect 97803 33412 97804 33452
rect 97844 33412 97845 33452
rect 97803 33403 97845 33412
rect 98187 33452 98229 33461
rect 98187 33412 98188 33452
rect 98228 33412 98229 33452
rect 98187 33403 98229 33412
rect 576 33284 99360 33308
rect 576 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 7112 33284
rect 7152 33244 7194 33284
rect 7234 33244 7276 33284
rect 7316 33244 7358 33284
rect 7398 33244 7440 33284
rect 7480 33244 11112 33284
rect 11152 33244 11194 33284
rect 11234 33244 11276 33284
rect 11316 33244 11358 33284
rect 11398 33244 11440 33284
rect 11480 33244 15112 33284
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15480 33244 19112 33284
rect 19152 33244 19194 33284
rect 19234 33244 19276 33284
rect 19316 33244 19358 33284
rect 19398 33244 19440 33284
rect 19480 33244 23112 33284
rect 23152 33244 23194 33284
rect 23234 33244 23276 33284
rect 23316 33244 23358 33284
rect 23398 33244 23440 33284
rect 23480 33244 27112 33284
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27480 33244 31112 33284
rect 31152 33244 31194 33284
rect 31234 33244 31276 33284
rect 31316 33244 31358 33284
rect 31398 33244 31440 33284
rect 31480 33244 35112 33284
rect 35152 33244 35194 33284
rect 35234 33244 35276 33284
rect 35316 33244 35358 33284
rect 35398 33244 35440 33284
rect 35480 33244 39112 33284
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39480 33244 43112 33284
rect 43152 33244 43194 33284
rect 43234 33244 43276 33284
rect 43316 33244 43358 33284
rect 43398 33244 43440 33284
rect 43480 33244 47112 33284
rect 47152 33244 47194 33284
rect 47234 33244 47276 33284
rect 47316 33244 47358 33284
rect 47398 33244 47440 33284
rect 47480 33244 51112 33284
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51480 33244 55112 33284
rect 55152 33244 55194 33284
rect 55234 33244 55276 33284
rect 55316 33244 55358 33284
rect 55398 33244 55440 33284
rect 55480 33244 59112 33284
rect 59152 33244 59194 33284
rect 59234 33244 59276 33284
rect 59316 33244 59358 33284
rect 59398 33244 59440 33284
rect 59480 33244 63112 33284
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63480 33244 67112 33284
rect 67152 33244 67194 33284
rect 67234 33244 67276 33284
rect 67316 33244 67358 33284
rect 67398 33244 67440 33284
rect 67480 33244 99360 33284
rect 576 33220 99360 33244
rect 74187 33116 74229 33125
rect 74187 33076 74188 33116
rect 74228 33076 74229 33116
rect 74187 33067 74229 33076
rect 77067 33116 77109 33125
rect 77067 33076 77068 33116
rect 77108 33076 77109 33116
rect 77067 33067 77109 33076
rect 78891 33116 78933 33125
rect 78891 33076 78892 33116
rect 78932 33076 78933 33116
rect 78891 33067 78933 33076
rect 86475 33116 86517 33125
rect 86475 33076 86476 33116
rect 86516 33076 86517 33116
rect 86475 33067 86517 33076
rect 90891 33116 90933 33125
rect 90891 33076 90892 33116
rect 90932 33076 90933 33116
rect 90891 33067 90933 33076
rect 92331 33116 92373 33125
rect 92331 33076 92332 33116
rect 92372 33076 92373 33116
rect 92331 33067 92373 33076
rect 94059 33116 94101 33125
rect 94059 33076 94060 33116
rect 94100 33076 94101 33116
rect 94059 33067 94101 33076
rect 74859 33032 74901 33041
rect 74859 32992 74860 33032
rect 74900 32992 74901 33032
rect 74859 32983 74901 32992
rect 76011 33032 76053 33041
rect 76011 32992 76012 33032
rect 76052 32992 76053 33032
rect 76011 32983 76053 32992
rect 83307 33032 83349 33041
rect 83307 32992 83308 33032
rect 83348 32992 83349 33032
rect 83307 32983 83349 32992
rect 84843 33032 84885 33041
rect 84843 32992 84844 33032
rect 84884 32992 84885 33032
rect 84843 32983 84885 32992
rect 88107 33032 88149 33041
rect 88107 32992 88108 33032
rect 88148 32992 88149 33032
rect 88107 32983 88149 32992
rect 92715 33032 92757 33041
rect 92715 32992 92716 33032
rect 92756 32992 92757 33032
rect 92715 32983 92757 32992
rect 94923 33032 94965 33041
rect 94923 32992 94924 33032
rect 94964 32992 94965 33032
rect 94923 32983 94965 32992
rect 96939 33032 96981 33041
rect 96939 32992 96940 33032
rect 96980 32992 96981 33032
rect 96939 32983 96981 32992
rect 90691 32959 90749 32960
rect 72643 32948 72701 32949
rect 72643 32908 72652 32948
rect 72692 32908 72701 32948
rect 72643 32907 72701 32908
rect 74371 32948 74429 32949
rect 74371 32908 74380 32948
rect 74420 32908 74429 32948
rect 74371 32907 74429 32908
rect 74659 32948 74717 32949
rect 74659 32908 74668 32948
rect 74708 32908 74717 32948
rect 74659 32907 74717 32908
rect 75811 32948 75869 32949
rect 75811 32908 75820 32948
rect 75860 32908 75869 32948
rect 75811 32907 75869 32908
rect 77251 32948 77309 32949
rect 77251 32908 77260 32948
rect 77300 32908 77309 32948
rect 77251 32907 77309 32908
rect 78691 32948 78749 32949
rect 78691 32908 78700 32948
rect 78740 32908 78749 32948
rect 78691 32907 78749 32908
rect 79371 32948 79413 32957
rect 79371 32908 79372 32948
rect 79412 32908 79413 32948
rect 79371 32899 79413 32908
rect 80611 32948 80669 32949
rect 80611 32908 80620 32948
rect 80660 32908 80669 32948
rect 80611 32907 80669 32908
rect 82051 32948 82109 32949
rect 82051 32908 82060 32948
rect 82100 32908 82109 32948
rect 82051 32907 82109 32908
rect 83107 32948 83165 32949
rect 83107 32908 83116 32948
rect 83156 32908 83165 32948
rect 83107 32907 83165 32908
rect 83595 32948 83637 32957
rect 83595 32908 83596 32948
rect 83636 32908 83637 32948
rect 83595 32899 83637 32908
rect 84643 32948 84701 32949
rect 84643 32908 84652 32948
rect 84692 32908 84701 32948
rect 84643 32907 84701 32908
rect 86275 32948 86333 32949
rect 86275 32908 86284 32948
rect 86324 32908 86333 32948
rect 86275 32907 86333 32908
rect 86955 32948 86997 32957
rect 86955 32908 86956 32948
rect 86996 32908 86997 32948
rect 86955 32899 86997 32908
rect 87907 32948 87965 32949
rect 87907 32908 87916 32948
rect 87956 32908 87965 32948
rect 87907 32907 87965 32908
rect 88395 32948 88437 32957
rect 88395 32908 88396 32948
rect 88436 32908 88437 32948
rect 88395 32899 88437 32908
rect 88963 32948 89021 32949
rect 88963 32908 88972 32948
rect 89012 32908 89021 32948
rect 88963 32907 89021 32908
rect 90027 32948 90069 32957
rect 90027 32908 90028 32948
rect 90068 32908 90069 32948
rect 90691 32919 90700 32959
rect 90740 32919 90749 32959
rect 90691 32918 90749 32919
rect 91083 32948 91125 32957
rect 90027 32899 90069 32908
rect 91083 32908 91084 32948
rect 91124 32908 91125 32948
rect 91083 32899 91125 32908
rect 92515 32948 92573 32949
rect 92515 32908 92524 32948
rect 92564 32908 92573 32948
rect 92515 32907 92573 32908
rect 93099 32948 93141 32957
rect 93099 32908 93100 32948
rect 93140 32908 93141 32948
rect 93099 32899 93141 32908
rect 93859 32948 93917 32949
rect 93859 32908 93868 32948
rect 93908 32908 93917 32948
rect 93859 32907 93917 32908
rect 95115 32948 95157 32957
rect 95115 32908 95116 32948
rect 95156 32908 95157 32948
rect 95115 32899 95157 32908
rect 96739 32948 96797 32949
rect 96739 32908 96748 32948
rect 96788 32908 96797 32948
rect 96739 32907 96797 32908
rect 98659 32948 98717 32949
rect 98659 32908 98668 32948
rect 98708 32908 98717 32948
rect 98659 32907 98717 32908
rect 80037 32877 80095 32878
rect 71491 32864 71549 32865
rect 71491 32824 71500 32864
rect 71540 32824 71549 32864
rect 71491 32823 71549 32824
rect 71595 32864 71637 32873
rect 71595 32824 71596 32864
rect 71636 32824 71637 32864
rect 71595 32815 71637 32824
rect 72355 32864 72413 32865
rect 72355 32824 72364 32864
rect 72404 32824 72413 32864
rect 72355 32823 72413 32824
rect 73027 32864 73085 32865
rect 73027 32824 73036 32864
rect 73076 32824 73085 32864
rect 73027 32823 73085 32824
rect 73603 32864 73661 32865
rect 73603 32824 73612 32864
rect 73652 32824 73661 32864
rect 73603 32823 73661 32824
rect 73987 32864 74045 32865
rect 73987 32824 73996 32864
rect 74036 32824 74045 32864
rect 73987 32823 74045 32824
rect 75139 32864 75197 32865
rect 75139 32824 75148 32864
rect 75188 32824 75197 32864
rect 75139 32823 75197 32824
rect 75427 32864 75485 32865
rect 75427 32824 75436 32864
rect 75476 32824 75485 32864
rect 75427 32823 75485 32824
rect 76203 32864 76245 32873
rect 76203 32824 76204 32864
rect 76244 32824 76245 32864
rect 76203 32815 76245 32824
rect 76291 32864 76349 32865
rect 76291 32824 76300 32864
rect 76340 32824 76349 32864
rect 76291 32823 76349 32824
rect 76579 32864 76637 32865
rect 76579 32824 76588 32864
rect 76628 32824 76637 32864
rect 76579 32823 76637 32824
rect 76867 32864 76925 32865
rect 76867 32824 76876 32864
rect 76916 32824 76925 32864
rect 76867 32823 76925 32824
rect 77443 32864 77501 32865
rect 77443 32824 77452 32864
rect 77492 32824 77501 32864
rect 77443 32823 77501 32824
rect 77547 32864 77589 32873
rect 77547 32824 77548 32864
rect 77588 32824 77589 32864
rect 77547 32815 77589 32824
rect 77827 32864 77885 32865
rect 77827 32824 77836 32864
rect 77876 32824 77885 32864
rect 77827 32823 77885 32824
rect 78115 32864 78173 32865
rect 78115 32824 78124 32864
rect 78164 32824 78173 32864
rect 78115 32823 78173 32824
rect 78315 32864 78357 32873
rect 78315 32824 78316 32864
rect 78356 32824 78357 32864
rect 78315 32815 78357 32824
rect 78403 32864 78461 32865
rect 78403 32824 78412 32864
rect 78452 32824 78461 32864
rect 78403 32823 78461 32824
rect 79075 32864 79133 32865
rect 79075 32824 79084 32864
rect 79124 32824 79133 32864
rect 79075 32823 79133 32824
rect 79459 32864 79517 32865
rect 79459 32824 79468 32864
rect 79508 32824 79517 32864
rect 79459 32823 79517 32824
rect 79659 32864 79701 32873
rect 79659 32824 79660 32864
rect 79700 32824 79701 32864
rect 79659 32815 79701 32824
rect 79747 32864 79805 32865
rect 79747 32824 79756 32864
rect 79796 32824 79805 32864
rect 80037 32837 80046 32877
rect 80086 32837 80095 32877
rect 91747 32877 91805 32878
rect 80037 32836 80095 32837
rect 80227 32864 80285 32865
rect 79747 32823 79805 32824
rect 80227 32824 80236 32864
rect 80276 32824 80285 32864
rect 80227 32823 80285 32824
rect 81003 32864 81045 32873
rect 81003 32824 81004 32864
rect 81044 32824 81045 32864
rect 81003 32815 81045 32824
rect 81091 32864 81149 32865
rect 81091 32824 81100 32864
rect 81140 32824 81149 32864
rect 81091 32823 81149 32824
rect 81379 32864 81437 32865
rect 81379 32824 81388 32864
rect 81428 32824 81437 32864
rect 81379 32823 81437 32824
rect 81667 32864 81725 32865
rect 81667 32824 81676 32864
rect 81716 32824 81725 32864
rect 81667 32823 81725 32824
rect 82243 32864 82301 32865
rect 82243 32824 82252 32864
rect 82292 32824 82301 32864
rect 82243 32823 82301 32824
rect 82347 32864 82389 32873
rect 82347 32824 82348 32864
rect 82388 32824 82389 32864
rect 82347 32815 82389 32824
rect 82627 32864 82685 32865
rect 82627 32824 82636 32864
rect 82676 32824 82685 32864
rect 82627 32823 82685 32824
rect 82915 32864 82973 32865
rect 82915 32824 82924 32864
rect 82964 32824 82973 32864
rect 82915 32823 82973 32824
rect 83491 32864 83549 32865
rect 83491 32824 83500 32864
rect 83540 32824 83549 32864
rect 83491 32823 83549 32824
rect 83787 32864 83829 32873
rect 83787 32824 83788 32864
rect 83828 32824 83829 32864
rect 83787 32815 83829 32824
rect 83875 32864 83933 32865
rect 83875 32824 83884 32864
rect 83924 32824 83933 32864
rect 83875 32823 83933 32824
rect 84163 32864 84221 32865
rect 84163 32824 84172 32864
rect 84212 32824 84221 32864
rect 84163 32823 84221 32824
rect 84451 32864 84509 32865
rect 84451 32824 84460 32864
rect 84500 32824 84509 32864
rect 84451 32823 84509 32824
rect 85027 32864 85085 32865
rect 85027 32824 85036 32864
rect 85076 32824 85085 32864
rect 85027 32823 85085 32824
rect 85131 32864 85173 32873
rect 85131 32824 85132 32864
rect 85172 32824 85173 32864
rect 85131 32815 85173 32824
rect 85411 32864 85469 32865
rect 85411 32824 85420 32864
rect 85460 32824 85469 32864
rect 85411 32823 85469 32824
rect 85699 32864 85757 32865
rect 85699 32824 85708 32864
rect 85748 32824 85757 32864
rect 85699 32823 85757 32824
rect 85987 32864 86045 32865
rect 85987 32824 85996 32864
rect 86036 32824 86045 32864
rect 85987 32823 86045 32824
rect 86659 32864 86717 32865
rect 86659 32824 86668 32864
rect 86708 32824 86717 32864
rect 86659 32823 86717 32824
rect 87043 32864 87101 32865
rect 87043 32824 87052 32864
rect 87092 32824 87101 32864
rect 87043 32823 87101 32824
rect 87243 32864 87285 32873
rect 87243 32824 87244 32864
rect 87284 32824 87285 32864
rect 87243 32815 87285 32824
rect 87331 32864 87389 32865
rect 87331 32824 87340 32864
rect 87380 32824 87389 32864
rect 87331 32823 87389 32824
rect 87619 32864 87677 32865
rect 87619 32824 87628 32864
rect 87668 32824 87677 32864
rect 87619 32823 87677 32824
rect 88291 32864 88349 32865
rect 88291 32824 88300 32864
rect 88340 32824 88349 32864
rect 88291 32823 88349 32824
rect 88587 32864 88629 32873
rect 88587 32824 88588 32864
rect 88628 32824 88629 32864
rect 88587 32815 88629 32824
rect 88675 32864 88733 32865
rect 88675 32824 88684 32864
rect 88724 32824 88733 32864
rect 88675 32823 88733 32824
rect 89443 32864 89501 32865
rect 89443 32824 89452 32864
rect 89492 32824 89501 32864
rect 89443 32823 89501 32824
rect 89643 32864 89685 32873
rect 89643 32824 89644 32864
rect 89684 32824 89685 32864
rect 89643 32815 89685 32824
rect 89731 32864 89789 32865
rect 89731 32824 89740 32864
rect 89780 32824 89789 32864
rect 89731 32823 89789 32824
rect 89923 32864 89981 32865
rect 89923 32824 89932 32864
rect 89972 32824 89981 32864
rect 89923 32823 89981 32824
rect 90307 32864 90365 32865
rect 90307 32824 90316 32864
rect 90356 32824 90365 32864
rect 90307 32823 90365 32824
rect 91171 32864 91229 32865
rect 91171 32824 91180 32864
rect 91220 32824 91229 32864
rect 91171 32823 91229 32824
rect 91371 32864 91413 32873
rect 91371 32824 91372 32864
rect 91412 32824 91413 32864
rect 91371 32815 91413 32824
rect 91459 32864 91517 32865
rect 91459 32824 91468 32864
rect 91508 32824 91517 32864
rect 91747 32837 91756 32877
rect 91796 32837 91805 32877
rect 91747 32836 91805 32837
rect 92035 32864 92093 32865
rect 91459 32823 91517 32824
rect 92035 32824 92044 32864
rect 92084 32824 92093 32864
rect 92035 32823 92093 32824
rect 92803 32864 92861 32865
rect 92803 32824 92812 32864
rect 92852 32824 92861 32864
rect 92803 32823 92861 32824
rect 92995 32864 93053 32865
rect 92995 32824 93004 32864
rect 93044 32824 93053 32864
rect 92995 32823 93053 32824
rect 93291 32864 93333 32873
rect 93291 32824 93292 32864
rect 93332 32824 93333 32864
rect 93291 32815 93333 32824
rect 93379 32864 93437 32865
rect 93379 32824 93388 32864
rect 93428 32824 93437 32864
rect 93379 32823 93437 32824
rect 93667 32864 93725 32865
rect 93667 32824 93676 32864
rect 93716 32824 93725 32864
rect 93667 32823 93725 32824
rect 94251 32864 94293 32873
rect 94251 32824 94252 32864
rect 94292 32824 94293 32864
rect 94251 32815 94293 32824
rect 94339 32864 94397 32865
rect 94339 32824 94348 32864
rect 94388 32824 94397 32864
rect 94339 32823 94397 32824
rect 94627 32864 94685 32865
rect 94627 32824 94636 32864
rect 94676 32824 94685 32864
rect 94627 32823 94685 32824
rect 94819 32864 94877 32865
rect 94819 32824 94828 32864
rect 94868 32824 94877 32864
rect 94819 32823 94877 32824
rect 95203 32864 95261 32865
rect 95203 32824 95212 32864
rect 95252 32824 95261 32864
rect 95203 32823 95261 32824
rect 95491 32864 95549 32865
rect 95491 32824 95500 32864
rect 95540 32824 95549 32864
rect 95491 32823 95549 32824
rect 95683 32864 95741 32865
rect 95683 32824 95692 32864
rect 95732 32824 95741 32864
rect 95683 32823 95741 32824
rect 95787 32864 95829 32873
rect 95787 32824 95788 32864
rect 95828 32824 95829 32864
rect 95787 32815 95829 32824
rect 96067 32864 96125 32865
rect 96067 32824 96076 32864
rect 96116 32824 96125 32864
rect 96067 32823 96125 32824
rect 96355 32864 96413 32865
rect 96355 32824 96364 32864
rect 96404 32824 96413 32864
rect 96355 32823 96413 32824
rect 97219 32864 97277 32865
rect 97219 32824 97228 32864
rect 97268 32824 97277 32864
rect 97219 32823 97277 32824
rect 97507 32864 97565 32865
rect 97507 32824 97516 32864
rect 97556 32824 97565 32864
rect 97507 32823 97565 32824
rect 97795 32864 97853 32865
rect 97795 32824 97804 32864
rect 97844 32824 97853 32864
rect 97795 32823 97853 32824
rect 98083 32864 98141 32865
rect 98083 32824 98092 32864
rect 98132 32824 98141 32864
rect 98083 32823 98141 32824
rect 98851 32864 98909 32865
rect 98851 32824 98860 32864
rect 98900 32824 98909 32864
rect 98851 32823 98909 32824
rect 99139 32864 99197 32865
rect 99139 32824 99148 32864
rect 99188 32824 99197 32864
rect 99139 32823 99197 32824
rect 85899 32780 85941 32789
rect 85899 32740 85900 32780
rect 85940 32740 85941 32780
rect 85899 32731 85941 32740
rect 93579 32780 93621 32789
rect 93579 32740 93580 32780
rect 93620 32740 93621 32780
rect 93579 32731 93621 32740
rect 94539 32780 94581 32789
rect 94539 32740 94540 32780
rect 94580 32740 94581 32780
rect 94539 32731 94581 32740
rect 95979 32780 96021 32789
rect 95979 32740 95980 32780
rect 96020 32740 96021 32780
rect 95979 32731 96021 32740
rect 72459 32696 72501 32705
rect 72459 32656 72460 32696
rect 72500 32656 72501 32696
rect 72459 32647 72501 32656
rect 72843 32696 72885 32705
rect 72843 32656 72844 32696
rect 72884 32656 72885 32696
rect 72843 32647 72885 32656
rect 73131 32696 73173 32705
rect 73131 32656 73132 32696
rect 73172 32656 73173 32696
rect 73131 32647 73173 32656
rect 73707 32696 73749 32705
rect 73707 32656 73708 32696
rect 73748 32656 73749 32696
rect 73707 32647 73749 32656
rect 73899 32696 73941 32705
rect 73899 32656 73900 32696
rect 73940 32656 73941 32696
rect 73899 32647 73941 32656
rect 75051 32696 75093 32705
rect 75051 32656 75052 32696
rect 75092 32656 75093 32696
rect 75051 32647 75093 32656
rect 75339 32696 75381 32705
rect 75339 32656 75340 32696
rect 75380 32656 75381 32696
rect 75339 32647 75381 32656
rect 76491 32696 76533 32705
rect 76491 32656 76492 32696
rect 76532 32656 76533 32696
rect 76491 32647 76533 32656
rect 76779 32696 76821 32705
rect 76779 32656 76780 32696
rect 76820 32656 76821 32696
rect 76779 32647 76821 32656
rect 77739 32696 77781 32705
rect 77739 32656 77740 32696
rect 77780 32656 77781 32696
rect 77739 32647 77781 32656
rect 78027 32696 78069 32705
rect 78027 32656 78028 32696
rect 78068 32656 78069 32696
rect 78027 32647 78069 32656
rect 79179 32696 79221 32705
rect 79179 32656 79180 32696
rect 79220 32656 79221 32696
rect 79179 32647 79221 32656
rect 79947 32696 79989 32705
rect 79947 32656 79948 32696
rect 79988 32656 79989 32696
rect 79947 32647 79989 32656
rect 80331 32696 80373 32705
rect 80331 32656 80332 32696
rect 80372 32656 80373 32696
rect 80331 32647 80373 32656
rect 80811 32696 80853 32705
rect 80811 32656 80812 32696
rect 80852 32656 80853 32696
rect 80811 32647 80853 32656
rect 81291 32696 81333 32705
rect 81291 32656 81292 32696
rect 81332 32656 81333 32696
rect 81291 32647 81333 32656
rect 81579 32696 81621 32705
rect 81579 32656 81580 32696
rect 81620 32656 81621 32696
rect 81579 32647 81621 32656
rect 81867 32696 81909 32705
rect 81867 32656 81868 32696
rect 81908 32656 81909 32696
rect 81867 32647 81909 32656
rect 82539 32696 82581 32705
rect 82539 32656 82540 32696
rect 82580 32656 82581 32696
rect 82539 32647 82581 32656
rect 82827 32696 82869 32705
rect 82827 32656 82828 32696
rect 82868 32656 82869 32696
rect 82827 32647 82869 32656
rect 84075 32696 84117 32705
rect 84075 32656 84076 32696
rect 84116 32656 84117 32696
rect 84075 32647 84117 32656
rect 84363 32696 84405 32705
rect 84363 32656 84364 32696
rect 84404 32656 84405 32696
rect 84363 32647 84405 32656
rect 85323 32696 85365 32705
rect 85323 32656 85324 32696
rect 85364 32656 85365 32696
rect 85323 32647 85365 32656
rect 85611 32696 85653 32705
rect 85611 32656 85612 32696
rect 85652 32656 85653 32696
rect 85611 32647 85653 32656
rect 86763 32696 86805 32705
rect 86763 32656 86764 32696
rect 86804 32656 86805 32696
rect 86763 32647 86805 32656
rect 87531 32696 87573 32705
rect 87531 32656 87532 32696
rect 87572 32656 87573 32696
rect 87531 32647 87573 32656
rect 89163 32696 89205 32705
rect 89163 32656 89164 32696
rect 89204 32656 89205 32696
rect 89163 32647 89205 32656
rect 89355 32696 89397 32705
rect 89355 32656 89356 32696
rect 89396 32656 89397 32696
rect 89355 32647 89397 32656
rect 90219 32696 90261 32705
rect 90219 32656 90220 32696
rect 90260 32656 90261 32696
rect 90219 32647 90261 32656
rect 91659 32696 91701 32705
rect 91659 32656 91660 32696
rect 91700 32656 91701 32696
rect 91659 32647 91701 32656
rect 91947 32696 91989 32705
rect 91947 32656 91948 32696
rect 91988 32656 91989 32696
rect 91947 32647 91989 32656
rect 95403 32696 95445 32705
rect 95403 32656 95404 32696
rect 95444 32656 95445 32696
rect 95403 32647 95445 32656
rect 96267 32696 96309 32705
rect 96267 32656 96268 32696
rect 96308 32656 96309 32696
rect 96267 32647 96309 32656
rect 97131 32696 97173 32705
rect 97131 32656 97132 32696
rect 97172 32656 97173 32696
rect 97131 32647 97173 32656
rect 97419 32696 97461 32705
rect 97419 32656 97420 32696
rect 97460 32656 97461 32696
rect 97419 32647 97461 32656
rect 97707 32696 97749 32705
rect 97707 32656 97708 32696
rect 97748 32656 97749 32696
rect 97707 32647 97749 32656
rect 97995 32696 98037 32705
rect 97995 32656 97996 32696
rect 98036 32656 98037 32696
rect 97995 32647 98037 32656
rect 98475 32696 98517 32705
rect 98475 32656 98476 32696
rect 98516 32656 98517 32696
rect 98475 32647 98517 32656
rect 98955 32696 98997 32705
rect 98955 32656 98956 32696
rect 98996 32656 98997 32696
rect 98955 32647 98997 32656
rect 99243 32696 99285 32705
rect 99243 32656 99244 32696
rect 99284 32656 99285 32696
rect 99243 32647 99285 32656
rect 576 32528 99360 32552
rect 576 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 8352 32528
rect 8392 32488 8434 32528
rect 8474 32488 8516 32528
rect 8556 32488 8598 32528
rect 8638 32488 8680 32528
rect 8720 32488 12352 32528
rect 12392 32488 12434 32528
rect 12474 32488 12516 32528
rect 12556 32488 12598 32528
rect 12638 32488 12680 32528
rect 12720 32488 16352 32528
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16720 32488 20352 32528
rect 20392 32488 20434 32528
rect 20474 32488 20516 32528
rect 20556 32488 20598 32528
rect 20638 32488 20680 32528
rect 20720 32488 24352 32528
rect 24392 32488 24434 32528
rect 24474 32488 24516 32528
rect 24556 32488 24598 32528
rect 24638 32488 24680 32528
rect 24720 32488 28352 32528
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28720 32488 32352 32528
rect 32392 32488 32434 32528
rect 32474 32488 32516 32528
rect 32556 32488 32598 32528
rect 32638 32488 32680 32528
rect 32720 32488 36352 32528
rect 36392 32488 36434 32528
rect 36474 32488 36516 32528
rect 36556 32488 36598 32528
rect 36638 32488 36680 32528
rect 36720 32488 40352 32528
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40720 32488 44352 32528
rect 44392 32488 44434 32528
rect 44474 32488 44516 32528
rect 44556 32488 44598 32528
rect 44638 32488 44680 32528
rect 44720 32488 48352 32528
rect 48392 32488 48434 32528
rect 48474 32488 48516 32528
rect 48556 32488 48598 32528
rect 48638 32488 48680 32528
rect 48720 32488 52352 32528
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52720 32488 56352 32528
rect 56392 32488 56434 32528
rect 56474 32488 56516 32528
rect 56556 32488 56598 32528
rect 56638 32488 56680 32528
rect 56720 32488 60352 32528
rect 60392 32488 60434 32528
rect 60474 32488 60516 32528
rect 60556 32488 60598 32528
rect 60638 32488 60680 32528
rect 60720 32488 64352 32528
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64720 32488 68352 32528
rect 68392 32488 68434 32528
rect 68474 32488 68516 32528
rect 68556 32488 68598 32528
rect 68638 32488 68680 32528
rect 68720 32488 99360 32528
rect 576 32464 99360 32488
rect 70731 32360 70773 32369
rect 70731 32320 70732 32360
rect 70772 32320 70773 32360
rect 70731 32311 70773 32320
rect 71403 32360 71445 32369
rect 71403 32320 71404 32360
rect 71444 32320 71445 32360
rect 71403 32311 71445 32320
rect 70915 32108 70973 32109
rect 70915 32068 70924 32108
rect 70964 32068 70973 32108
rect 70915 32067 70973 32068
rect 71203 32108 71261 32109
rect 71203 32068 71212 32108
rect 71252 32068 71261 32108
rect 71203 32067 71261 32068
rect 70731 31940 70773 31949
rect 70731 31900 70732 31940
rect 70772 31900 70773 31940
rect 70731 31891 70773 31900
rect 576 31772 71520 31796
rect 576 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 7112 31772
rect 7152 31732 7194 31772
rect 7234 31732 7276 31772
rect 7316 31732 7358 31772
rect 7398 31732 7440 31772
rect 7480 31732 11112 31772
rect 11152 31732 11194 31772
rect 11234 31732 11276 31772
rect 11316 31732 11358 31772
rect 11398 31732 11440 31772
rect 11480 31732 15112 31772
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15480 31732 19112 31772
rect 19152 31732 19194 31772
rect 19234 31732 19276 31772
rect 19316 31732 19358 31772
rect 19398 31732 19440 31772
rect 19480 31732 23112 31772
rect 23152 31732 23194 31772
rect 23234 31732 23276 31772
rect 23316 31732 23358 31772
rect 23398 31732 23440 31772
rect 23480 31732 27112 31772
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27480 31732 31112 31772
rect 31152 31732 31194 31772
rect 31234 31732 31276 31772
rect 31316 31732 31358 31772
rect 31398 31732 31440 31772
rect 31480 31732 35112 31772
rect 35152 31732 35194 31772
rect 35234 31732 35276 31772
rect 35316 31732 35358 31772
rect 35398 31732 35440 31772
rect 35480 31732 39112 31772
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39480 31732 43112 31772
rect 43152 31732 43194 31772
rect 43234 31732 43276 31772
rect 43316 31732 43358 31772
rect 43398 31732 43440 31772
rect 43480 31732 47112 31772
rect 47152 31732 47194 31772
rect 47234 31732 47276 31772
rect 47316 31732 47358 31772
rect 47398 31732 47440 31772
rect 47480 31732 51112 31772
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51480 31732 55112 31772
rect 55152 31732 55194 31772
rect 55234 31732 55276 31772
rect 55316 31732 55358 31772
rect 55398 31732 55440 31772
rect 55480 31732 59112 31772
rect 59152 31732 59194 31772
rect 59234 31732 59276 31772
rect 59316 31732 59358 31772
rect 59398 31732 59440 31772
rect 59480 31732 63112 31772
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63480 31732 67112 31772
rect 67152 31732 67194 31772
rect 67234 31732 67276 31772
rect 67316 31732 67358 31772
rect 67398 31732 67440 31772
rect 67480 31732 71520 31772
rect 576 31708 71520 31732
rect 70827 31604 70869 31613
rect 70827 31564 70828 31604
rect 70868 31564 70869 31604
rect 70827 31555 70869 31564
rect 71115 31520 71157 31529
rect 71115 31480 71116 31520
rect 71156 31480 71157 31520
rect 71115 31471 71157 31480
rect 70627 31436 70685 31437
rect 70627 31396 70636 31436
rect 70676 31396 70685 31436
rect 70627 31395 70685 31396
rect 71011 31352 71069 31353
rect 71011 31312 71020 31352
rect 71060 31312 71069 31352
rect 71011 31311 71069 31312
rect 576 31016 71520 31040
rect 576 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 8352 31016
rect 8392 30976 8434 31016
rect 8474 30976 8516 31016
rect 8556 30976 8598 31016
rect 8638 30976 8680 31016
rect 8720 30976 12352 31016
rect 12392 30976 12434 31016
rect 12474 30976 12516 31016
rect 12556 30976 12598 31016
rect 12638 30976 12680 31016
rect 12720 30976 16352 31016
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16720 30976 20352 31016
rect 20392 30976 20434 31016
rect 20474 30976 20516 31016
rect 20556 30976 20598 31016
rect 20638 30976 20680 31016
rect 20720 30976 24352 31016
rect 24392 30976 24434 31016
rect 24474 30976 24516 31016
rect 24556 30976 24598 31016
rect 24638 30976 24680 31016
rect 24720 30976 28352 31016
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28720 30976 32352 31016
rect 32392 30976 32434 31016
rect 32474 30976 32516 31016
rect 32556 30976 32598 31016
rect 32638 30976 32680 31016
rect 32720 30976 36352 31016
rect 36392 30976 36434 31016
rect 36474 30976 36516 31016
rect 36556 30976 36598 31016
rect 36638 30976 36680 31016
rect 36720 30976 40352 31016
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40720 30976 44352 31016
rect 44392 30976 44434 31016
rect 44474 30976 44516 31016
rect 44556 30976 44598 31016
rect 44638 30976 44680 31016
rect 44720 30976 48352 31016
rect 48392 30976 48434 31016
rect 48474 30976 48516 31016
rect 48556 30976 48598 31016
rect 48638 30976 48680 31016
rect 48720 30976 52352 31016
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52720 30976 56352 31016
rect 56392 30976 56434 31016
rect 56474 30976 56516 31016
rect 56556 30976 56598 31016
rect 56638 30976 56680 31016
rect 56720 30976 60352 31016
rect 60392 30976 60434 31016
rect 60474 30976 60516 31016
rect 60556 30976 60598 31016
rect 60638 30976 60680 31016
rect 60720 30976 64352 31016
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64720 30976 68352 31016
rect 68392 30976 68434 31016
rect 68474 30976 68516 31016
rect 68556 30976 68598 31016
rect 68638 30976 68680 31016
rect 68720 30976 71520 31016
rect 576 30952 71520 30976
rect 576 30260 71520 30284
rect 576 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 7112 30260
rect 7152 30220 7194 30260
rect 7234 30220 7276 30260
rect 7316 30220 7358 30260
rect 7398 30220 7440 30260
rect 7480 30220 11112 30260
rect 11152 30220 11194 30260
rect 11234 30220 11276 30260
rect 11316 30220 11358 30260
rect 11398 30220 11440 30260
rect 11480 30220 15112 30260
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15480 30220 19112 30260
rect 19152 30220 19194 30260
rect 19234 30220 19276 30260
rect 19316 30220 19358 30260
rect 19398 30220 19440 30260
rect 19480 30220 23112 30260
rect 23152 30220 23194 30260
rect 23234 30220 23276 30260
rect 23316 30220 23358 30260
rect 23398 30220 23440 30260
rect 23480 30220 27112 30260
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27480 30220 31112 30260
rect 31152 30220 31194 30260
rect 31234 30220 31276 30260
rect 31316 30220 31358 30260
rect 31398 30220 31440 30260
rect 31480 30220 35112 30260
rect 35152 30220 35194 30260
rect 35234 30220 35276 30260
rect 35316 30220 35358 30260
rect 35398 30220 35440 30260
rect 35480 30220 39112 30260
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39480 30220 43112 30260
rect 43152 30220 43194 30260
rect 43234 30220 43276 30260
rect 43316 30220 43358 30260
rect 43398 30220 43440 30260
rect 43480 30220 47112 30260
rect 47152 30220 47194 30260
rect 47234 30220 47276 30260
rect 47316 30220 47358 30260
rect 47398 30220 47440 30260
rect 47480 30220 51112 30260
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51480 30220 55112 30260
rect 55152 30220 55194 30260
rect 55234 30220 55276 30260
rect 55316 30220 55358 30260
rect 55398 30220 55440 30260
rect 55480 30220 59112 30260
rect 59152 30220 59194 30260
rect 59234 30220 59276 30260
rect 59316 30220 59358 30260
rect 59398 30220 59440 30260
rect 59480 30220 63112 30260
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63480 30220 67112 30260
rect 67152 30220 67194 30260
rect 67234 30220 67276 30260
rect 67316 30220 67358 30260
rect 67398 30220 67440 30260
rect 67480 30220 71520 30260
rect 576 30196 71520 30220
rect 576 29504 71520 29528
rect 576 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 8352 29504
rect 8392 29464 8434 29504
rect 8474 29464 8516 29504
rect 8556 29464 8598 29504
rect 8638 29464 8680 29504
rect 8720 29464 12352 29504
rect 12392 29464 12434 29504
rect 12474 29464 12516 29504
rect 12556 29464 12598 29504
rect 12638 29464 12680 29504
rect 12720 29464 16352 29504
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16720 29464 20352 29504
rect 20392 29464 20434 29504
rect 20474 29464 20516 29504
rect 20556 29464 20598 29504
rect 20638 29464 20680 29504
rect 20720 29464 24352 29504
rect 24392 29464 24434 29504
rect 24474 29464 24516 29504
rect 24556 29464 24598 29504
rect 24638 29464 24680 29504
rect 24720 29464 28352 29504
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28720 29464 32352 29504
rect 32392 29464 32434 29504
rect 32474 29464 32516 29504
rect 32556 29464 32598 29504
rect 32638 29464 32680 29504
rect 32720 29464 36352 29504
rect 36392 29464 36434 29504
rect 36474 29464 36516 29504
rect 36556 29464 36598 29504
rect 36638 29464 36680 29504
rect 36720 29464 40352 29504
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40720 29464 44352 29504
rect 44392 29464 44434 29504
rect 44474 29464 44516 29504
rect 44556 29464 44598 29504
rect 44638 29464 44680 29504
rect 44720 29464 48352 29504
rect 48392 29464 48434 29504
rect 48474 29464 48516 29504
rect 48556 29464 48598 29504
rect 48638 29464 48680 29504
rect 48720 29464 52352 29504
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52720 29464 56352 29504
rect 56392 29464 56434 29504
rect 56474 29464 56516 29504
rect 56556 29464 56598 29504
rect 56638 29464 56680 29504
rect 56720 29464 60352 29504
rect 60392 29464 60434 29504
rect 60474 29464 60516 29504
rect 60556 29464 60598 29504
rect 60638 29464 60680 29504
rect 60720 29464 64352 29504
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64720 29464 68352 29504
rect 68392 29464 68434 29504
rect 68474 29464 68516 29504
rect 68556 29464 68598 29504
rect 68638 29464 68680 29504
rect 68720 29464 71520 29504
rect 576 29440 71520 29464
rect 576 28748 71520 28772
rect 576 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 7112 28748
rect 7152 28708 7194 28748
rect 7234 28708 7276 28748
rect 7316 28708 7358 28748
rect 7398 28708 7440 28748
rect 7480 28708 11112 28748
rect 11152 28708 11194 28748
rect 11234 28708 11276 28748
rect 11316 28708 11358 28748
rect 11398 28708 11440 28748
rect 11480 28708 15112 28748
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15480 28708 19112 28748
rect 19152 28708 19194 28748
rect 19234 28708 19276 28748
rect 19316 28708 19358 28748
rect 19398 28708 19440 28748
rect 19480 28708 23112 28748
rect 23152 28708 23194 28748
rect 23234 28708 23276 28748
rect 23316 28708 23358 28748
rect 23398 28708 23440 28748
rect 23480 28708 27112 28748
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27480 28708 31112 28748
rect 31152 28708 31194 28748
rect 31234 28708 31276 28748
rect 31316 28708 31358 28748
rect 31398 28708 31440 28748
rect 31480 28708 35112 28748
rect 35152 28708 35194 28748
rect 35234 28708 35276 28748
rect 35316 28708 35358 28748
rect 35398 28708 35440 28748
rect 35480 28708 39112 28748
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39480 28708 43112 28748
rect 43152 28708 43194 28748
rect 43234 28708 43276 28748
rect 43316 28708 43358 28748
rect 43398 28708 43440 28748
rect 43480 28708 47112 28748
rect 47152 28708 47194 28748
rect 47234 28708 47276 28748
rect 47316 28708 47358 28748
rect 47398 28708 47440 28748
rect 47480 28708 51112 28748
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51480 28708 55112 28748
rect 55152 28708 55194 28748
rect 55234 28708 55276 28748
rect 55316 28708 55358 28748
rect 55398 28708 55440 28748
rect 55480 28708 59112 28748
rect 59152 28708 59194 28748
rect 59234 28708 59276 28748
rect 59316 28708 59358 28748
rect 59398 28708 59440 28748
rect 59480 28708 63112 28748
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63480 28708 67112 28748
rect 67152 28708 67194 28748
rect 67234 28708 67276 28748
rect 67316 28708 67358 28748
rect 67398 28708 67440 28748
rect 67480 28708 71520 28748
rect 576 28684 71520 28708
rect 576 27992 71520 28016
rect 576 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 8352 27992
rect 8392 27952 8434 27992
rect 8474 27952 8516 27992
rect 8556 27952 8598 27992
rect 8638 27952 8680 27992
rect 8720 27952 12352 27992
rect 12392 27952 12434 27992
rect 12474 27952 12516 27992
rect 12556 27952 12598 27992
rect 12638 27952 12680 27992
rect 12720 27952 16352 27992
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16720 27952 20352 27992
rect 20392 27952 20434 27992
rect 20474 27952 20516 27992
rect 20556 27952 20598 27992
rect 20638 27952 20680 27992
rect 20720 27952 24352 27992
rect 24392 27952 24434 27992
rect 24474 27952 24516 27992
rect 24556 27952 24598 27992
rect 24638 27952 24680 27992
rect 24720 27952 28352 27992
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28720 27952 32352 27992
rect 32392 27952 32434 27992
rect 32474 27952 32516 27992
rect 32556 27952 32598 27992
rect 32638 27952 32680 27992
rect 32720 27952 36352 27992
rect 36392 27952 36434 27992
rect 36474 27952 36516 27992
rect 36556 27952 36598 27992
rect 36638 27952 36680 27992
rect 36720 27952 40352 27992
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40720 27952 44352 27992
rect 44392 27952 44434 27992
rect 44474 27952 44516 27992
rect 44556 27952 44598 27992
rect 44638 27952 44680 27992
rect 44720 27952 48352 27992
rect 48392 27952 48434 27992
rect 48474 27952 48516 27992
rect 48556 27952 48598 27992
rect 48638 27952 48680 27992
rect 48720 27952 52352 27992
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52720 27952 56352 27992
rect 56392 27952 56434 27992
rect 56474 27952 56516 27992
rect 56556 27952 56598 27992
rect 56638 27952 56680 27992
rect 56720 27952 60352 27992
rect 60392 27952 60434 27992
rect 60474 27952 60516 27992
rect 60556 27952 60598 27992
rect 60638 27952 60680 27992
rect 60720 27952 64352 27992
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64720 27952 68352 27992
rect 68392 27952 68434 27992
rect 68474 27952 68516 27992
rect 68556 27952 68598 27992
rect 68638 27952 68680 27992
rect 68720 27952 71520 27992
rect 576 27928 71520 27952
rect 69955 27656 70013 27657
rect 69955 27616 69964 27656
rect 70004 27616 70013 27656
rect 69955 27615 70013 27616
rect 70147 27656 70205 27657
rect 70147 27616 70156 27656
rect 70196 27616 70205 27656
rect 70147 27615 70205 27616
rect 70915 27656 70973 27657
rect 70915 27616 70924 27656
rect 70964 27616 70973 27656
rect 70915 27615 70973 27616
rect 70531 27572 70589 27573
rect 70531 27532 70540 27572
rect 70580 27532 70589 27572
rect 70531 27531 70589 27532
rect 71203 27572 71261 27573
rect 71203 27532 71212 27572
rect 71252 27532 71261 27572
rect 71203 27531 71261 27532
rect 70347 27488 70389 27497
rect 70347 27448 70348 27488
rect 70388 27448 70389 27488
rect 70347 27439 70389 27448
rect 71019 27404 71061 27413
rect 71019 27364 71020 27404
rect 71060 27364 71061 27404
rect 71019 27355 71061 27364
rect 71403 27404 71445 27413
rect 71403 27364 71404 27404
rect 71444 27364 71445 27404
rect 71403 27355 71445 27364
rect 576 27236 71520 27260
rect 576 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 7112 27236
rect 7152 27196 7194 27236
rect 7234 27196 7276 27236
rect 7316 27196 7358 27236
rect 7398 27196 7440 27236
rect 7480 27196 11112 27236
rect 11152 27196 11194 27236
rect 11234 27196 11276 27236
rect 11316 27196 11358 27236
rect 11398 27196 11440 27236
rect 11480 27196 15112 27236
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15480 27196 19112 27236
rect 19152 27196 19194 27236
rect 19234 27196 19276 27236
rect 19316 27196 19358 27236
rect 19398 27196 19440 27236
rect 19480 27196 23112 27236
rect 23152 27196 23194 27236
rect 23234 27196 23276 27236
rect 23316 27196 23358 27236
rect 23398 27196 23440 27236
rect 23480 27196 27112 27236
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27480 27196 31112 27236
rect 31152 27196 31194 27236
rect 31234 27196 31276 27236
rect 31316 27196 31358 27236
rect 31398 27196 31440 27236
rect 31480 27196 35112 27236
rect 35152 27196 35194 27236
rect 35234 27196 35276 27236
rect 35316 27196 35358 27236
rect 35398 27196 35440 27236
rect 35480 27196 39112 27236
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39480 27196 43112 27236
rect 43152 27196 43194 27236
rect 43234 27196 43276 27236
rect 43316 27196 43358 27236
rect 43398 27196 43440 27236
rect 43480 27196 47112 27236
rect 47152 27196 47194 27236
rect 47234 27196 47276 27236
rect 47316 27196 47358 27236
rect 47398 27196 47440 27236
rect 47480 27196 51112 27236
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51480 27196 55112 27236
rect 55152 27196 55194 27236
rect 55234 27196 55276 27236
rect 55316 27196 55358 27236
rect 55398 27196 55440 27236
rect 55480 27196 59112 27236
rect 59152 27196 59194 27236
rect 59234 27196 59276 27236
rect 59316 27196 59358 27236
rect 59398 27196 59440 27236
rect 59480 27196 63112 27236
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63480 27196 67112 27236
rect 67152 27196 67194 27236
rect 67234 27196 67276 27236
rect 67316 27196 67358 27236
rect 67398 27196 67440 27236
rect 67480 27196 71520 27236
rect 576 27172 71520 27196
rect 69763 26900 69821 26901
rect 69763 26860 69772 26900
rect 69812 26860 69821 26900
rect 69763 26859 69821 26860
rect 70339 26900 70397 26901
rect 70339 26860 70348 26900
rect 70388 26860 70397 26900
rect 70339 26859 70397 26860
rect 70723 26900 70781 26901
rect 70723 26860 70732 26900
rect 70772 26860 70781 26900
rect 70723 26859 70781 26860
rect 71107 26900 71165 26901
rect 71107 26860 71116 26900
rect 71156 26860 71165 26900
rect 71107 26859 71165 26860
rect 69963 26648 70005 26657
rect 69963 26608 69964 26648
rect 70004 26608 70005 26648
rect 69963 26599 70005 26608
rect 70539 26648 70581 26657
rect 70539 26608 70540 26648
rect 70580 26608 70581 26648
rect 70539 26599 70581 26608
rect 70923 26648 70965 26657
rect 70923 26608 70924 26648
rect 70964 26608 70965 26648
rect 70923 26599 70965 26608
rect 71307 26648 71349 26657
rect 71307 26608 71308 26648
rect 71348 26608 71349 26648
rect 71307 26599 71349 26608
rect 576 26480 71520 26504
rect 576 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 8352 26480
rect 8392 26440 8434 26480
rect 8474 26440 8516 26480
rect 8556 26440 8598 26480
rect 8638 26440 8680 26480
rect 8720 26440 12352 26480
rect 12392 26440 12434 26480
rect 12474 26440 12516 26480
rect 12556 26440 12598 26480
rect 12638 26440 12680 26480
rect 12720 26440 16352 26480
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16720 26440 20352 26480
rect 20392 26440 20434 26480
rect 20474 26440 20516 26480
rect 20556 26440 20598 26480
rect 20638 26440 20680 26480
rect 20720 26440 24352 26480
rect 24392 26440 24434 26480
rect 24474 26440 24516 26480
rect 24556 26440 24598 26480
rect 24638 26440 24680 26480
rect 24720 26440 28352 26480
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28720 26440 32352 26480
rect 32392 26440 32434 26480
rect 32474 26440 32516 26480
rect 32556 26440 32598 26480
rect 32638 26440 32680 26480
rect 32720 26440 36352 26480
rect 36392 26440 36434 26480
rect 36474 26440 36516 26480
rect 36556 26440 36598 26480
rect 36638 26440 36680 26480
rect 36720 26440 40352 26480
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40720 26440 44352 26480
rect 44392 26440 44434 26480
rect 44474 26440 44516 26480
rect 44556 26440 44598 26480
rect 44638 26440 44680 26480
rect 44720 26440 48352 26480
rect 48392 26440 48434 26480
rect 48474 26440 48516 26480
rect 48556 26440 48598 26480
rect 48638 26440 48680 26480
rect 48720 26440 52352 26480
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52720 26440 56352 26480
rect 56392 26440 56434 26480
rect 56474 26440 56516 26480
rect 56556 26440 56598 26480
rect 56638 26440 56680 26480
rect 56720 26440 60352 26480
rect 60392 26440 60434 26480
rect 60474 26440 60516 26480
rect 60556 26440 60598 26480
rect 60638 26440 60680 26480
rect 60720 26440 64352 26480
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64720 26440 68352 26480
rect 68392 26440 68434 26480
rect 68474 26440 68516 26480
rect 68556 26440 68598 26480
rect 68638 26440 68680 26480
rect 68720 26440 71520 26480
rect 576 26416 71520 26440
rect 71019 26312 71061 26321
rect 71019 26272 71020 26312
rect 71060 26272 71061 26312
rect 71019 26263 71061 26272
rect 71403 26312 71445 26321
rect 71403 26272 71404 26312
rect 71444 26272 71445 26312
rect 71403 26263 71445 26272
rect 70915 26144 70973 26145
rect 70915 26104 70924 26144
rect 70964 26104 70973 26144
rect 70915 26103 70973 26104
rect 71299 26144 71357 26145
rect 71299 26104 71308 26144
rect 71348 26104 71357 26144
rect 71299 26103 71357 26104
rect 576 25724 99360 25748
rect 576 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 7112 25724
rect 7152 25684 7194 25724
rect 7234 25684 7276 25724
rect 7316 25684 7358 25724
rect 7398 25684 7440 25724
rect 7480 25684 11112 25724
rect 11152 25684 11194 25724
rect 11234 25684 11276 25724
rect 11316 25684 11358 25724
rect 11398 25684 11440 25724
rect 11480 25684 15112 25724
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15480 25684 19112 25724
rect 19152 25684 19194 25724
rect 19234 25684 19276 25724
rect 19316 25684 19358 25724
rect 19398 25684 19440 25724
rect 19480 25684 23112 25724
rect 23152 25684 23194 25724
rect 23234 25684 23276 25724
rect 23316 25684 23358 25724
rect 23398 25684 23440 25724
rect 23480 25684 27112 25724
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27480 25684 31112 25724
rect 31152 25684 31194 25724
rect 31234 25684 31276 25724
rect 31316 25684 31358 25724
rect 31398 25684 31440 25724
rect 31480 25684 35112 25724
rect 35152 25684 35194 25724
rect 35234 25684 35276 25724
rect 35316 25684 35358 25724
rect 35398 25684 35440 25724
rect 35480 25684 39112 25724
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39480 25684 43112 25724
rect 43152 25684 43194 25724
rect 43234 25684 43276 25724
rect 43316 25684 43358 25724
rect 43398 25684 43440 25724
rect 43480 25684 47112 25724
rect 47152 25684 47194 25724
rect 47234 25684 47276 25724
rect 47316 25684 47358 25724
rect 47398 25684 47440 25724
rect 47480 25684 51112 25724
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51480 25684 55112 25724
rect 55152 25684 55194 25724
rect 55234 25684 55276 25724
rect 55316 25684 55358 25724
rect 55398 25684 55440 25724
rect 55480 25684 59112 25724
rect 59152 25684 59194 25724
rect 59234 25684 59276 25724
rect 59316 25684 59358 25724
rect 59398 25684 59440 25724
rect 59480 25684 63112 25724
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63480 25684 67112 25724
rect 67152 25684 67194 25724
rect 67234 25684 67276 25724
rect 67316 25684 67358 25724
rect 67398 25684 67440 25724
rect 67480 25684 99360 25724
rect 576 25660 99360 25684
rect 72747 25556 72789 25565
rect 72747 25516 72748 25556
rect 72788 25516 72789 25556
rect 72747 25507 72789 25516
rect 73131 25556 73173 25565
rect 73131 25516 73132 25556
rect 73172 25516 73173 25556
rect 73131 25507 73173 25516
rect 73515 25556 73557 25565
rect 73515 25516 73516 25556
rect 73556 25516 73557 25556
rect 73515 25507 73557 25516
rect 74091 25556 74133 25565
rect 74091 25516 74092 25556
rect 74132 25516 74133 25556
rect 74091 25507 74133 25516
rect 75723 25556 75765 25565
rect 75723 25516 75724 25556
rect 75764 25516 75765 25556
rect 75723 25507 75765 25516
rect 75915 25556 75957 25565
rect 75915 25516 75916 25556
rect 75956 25516 75957 25556
rect 75915 25507 75957 25516
rect 76203 25556 76245 25565
rect 76203 25516 76204 25556
rect 76244 25516 76245 25556
rect 76203 25507 76245 25516
rect 76875 25556 76917 25565
rect 76875 25516 76876 25556
rect 76916 25516 76917 25556
rect 76875 25507 76917 25516
rect 77163 25556 77205 25565
rect 77163 25516 77164 25556
rect 77204 25516 77205 25556
rect 77163 25507 77205 25516
rect 77931 25556 77973 25565
rect 77931 25516 77932 25556
rect 77972 25516 77973 25556
rect 77931 25507 77973 25516
rect 78219 25556 78261 25565
rect 78219 25516 78220 25556
rect 78260 25516 78261 25556
rect 78219 25507 78261 25516
rect 78507 25556 78549 25565
rect 78507 25516 78508 25556
rect 78548 25516 78549 25556
rect 78507 25507 78549 25516
rect 78795 25556 78837 25565
rect 78795 25516 78796 25556
rect 78836 25516 78837 25556
rect 78795 25507 78837 25516
rect 79179 25556 79221 25565
rect 79179 25516 79180 25556
rect 79220 25516 79221 25556
rect 79179 25507 79221 25516
rect 79563 25556 79605 25565
rect 79563 25516 79564 25556
rect 79604 25516 79605 25556
rect 79563 25507 79605 25516
rect 79755 25556 79797 25565
rect 79755 25516 79756 25556
rect 79796 25516 79797 25556
rect 79755 25507 79797 25516
rect 80139 25556 80181 25565
rect 80139 25516 80140 25556
rect 80180 25516 80181 25556
rect 80139 25507 80181 25516
rect 80331 25556 80373 25565
rect 80331 25516 80332 25556
rect 80372 25516 80373 25556
rect 80331 25507 80373 25516
rect 80811 25556 80853 25565
rect 80811 25516 80812 25556
rect 80852 25516 80853 25556
rect 80811 25507 80853 25516
rect 81195 25556 81237 25565
rect 81195 25516 81196 25556
rect 81236 25516 81237 25556
rect 81195 25507 81237 25516
rect 81579 25556 81621 25565
rect 81579 25516 81580 25556
rect 81620 25516 81621 25556
rect 81579 25507 81621 25516
rect 82059 25556 82101 25565
rect 82059 25516 82060 25556
rect 82100 25516 82101 25556
rect 82059 25507 82101 25516
rect 82347 25556 82389 25565
rect 82347 25516 82348 25556
rect 82388 25516 82389 25556
rect 82347 25507 82389 25516
rect 82731 25556 82773 25565
rect 82731 25516 82732 25556
rect 82772 25516 82773 25556
rect 82731 25507 82773 25516
rect 83115 25556 83157 25565
rect 83115 25516 83116 25556
rect 83156 25516 83157 25556
rect 83115 25507 83157 25516
rect 83979 25556 84021 25565
rect 83979 25516 83980 25556
rect 84020 25516 84021 25556
rect 83979 25507 84021 25516
rect 84267 25556 84309 25565
rect 84267 25516 84268 25556
rect 84308 25516 84309 25556
rect 84267 25507 84309 25516
rect 84555 25556 84597 25565
rect 84555 25516 84556 25556
rect 84596 25516 84597 25556
rect 84555 25507 84597 25516
rect 84843 25556 84885 25565
rect 84843 25516 84844 25556
rect 84884 25516 84885 25556
rect 84843 25507 84885 25516
rect 85227 25556 85269 25565
rect 85227 25516 85228 25556
rect 85268 25516 85269 25556
rect 85227 25507 85269 25516
rect 85611 25556 85653 25565
rect 85611 25516 85612 25556
rect 85652 25516 85653 25556
rect 85611 25507 85653 25516
rect 85995 25556 86037 25565
rect 85995 25516 85996 25556
rect 86036 25516 86037 25556
rect 85995 25507 86037 25516
rect 86379 25556 86421 25565
rect 86379 25516 86380 25556
rect 86420 25516 86421 25556
rect 86379 25507 86421 25516
rect 87531 25556 87573 25565
rect 87531 25516 87532 25556
rect 87572 25516 87573 25556
rect 87531 25507 87573 25516
rect 87819 25556 87861 25565
rect 87819 25516 87820 25556
rect 87860 25516 87861 25556
rect 87819 25507 87861 25516
rect 88107 25556 88149 25565
rect 88107 25516 88108 25556
rect 88148 25516 88149 25556
rect 88107 25507 88149 25516
rect 88395 25556 88437 25565
rect 88395 25516 88396 25556
rect 88436 25516 88437 25556
rect 88395 25507 88437 25516
rect 88779 25556 88821 25565
rect 88779 25516 88780 25556
rect 88820 25516 88821 25556
rect 88779 25507 88821 25516
rect 89163 25556 89205 25565
rect 89163 25516 89164 25556
rect 89204 25516 89205 25556
rect 89163 25507 89205 25516
rect 89931 25556 89973 25565
rect 89931 25516 89932 25556
rect 89972 25516 89973 25556
rect 89931 25507 89973 25516
rect 90219 25556 90261 25565
rect 90219 25516 90220 25556
rect 90260 25516 90261 25556
rect 90219 25507 90261 25516
rect 90507 25556 90549 25565
rect 90507 25516 90508 25556
rect 90548 25516 90549 25556
rect 90507 25507 90549 25516
rect 90795 25556 90837 25565
rect 90795 25516 90796 25556
rect 90836 25516 90837 25556
rect 90795 25507 90837 25516
rect 91179 25556 91221 25565
rect 91179 25516 91180 25556
rect 91220 25516 91221 25556
rect 91179 25507 91221 25516
rect 91563 25556 91605 25565
rect 91563 25516 91564 25556
rect 91604 25516 91605 25556
rect 91563 25507 91605 25516
rect 92043 25556 92085 25565
rect 92043 25516 92044 25556
rect 92084 25516 92085 25556
rect 92043 25507 92085 25516
rect 92811 25556 92853 25565
rect 92811 25516 92812 25556
rect 92852 25516 92853 25556
rect 92811 25507 92853 25516
rect 93195 25556 93237 25565
rect 93195 25516 93196 25556
rect 93236 25516 93237 25556
rect 93195 25507 93237 25516
rect 93579 25556 93621 25565
rect 93579 25516 93580 25556
rect 93620 25516 93621 25556
rect 93579 25507 93621 25516
rect 94059 25556 94101 25565
rect 94059 25516 94060 25556
rect 94100 25516 94101 25556
rect 94059 25507 94101 25516
rect 94347 25556 94389 25565
rect 94347 25516 94348 25556
rect 94388 25516 94389 25556
rect 94347 25507 94389 25516
rect 94827 25556 94869 25565
rect 94827 25516 94828 25556
rect 94868 25516 94869 25556
rect 94827 25507 94869 25516
rect 95211 25556 95253 25565
rect 95211 25516 95212 25556
rect 95252 25516 95253 25556
rect 95211 25507 95253 25516
rect 96075 25556 96117 25565
rect 96075 25516 96076 25556
rect 96116 25516 96117 25556
rect 96075 25507 96117 25516
rect 96363 25556 96405 25565
rect 96363 25516 96364 25556
rect 96404 25516 96405 25556
rect 96363 25507 96405 25516
rect 96843 25556 96885 25565
rect 96843 25516 96844 25556
rect 96884 25516 96885 25556
rect 96843 25507 96885 25516
rect 97227 25556 97269 25565
rect 97227 25516 97228 25556
rect 97268 25516 97269 25556
rect 97227 25507 97269 25516
rect 97419 25556 97461 25565
rect 97419 25516 97420 25556
rect 97460 25516 97461 25556
rect 97419 25507 97461 25516
rect 97707 25556 97749 25565
rect 97707 25516 97708 25556
rect 97748 25516 97749 25556
rect 97707 25507 97749 25516
rect 98091 25556 98133 25565
rect 98091 25516 98092 25556
rect 98132 25516 98133 25556
rect 98091 25507 98133 25516
rect 98379 25556 98421 25565
rect 98379 25516 98380 25556
rect 98420 25516 98421 25556
rect 98379 25507 98421 25516
rect 98763 25556 98805 25565
rect 98763 25516 98764 25556
rect 98804 25516 98805 25556
rect 98763 25507 98805 25516
rect 74667 25472 74709 25481
rect 74667 25432 74668 25472
rect 74708 25432 74709 25472
rect 74667 25423 74709 25432
rect 75243 25472 75285 25481
rect 75243 25432 75244 25472
rect 75284 25432 75285 25472
rect 75243 25423 75285 25432
rect 76491 25472 76533 25481
rect 76491 25432 76492 25472
rect 76532 25432 76533 25472
rect 76491 25423 76533 25432
rect 77739 25472 77781 25481
rect 77739 25432 77740 25472
rect 77780 25432 77781 25472
rect 77739 25423 77781 25432
rect 83787 25472 83829 25481
rect 83787 25432 83788 25472
rect 83828 25432 83829 25472
rect 83787 25423 83829 25432
rect 87339 25472 87381 25481
rect 87339 25432 87340 25472
rect 87380 25432 87381 25472
rect 87339 25423 87381 25432
rect 89739 25472 89781 25481
rect 89739 25432 89740 25472
rect 89780 25432 89781 25472
rect 89739 25423 89781 25432
rect 72931 25388 72989 25389
rect 72931 25348 72940 25388
rect 72980 25348 72989 25388
rect 72931 25347 72989 25348
rect 73315 25388 73373 25389
rect 73315 25348 73324 25388
rect 73364 25348 73373 25388
rect 73315 25347 73373 25348
rect 73891 25388 73949 25389
rect 73891 25348 73900 25388
rect 73940 25348 73949 25388
rect 73891 25347 73949 25348
rect 74467 25388 74525 25389
rect 74467 25348 74476 25388
rect 74516 25348 74525 25388
rect 74467 25347 74525 25348
rect 74851 25388 74909 25389
rect 74851 25348 74860 25388
rect 74900 25348 74909 25388
rect 74851 25347 74909 25348
rect 75043 25388 75101 25389
rect 75043 25348 75052 25388
rect 75092 25348 75101 25388
rect 75043 25347 75101 25348
rect 75523 25388 75581 25389
rect 75523 25348 75532 25388
rect 75572 25348 75581 25388
rect 75523 25347 75581 25348
rect 77539 25388 77597 25389
rect 77539 25348 77548 25388
rect 77588 25348 77597 25388
rect 77539 25347 77597 25348
rect 83587 25388 83645 25389
rect 83587 25348 83596 25388
rect 83636 25348 83645 25388
rect 83587 25347 83645 25348
rect 87139 25388 87197 25389
rect 87139 25348 87148 25388
rect 87188 25348 87197 25388
rect 87139 25347 87197 25348
rect 89539 25388 89597 25389
rect 89539 25348 89548 25388
rect 89588 25348 89597 25388
rect 89539 25347 89597 25348
rect 95683 25388 95741 25389
rect 95683 25348 95692 25388
rect 95732 25348 95741 25388
rect 95683 25347 95741 25348
rect 98563 25388 98621 25389
rect 98563 25348 98572 25388
rect 98612 25348 98621 25388
rect 98563 25347 98621 25348
rect 643 25304 701 25305
rect 643 25264 652 25304
rect 692 25264 701 25304
rect 643 25263 701 25264
rect 835 25304 893 25305
rect 835 25264 844 25304
rect 884 25264 893 25304
rect 835 25263 893 25264
rect 72643 25304 72701 25305
rect 72643 25264 72652 25304
rect 72692 25264 72701 25304
rect 72643 25263 72701 25264
rect 76003 25304 76061 25305
rect 76003 25264 76012 25304
rect 76052 25264 76061 25304
rect 76003 25263 76061 25264
rect 76291 25304 76349 25305
rect 76291 25264 76300 25304
rect 76340 25264 76349 25304
rect 76291 25263 76349 25264
rect 76579 25304 76637 25305
rect 76579 25264 76588 25304
rect 76628 25264 76637 25304
rect 76579 25263 76637 25264
rect 76771 25304 76829 25305
rect 76771 25264 76780 25304
rect 76820 25264 76829 25304
rect 76771 25263 76829 25264
rect 77059 25304 77117 25305
rect 77059 25264 77068 25304
rect 77108 25264 77117 25304
rect 77059 25263 77117 25264
rect 78019 25304 78077 25305
rect 78019 25264 78028 25304
rect 78068 25264 78077 25304
rect 78019 25263 78077 25264
rect 78307 25304 78365 25305
rect 78307 25264 78316 25304
rect 78356 25264 78365 25304
rect 78307 25263 78365 25264
rect 78595 25304 78653 25305
rect 78595 25264 78604 25304
rect 78644 25264 78653 25304
rect 78595 25263 78653 25264
rect 78883 25304 78941 25305
rect 78883 25264 78892 25304
rect 78932 25264 78941 25304
rect 79843 25304 79901 25305
rect 78883 25263 78941 25264
rect 79070 25293 79112 25302
rect 79070 25253 79071 25293
rect 79111 25253 79112 25293
rect 79070 25244 79112 25253
rect 79459 25293 79517 25294
rect 79459 25253 79468 25293
rect 79508 25253 79517 25293
rect 79843 25264 79852 25304
rect 79892 25264 79901 25304
rect 79843 25263 79901 25264
rect 80035 25304 80093 25305
rect 80035 25264 80044 25304
rect 80084 25264 80093 25304
rect 80035 25263 80093 25264
rect 80419 25304 80477 25305
rect 80419 25264 80428 25304
rect 80468 25264 80477 25304
rect 81475 25304 81533 25305
rect 80419 25263 80477 25264
rect 80707 25293 80765 25294
rect 79459 25252 79517 25253
rect 80707 25253 80716 25293
rect 80756 25253 80765 25293
rect 80707 25252 80765 25253
rect 81091 25293 81149 25294
rect 81091 25253 81100 25293
rect 81140 25253 81149 25293
rect 81475 25264 81484 25304
rect 81524 25264 81533 25304
rect 81475 25263 81533 25264
rect 81955 25304 82013 25305
rect 81955 25264 81964 25304
rect 82004 25264 82013 25304
rect 82627 25304 82685 25305
rect 81955 25263 82013 25264
rect 82243 25293 82301 25294
rect 81091 25252 81149 25253
rect 82243 25253 82252 25293
rect 82292 25253 82301 25293
rect 82627 25264 82636 25304
rect 82676 25264 82685 25304
rect 82627 25263 82685 25264
rect 83203 25304 83261 25305
rect 83203 25264 83212 25304
rect 83252 25264 83261 25304
rect 83203 25263 83261 25264
rect 84067 25304 84125 25305
rect 84067 25264 84076 25304
rect 84116 25264 84125 25304
rect 84067 25263 84125 25264
rect 84355 25304 84413 25305
rect 84355 25264 84364 25304
rect 84404 25264 84413 25304
rect 84355 25263 84413 25264
rect 84643 25304 84701 25305
rect 84643 25264 84652 25304
rect 84692 25264 84701 25304
rect 84643 25263 84701 25264
rect 84931 25304 84989 25305
rect 84931 25264 84940 25304
rect 84980 25264 84989 25304
rect 84931 25263 84989 25264
rect 85123 25304 85181 25305
rect 85123 25264 85132 25304
rect 85172 25264 85181 25304
rect 85123 25263 85181 25264
rect 85507 25304 85565 25305
rect 85507 25264 85516 25304
rect 85556 25264 85565 25304
rect 85507 25263 85565 25264
rect 85891 25304 85949 25305
rect 85891 25264 85900 25304
rect 85940 25264 85949 25304
rect 85891 25263 85949 25264
rect 86467 25304 86525 25305
rect 86467 25264 86476 25304
rect 86516 25264 86525 25304
rect 86467 25263 86525 25264
rect 86755 25304 86813 25305
rect 86755 25264 86764 25304
rect 86804 25264 86813 25304
rect 86755 25263 86813 25264
rect 86947 25304 87005 25305
rect 86947 25264 86956 25304
rect 86996 25264 87005 25304
rect 86947 25263 87005 25264
rect 87619 25304 87677 25305
rect 87619 25264 87628 25304
rect 87668 25264 87677 25304
rect 87619 25263 87677 25264
rect 87907 25304 87965 25305
rect 87907 25264 87916 25304
rect 87956 25264 87965 25304
rect 87907 25263 87965 25264
rect 88195 25304 88253 25305
rect 88195 25264 88204 25304
rect 88244 25264 88253 25304
rect 88195 25263 88253 25264
rect 88483 25304 88541 25305
rect 88483 25264 88492 25304
rect 88532 25264 88541 25304
rect 88483 25263 88541 25264
rect 88675 25304 88733 25305
rect 88675 25264 88684 25304
rect 88724 25264 88733 25304
rect 88675 25263 88733 25264
rect 89059 25304 89117 25305
rect 89059 25264 89068 25304
rect 89108 25264 89117 25304
rect 89059 25263 89117 25264
rect 90019 25304 90077 25305
rect 90019 25264 90028 25304
rect 90068 25264 90077 25304
rect 90019 25263 90077 25264
rect 90307 25304 90365 25305
rect 90307 25264 90316 25304
rect 90356 25264 90365 25304
rect 90307 25263 90365 25264
rect 90595 25304 90653 25305
rect 90595 25264 90604 25304
rect 90644 25264 90653 25304
rect 90595 25263 90653 25264
rect 90883 25304 90941 25305
rect 90883 25264 90892 25304
rect 90932 25264 90941 25304
rect 90883 25263 90941 25264
rect 91267 25304 91325 25305
rect 91267 25264 91276 25304
rect 91316 25264 91325 25304
rect 91939 25304 91997 25305
rect 91267 25263 91325 25264
rect 91454 25293 91496 25302
rect 82243 25252 82301 25253
rect 91454 25253 91455 25293
rect 91495 25253 91496 25293
rect 91939 25264 91948 25304
rect 91988 25264 91997 25304
rect 91939 25263 91997 25264
rect 92323 25304 92381 25305
rect 92323 25264 92332 25304
rect 92372 25264 92381 25304
rect 92323 25263 92381 25264
rect 92515 25304 92573 25305
rect 92515 25264 92524 25304
rect 92564 25264 92573 25304
rect 92515 25263 92573 25264
rect 92899 25304 92957 25305
rect 92899 25264 92908 25304
rect 92948 25264 92957 25304
rect 93667 25304 93725 25305
rect 92899 25263 92957 25264
rect 93086 25293 93128 25302
rect 91454 25244 91496 25253
rect 93086 25253 93087 25293
rect 93127 25253 93128 25293
rect 93667 25264 93676 25304
rect 93716 25264 93725 25304
rect 93667 25263 93725 25264
rect 93955 25304 94013 25305
rect 93955 25264 93964 25304
rect 94004 25264 94013 25304
rect 94915 25304 94973 25305
rect 93955 25263 94013 25264
rect 94243 25293 94301 25294
rect 93086 25244 93128 25253
rect 94243 25253 94252 25293
rect 94292 25253 94301 25293
rect 94915 25264 94924 25304
rect 94964 25264 94973 25304
rect 94915 25263 94973 25264
rect 95299 25304 95357 25305
rect 95299 25264 95308 25304
rect 95348 25264 95357 25304
rect 95299 25263 95357 25264
rect 96163 25304 96221 25305
rect 96163 25264 96172 25304
rect 96212 25264 96221 25304
rect 96163 25263 96221 25264
rect 96451 25304 96509 25305
rect 96451 25264 96460 25304
rect 96500 25264 96509 25304
rect 96451 25263 96509 25264
rect 96739 25304 96797 25305
rect 96739 25264 96748 25304
rect 96788 25264 96797 25304
rect 97507 25304 97565 25305
rect 96739 25263 96797 25264
rect 97118 25293 97176 25294
rect 94243 25252 94301 25253
rect 97118 25253 97127 25293
rect 97167 25253 97176 25293
rect 97507 25264 97516 25304
rect 97556 25264 97565 25304
rect 97507 25263 97565 25264
rect 97795 25304 97853 25305
rect 97795 25264 97804 25304
rect 97844 25264 97853 25304
rect 97795 25263 97853 25264
rect 97987 25304 98045 25305
rect 97987 25264 97996 25304
rect 98036 25264 98045 25304
rect 97987 25263 98045 25264
rect 98851 25304 98909 25305
rect 98851 25264 98860 25304
rect 98900 25264 98909 25304
rect 98851 25263 98909 25264
rect 97118 25252 97176 25253
rect 74283 25136 74325 25145
rect 74283 25096 74284 25136
rect 74324 25096 74325 25136
rect 74283 25087 74325 25096
rect 95883 25136 95925 25145
rect 95883 25096 95884 25136
rect 95924 25096 95925 25136
rect 95883 25087 95925 25096
rect 576 24968 99360 24992
rect 576 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 8352 24968
rect 8392 24928 8434 24968
rect 8474 24928 8516 24968
rect 8556 24928 8598 24968
rect 8638 24928 8680 24968
rect 8720 24928 12352 24968
rect 12392 24928 12434 24968
rect 12474 24928 12516 24968
rect 12556 24928 12598 24968
rect 12638 24928 12680 24968
rect 12720 24928 16352 24968
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16720 24928 20352 24968
rect 20392 24928 20434 24968
rect 20474 24928 20516 24968
rect 20556 24928 20598 24968
rect 20638 24928 20680 24968
rect 20720 24928 24352 24968
rect 24392 24928 24434 24968
rect 24474 24928 24516 24968
rect 24556 24928 24598 24968
rect 24638 24928 24680 24968
rect 24720 24928 28352 24968
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28720 24928 32352 24968
rect 32392 24928 32434 24968
rect 32474 24928 32516 24968
rect 32556 24928 32598 24968
rect 32638 24928 32680 24968
rect 32720 24928 36352 24968
rect 36392 24928 36434 24968
rect 36474 24928 36516 24968
rect 36556 24928 36598 24968
rect 36638 24928 36680 24968
rect 36720 24928 40352 24968
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40720 24928 44352 24968
rect 44392 24928 44434 24968
rect 44474 24928 44516 24968
rect 44556 24928 44598 24968
rect 44638 24928 44680 24968
rect 44720 24928 48352 24968
rect 48392 24928 48434 24968
rect 48474 24928 48516 24968
rect 48556 24928 48598 24968
rect 48638 24928 48680 24968
rect 48720 24928 52352 24968
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52720 24928 56352 24968
rect 56392 24928 56434 24968
rect 56474 24928 56516 24968
rect 56556 24928 56598 24968
rect 56638 24928 56680 24968
rect 56720 24928 60352 24968
rect 60392 24928 60434 24968
rect 60474 24928 60516 24968
rect 60556 24928 60598 24968
rect 60638 24928 60680 24968
rect 60720 24928 64352 24968
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64720 24928 68352 24968
rect 68392 24928 68434 24968
rect 68474 24928 68516 24968
rect 68556 24928 68598 24968
rect 68638 24928 68680 24968
rect 68720 24928 99360 24968
rect 576 24904 99360 24928
rect 73323 24800 73365 24809
rect 73323 24760 73324 24800
rect 73364 24760 73365 24800
rect 73323 24751 73365 24760
rect 73515 24800 73557 24809
rect 73515 24760 73516 24800
rect 73556 24760 73557 24800
rect 73515 24751 73557 24760
rect 73995 24800 74037 24809
rect 73995 24760 73996 24800
rect 74036 24760 74037 24800
rect 73995 24751 74037 24760
rect 74859 24800 74901 24809
rect 74859 24760 74860 24800
rect 74900 24760 74901 24800
rect 74859 24751 74901 24760
rect 75435 24800 75477 24809
rect 75435 24760 75436 24800
rect 75476 24760 75477 24800
rect 75435 24751 75477 24760
rect 75627 24800 75669 24809
rect 75627 24760 75628 24800
rect 75668 24760 75669 24800
rect 75627 24751 75669 24760
rect 76203 24800 76245 24809
rect 76203 24760 76204 24800
rect 76244 24760 76245 24800
rect 76203 24751 76245 24760
rect 76587 24800 76629 24809
rect 76587 24760 76588 24800
rect 76628 24760 76629 24800
rect 76587 24751 76629 24760
rect 77067 24800 77109 24809
rect 77067 24760 77068 24800
rect 77108 24760 77109 24800
rect 77067 24751 77109 24760
rect 77451 24800 77493 24809
rect 77451 24760 77452 24800
rect 77492 24760 77493 24800
rect 77451 24751 77493 24760
rect 78027 24800 78069 24809
rect 78027 24760 78028 24800
rect 78068 24760 78069 24800
rect 78027 24751 78069 24760
rect 78411 24800 78453 24809
rect 78411 24760 78412 24800
rect 78452 24760 78453 24800
rect 78411 24751 78453 24760
rect 78795 24800 78837 24809
rect 78795 24760 78796 24800
rect 78836 24760 78837 24800
rect 78795 24751 78837 24760
rect 79179 24800 79221 24809
rect 79179 24760 79180 24800
rect 79220 24760 79221 24800
rect 79179 24751 79221 24760
rect 79563 24800 79605 24809
rect 79563 24760 79564 24800
rect 79604 24760 79605 24800
rect 79563 24751 79605 24760
rect 79947 24800 79989 24809
rect 79947 24760 79948 24800
rect 79988 24760 79989 24800
rect 79947 24751 79989 24760
rect 81195 24800 81237 24809
rect 81195 24760 81196 24800
rect 81236 24760 81237 24800
rect 81195 24751 81237 24760
rect 81579 24800 81621 24809
rect 81579 24760 81580 24800
rect 81620 24760 81621 24800
rect 81579 24751 81621 24760
rect 81963 24800 82005 24809
rect 81963 24760 81964 24800
rect 82004 24760 82005 24800
rect 81963 24751 82005 24760
rect 82347 24800 82389 24809
rect 82347 24760 82348 24800
rect 82388 24760 82389 24800
rect 82347 24751 82389 24760
rect 83115 24800 83157 24809
rect 83115 24760 83116 24800
rect 83156 24760 83157 24800
rect 83115 24751 83157 24760
rect 83499 24800 83541 24809
rect 83499 24760 83500 24800
rect 83540 24760 83541 24800
rect 83499 24751 83541 24760
rect 83883 24800 83925 24809
rect 83883 24760 83884 24800
rect 83924 24760 83925 24800
rect 83883 24751 83925 24760
rect 84459 24800 84501 24809
rect 84459 24760 84460 24800
rect 84500 24760 84501 24800
rect 84459 24751 84501 24760
rect 84843 24800 84885 24809
rect 84843 24760 84844 24800
rect 84884 24760 84885 24800
rect 84843 24751 84885 24760
rect 85515 24800 85557 24809
rect 85515 24760 85516 24800
rect 85556 24760 85557 24800
rect 85515 24751 85557 24760
rect 86283 24800 86325 24809
rect 86283 24760 86284 24800
rect 86324 24760 86325 24800
rect 86283 24751 86325 24760
rect 87147 24800 87189 24809
rect 87147 24760 87148 24800
rect 87188 24760 87189 24800
rect 87147 24751 87189 24760
rect 87531 24800 87573 24809
rect 87531 24760 87532 24800
rect 87572 24760 87573 24800
rect 87531 24751 87573 24760
rect 88299 24800 88341 24809
rect 88299 24760 88300 24800
rect 88340 24760 88341 24800
rect 88299 24751 88341 24760
rect 88683 24800 88725 24809
rect 88683 24760 88684 24800
rect 88724 24760 88725 24800
rect 88683 24751 88725 24760
rect 89451 24800 89493 24809
rect 89451 24760 89452 24800
rect 89492 24760 89493 24800
rect 89451 24751 89493 24760
rect 89931 24800 89973 24809
rect 89931 24760 89932 24800
rect 89972 24760 89973 24800
rect 89931 24751 89973 24760
rect 90315 24800 90357 24809
rect 90315 24760 90316 24800
rect 90356 24760 90357 24800
rect 90315 24751 90357 24760
rect 90699 24800 90741 24809
rect 90699 24760 90700 24800
rect 90740 24760 90741 24800
rect 90699 24751 90741 24760
rect 91179 24800 91221 24809
rect 91179 24760 91180 24800
rect 91220 24760 91221 24800
rect 91179 24751 91221 24760
rect 91851 24800 91893 24809
rect 91851 24760 91852 24800
rect 91892 24760 91893 24800
rect 91851 24751 91893 24760
rect 92139 24800 92181 24809
rect 92139 24760 92140 24800
rect 92180 24760 92181 24800
rect 92139 24751 92181 24760
rect 92907 24800 92949 24809
rect 92907 24760 92908 24800
rect 92948 24760 92949 24800
rect 92907 24751 92949 24760
rect 93291 24800 93333 24809
rect 93291 24760 93292 24800
rect 93332 24760 93333 24800
rect 93291 24751 93333 24760
rect 93963 24800 94005 24809
rect 93963 24760 93964 24800
rect 94004 24760 94005 24800
rect 93963 24751 94005 24760
rect 94347 24800 94389 24809
rect 94347 24760 94348 24800
rect 94388 24760 94389 24800
rect 94347 24751 94389 24760
rect 94731 24800 94773 24809
rect 94731 24760 94732 24800
rect 94772 24760 94773 24800
rect 94731 24751 94773 24760
rect 95115 24800 95157 24809
rect 95115 24760 95116 24800
rect 95156 24760 95157 24800
rect 95115 24751 95157 24760
rect 95595 24800 95637 24809
rect 95595 24760 95596 24800
rect 95636 24760 95637 24800
rect 95595 24751 95637 24760
rect 95979 24800 96021 24809
rect 95979 24760 95980 24800
rect 96020 24760 96021 24800
rect 95979 24751 96021 24760
rect 96171 24800 96213 24809
rect 96171 24760 96172 24800
rect 96212 24760 96213 24800
rect 96171 24751 96213 24760
rect 96555 24800 96597 24809
rect 96555 24760 96556 24800
rect 96596 24760 96597 24800
rect 96555 24751 96597 24760
rect 96939 24800 96981 24809
rect 96939 24760 96940 24800
rect 96980 24760 96981 24800
rect 96939 24751 96981 24760
rect 97323 24800 97365 24809
rect 97323 24760 97324 24800
rect 97364 24760 97365 24800
rect 97323 24751 97365 24760
rect 97707 24800 97749 24809
rect 97707 24760 97708 24800
rect 97748 24760 97749 24800
rect 97707 24751 97749 24760
rect 98091 24800 98133 24809
rect 98091 24760 98092 24800
rect 98132 24760 98133 24800
rect 98091 24751 98133 24760
rect 643 24632 701 24633
rect 643 24592 652 24632
rect 692 24592 701 24632
rect 643 24591 701 24592
rect 835 24632 893 24633
rect 835 24592 844 24632
rect 884 24592 893 24632
rect 835 24591 893 24592
rect 73219 24632 73277 24633
rect 73219 24592 73228 24632
rect 73268 24592 73277 24632
rect 73219 24591 73277 24592
rect 73603 24632 73661 24633
rect 73603 24592 73612 24632
rect 73652 24592 73661 24632
rect 73603 24591 73661 24592
rect 75715 24632 75773 24633
rect 75715 24592 75724 24632
rect 75764 24592 75773 24632
rect 75715 24591 75773 24592
rect 80419 24632 80477 24633
rect 80419 24592 80428 24632
rect 80468 24592 80477 24632
rect 80419 24591 80477 24592
rect 80611 24632 80669 24633
rect 80611 24592 80620 24632
rect 80660 24592 80669 24632
rect 80611 24591 80669 24592
rect 87723 24632 87765 24641
rect 87723 24592 87724 24632
rect 87764 24592 87765 24632
rect 87723 24583 87765 24592
rect 87811 24632 87869 24633
rect 87811 24592 87820 24632
rect 87860 24592 87869 24632
rect 87811 24591 87869 24592
rect 73795 24548 73853 24549
rect 73795 24508 73804 24548
rect 73844 24508 73853 24548
rect 73795 24507 73853 24508
rect 74179 24548 74237 24549
rect 74179 24508 74188 24548
rect 74228 24508 74237 24548
rect 74179 24507 74237 24508
rect 74659 24548 74717 24549
rect 74659 24508 74668 24548
rect 74708 24508 74717 24548
rect 74659 24507 74717 24508
rect 75235 24548 75293 24549
rect 75235 24508 75244 24548
rect 75284 24508 75293 24548
rect 75235 24507 75293 24508
rect 76003 24548 76061 24549
rect 76003 24508 76012 24548
rect 76052 24508 76061 24548
rect 76003 24507 76061 24508
rect 76387 24548 76445 24549
rect 76387 24508 76396 24548
rect 76436 24508 76445 24548
rect 76387 24507 76445 24508
rect 76867 24548 76925 24549
rect 76867 24508 76876 24548
rect 76916 24508 76925 24548
rect 76867 24507 76925 24508
rect 77251 24548 77309 24549
rect 77251 24508 77260 24548
rect 77300 24508 77309 24548
rect 77251 24507 77309 24508
rect 77635 24548 77693 24549
rect 77635 24508 77644 24548
rect 77684 24508 77693 24548
rect 77635 24507 77693 24508
rect 78211 24548 78269 24549
rect 78211 24508 78220 24548
rect 78260 24508 78269 24548
rect 78211 24507 78269 24508
rect 78595 24548 78653 24549
rect 78595 24508 78604 24548
rect 78644 24508 78653 24548
rect 78595 24507 78653 24508
rect 78979 24548 79037 24549
rect 78979 24508 78988 24548
rect 79028 24508 79037 24548
rect 78979 24507 79037 24508
rect 79363 24548 79421 24549
rect 79363 24508 79372 24548
rect 79412 24508 79421 24548
rect 79363 24507 79421 24508
rect 79747 24548 79805 24549
rect 79747 24508 79756 24548
rect 79796 24508 79805 24548
rect 79747 24507 79805 24508
rect 80131 24548 80189 24549
rect 80131 24508 80140 24548
rect 80180 24508 80189 24548
rect 80131 24507 80189 24508
rect 80995 24548 81053 24549
rect 80995 24508 81004 24548
rect 81044 24508 81053 24548
rect 80995 24507 81053 24508
rect 81379 24548 81437 24549
rect 81379 24508 81388 24548
rect 81428 24508 81437 24548
rect 81379 24507 81437 24508
rect 81763 24548 81821 24549
rect 81763 24508 81772 24548
rect 81812 24508 81821 24548
rect 81763 24507 81821 24508
rect 82147 24548 82205 24549
rect 82147 24508 82156 24548
rect 82196 24508 82205 24548
rect 82147 24507 82205 24508
rect 82531 24548 82589 24549
rect 82531 24508 82540 24548
rect 82580 24508 82589 24548
rect 82531 24507 82589 24508
rect 82915 24548 82973 24549
rect 82915 24508 82924 24548
rect 82964 24508 82973 24548
rect 82915 24507 82973 24508
rect 83299 24548 83357 24549
rect 83299 24508 83308 24548
rect 83348 24508 83357 24548
rect 83299 24507 83357 24508
rect 83683 24548 83741 24549
rect 83683 24508 83692 24548
rect 83732 24508 83741 24548
rect 83683 24507 83741 24508
rect 84067 24548 84125 24549
rect 84067 24508 84076 24548
rect 84116 24508 84125 24548
rect 84067 24507 84125 24508
rect 84643 24548 84701 24549
rect 84643 24508 84652 24548
rect 84692 24508 84701 24548
rect 84643 24507 84701 24508
rect 85027 24548 85085 24549
rect 85027 24508 85036 24548
rect 85076 24508 85085 24548
rect 85027 24507 85085 24508
rect 85315 24548 85373 24549
rect 85315 24508 85324 24548
rect 85364 24508 85373 24548
rect 85315 24507 85373 24508
rect 86083 24548 86141 24549
rect 86083 24508 86092 24548
rect 86132 24508 86141 24548
rect 86083 24507 86141 24508
rect 86563 24548 86621 24549
rect 86563 24508 86572 24548
rect 86612 24508 86621 24548
rect 86563 24507 86621 24508
rect 86947 24548 87005 24549
rect 86947 24508 86956 24548
rect 86996 24508 87005 24548
rect 86947 24507 87005 24508
rect 87331 24548 87389 24549
rect 87331 24508 87340 24548
rect 87380 24508 87389 24548
rect 87331 24507 87389 24508
rect 88099 24548 88157 24549
rect 88099 24508 88108 24548
rect 88148 24508 88157 24548
rect 88099 24507 88157 24508
rect 88483 24548 88541 24549
rect 88483 24508 88492 24548
rect 88532 24508 88541 24548
rect 88483 24507 88541 24508
rect 88867 24548 88925 24549
rect 88867 24508 88876 24548
rect 88916 24508 88925 24548
rect 88867 24507 88925 24508
rect 89251 24548 89309 24549
rect 89251 24508 89260 24548
rect 89300 24508 89309 24548
rect 89251 24507 89309 24508
rect 89731 24548 89789 24549
rect 89731 24508 89740 24548
rect 89780 24508 89789 24548
rect 89731 24507 89789 24508
rect 90115 24548 90173 24549
rect 90115 24508 90124 24548
rect 90164 24508 90173 24548
rect 90115 24507 90173 24508
rect 90499 24548 90557 24549
rect 90499 24508 90508 24548
rect 90548 24508 90557 24548
rect 90499 24507 90557 24508
rect 90979 24548 91037 24549
rect 90979 24508 90988 24548
rect 91028 24508 91037 24548
rect 90979 24507 91037 24508
rect 91651 24548 91709 24549
rect 91651 24508 91660 24548
rect 91700 24508 91709 24548
rect 91651 24507 91709 24508
rect 92323 24548 92381 24549
rect 92323 24508 92332 24548
rect 92372 24508 92381 24548
rect 92323 24507 92381 24508
rect 92707 24548 92765 24549
rect 92707 24508 92716 24548
rect 92756 24508 92765 24548
rect 92707 24507 92765 24508
rect 93091 24548 93149 24549
rect 93091 24508 93100 24548
rect 93140 24508 93149 24548
rect 93091 24507 93149 24508
rect 93475 24548 93533 24549
rect 93475 24508 93484 24548
rect 93524 24508 93533 24548
rect 93475 24507 93533 24508
rect 93763 24548 93821 24549
rect 93763 24508 93772 24548
rect 93812 24508 93821 24548
rect 93763 24507 93821 24508
rect 94147 24548 94205 24549
rect 94147 24508 94156 24548
rect 94196 24508 94205 24548
rect 94147 24507 94205 24508
rect 94531 24548 94589 24549
rect 94531 24508 94540 24548
rect 94580 24508 94589 24548
rect 94531 24507 94589 24508
rect 94915 24548 94973 24549
rect 94915 24508 94924 24548
rect 94964 24508 94973 24548
rect 94915 24507 94973 24508
rect 95395 24548 95453 24549
rect 95395 24508 95404 24548
rect 95444 24508 95453 24548
rect 95395 24507 95453 24508
rect 95779 24548 95837 24549
rect 95779 24508 95788 24548
rect 95828 24508 95837 24548
rect 95779 24507 95837 24508
rect 96355 24548 96413 24549
rect 96355 24508 96364 24548
rect 96404 24508 96413 24548
rect 96355 24507 96413 24508
rect 96739 24548 96797 24549
rect 96739 24508 96748 24548
rect 96788 24508 96797 24548
rect 96739 24507 96797 24508
rect 97123 24548 97181 24549
rect 97123 24508 97132 24548
rect 97172 24508 97181 24548
rect 97123 24507 97181 24508
rect 97507 24548 97565 24549
rect 97507 24508 97516 24548
rect 97556 24508 97565 24548
rect 97507 24507 97565 24508
rect 97891 24548 97949 24549
rect 97891 24508 97900 24548
rect 97940 24508 97949 24548
rect 97891 24507 97949 24508
rect 98275 24548 98333 24549
rect 98275 24508 98284 24548
rect 98324 24508 98333 24548
rect 98275 24507 98333 24508
rect 77835 24464 77877 24473
rect 77835 24424 77836 24464
rect 77876 24424 77877 24464
rect 77835 24415 77877 24424
rect 84267 24464 84309 24473
rect 84267 24424 84268 24464
rect 84308 24424 84309 24464
rect 84267 24415 84309 24424
rect 86763 24464 86805 24473
rect 86763 24424 86764 24464
rect 86804 24424 86805 24464
rect 86763 24415 86805 24424
rect 89067 24464 89109 24473
rect 89067 24424 89068 24464
rect 89108 24424 89109 24464
rect 89067 24415 89109 24424
rect 92523 24464 92565 24473
rect 92523 24424 92524 24464
rect 92564 24424 92565 24464
rect 92523 24415 92565 24424
rect 74379 24380 74421 24389
rect 74379 24340 74380 24380
rect 74420 24340 74421 24380
rect 74379 24331 74421 24340
rect 80811 24380 80853 24389
rect 80811 24340 80812 24380
rect 80852 24340 80853 24380
rect 80811 24331 80853 24340
rect 576 24212 99516 24236
rect 576 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 7112 24212
rect 7152 24172 7194 24212
rect 7234 24172 7276 24212
rect 7316 24172 7358 24212
rect 7398 24172 7440 24212
rect 7480 24172 11112 24212
rect 11152 24172 11194 24212
rect 11234 24172 11276 24212
rect 11316 24172 11358 24212
rect 11398 24172 11440 24212
rect 11480 24172 15112 24212
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15480 24172 19112 24212
rect 19152 24172 19194 24212
rect 19234 24172 19276 24212
rect 19316 24172 19358 24212
rect 19398 24172 19440 24212
rect 19480 24172 23112 24212
rect 23152 24172 23194 24212
rect 23234 24172 23276 24212
rect 23316 24172 23358 24212
rect 23398 24172 23440 24212
rect 23480 24172 27112 24212
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27480 24172 31112 24212
rect 31152 24172 31194 24212
rect 31234 24172 31276 24212
rect 31316 24172 31358 24212
rect 31398 24172 31440 24212
rect 31480 24172 35112 24212
rect 35152 24172 35194 24212
rect 35234 24172 35276 24212
rect 35316 24172 35358 24212
rect 35398 24172 35440 24212
rect 35480 24172 39112 24212
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39480 24172 43112 24212
rect 43152 24172 43194 24212
rect 43234 24172 43276 24212
rect 43316 24172 43358 24212
rect 43398 24172 43440 24212
rect 43480 24172 47112 24212
rect 47152 24172 47194 24212
rect 47234 24172 47276 24212
rect 47316 24172 47358 24212
rect 47398 24172 47440 24212
rect 47480 24172 51112 24212
rect 51152 24172 51194 24212
rect 51234 24172 51276 24212
rect 51316 24172 51358 24212
rect 51398 24172 51440 24212
rect 51480 24172 55112 24212
rect 55152 24172 55194 24212
rect 55234 24172 55276 24212
rect 55316 24172 55358 24212
rect 55398 24172 55440 24212
rect 55480 24172 59112 24212
rect 59152 24172 59194 24212
rect 59234 24172 59276 24212
rect 59316 24172 59358 24212
rect 59398 24172 59440 24212
rect 59480 24172 63112 24212
rect 63152 24172 63194 24212
rect 63234 24172 63276 24212
rect 63316 24172 63358 24212
rect 63398 24172 63440 24212
rect 63480 24172 67112 24212
rect 67152 24172 67194 24212
rect 67234 24172 67276 24212
rect 67316 24172 67358 24212
rect 67398 24172 67440 24212
rect 67480 24172 71112 24212
rect 71152 24172 71194 24212
rect 71234 24172 71276 24212
rect 71316 24172 71358 24212
rect 71398 24172 71440 24212
rect 71480 24172 75112 24212
rect 75152 24172 75194 24212
rect 75234 24172 75276 24212
rect 75316 24172 75358 24212
rect 75398 24172 75440 24212
rect 75480 24172 79112 24212
rect 79152 24172 79194 24212
rect 79234 24172 79276 24212
rect 79316 24172 79358 24212
rect 79398 24172 79440 24212
rect 79480 24172 83112 24212
rect 83152 24172 83194 24212
rect 83234 24172 83276 24212
rect 83316 24172 83358 24212
rect 83398 24172 83440 24212
rect 83480 24172 87112 24212
rect 87152 24172 87194 24212
rect 87234 24172 87276 24212
rect 87316 24172 87358 24212
rect 87398 24172 87440 24212
rect 87480 24172 91112 24212
rect 91152 24172 91194 24212
rect 91234 24172 91276 24212
rect 91316 24172 91358 24212
rect 91398 24172 91440 24212
rect 91480 24172 95112 24212
rect 95152 24172 95194 24212
rect 95234 24172 95276 24212
rect 95316 24172 95358 24212
rect 95398 24172 95440 24212
rect 95480 24172 99112 24212
rect 99152 24172 99194 24212
rect 99234 24172 99276 24212
rect 99316 24172 99358 24212
rect 99398 24172 99440 24212
rect 99480 24172 99516 24212
rect 576 24148 99516 24172
rect 81867 24044 81909 24053
rect 81867 24004 81868 24044
rect 81908 24004 81909 24044
rect 81867 23995 81909 24004
rect 80139 23960 80181 23969
rect 80139 23920 80140 23960
rect 80180 23920 80181 23960
rect 80139 23911 80181 23920
rect 82635 23960 82677 23969
rect 82635 23920 82636 23960
rect 82676 23920 82677 23960
rect 82635 23911 82677 23920
rect 85131 23960 85173 23969
rect 85131 23920 85132 23960
rect 85172 23920 85173 23960
rect 85131 23911 85173 23920
rect 85899 23960 85941 23969
rect 85899 23920 85900 23960
rect 85940 23920 85941 23960
rect 85899 23911 85941 23920
rect 86667 23960 86709 23969
rect 86667 23920 86668 23960
rect 86708 23920 86709 23960
rect 86667 23911 86709 23920
rect 87915 23960 87957 23969
rect 87915 23920 87916 23960
rect 87956 23920 87957 23960
rect 87915 23911 87957 23920
rect 89067 23960 89109 23969
rect 89067 23920 89068 23960
rect 89108 23920 89109 23960
rect 89067 23911 89109 23920
rect 91467 23960 91509 23969
rect 91467 23920 91468 23960
rect 91508 23920 91509 23960
rect 91467 23911 91509 23920
rect 92427 23960 92469 23969
rect 92427 23920 92428 23960
rect 92468 23920 92469 23960
rect 92427 23911 92469 23920
rect 93579 23960 93621 23969
rect 93579 23920 93580 23960
rect 93620 23920 93621 23960
rect 93579 23911 93621 23920
rect 80323 23876 80381 23877
rect 80323 23836 80332 23876
rect 80372 23836 80381 23876
rect 80323 23835 80381 23836
rect 81667 23876 81725 23877
rect 81667 23836 81676 23876
rect 81716 23836 81725 23876
rect 81667 23835 81725 23836
rect 82435 23876 82493 23877
rect 82435 23836 82444 23876
rect 82484 23836 82493 23876
rect 82435 23835 82493 23836
rect 84931 23876 84989 23877
rect 84931 23836 84940 23876
rect 84980 23836 84989 23876
rect 84931 23835 84989 23836
rect 85699 23876 85757 23877
rect 85699 23836 85708 23876
rect 85748 23836 85757 23876
rect 85699 23835 85757 23836
rect 86467 23876 86525 23877
rect 86467 23836 86476 23876
rect 86516 23836 86525 23876
rect 86467 23835 86525 23836
rect 87715 23876 87773 23877
rect 87715 23836 87724 23876
rect 87764 23836 87773 23876
rect 87715 23835 87773 23836
rect 88867 23876 88925 23877
rect 88867 23836 88876 23876
rect 88916 23836 88925 23876
rect 88867 23835 88925 23836
rect 91267 23876 91325 23877
rect 91267 23836 91276 23876
rect 91316 23836 91325 23876
rect 91267 23835 91325 23836
rect 93379 23876 93437 23877
rect 93379 23836 93388 23876
rect 93428 23836 93437 23876
rect 93379 23835 93437 23836
rect 643 23792 701 23793
rect 643 23752 652 23792
rect 692 23752 701 23792
rect 643 23751 701 23752
rect 835 23792 893 23793
rect 835 23752 844 23792
rect 884 23752 893 23792
rect 835 23751 893 23752
rect 92323 23792 92381 23793
rect 92323 23752 92332 23792
rect 92372 23752 92381 23792
rect 92323 23751 92381 23752
rect 576 23456 99360 23480
rect 576 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 8352 23456
rect 8392 23416 8434 23456
rect 8474 23416 8516 23456
rect 8556 23416 8598 23456
rect 8638 23416 8680 23456
rect 8720 23416 12352 23456
rect 12392 23416 12434 23456
rect 12474 23416 12516 23456
rect 12556 23416 12598 23456
rect 12638 23416 12680 23456
rect 12720 23416 16352 23456
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16720 23416 20352 23456
rect 20392 23416 20434 23456
rect 20474 23416 20516 23456
rect 20556 23416 20598 23456
rect 20638 23416 20680 23456
rect 20720 23416 24352 23456
rect 24392 23416 24434 23456
rect 24474 23416 24516 23456
rect 24556 23416 24598 23456
rect 24638 23416 24680 23456
rect 24720 23416 28352 23456
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28720 23416 32352 23456
rect 32392 23416 32434 23456
rect 32474 23416 32516 23456
rect 32556 23416 32598 23456
rect 32638 23416 32680 23456
rect 32720 23416 36352 23456
rect 36392 23416 36434 23456
rect 36474 23416 36516 23456
rect 36556 23416 36598 23456
rect 36638 23416 36680 23456
rect 36720 23416 40352 23456
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40720 23416 44352 23456
rect 44392 23416 44434 23456
rect 44474 23416 44516 23456
rect 44556 23416 44598 23456
rect 44638 23416 44680 23456
rect 44720 23416 48352 23456
rect 48392 23416 48434 23456
rect 48474 23416 48516 23456
rect 48556 23416 48598 23456
rect 48638 23416 48680 23456
rect 48720 23416 52352 23456
rect 52392 23416 52434 23456
rect 52474 23416 52516 23456
rect 52556 23416 52598 23456
rect 52638 23416 52680 23456
rect 52720 23416 56352 23456
rect 56392 23416 56434 23456
rect 56474 23416 56516 23456
rect 56556 23416 56598 23456
rect 56638 23416 56680 23456
rect 56720 23416 60352 23456
rect 60392 23416 60434 23456
rect 60474 23416 60516 23456
rect 60556 23416 60598 23456
rect 60638 23416 60680 23456
rect 60720 23416 64352 23456
rect 64392 23416 64434 23456
rect 64474 23416 64516 23456
rect 64556 23416 64598 23456
rect 64638 23416 64680 23456
rect 64720 23416 68352 23456
rect 68392 23416 68434 23456
rect 68474 23416 68516 23456
rect 68556 23416 68598 23456
rect 68638 23416 68680 23456
rect 68720 23416 72352 23456
rect 72392 23416 72434 23456
rect 72474 23416 72516 23456
rect 72556 23416 72598 23456
rect 72638 23416 72680 23456
rect 72720 23416 76352 23456
rect 76392 23416 76434 23456
rect 76474 23416 76516 23456
rect 76556 23416 76598 23456
rect 76638 23416 76680 23456
rect 76720 23416 80352 23456
rect 80392 23416 80434 23456
rect 80474 23416 80516 23456
rect 80556 23416 80598 23456
rect 80638 23416 80680 23456
rect 80720 23416 84352 23456
rect 84392 23416 84434 23456
rect 84474 23416 84516 23456
rect 84556 23416 84598 23456
rect 84638 23416 84680 23456
rect 84720 23416 88352 23456
rect 88392 23416 88434 23456
rect 88474 23416 88516 23456
rect 88556 23416 88598 23456
rect 88638 23416 88680 23456
rect 88720 23416 92352 23456
rect 92392 23416 92434 23456
rect 92474 23416 92516 23456
rect 92556 23416 92598 23456
rect 92638 23416 92680 23456
rect 92720 23416 96352 23456
rect 96392 23416 96434 23456
rect 96474 23416 96516 23456
rect 96556 23416 96598 23456
rect 96638 23416 96680 23456
rect 96720 23416 99360 23456
rect 576 23392 99360 23416
rect 643 23120 701 23121
rect 643 23080 652 23120
rect 692 23080 701 23120
rect 643 23079 701 23080
rect 835 23120 893 23121
rect 835 23080 844 23120
rect 884 23080 893 23120
rect 835 23079 893 23080
rect 576 22700 99516 22724
rect 576 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 7112 22700
rect 7152 22660 7194 22700
rect 7234 22660 7276 22700
rect 7316 22660 7358 22700
rect 7398 22660 7440 22700
rect 7480 22660 11112 22700
rect 11152 22660 11194 22700
rect 11234 22660 11276 22700
rect 11316 22660 11358 22700
rect 11398 22660 11440 22700
rect 11480 22660 15112 22700
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15480 22660 19112 22700
rect 19152 22660 19194 22700
rect 19234 22660 19276 22700
rect 19316 22660 19358 22700
rect 19398 22660 19440 22700
rect 19480 22660 23112 22700
rect 23152 22660 23194 22700
rect 23234 22660 23276 22700
rect 23316 22660 23358 22700
rect 23398 22660 23440 22700
rect 23480 22660 27112 22700
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27480 22660 31112 22700
rect 31152 22660 31194 22700
rect 31234 22660 31276 22700
rect 31316 22660 31358 22700
rect 31398 22660 31440 22700
rect 31480 22660 35112 22700
rect 35152 22660 35194 22700
rect 35234 22660 35276 22700
rect 35316 22660 35358 22700
rect 35398 22660 35440 22700
rect 35480 22660 39112 22700
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39480 22660 43112 22700
rect 43152 22660 43194 22700
rect 43234 22660 43276 22700
rect 43316 22660 43358 22700
rect 43398 22660 43440 22700
rect 43480 22660 47112 22700
rect 47152 22660 47194 22700
rect 47234 22660 47276 22700
rect 47316 22660 47358 22700
rect 47398 22660 47440 22700
rect 47480 22660 51112 22700
rect 51152 22660 51194 22700
rect 51234 22660 51276 22700
rect 51316 22660 51358 22700
rect 51398 22660 51440 22700
rect 51480 22660 55112 22700
rect 55152 22660 55194 22700
rect 55234 22660 55276 22700
rect 55316 22660 55358 22700
rect 55398 22660 55440 22700
rect 55480 22660 59112 22700
rect 59152 22660 59194 22700
rect 59234 22660 59276 22700
rect 59316 22660 59358 22700
rect 59398 22660 59440 22700
rect 59480 22660 63112 22700
rect 63152 22660 63194 22700
rect 63234 22660 63276 22700
rect 63316 22660 63358 22700
rect 63398 22660 63440 22700
rect 63480 22660 67112 22700
rect 67152 22660 67194 22700
rect 67234 22660 67276 22700
rect 67316 22660 67358 22700
rect 67398 22660 67440 22700
rect 67480 22660 71112 22700
rect 71152 22660 71194 22700
rect 71234 22660 71276 22700
rect 71316 22660 71358 22700
rect 71398 22660 71440 22700
rect 71480 22660 75112 22700
rect 75152 22660 75194 22700
rect 75234 22660 75276 22700
rect 75316 22660 75358 22700
rect 75398 22660 75440 22700
rect 75480 22660 79112 22700
rect 79152 22660 79194 22700
rect 79234 22660 79276 22700
rect 79316 22660 79358 22700
rect 79398 22660 79440 22700
rect 79480 22660 83112 22700
rect 83152 22660 83194 22700
rect 83234 22660 83276 22700
rect 83316 22660 83358 22700
rect 83398 22660 83440 22700
rect 83480 22660 87112 22700
rect 87152 22660 87194 22700
rect 87234 22660 87276 22700
rect 87316 22660 87358 22700
rect 87398 22660 87440 22700
rect 87480 22660 91112 22700
rect 91152 22660 91194 22700
rect 91234 22660 91276 22700
rect 91316 22660 91358 22700
rect 91398 22660 91440 22700
rect 91480 22660 95112 22700
rect 95152 22660 95194 22700
rect 95234 22660 95276 22700
rect 95316 22660 95358 22700
rect 95398 22660 95440 22700
rect 95480 22660 99112 22700
rect 99152 22660 99194 22700
rect 99234 22660 99276 22700
rect 99316 22660 99358 22700
rect 99398 22660 99440 22700
rect 99480 22660 99516 22700
rect 576 22636 99516 22660
rect 651 22448 693 22457
rect 651 22408 652 22448
rect 692 22408 693 22448
rect 651 22399 693 22408
rect 576 21944 99360 21968
rect 576 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 8352 21944
rect 8392 21904 8434 21944
rect 8474 21904 8516 21944
rect 8556 21904 8598 21944
rect 8638 21904 8680 21944
rect 8720 21904 12352 21944
rect 12392 21904 12434 21944
rect 12474 21904 12516 21944
rect 12556 21904 12598 21944
rect 12638 21904 12680 21944
rect 12720 21904 16352 21944
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16720 21904 20352 21944
rect 20392 21904 20434 21944
rect 20474 21904 20516 21944
rect 20556 21904 20598 21944
rect 20638 21904 20680 21944
rect 20720 21904 24352 21944
rect 24392 21904 24434 21944
rect 24474 21904 24516 21944
rect 24556 21904 24598 21944
rect 24638 21904 24680 21944
rect 24720 21904 28352 21944
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28720 21904 32352 21944
rect 32392 21904 32434 21944
rect 32474 21904 32516 21944
rect 32556 21904 32598 21944
rect 32638 21904 32680 21944
rect 32720 21904 36352 21944
rect 36392 21904 36434 21944
rect 36474 21904 36516 21944
rect 36556 21904 36598 21944
rect 36638 21904 36680 21944
rect 36720 21904 40352 21944
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40720 21904 44352 21944
rect 44392 21904 44434 21944
rect 44474 21904 44516 21944
rect 44556 21904 44598 21944
rect 44638 21904 44680 21944
rect 44720 21904 48352 21944
rect 48392 21904 48434 21944
rect 48474 21904 48516 21944
rect 48556 21904 48598 21944
rect 48638 21904 48680 21944
rect 48720 21904 52352 21944
rect 52392 21904 52434 21944
rect 52474 21904 52516 21944
rect 52556 21904 52598 21944
rect 52638 21904 52680 21944
rect 52720 21904 56352 21944
rect 56392 21904 56434 21944
rect 56474 21904 56516 21944
rect 56556 21904 56598 21944
rect 56638 21904 56680 21944
rect 56720 21904 60352 21944
rect 60392 21904 60434 21944
rect 60474 21904 60516 21944
rect 60556 21904 60598 21944
rect 60638 21904 60680 21944
rect 60720 21904 64352 21944
rect 64392 21904 64434 21944
rect 64474 21904 64516 21944
rect 64556 21904 64598 21944
rect 64638 21904 64680 21944
rect 64720 21904 68352 21944
rect 68392 21904 68434 21944
rect 68474 21904 68516 21944
rect 68556 21904 68598 21944
rect 68638 21904 68680 21944
rect 68720 21904 72352 21944
rect 72392 21904 72434 21944
rect 72474 21904 72516 21944
rect 72556 21904 72598 21944
rect 72638 21904 72680 21944
rect 72720 21904 76352 21944
rect 76392 21904 76434 21944
rect 76474 21904 76516 21944
rect 76556 21904 76598 21944
rect 76638 21904 76680 21944
rect 76720 21904 80352 21944
rect 80392 21904 80434 21944
rect 80474 21904 80516 21944
rect 80556 21904 80598 21944
rect 80638 21904 80680 21944
rect 80720 21904 84352 21944
rect 84392 21904 84434 21944
rect 84474 21904 84516 21944
rect 84556 21904 84598 21944
rect 84638 21904 84680 21944
rect 84720 21904 88352 21944
rect 88392 21904 88434 21944
rect 88474 21904 88516 21944
rect 88556 21904 88598 21944
rect 88638 21904 88680 21944
rect 88720 21904 92352 21944
rect 92392 21904 92434 21944
rect 92474 21904 92516 21944
rect 92556 21904 92598 21944
rect 92638 21904 92680 21944
rect 92720 21904 96352 21944
rect 96392 21904 96434 21944
rect 96474 21904 96516 21944
rect 96556 21904 96598 21944
rect 96638 21904 96680 21944
rect 96720 21904 99360 21944
rect 576 21880 99360 21904
rect 576 21188 99516 21212
rect 576 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 7112 21188
rect 7152 21148 7194 21188
rect 7234 21148 7276 21188
rect 7316 21148 7358 21188
rect 7398 21148 7440 21188
rect 7480 21148 11112 21188
rect 11152 21148 11194 21188
rect 11234 21148 11276 21188
rect 11316 21148 11358 21188
rect 11398 21148 11440 21188
rect 11480 21148 15112 21188
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15480 21148 19112 21188
rect 19152 21148 19194 21188
rect 19234 21148 19276 21188
rect 19316 21148 19358 21188
rect 19398 21148 19440 21188
rect 19480 21148 23112 21188
rect 23152 21148 23194 21188
rect 23234 21148 23276 21188
rect 23316 21148 23358 21188
rect 23398 21148 23440 21188
rect 23480 21148 27112 21188
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27480 21148 31112 21188
rect 31152 21148 31194 21188
rect 31234 21148 31276 21188
rect 31316 21148 31358 21188
rect 31398 21148 31440 21188
rect 31480 21148 35112 21188
rect 35152 21148 35194 21188
rect 35234 21148 35276 21188
rect 35316 21148 35358 21188
rect 35398 21148 35440 21188
rect 35480 21148 39112 21188
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39480 21148 43112 21188
rect 43152 21148 43194 21188
rect 43234 21148 43276 21188
rect 43316 21148 43358 21188
rect 43398 21148 43440 21188
rect 43480 21148 47112 21188
rect 47152 21148 47194 21188
rect 47234 21148 47276 21188
rect 47316 21148 47358 21188
rect 47398 21148 47440 21188
rect 47480 21148 51112 21188
rect 51152 21148 51194 21188
rect 51234 21148 51276 21188
rect 51316 21148 51358 21188
rect 51398 21148 51440 21188
rect 51480 21148 55112 21188
rect 55152 21148 55194 21188
rect 55234 21148 55276 21188
rect 55316 21148 55358 21188
rect 55398 21148 55440 21188
rect 55480 21148 59112 21188
rect 59152 21148 59194 21188
rect 59234 21148 59276 21188
rect 59316 21148 59358 21188
rect 59398 21148 59440 21188
rect 59480 21148 63112 21188
rect 63152 21148 63194 21188
rect 63234 21148 63276 21188
rect 63316 21148 63358 21188
rect 63398 21148 63440 21188
rect 63480 21148 67112 21188
rect 67152 21148 67194 21188
rect 67234 21148 67276 21188
rect 67316 21148 67358 21188
rect 67398 21148 67440 21188
rect 67480 21148 71112 21188
rect 71152 21148 71194 21188
rect 71234 21148 71276 21188
rect 71316 21148 71358 21188
rect 71398 21148 71440 21188
rect 71480 21148 75112 21188
rect 75152 21148 75194 21188
rect 75234 21148 75276 21188
rect 75316 21148 75358 21188
rect 75398 21148 75440 21188
rect 75480 21148 79112 21188
rect 79152 21148 79194 21188
rect 79234 21148 79276 21188
rect 79316 21148 79358 21188
rect 79398 21148 79440 21188
rect 79480 21148 83112 21188
rect 83152 21148 83194 21188
rect 83234 21148 83276 21188
rect 83316 21148 83358 21188
rect 83398 21148 83440 21188
rect 83480 21148 87112 21188
rect 87152 21148 87194 21188
rect 87234 21148 87276 21188
rect 87316 21148 87358 21188
rect 87398 21148 87440 21188
rect 87480 21148 91112 21188
rect 91152 21148 91194 21188
rect 91234 21148 91276 21188
rect 91316 21148 91358 21188
rect 91398 21148 91440 21188
rect 91480 21148 95112 21188
rect 95152 21148 95194 21188
rect 95234 21148 95276 21188
rect 95316 21148 95358 21188
rect 95398 21148 95440 21188
rect 95480 21148 99112 21188
rect 99152 21148 99194 21188
rect 99234 21148 99276 21188
rect 99316 21148 99358 21188
rect 99398 21148 99440 21188
rect 99480 21148 99516 21188
rect 576 21124 99516 21148
rect 651 20936 693 20945
rect 651 20896 652 20936
rect 692 20896 693 20936
rect 651 20887 693 20896
rect 576 20432 99360 20456
rect 576 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 8352 20432
rect 8392 20392 8434 20432
rect 8474 20392 8516 20432
rect 8556 20392 8598 20432
rect 8638 20392 8680 20432
rect 8720 20392 12352 20432
rect 12392 20392 12434 20432
rect 12474 20392 12516 20432
rect 12556 20392 12598 20432
rect 12638 20392 12680 20432
rect 12720 20392 16352 20432
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16720 20392 20352 20432
rect 20392 20392 20434 20432
rect 20474 20392 20516 20432
rect 20556 20392 20598 20432
rect 20638 20392 20680 20432
rect 20720 20392 24352 20432
rect 24392 20392 24434 20432
rect 24474 20392 24516 20432
rect 24556 20392 24598 20432
rect 24638 20392 24680 20432
rect 24720 20392 28352 20432
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28720 20392 32352 20432
rect 32392 20392 32434 20432
rect 32474 20392 32516 20432
rect 32556 20392 32598 20432
rect 32638 20392 32680 20432
rect 32720 20392 36352 20432
rect 36392 20392 36434 20432
rect 36474 20392 36516 20432
rect 36556 20392 36598 20432
rect 36638 20392 36680 20432
rect 36720 20392 40352 20432
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40720 20392 44352 20432
rect 44392 20392 44434 20432
rect 44474 20392 44516 20432
rect 44556 20392 44598 20432
rect 44638 20392 44680 20432
rect 44720 20392 48352 20432
rect 48392 20392 48434 20432
rect 48474 20392 48516 20432
rect 48556 20392 48598 20432
rect 48638 20392 48680 20432
rect 48720 20392 52352 20432
rect 52392 20392 52434 20432
rect 52474 20392 52516 20432
rect 52556 20392 52598 20432
rect 52638 20392 52680 20432
rect 52720 20392 56352 20432
rect 56392 20392 56434 20432
rect 56474 20392 56516 20432
rect 56556 20392 56598 20432
rect 56638 20392 56680 20432
rect 56720 20392 60352 20432
rect 60392 20392 60434 20432
rect 60474 20392 60516 20432
rect 60556 20392 60598 20432
rect 60638 20392 60680 20432
rect 60720 20392 64352 20432
rect 64392 20392 64434 20432
rect 64474 20392 64516 20432
rect 64556 20392 64598 20432
rect 64638 20392 64680 20432
rect 64720 20392 68352 20432
rect 68392 20392 68434 20432
rect 68474 20392 68516 20432
rect 68556 20392 68598 20432
rect 68638 20392 68680 20432
rect 68720 20392 72352 20432
rect 72392 20392 72434 20432
rect 72474 20392 72516 20432
rect 72556 20392 72598 20432
rect 72638 20392 72680 20432
rect 72720 20392 76352 20432
rect 76392 20392 76434 20432
rect 76474 20392 76516 20432
rect 76556 20392 76598 20432
rect 76638 20392 76680 20432
rect 76720 20392 80352 20432
rect 80392 20392 80434 20432
rect 80474 20392 80516 20432
rect 80556 20392 80598 20432
rect 80638 20392 80680 20432
rect 80720 20392 84352 20432
rect 84392 20392 84434 20432
rect 84474 20392 84516 20432
rect 84556 20392 84598 20432
rect 84638 20392 84680 20432
rect 84720 20392 88352 20432
rect 88392 20392 88434 20432
rect 88474 20392 88516 20432
rect 88556 20392 88598 20432
rect 88638 20392 88680 20432
rect 88720 20392 92352 20432
rect 92392 20392 92434 20432
rect 92474 20392 92516 20432
rect 92556 20392 92598 20432
rect 92638 20392 92680 20432
rect 92720 20392 96352 20432
rect 96392 20392 96434 20432
rect 96474 20392 96516 20432
rect 96556 20392 96598 20432
rect 96638 20392 96680 20432
rect 96720 20392 99360 20432
rect 576 20368 99360 20392
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 576 19676 99516 19700
rect 576 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 7112 19676
rect 7152 19636 7194 19676
rect 7234 19636 7276 19676
rect 7316 19636 7358 19676
rect 7398 19636 7440 19676
rect 7480 19636 11112 19676
rect 11152 19636 11194 19676
rect 11234 19636 11276 19676
rect 11316 19636 11358 19676
rect 11398 19636 11440 19676
rect 11480 19636 15112 19676
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15480 19636 19112 19676
rect 19152 19636 19194 19676
rect 19234 19636 19276 19676
rect 19316 19636 19358 19676
rect 19398 19636 19440 19676
rect 19480 19636 23112 19676
rect 23152 19636 23194 19676
rect 23234 19636 23276 19676
rect 23316 19636 23358 19676
rect 23398 19636 23440 19676
rect 23480 19636 27112 19676
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27480 19636 31112 19676
rect 31152 19636 31194 19676
rect 31234 19636 31276 19676
rect 31316 19636 31358 19676
rect 31398 19636 31440 19676
rect 31480 19636 35112 19676
rect 35152 19636 35194 19676
rect 35234 19636 35276 19676
rect 35316 19636 35358 19676
rect 35398 19636 35440 19676
rect 35480 19636 39112 19676
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39480 19636 43112 19676
rect 43152 19636 43194 19676
rect 43234 19636 43276 19676
rect 43316 19636 43358 19676
rect 43398 19636 43440 19676
rect 43480 19636 47112 19676
rect 47152 19636 47194 19676
rect 47234 19636 47276 19676
rect 47316 19636 47358 19676
rect 47398 19636 47440 19676
rect 47480 19636 51112 19676
rect 51152 19636 51194 19676
rect 51234 19636 51276 19676
rect 51316 19636 51358 19676
rect 51398 19636 51440 19676
rect 51480 19636 55112 19676
rect 55152 19636 55194 19676
rect 55234 19636 55276 19676
rect 55316 19636 55358 19676
rect 55398 19636 55440 19676
rect 55480 19636 59112 19676
rect 59152 19636 59194 19676
rect 59234 19636 59276 19676
rect 59316 19636 59358 19676
rect 59398 19636 59440 19676
rect 59480 19636 63112 19676
rect 63152 19636 63194 19676
rect 63234 19636 63276 19676
rect 63316 19636 63358 19676
rect 63398 19636 63440 19676
rect 63480 19636 67112 19676
rect 67152 19636 67194 19676
rect 67234 19636 67276 19676
rect 67316 19636 67358 19676
rect 67398 19636 67440 19676
rect 67480 19636 71112 19676
rect 71152 19636 71194 19676
rect 71234 19636 71276 19676
rect 71316 19636 71358 19676
rect 71398 19636 71440 19676
rect 71480 19636 75112 19676
rect 75152 19636 75194 19676
rect 75234 19636 75276 19676
rect 75316 19636 75358 19676
rect 75398 19636 75440 19676
rect 75480 19636 79112 19676
rect 79152 19636 79194 19676
rect 79234 19636 79276 19676
rect 79316 19636 79358 19676
rect 79398 19636 79440 19676
rect 79480 19636 83112 19676
rect 83152 19636 83194 19676
rect 83234 19636 83276 19676
rect 83316 19636 83358 19676
rect 83398 19636 83440 19676
rect 83480 19636 87112 19676
rect 87152 19636 87194 19676
rect 87234 19636 87276 19676
rect 87316 19636 87358 19676
rect 87398 19636 87440 19676
rect 87480 19636 91112 19676
rect 91152 19636 91194 19676
rect 91234 19636 91276 19676
rect 91316 19636 91358 19676
rect 91398 19636 91440 19676
rect 91480 19636 95112 19676
rect 95152 19636 95194 19676
rect 95234 19636 95276 19676
rect 95316 19636 95358 19676
rect 95398 19636 95440 19676
rect 95480 19636 99112 19676
rect 99152 19636 99194 19676
rect 99234 19636 99276 19676
rect 99316 19636 99358 19676
rect 99398 19636 99440 19676
rect 99480 19636 99516 19676
rect 576 19612 99516 19636
rect 651 19424 693 19433
rect 651 19384 652 19424
rect 692 19384 693 19424
rect 651 19375 693 19384
rect 576 18920 99360 18944
rect 576 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 8352 18920
rect 8392 18880 8434 18920
rect 8474 18880 8516 18920
rect 8556 18880 8598 18920
rect 8638 18880 8680 18920
rect 8720 18880 12352 18920
rect 12392 18880 12434 18920
rect 12474 18880 12516 18920
rect 12556 18880 12598 18920
rect 12638 18880 12680 18920
rect 12720 18880 16352 18920
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16720 18880 20352 18920
rect 20392 18880 20434 18920
rect 20474 18880 20516 18920
rect 20556 18880 20598 18920
rect 20638 18880 20680 18920
rect 20720 18880 24352 18920
rect 24392 18880 24434 18920
rect 24474 18880 24516 18920
rect 24556 18880 24598 18920
rect 24638 18880 24680 18920
rect 24720 18880 28352 18920
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28720 18880 32352 18920
rect 32392 18880 32434 18920
rect 32474 18880 32516 18920
rect 32556 18880 32598 18920
rect 32638 18880 32680 18920
rect 32720 18880 36352 18920
rect 36392 18880 36434 18920
rect 36474 18880 36516 18920
rect 36556 18880 36598 18920
rect 36638 18880 36680 18920
rect 36720 18880 40352 18920
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40720 18880 44352 18920
rect 44392 18880 44434 18920
rect 44474 18880 44516 18920
rect 44556 18880 44598 18920
rect 44638 18880 44680 18920
rect 44720 18880 48352 18920
rect 48392 18880 48434 18920
rect 48474 18880 48516 18920
rect 48556 18880 48598 18920
rect 48638 18880 48680 18920
rect 48720 18880 52352 18920
rect 52392 18880 52434 18920
rect 52474 18880 52516 18920
rect 52556 18880 52598 18920
rect 52638 18880 52680 18920
rect 52720 18880 56352 18920
rect 56392 18880 56434 18920
rect 56474 18880 56516 18920
rect 56556 18880 56598 18920
rect 56638 18880 56680 18920
rect 56720 18880 60352 18920
rect 60392 18880 60434 18920
rect 60474 18880 60516 18920
rect 60556 18880 60598 18920
rect 60638 18880 60680 18920
rect 60720 18880 64352 18920
rect 64392 18880 64434 18920
rect 64474 18880 64516 18920
rect 64556 18880 64598 18920
rect 64638 18880 64680 18920
rect 64720 18880 68352 18920
rect 68392 18880 68434 18920
rect 68474 18880 68516 18920
rect 68556 18880 68598 18920
rect 68638 18880 68680 18920
rect 68720 18880 72352 18920
rect 72392 18880 72434 18920
rect 72474 18880 72516 18920
rect 72556 18880 72598 18920
rect 72638 18880 72680 18920
rect 72720 18880 76352 18920
rect 76392 18880 76434 18920
rect 76474 18880 76516 18920
rect 76556 18880 76598 18920
rect 76638 18880 76680 18920
rect 76720 18880 80352 18920
rect 80392 18880 80434 18920
rect 80474 18880 80516 18920
rect 80556 18880 80598 18920
rect 80638 18880 80680 18920
rect 80720 18880 84352 18920
rect 84392 18880 84434 18920
rect 84474 18880 84516 18920
rect 84556 18880 84598 18920
rect 84638 18880 84680 18920
rect 84720 18880 88352 18920
rect 88392 18880 88434 18920
rect 88474 18880 88516 18920
rect 88556 18880 88598 18920
rect 88638 18880 88680 18920
rect 88720 18880 92352 18920
rect 92392 18880 92434 18920
rect 92474 18880 92516 18920
rect 92556 18880 92598 18920
rect 92638 18880 92680 18920
rect 92720 18880 96352 18920
rect 96392 18880 96434 18920
rect 96474 18880 96516 18920
rect 96556 18880 96598 18920
rect 96638 18880 96680 18920
rect 96720 18880 99360 18920
rect 576 18856 99360 18880
rect 651 18416 693 18425
rect 651 18376 652 18416
rect 692 18376 693 18416
rect 651 18367 693 18376
rect 576 18164 99516 18188
rect 576 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 7112 18164
rect 7152 18124 7194 18164
rect 7234 18124 7276 18164
rect 7316 18124 7358 18164
rect 7398 18124 7440 18164
rect 7480 18124 11112 18164
rect 11152 18124 11194 18164
rect 11234 18124 11276 18164
rect 11316 18124 11358 18164
rect 11398 18124 11440 18164
rect 11480 18124 15112 18164
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15480 18124 19112 18164
rect 19152 18124 19194 18164
rect 19234 18124 19276 18164
rect 19316 18124 19358 18164
rect 19398 18124 19440 18164
rect 19480 18124 23112 18164
rect 23152 18124 23194 18164
rect 23234 18124 23276 18164
rect 23316 18124 23358 18164
rect 23398 18124 23440 18164
rect 23480 18124 27112 18164
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27480 18124 31112 18164
rect 31152 18124 31194 18164
rect 31234 18124 31276 18164
rect 31316 18124 31358 18164
rect 31398 18124 31440 18164
rect 31480 18124 35112 18164
rect 35152 18124 35194 18164
rect 35234 18124 35276 18164
rect 35316 18124 35358 18164
rect 35398 18124 35440 18164
rect 35480 18124 39112 18164
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39480 18124 43112 18164
rect 43152 18124 43194 18164
rect 43234 18124 43276 18164
rect 43316 18124 43358 18164
rect 43398 18124 43440 18164
rect 43480 18124 47112 18164
rect 47152 18124 47194 18164
rect 47234 18124 47276 18164
rect 47316 18124 47358 18164
rect 47398 18124 47440 18164
rect 47480 18124 51112 18164
rect 51152 18124 51194 18164
rect 51234 18124 51276 18164
rect 51316 18124 51358 18164
rect 51398 18124 51440 18164
rect 51480 18124 55112 18164
rect 55152 18124 55194 18164
rect 55234 18124 55276 18164
rect 55316 18124 55358 18164
rect 55398 18124 55440 18164
rect 55480 18124 59112 18164
rect 59152 18124 59194 18164
rect 59234 18124 59276 18164
rect 59316 18124 59358 18164
rect 59398 18124 59440 18164
rect 59480 18124 63112 18164
rect 63152 18124 63194 18164
rect 63234 18124 63276 18164
rect 63316 18124 63358 18164
rect 63398 18124 63440 18164
rect 63480 18124 67112 18164
rect 67152 18124 67194 18164
rect 67234 18124 67276 18164
rect 67316 18124 67358 18164
rect 67398 18124 67440 18164
rect 67480 18124 71112 18164
rect 71152 18124 71194 18164
rect 71234 18124 71276 18164
rect 71316 18124 71358 18164
rect 71398 18124 71440 18164
rect 71480 18124 75112 18164
rect 75152 18124 75194 18164
rect 75234 18124 75276 18164
rect 75316 18124 75358 18164
rect 75398 18124 75440 18164
rect 75480 18124 79112 18164
rect 79152 18124 79194 18164
rect 79234 18124 79276 18164
rect 79316 18124 79358 18164
rect 79398 18124 79440 18164
rect 79480 18124 83112 18164
rect 83152 18124 83194 18164
rect 83234 18124 83276 18164
rect 83316 18124 83358 18164
rect 83398 18124 83440 18164
rect 83480 18124 87112 18164
rect 87152 18124 87194 18164
rect 87234 18124 87276 18164
rect 87316 18124 87358 18164
rect 87398 18124 87440 18164
rect 87480 18124 91112 18164
rect 91152 18124 91194 18164
rect 91234 18124 91276 18164
rect 91316 18124 91358 18164
rect 91398 18124 91440 18164
rect 91480 18124 95112 18164
rect 95152 18124 95194 18164
rect 95234 18124 95276 18164
rect 95316 18124 95358 18164
rect 95398 18124 95440 18164
rect 95480 18124 99112 18164
rect 99152 18124 99194 18164
rect 99234 18124 99276 18164
rect 99316 18124 99358 18164
rect 99398 18124 99440 18164
rect 99480 18124 99516 18164
rect 576 18100 99516 18124
rect 651 17912 693 17921
rect 651 17872 652 17912
rect 692 17872 693 17912
rect 651 17863 693 17872
rect 576 17408 99360 17432
rect 576 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 8352 17408
rect 8392 17368 8434 17408
rect 8474 17368 8516 17408
rect 8556 17368 8598 17408
rect 8638 17368 8680 17408
rect 8720 17368 12352 17408
rect 12392 17368 12434 17408
rect 12474 17368 12516 17408
rect 12556 17368 12598 17408
rect 12638 17368 12680 17408
rect 12720 17368 16352 17408
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16720 17368 20352 17408
rect 20392 17368 20434 17408
rect 20474 17368 20516 17408
rect 20556 17368 20598 17408
rect 20638 17368 20680 17408
rect 20720 17368 24352 17408
rect 24392 17368 24434 17408
rect 24474 17368 24516 17408
rect 24556 17368 24598 17408
rect 24638 17368 24680 17408
rect 24720 17368 28352 17408
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28720 17368 32352 17408
rect 32392 17368 32434 17408
rect 32474 17368 32516 17408
rect 32556 17368 32598 17408
rect 32638 17368 32680 17408
rect 32720 17368 36352 17408
rect 36392 17368 36434 17408
rect 36474 17368 36516 17408
rect 36556 17368 36598 17408
rect 36638 17368 36680 17408
rect 36720 17368 40352 17408
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40720 17368 44352 17408
rect 44392 17368 44434 17408
rect 44474 17368 44516 17408
rect 44556 17368 44598 17408
rect 44638 17368 44680 17408
rect 44720 17368 48352 17408
rect 48392 17368 48434 17408
rect 48474 17368 48516 17408
rect 48556 17368 48598 17408
rect 48638 17368 48680 17408
rect 48720 17368 52352 17408
rect 52392 17368 52434 17408
rect 52474 17368 52516 17408
rect 52556 17368 52598 17408
rect 52638 17368 52680 17408
rect 52720 17368 56352 17408
rect 56392 17368 56434 17408
rect 56474 17368 56516 17408
rect 56556 17368 56598 17408
rect 56638 17368 56680 17408
rect 56720 17368 60352 17408
rect 60392 17368 60434 17408
rect 60474 17368 60516 17408
rect 60556 17368 60598 17408
rect 60638 17368 60680 17408
rect 60720 17368 64352 17408
rect 64392 17368 64434 17408
rect 64474 17368 64516 17408
rect 64556 17368 64598 17408
rect 64638 17368 64680 17408
rect 64720 17368 68352 17408
rect 68392 17368 68434 17408
rect 68474 17368 68516 17408
rect 68556 17368 68598 17408
rect 68638 17368 68680 17408
rect 68720 17368 72352 17408
rect 72392 17368 72434 17408
rect 72474 17368 72516 17408
rect 72556 17368 72598 17408
rect 72638 17368 72680 17408
rect 72720 17368 76352 17408
rect 76392 17368 76434 17408
rect 76474 17368 76516 17408
rect 76556 17368 76598 17408
rect 76638 17368 76680 17408
rect 76720 17368 80352 17408
rect 80392 17368 80434 17408
rect 80474 17368 80516 17408
rect 80556 17368 80598 17408
rect 80638 17368 80680 17408
rect 80720 17368 84352 17408
rect 84392 17368 84434 17408
rect 84474 17368 84516 17408
rect 84556 17368 84598 17408
rect 84638 17368 84680 17408
rect 84720 17368 88352 17408
rect 88392 17368 88434 17408
rect 88474 17368 88516 17408
rect 88556 17368 88598 17408
rect 88638 17368 88680 17408
rect 88720 17368 92352 17408
rect 92392 17368 92434 17408
rect 92474 17368 92516 17408
rect 92556 17368 92598 17408
rect 92638 17368 92680 17408
rect 92720 17368 96352 17408
rect 96392 17368 96434 17408
rect 96474 17368 96516 17408
rect 96556 17368 96598 17408
rect 96638 17368 96680 17408
rect 96720 17368 99360 17408
rect 576 17344 99360 17368
rect 86563 17072 86621 17073
rect 86563 17032 86572 17072
rect 86612 17032 86621 17072
rect 86563 17031 86621 17032
rect 86755 17072 86813 17073
rect 86755 17032 86764 17072
rect 86804 17032 86813 17072
rect 86755 17031 86813 17032
rect 80419 16988 80477 16989
rect 80419 16948 80428 16988
rect 80468 16948 80477 16988
rect 80419 16947 80477 16948
rect 86179 16988 86237 16989
rect 86179 16948 86188 16988
rect 86228 16948 86237 16988
rect 86179 16947 86237 16948
rect 651 16904 693 16913
rect 651 16864 652 16904
rect 692 16864 693 16904
rect 651 16855 693 16864
rect 80619 16820 80661 16829
rect 80619 16780 80620 16820
rect 80660 16780 80661 16820
rect 80619 16771 80661 16780
rect 86379 16820 86421 16829
rect 86379 16780 86380 16820
rect 86420 16780 86421 16820
rect 86379 16771 86421 16780
rect 576 16652 99516 16676
rect 576 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 7112 16652
rect 7152 16612 7194 16652
rect 7234 16612 7276 16652
rect 7316 16612 7358 16652
rect 7398 16612 7440 16652
rect 7480 16612 11112 16652
rect 11152 16612 11194 16652
rect 11234 16612 11276 16652
rect 11316 16612 11358 16652
rect 11398 16612 11440 16652
rect 11480 16612 15112 16652
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15480 16612 19112 16652
rect 19152 16612 19194 16652
rect 19234 16612 19276 16652
rect 19316 16612 19358 16652
rect 19398 16612 19440 16652
rect 19480 16612 23112 16652
rect 23152 16612 23194 16652
rect 23234 16612 23276 16652
rect 23316 16612 23358 16652
rect 23398 16612 23440 16652
rect 23480 16612 27112 16652
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27480 16612 31112 16652
rect 31152 16612 31194 16652
rect 31234 16612 31276 16652
rect 31316 16612 31358 16652
rect 31398 16612 31440 16652
rect 31480 16612 35112 16652
rect 35152 16612 35194 16652
rect 35234 16612 35276 16652
rect 35316 16612 35358 16652
rect 35398 16612 35440 16652
rect 35480 16612 39112 16652
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39480 16612 43112 16652
rect 43152 16612 43194 16652
rect 43234 16612 43276 16652
rect 43316 16612 43358 16652
rect 43398 16612 43440 16652
rect 43480 16612 47112 16652
rect 47152 16612 47194 16652
rect 47234 16612 47276 16652
rect 47316 16612 47358 16652
rect 47398 16612 47440 16652
rect 47480 16612 51112 16652
rect 51152 16612 51194 16652
rect 51234 16612 51276 16652
rect 51316 16612 51358 16652
rect 51398 16612 51440 16652
rect 51480 16612 55112 16652
rect 55152 16612 55194 16652
rect 55234 16612 55276 16652
rect 55316 16612 55358 16652
rect 55398 16612 55440 16652
rect 55480 16612 59112 16652
rect 59152 16612 59194 16652
rect 59234 16612 59276 16652
rect 59316 16612 59358 16652
rect 59398 16612 59440 16652
rect 59480 16612 63112 16652
rect 63152 16612 63194 16652
rect 63234 16612 63276 16652
rect 63316 16612 63358 16652
rect 63398 16612 63440 16652
rect 63480 16612 67112 16652
rect 67152 16612 67194 16652
rect 67234 16612 67276 16652
rect 67316 16612 67358 16652
rect 67398 16612 67440 16652
rect 67480 16612 71112 16652
rect 71152 16612 71194 16652
rect 71234 16612 71276 16652
rect 71316 16612 71358 16652
rect 71398 16612 71440 16652
rect 71480 16612 75112 16652
rect 75152 16612 75194 16652
rect 75234 16612 75276 16652
rect 75316 16612 75358 16652
rect 75398 16612 75440 16652
rect 75480 16612 79112 16652
rect 79152 16612 79194 16652
rect 79234 16612 79276 16652
rect 79316 16612 79358 16652
rect 79398 16612 79440 16652
rect 79480 16612 83112 16652
rect 83152 16612 83194 16652
rect 83234 16612 83276 16652
rect 83316 16612 83358 16652
rect 83398 16612 83440 16652
rect 83480 16612 87112 16652
rect 87152 16612 87194 16652
rect 87234 16612 87276 16652
rect 87316 16612 87358 16652
rect 87398 16612 87440 16652
rect 87480 16612 91112 16652
rect 91152 16612 91194 16652
rect 91234 16612 91276 16652
rect 91316 16612 91358 16652
rect 91398 16612 91440 16652
rect 91480 16612 95112 16652
rect 95152 16612 95194 16652
rect 95234 16612 95276 16652
rect 95316 16612 95358 16652
rect 95398 16612 95440 16652
rect 95480 16612 99112 16652
rect 99152 16612 99194 16652
rect 99234 16612 99276 16652
rect 99316 16612 99358 16652
rect 99398 16612 99440 16652
rect 99480 16612 99516 16652
rect 576 16588 99516 16612
rect 651 16400 693 16409
rect 651 16360 652 16400
rect 692 16360 693 16400
rect 651 16351 693 16360
rect 74475 16400 74517 16409
rect 74475 16360 74476 16400
rect 74516 16360 74517 16400
rect 74475 16351 74517 16360
rect 81579 16400 81621 16409
rect 81579 16360 81580 16400
rect 81620 16360 81621 16400
rect 81579 16351 81621 16360
rect 83115 16400 83157 16409
rect 83115 16360 83116 16400
rect 83156 16360 83157 16400
rect 83115 16351 83157 16360
rect 73891 16316 73949 16317
rect 73891 16276 73900 16316
rect 73940 16276 73949 16316
rect 73891 16275 73949 16276
rect 74275 16316 74333 16317
rect 74275 16276 74284 16316
rect 74324 16276 74333 16316
rect 74275 16275 74333 16276
rect 76771 16316 76829 16317
rect 76771 16276 76780 16316
rect 76820 16276 76829 16316
rect 76771 16275 76829 16276
rect 77155 16316 77213 16317
rect 77155 16276 77164 16316
rect 77204 16276 77213 16316
rect 77155 16275 77213 16276
rect 80515 16316 80573 16317
rect 80515 16276 80524 16316
rect 80564 16276 80573 16316
rect 80515 16275 80573 16276
rect 81187 16316 81245 16317
rect 81187 16276 81196 16316
rect 81236 16276 81245 16316
rect 81187 16275 81245 16276
rect 81763 16316 81821 16317
rect 81763 16276 81772 16316
rect 81812 16276 81821 16316
rect 81763 16275 81821 16276
rect 82147 16316 82205 16317
rect 82147 16276 82156 16316
rect 82196 16276 82205 16316
rect 82147 16275 82205 16276
rect 82531 16316 82589 16317
rect 82531 16276 82540 16316
rect 82580 16276 82589 16316
rect 82531 16275 82589 16276
rect 83299 16316 83357 16317
rect 83299 16276 83308 16316
rect 83348 16276 83357 16316
rect 83299 16275 83357 16276
rect 83779 16316 83837 16317
rect 83779 16276 83788 16316
rect 83828 16276 83837 16316
rect 83779 16275 83837 16276
rect 84643 16316 84701 16317
rect 84643 16276 84652 16316
rect 84692 16276 84701 16316
rect 84643 16275 84701 16276
rect 86563 16316 86621 16317
rect 86563 16276 86572 16316
rect 86612 16276 86621 16316
rect 86563 16275 86621 16276
rect 87427 16316 87485 16317
rect 87427 16276 87436 16316
rect 87476 16276 87485 16316
rect 87427 16275 87485 16276
rect 88195 16316 88253 16317
rect 88195 16276 88204 16316
rect 88244 16276 88253 16316
rect 88195 16275 88253 16276
rect 89347 16316 89405 16317
rect 89347 16276 89356 16316
rect 89396 16276 89405 16316
rect 89347 16275 89405 16276
rect 90595 16316 90653 16317
rect 90595 16276 90604 16316
rect 90644 16276 90653 16316
rect 90595 16275 90653 16276
rect 92227 16316 92285 16317
rect 92227 16276 92236 16316
rect 92276 16276 92285 16316
rect 92227 16275 92285 16276
rect 92419 16316 92477 16317
rect 92419 16276 92428 16316
rect 92468 16276 92477 16316
rect 92419 16275 92477 16276
rect 94051 16316 94109 16317
rect 94051 16276 94060 16316
rect 94100 16276 94109 16316
rect 94051 16275 94109 16276
rect 95587 16316 95645 16317
rect 95587 16276 95596 16316
rect 95636 16276 95645 16316
rect 95587 16275 95645 16276
rect 90979 16232 91037 16233
rect 90979 16192 90988 16232
rect 91028 16192 91037 16232
rect 90979 16191 91037 16192
rect 74091 16064 74133 16073
rect 74091 16024 74092 16064
rect 74132 16024 74133 16064
rect 74091 16015 74133 16024
rect 76971 16064 77013 16073
rect 76971 16024 76972 16064
rect 77012 16024 77013 16064
rect 76971 16015 77013 16024
rect 77355 16064 77397 16073
rect 77355 16024 77356 16064
rect 77396 16024 77397 16064
rect 77355 16015 77397 16024
rect 80331 16064 80373 16073
rect 80331 16024 80332 16064
rect 80372 16024 80373 16064
rect 80331 16015 80373 16024
rect 81387 16064 81429 16073
rect 81387 16024 81388 16064
rect 81428 16024 81429 16064
rect 81387 16015 81429 16024
rect 81963 16064 82005 16073
rect 81963 16024 81964 16064
rect 82004 16024 82005 16064
rect 81963 16015 82005 16024
rect 82731 16064 82773 16073
rect 82731 16024 82732 16064
rect 82772 16024 82773 16064
rect 82731 16015 82773 16024
rect 83979 16064 84021 16073
rect 83979 16024 83980 16064
rect 84020 16024 84021 16064
rect 83979 16015 84021 16024
rect 84843 16064 84885 16073
rect 84843 16024 84844 16064
rect 84884 16024 84885 16064
rect 84843 16015 84885 16024
rect 86379 16064 86421 16073
rect 86379 16024 86380 16064
rect 86420 16024 86421 16064
rect 86379 16015 86421 16024
rect 87627 16064 87669 16073
rect 87627 16024 87628 16064
rect 87668 16024 87669 16064
rect 87627 16015 87669 16024
rect 88011 16064 88053 16073
rect 88011 16024 88012 16064
rect 88052 16024 88053 16064
rect 88011 16015 88053 16024
rect 89163 16064 89205 16073
rect 89163 16024 89164 16064
rect 89204 16024 89205 16064
rect 89163 16015 89205 16024
rect 90795 16064 90837 16073
rect 90795 16024 90796 16064
rect 90836 16024 90837 16064
rect 90795 16015 90837 16024
rect 91083 16064 91125 16073
rect 91083 16024 91084 16064
rect 91124 16024 91125 16064
rect 91083 16015 91125 16024
rect 92043 16064 92085 16073
rect 92043 16024 92044 16064
rect 92084 16024 92085 16064
rect 92043 16015 92085 16024
rect 92619 16064 92661 16073
rect 92619 16024 92620 16064
rect 92660 16024 92661 16064
rect 92619 16015 92661 16024
rect 93867 16064 93909 16073
rect 93867 16024 93868 16064
rect 93908 16024 93909 16064
rect 93867 16015 93909 16024
rect 95787 16064 95829 16073
rect 95787 16024 95788 16064
rect 95828 16024 95829 16064
rect 95787 16015 95829 16024
rect 576 15896 99360 15920
rect 576 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 8352 15896
rect 8392 15856 8434 15896
rect 8474 15856 8516 15896
rect 8556 15856 8598 15896
rect 8638 15856 8680 15896
rect 8720 15856 12352 15896
rect 12392 15856 12434 15896
rect 12474 15856 12516 15896
rect 12556 15856 12598 15896
rect 12638 15856 12680 15896
rect 12720 15856 16352 15896
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16720 15856 20352 15896
rect 20392 15856 20434 15896
rect 20474 15856 20516 15896
rect 20556 15856 20598 15896
rect 20638 15856 20680 15896
rect 20720 15856 24352 15896
rect 24392 15856 24434 15896
rect 24474 15856 24516 15896
rect 24556 15856 24598 15896
rect 24638 15856 24680 15896
rect 24720 15856 28352 15896
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28720 15856 32352 15896
rect 32392 15856 32434 15896
rect 32474 15856 32516 15896
rect 32556 15856 32598 15896
rect 32638 15856 32680 15896
rect 32720 15856 36352 15896
rect 36392 15856 36434 15896
rect 36474 15856 36516 15896
rect 36556 15856 36598 15896
rect 36638 15856 36680 15896
rect 36720 15856 40352 15896
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40720 15856 44352 15896
rect 44392 15856 44434 15896
rect 44474 15856 44516 15896
rect 44556 15856 44598 15896
rect 44638 15856 44680 15896
rect 44720 15856 48352 15896
rect 48392 15856 48434 15896
rect 48474 15856 48516 15896
rect 48556 15856 48598 15896
rect 48638 15856 48680 15896
rect 48720 15856 52352 15896
rect 52392 15856 52434 15896
rect 52474 15856 52516 15896
rect 52556 15856 52598 15896
rect 52638 15856 52680 15896
rect 52720 15856 56352 15896
rect 56392 15856 56434 15896
rect 56474 15856 56516 15896
rect 56556 15856 56598 15896
rect 56638 15856 56680 15896
rect 56720 15856 60352 15896
rect 60392 15856 60434 15896
rect 60474 15856 60516 15896
rect 60556 15856 60598 15896
rect 60638 15856 60680 15896
rect 60720 15856 64352 15896
rect 64392 15856 64434 15896
rect 64474 15856 64516 15896
rect 64556 15856 64598 15896
rect 64638 15856 64680 15896
rect 64720 15856 68352 15896
rect 68392 15856 68434 15896
rect 68474 15856 68516 15896
rect 68556 15856 68598 15896
rect 68638 15856 68680 15896
rect 68720 15856 72352 15896
rect 72392 15856 72434 15896
rect 72474 15856 72516 15896
rect 72556 15856 72598 15896
rect 72638 15856 72680 15896
rect 72720 15856 76352 15896
rect 76392 15856 76434 15896
rect 76474 15856 76516 15896
rect 76556 15856 76598 15896
rect 76638 15856 76680 15896
rect 76720 15856 80352 15896
rect 80392 15856 80434 15896
rect 80474 15856 80516 15896
rect 80556 15856 80598 15896
rect 80638 15856 80680 15896
rect 80720 15856 84352 15896
rect 84392 15856 84434 15896
rect 84474 15856 84516 15896
rect 84556 15856 84598 15896
rect 84638 15856 84680 15896
rect 84720 15856 88352 15896
rect 88392 15856 88434 15896
rect 88474 15856 88516 15896
rect 88556 15856 88598 15896
rect 88638 15856 88680 15896
rect 88720 15856 92352 15896
rect 92392 15856 92434 15896
rect 92474 15856 92516 15896
rect 92556 15856 92598 15896
rect 92638 15856 92680 15896
rect 92720 15856 96352 15896
rect 96392 15856 96434 15896
rect 96474 15856 96516 15896
rect 96556 15856 96598 15896
rect 96638 15856 96680 15896
rect 96720 15856 99360 15896
rect 576 15832 99360 15856
rect 81763 15560 81821 15561
rect 81763 15520 81772 15560
rect 81812 15520 81821 15560
rect 81763 15519 81821 15520
rect 83875 15560 83933 15561
rect 83875 15520 83884 15560
rect 83924 15520 83933 15560
rect 83875 15519 83933 15520
rect 87427 15560 87485 15561
rect 87427 15520 87436 15560
rect 87476 15520 87485 15560
rect 87427 15519 87485 15520
rect 98563 15560 98621 15561
rect 98563 15520 98572 15560
rect 98612 15520 98621 15560
rect 98563 15519 98621 15520
rect 835 15476 893 15477
rect 835 15436 844 15476
rect 884 15436 893 15476
rect 835 15435 893 15436
rect 73699 15476 73757 15477
rect 73699 15436 73708 15476
rect 73748 15436 73757 15476
rect 73699 15435 73757 15436
rect 74275 15476 74333 15477
rect 74275 15436 74284 15476
rect 74324 15436 74333 15476
rect 74275 15435 74333 15436
rect 74851 15476 74909 15477
rect 74851 15436 74860 15476
rect 74900 15436 74909 15476
rect 74851 15435 74909 15436
rect 75331 15476 75389 15477
rect 75331 15436 75340 15476
rect 75380 15436 75389 15476
rect 75331 15435 75389 15436
rect 75811 15476 75869 15477
rect 75811 15436 75820 15476
rect 75860 15436 75869 15476
rect 75811 15435 75869 15436
rect 76195 15476 76253 15477
rect 76195 15436 76204 15476
rect 76244 15436 76253 15476
rect 76195 15435 76253 15436
rect 76579 15476 76637 15477
rect 76579 15436 76588 15476
rect 76628 15436 76637 15476
rect 76579 15435 76637 15436
rect 76963 15476 77021 15477
rect 76963 15436 76972 15476
rect 77012 15436 77021 15476
rect 76963 15435 77021 15436
rect 77347 15476 77405 15477
rect 77347 15436 77356 15476
rect 77396 15436 77405 15476
rect 77347 15435 77405 15436
rect 77731 15476 77789 15477
rect 77731 15436 77740 15476
rect 77780 15436 77789 15476
rect 77731 15435 77789 15436
rect 78115 15476 78173 15477
rect 78115 15436 78124 15476
rect 78164 15436 78173 15476
rect 78115 15435 78173 15436
rect 78595 15476 78653 15477
rect 78595 15436 78604 15476
rect 78644 15436 78653 15476
rect 79363 15476 79421 15477
rect 78595 15435 78653 15436
rect 79170 15465 79228 15466
rect 79170 15425 79179 15465
rect 79219 15425 79228 15465
rect 79363 15436 79372 15476
rect 79412 15436 79421 15476
rect 79363 15435 79421 15436
rect 79747 15476 79805 15477
rect 79747 15436 79756 15476
rect 79796 15436 79805 15476
rect 79747 15435 79805 15436
rect 80227 15476 80285 15477
rect 80227 15436 80236 15476
rect 80276 15436 80285 15476
rect 80227 15435 80285 15436
rect 80707 15476 80765 15477
rect 80707 15436 80716 15476
rect 80756 15436 80765 15476
rect 80707 15435 80765 15436
rect 81091 15476 81149 15477
rect 81091 15436 81100 15476
rect 81140 15436 81149 15476
rect 81091 15435 81149 15436
rect 83011 15476 83069 15477
rect 83011 15436 83020 15476
rect 83060 15436 83069 15476
rect 83011 15435 83069 15436
rect 83395 15476 83453 15477
rect 83395 15436 83404 15476
rect 83444 15436 83453 15476
rect 83395 15435 83453 15436
rect 84163 15476 84221 15477
rect 84163 15436 84172 15476
rect 84212 15436 84221 15476
rect 84163 15435 84221 15436
rect 84547 15476 84605 15477
rect 84547 15436 84556 15476
rect 84596 15436 84605 15476
rect 84547 15435 84605 15436
rect 85027 15476 85085 15477
rect 85027 15436 85036 15476
rect 85076 15436 85085 15476
rect 85027 15435 85085 15436
rect 85411 15476 85469 15477
rect 85411 15436 85420 15476
rect 85460 15436 85469 15476
rect 85411 15435 85469 15436
rect 85795 15476 85853 15477
rect 85795 15436 85804 15476
rect 85844 15436 85853 15476
rect 85795 15435 85853 15436
rect 86179 15476 86237 15477
rect 86179 15436 86188 15476
rect 86228 15436 86237 15476
rect 86179 15435 86237 15436
rect 86563 15476 86621 15477
rect 86563 15436 86572 15476
rect 86612 15436 86621 15476
rect 86563 15435 86621 15436
rect 87043 15476 87101 15477
rect 87043 15436 87052 15476
rect 87092 15436 87101 15476
rect 87043 15435 87101 15436
rect 87907 15476 87965 15477
rect 87907 15436 87916 15476
rect 87956 15436 87965 15476
rect 87907 15435 87965 15436
rect 88291 15476 88349 15477
rect 88291 15436 88300 15476
rect 88340 15436 88349 15476
rect 88291 15435 88349 15436
rect 88675 15476 88733 15477
rect 88675 15436 88684 15476
rect 88724 15436 88733 15476
rect 88675 15435 88733 15436
rect 89059 15476 89117 15477
rect 89059 15436 89068 15476
rect 89108 15436 89117 15476
rect 89059 15435 89117 15436
rect 89443 15476 89501 15477
rect 89443 15436 89452 15476
rect 89492 15436 89501 15476
rect 89443 15435 89501 15436
rect 89827 15476 89885 15477
rect 89827 15436 89836 15476
rect 89876 15436 89885 15476
rect 89827 15435 89885 15436
rect 90499 15476 90557 15477
rect 90499 15436 90508 15476
rect 90548 15436 90557 15476
rect 90499 15435 90557 15436
rect 91075 15476 91133 15477
rect 91075 15436 91084 15476
rect 91124 15436 91133 15476
rect 91075 15435 91133 15436
rect 91459 15476 91517 15477
rect 91459 15436 91468 15476
rect 91508 15436 91517 15476
rect 91459 15435 91517 15436
rect 91939 15476 91997 15477
rect 91939 15436 91948 15476
rect 91988 15436 91997 15476
rect 91939 15435 91997 15436
rect 92515 15476 92573 15477
rect 92515 15436 92524 15476
rect 92564 15436 92573 15476
rect 92515 15435 92573 15436
rect 92707 15476 92765 15477
rect 92707 15436 92716 15476
rect 92756 15436 92765 15476
rect 92707 15435 92765 15436
rect 93379 15476 93437 15477
rect 93379 15436 93388 15476
rect 93428 15436 93437 15476
rect 93379 15435 93437 15436
rect 93763 15476 93821 15477
rect 93763 15436 93772 15476
rect 93812 15436 93821 15476
rect 93763 15435 93821 15436
rect 94243 15476 94301 15477
rect 94243 15436 94252 15476
rect 94292 15436 94301 15476
rect 94243 15435 94301 15436
rect 94627 15476 94685 15477
rect 94627 15436 94636 15476
rect 94676 15436 94685 15476
rect 94627 15435 94685 15436
rect 95011 15476 95069 15477
rect 95011 15436 95020 15476
rect 95060 15436 95069 15476
rect 95011 15435 95069 15436
rect 95683 15476 95741 15477
rect 95683 15436 95692 15476
rect 95732 15436 95741 15476
rect 95683 15435 95741 15436
rect 96067 15476 96125 15477
rect 96067 15436 96076 15476
rect 96116 15436 96125 15476
rect 96067 15435 96125 15436
rect 96451 15476 96509 15477
rect 96451 15436 96460 15476
rect 96500 15436 96509 15476
rect 96451 15435 96509 15436
rect 96835 15476 96893 15477
rect 96835 15436 96844 15476
rect 96884 15436 96893 15476
rect 96835 15435 96893 15436
rect 97219 15476 97277 15477
rect 97219 15436 97228 15476
rect 97268 15436 97277 15476
rect 97219 15435 97277 15436
rect 97603 15476 97661 15477
rect 97603 15436 97612 15476
rect 97652 15436 97661 15476
rect 97603 15435 97661 15436
rect 97987 15476 98045 15477
rect 97987 15436 97996 15476
rect 98036 15436 98045 15476
rect 97987 15435 98045 15436
rect 98371 15476 98429 15477
rect 98371 15436 98380 15476
rect 98420 15436 98429 15476
rect 98371 15435 98429 15436
rect 79170 15424 79228 15425
rect 74091 15392 74133 15401
rect 74091 15352 74092 15392
rect 74132 15352 74133 15392
rect 74091 15343 74133 15352
rect 78795 15392 78837 15401
rect 78795 15352 78796 15392
rect 78836 15352 78837 15392
rect 78795 15343 78837 15352
rect 95499 15392 95541 15401
rect 95499 15352 95500 15392
rect 95540 15352 95541 15392
rect 95499 15343 95541 15352
rect 651 15308 693 15317
rect 651 15268 652 15308
rect 692 15268 693 15308
rect 651 15259 693 15268
rect 73899 15308 73941 15317
rect 73899 15268 73900 15308
rect 73940 15268 73941 15308
rect 73899 15259 73941 15268
rect 75051 15308 75093 15317
rect 75051 15268 75052 15308
rect 75092 15268 75093 15308
rect 75051 15259 75093 15268
rect 75531 15308 75573 15317
rect 75531 15268 75532 15308
rect 75572 15268 75573 15308
rect 75531 15259 75573 15268
rect 76011 15308 76053 15317
rect 76011 15268 76012 15308
rect 76052 15268 76053 15308
rect 76011 15259 76053 15268
rect 76395 15308 76437 15317
rect 76395 15268 76396 15308
rect 76436 15268 76437 15308
rect 76395 15259 76437 15268
rect 76779 15308 76821 15317
rect 76779 15268 76780 15308
rect 76820 15268 76821 15308
rect 76779 15259 76821 15268
rect 77163 15308 77205 15317
rect 77163 15268 77164 15308
rect 77204 15268 77205 15308
rect 77163 15259 77205 15268
rect 77547 15308 77589 15317
rect 77547 15268 77548 15308
rect 77588 15268 77589 15308
rect 77547 15259 77589 15268
rect 77931 15308 77973 15317
rect 77931 15268 77932 15308
rect 77972 15268 77973 15308
rect 77931 15259 77973 15268
rect 78315 15308 78357 15317
rect 78315 15268 78316 15308
rect 78356 15268 78357 15308
rect 78315 15259 78357 15268
rect 78987 15308 79029 15317
rect 78987 15268 78988 15308
rect 79028 15268 79029 15308
rect 78987 15259 79029 15268
rect 79563 15308 79605 15317
rect 79563 15268 79564 15308
rect 79604 15268 79605 15308
rect 79563 15259 79605 15268
rect 79947 15308 79989 15317
rect 79947 15268 79948 15308
rect 79988 15268 79989 15308
rect 79947 15259 79989 15268
rect 80427 15308 80469 15317
rect 80427 15268 80428 15308
rect 80468 15268 80469 15308
rect 80427 15259 80469 15268
rect 80907 15308 80949 15317
rect 80907 15268 80908 15308
rect 80948 15268 80949 15308
rect 80907 15259 80949 15268
rect 81291 15308 81333 15317
rect 81291 15268 81292 15308
rect 81332 15268 81333 15308
rect 81291 15259 81333 15268
rect 81867 15308 81909 15317
rect 81867 15268 81868 15308
rect 81908 15268 81909 15308
rect 81867 15259 81909 15268
rect 83211 15308 83253 15317
rect 83211 15268 83212 15308
rect 83252 15268 83253 15308
rect 83211 15259 83253 15268
rect 83595 15308 83637 15317
rect 83595 15268 83596 15308
rect 83636 15268 83637 15308
rect 83595 15259 83637 15268
rect 83979 15308 84021 15317
rect 83979 15268 83980 15308
rect 84020 15268 84021 15308
rect 83979 15259 84021 15268
rect 84363 15308 84405 15317
rect 84363 15268 84364 15308
rect 84404 15268 84405 15308
rect 84363 15259 84405 15268
rect 84747 15308 84789 15317
rect 84747 15268 84748 15308
rect 84788 15268 84789 15308
rect 84747 15259 84789 15268
rect 85227 15308 85269 15317
rect 85227 15268 85228 15308
rect 85268 15268 85269 15308
rect 85227 15259 85269 15268
rect 85611 15308 85653 15317
rect 85611 15268 85612 15308
rect 85652 15268 85653 15308
rect 85611 15259 85653 15268
rect 85995 15308 86037 15317
rect 85995 15268 85996 15308
rect 86036 15268 86037 15308
rect 85995 15259 86037 15268
rect 86379 15308 86421 15317
rect 86379 15268 86380 15308
rect 86420 15268 86421 15308
rect 86379 15259 86421 15268
rect 86763 15308 86805 15317
rect 86763 15268 86764 15308
rect 86804 15268 86805 15308
rect 86763 15259 86805 15268
rect 87243 15308 87285 15317
rect 87243 15268 87244 15308
rect 87284 15268 87285 15308
rect 87243 15259 87285 15268
rect 87531 15308 87573 15317
rect 87531 15268 87532 15308
rect 87572 15268 87573 15308
rect 87531 15259 87573 15268
rect 88107 15308 88149 15317
rect 88107 15268 88108 15308
rect 88148 15268 88149 15308
rect 88107 15259 88149 15268
rect 88491 15308 88533 15317
rect 88491 15268 88492 15308
rect 88532 15268 88533 15308
rect 88491 15259 88533 15268
rect 88875 15308 88917 15317
rect 88875 15268 88876 15308
rect 88916 15268 88917 15308
rect 88875 15259 88917 15268
rect 89259 15308 89301 15317
rect 89259 15268 89260 15308
rect 89300 15268 89301 15308
rect 89259 15259 89301 15268
rect 89643 15308 89685 15317
rect 89643 15268 89644 15308
rect 89684 15268 89685 15308
rect 89643 15259 89685 15268
rect 90027 15308 90069 15317
rect 90027 15268 90028 15308
rect 90068 15268 90069 15308
rect 90027 15259 90069 15268
rect 90699 15308 90741 15317
rect 90699 15268 90700 15308
rect 90740 15268 90741 15308
rect 90699 15259 90741 15268
rect 90891 15308 90933 15317
rect 90891 15268 90892 15308
rect 90932 15268 90933 15308
rect 90891 15259 90933 15268
rect 91659 15308 91701 15317
rect 91659 15268 91660 15308
rect 91700 15268 91701 15308
rect 91659 15259 91701 15268
rect 92139 15308 92181 15317
rect 92139 15268 92140 15308
rect 92180 15268 92181 15308
rect 92139 15259 92181 15268
rect 92331 15308 92373 15317
rect 92331 15268 92332 15308
rect 92372 15268 92373 15308
rect 92331 15259 92373 15268
rect 92907 15308 92949 15317
rect 92907 15268 92908 15308
rect 92948 15268 92949 15308
rect 92907 15259 92949 15268
rect 93579 15308 93621 15317
rect 93579 15268 93580 15308
rect 93620 15268 93621 15308
rect 93579 15259 93621 15268
rect 93963 15308 94005 15317
rect 93963 15268 93964 15308
rect 94004 15268 94005 15308
rect 93963 15259 94005 15268
rect 94443 15308 94485 15317
rect 94443 15268 94444 15308
rect 94484 15268 94485 15308
rect 94443 15259 94485 15268
rect 94827 15308 94869 15317
rect 94827 15268 94828 15308
rect 94868 15268 94869 15308
rect 94827 15259 94869 15268
rect 95211 15308 95253 15317
rect 95211 15268 95212 15308
rect 95252 15268 95253 15308
rect 95211 15259 95253 15268
rect 95883 15308 95925 15317
rect 95883 15268 95884 15308
rect 95924 15268 95925 15308
rect 95883 15259 95925 15268
rect 96267 15308 96309 15317
rect 96267 15268 96268 15308
rect 96308 15268 96309 15308
rect 96267 15259 96309 15268
rect 96651 15308 96693 15317
rect 96651 15268 96652 15308
rect 96692 15268 96693 15308
rect 96651 15259 96693 15268
rect 97035 15308 97077 15317
rect 97035 15268 97036 15308
rect 97076 15268 97077 15308
rect 97035 15259 97077 15268
rect 97419 15308 97461 15317
rect 97419 15268 97420 15308
rect 97460 15268 97461 15308
rect 97419 15259 97461 15268
rect 97803 15308 97845 15317
rect 97803 15268 97804 15308
rect 97844 15268 97845 15308
rect 97803 15259 97845 15268
rect 98187 15308 98229 15317
rect 98187 15268 98188 15308
rect 98228 15268 98229 15308
rect 98187 15259 98229 15268
rect 98667 15308 98709 15317
rect 98667 15268 98668 15308
rect 98708 15268 98709 15308
rect 98667 15259 98709 15268
rect 576 15140 99360 15164
rect 576 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 7112 15140
rect 7152 15100 7194 15140
rect 7234 15100 7276 15140
rect 7316 15100 7358 15140
rect 7398 15100 7440 15140
rect 7480 15100 11112 15140
rect 11152 15100 11194 15140
rect 11234 15100 11276 15140
rect 11316 15100 11358 15140
rect 11398 15100 11440 15140
rect 11480 15100 15112 15140
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15480 15100 19112 15140
rect 19152 15100 19194 15140
rect 19234 15100 19276 15140
rect 19316 15100 19358 15140
rect 19398 15100 19440 15140
rect 19480 15100 23112 15140
rect 23152 15100 23194 15140
rect 23234 15100 23276 15140
rect 23316 15100 23358 15140
rect 23398 15100 23440 15140
rect 23480 15100 27112 15140
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27480 15100 31112 15140
rect 31152 15100 31194 15140
rect 31234 15100 31276 15140
rect 31316 15100 31358 15140
rect 31398 15100 31440 15140
rect 31480 15100 35112 15140
rect 35152 15100 35194 15140
rect 35234 15100 35276 15140
rect 35316 15100 35358 15140
rect 35398 15100 35440 15140
rect 35480 15100 39112 15140
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39480 15100 43112 15140
rect 43152 15100 43194 15140
rect 43234 15100 43276 15140
rect 43316 15100 43358 15140
rect 43398 15100 43440 15140
rect 43480 15100 47112 15140
rect 47152 15100 47194 15140
rect 47234 15100 47276 15140
rect 47316 15100 47358 15140
rect 47398 15100 47440 15140
rect 47480 15100 51112 15140
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51480 15100 55112 15140
rect 55152 15100 55194 15140
rect 55234 15100 55276 15140
rect 55316 15100 55358 15140
rect 55398 15100 55440 15140
rect 55480 15100 59112 15140
rect 59152 15100 59194 15140
rect 59234 15100 59276 15140
rect 59316 15100 59358 15140
rect 59398 15100 59440 15140
rect 59480 15100 63112 15140
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63480 15100 67112 15140
rect 67152 15100 67194 15140
rect 67234 15100 67276 15140
rect 67316 15100 67358 15140
rect 67398 15100 67440 15140
rect 67480 15100 99360 15140
rect 576 15076 99360 15100
rect 1419 14972 1461 14981
rect 1419 14932 1420 14972
rect 1460 14932 1461 14972
rect 1419 14923 1461 14932
rect 73707 14888 73749 14897
rect 73707 14848 73708 14888
rect 73748 14848 73749 14888
rect 73707 14839 73749 14848
rect 835 14804 893 14805
rect 835 14764 844 14804
rect 884 14764 893 14804
rect 835 14763 893 14764
rect 1603 14804 1661 14805
rect 1603 14764 1612 14804
rect 1652 14764 1661 14804
rect 1603 14763 1661 14764
rect 1987 14804 2045 14805
rect 1987 14764 1996 14804
rect 2036 14764 2045 14804
rect 1987 14763 2045 14764
rect 73027 14804 73085 14805
rect 73027 14764 73036 14804
rect 73076 14764 73085 14804
rect 73027 14763 73085 14764
rect 73507 14804 73565 14805
rect 73507 14764 73516 14804
rect 73556 14764 73565 14804
rect 73507 14763 73565 14764
rect 74467 14804 74525 14805
rect 74467 14764 74476 14804
rect 74516 14764 74525 14804
rect 74467 14763 74525 14764
rect 78883 14804 78941 14805
rect 78883 14764 78892 14804
rect 78932 14764 78941 14804
rect 78883 14763 78941 14764
rect 82243 14804 82301 14805
rect 82243 14764 82252 14804
rect 82292 14764 82301 14804
rect 82243 14763 82301 14764
rect 91075 14804 91133 14805
rect 91075 14764 91084 14804
rect 91124 14764 91133 14804
rect 91075 14763 91133 14764
rect 92995 14804 93053 14805
rect 92995 14764 93004 14804
rect 93044 14764 93053 14804
rect 92995 14763 93053 14764
rect 96835 14804 96893 14805
rect 96835 14764 96844 14804
rect 96884 14764 96893 14804
rect 96835 14763 96893 14764
rect 98755 14804 98813 14805
rect 98755 14764 98764 14804
rect 98804 14764 98813 14804
rect 98755 14763 98813 14764
rect 92419 14733 92477 14734
rect 72739 14720 72797 14721
rect 72739 14680 72748 14720
rect 72788 14680 72797 14720
rect 72739 14679 72797 14680
rect 73891 14720 73949 14721
rect 73891 14680 73900 14720
rect 73940 14680 73949 14720
rect 73891 14679 73949 14680
rect 74179 14720 74237 14721
rect 74179 14680 74188 14720
rect 74228 14680 74237 14720
rect 74179 14679 74237 14680
rect 74851 14720 74909 14721
rect 74851 14680 74860 14720
rect 74900 14680 74909 14720
rect 74851 14679 74909 14680
rect 75331 14720 75389 14721
rect 75331 14680 75340 14720
rect 75380 14680 75389 14720
rect 75331 14679 75389 14680
rect 75811 14720 75869 14721
rect 75811 14680 75820 14720
rect 75860 14680 75869 14720
rect 75811 14679 75869 14680
rect 76099 14720 76157 14721
rect 76099 14680 76108 14720
rect 76148 14680 76157 14720
rect 76099 14679 76157 14680
rect 76579 14720 76637 14721
rect 76579 14680 76588 14720
rect 76628 14680 76637 14720
rect 76579 14679 76637 14680
rect 76963 14720 77021 14721
rect 76963 14680 76972 14720
rect 77012 14680 77021 14720
rect 76963 14679 77021 14680
rect 77347 14720 77405 14721
rect 77347 14680 77356 14720
rect 77396 14680 77405 14720
rect 77347 14679 77405 14680
rect 77827 14720 77885 14721
rect 77827 14680 77836 14720
rect 77876 14680 77885 14720
rect 77827 14679 77885 14680
rect 78115 14720 78173 14721
rect 78115 14680 78124 14720
rect 78164 14680 78173 14720
rect 78115 14679 78173 14680
rect 78691 14720 78749 14721
rect 78691 14680 78700 14720
rect 78740 14680 78749 14720
rect 78691 14679 78749 14680
rect 79363 14720 79421 14721
rect 79363 14680 79372 14720
rect 79412 14680 79421 14720
rect 79363 14679 79421 14680
rect 79651 14720 79709 14721
rect 79651 14680 79660 14720
rect 79700 14680 79709 14720
rect 79651 14679 79709 14680
rect 80131 14720 80189 14721
rect 80131 14680 80140 14720
rect 80180 14680 80189 14720
rect 80131 14679 80189 14680
rect 80419 14720 80477 14721
rect 80419 14680 80428 14720
rect 80468 14680 80477 14720
rect 80419 14679 80477 14680
rect 80803 14720 80861 14721
rect 80803 14680 80812 14720
rect 80852 14680 80861 14720
rect 80803 14679 80861 14680
rect 80995 14720 81053 14721
rect 80995 14680 81004 14720
rect 81044 14680 81053 14720
rect 80995 14679 81053 14680
rect 81379 14720 81437 14721
rect 81379 14680 81388 14720
rect 81428 14680 81437 14720
rect 81379 14679 81437 14680
rect 81955 14720 82013 14721
rect 81955 14680 81964 14720
rect 82004 14680 82013 14720
rect 81955 14679 82013 14680
rect 82627 14720 82685 14721
rect 82627 14680 82636 14720
rect 82676 14680 82685 14720
rect 82627 14679 82685 14680
rect 83011 14720 83069 14721
rect 83011 14680 83020 14720
rect 83060 14680 83069 14720
rect 83011 14679 83069 14680
rect 83395 14720 83453 14721
rect 83395 14680 83404 14720
rect 83444 14680 83453 14720
rect 83395 14679 83453 14680
rect 83779 14720 83837 14721
rect 83779 14680 83788 14720
rect 83828 14680 83837 14720
rect 83779 14679 83837 14680
rect 84547 14720 84605 14721
rect 84547 14680 84556 14720
rect 84596 14680 84605 14720
rect 84547 14679 84605 14680
rect 85027 14720 85085 14721
rect 85027 14680 85036 14720
rect 85076 14680 85085 14720
rect 85027 14679 85085 14680
rect 85411 14720 85469 14721
rect 85411 14680 85420 14720
rect 85460 14680 85469 14720
rect 85411 14679 85469 14680
rect 85795 14720 85853 14721
rect 85795 14680 85804 14720
rect 85844 14680 85853 14720
rect 85795 14679 85853 14680
rect 86371 14720 86429 14721
rect 86371 14680 86380 14720
rect 86420 14680 86429 14720
rect 86371 14679 86429 14680
rect 86755 14720 86813 14721
rect 86755 14680 86764 14720
rect 86804 14680 86813 14720
rect 86755 14679 86813 14680
rect 87043 14720 87101 14721
rect 87043 14680 87052 14720
rect 87092 14680 87101 14720
rect 87043 14679 87101 14680
rect 87907 14720 87965 14721
rect 87907 14680 87916 14720
rect 87956 14680 87965 14720
rect 87907 14679 87965 14680
rect 88195 14720 88253 14721
rect 88195 14680 88204 14720
rect 88244 14680 88253 14720
rect 88195 14679 88253 14680
rect 88579 14720 88637 14721
rect 88579 14680 88588 14720
rect 88628 14680 88637 14720
rect 88579 14679 88637 14680
rect 88963 14720 89021 14721
rect 88963 14680 88972 14720
rect 89012 14680 89021 14720
rect 88963 14679 89021 14680
rect 89635 14720 89693 14721
rect 89635 14680 89644 14720
rect 89684 14680 89693 14720
rect 89635 14679 89693 14680
rect 90019 14720 90077 14721
rect 90019 14680 90028 14720
rect 90068 14680 90077 14720
rect 90019 14679 90077 14680
rect 90211 14720 90269 14721
rect 90211 14680 90220 14720
rect 90260 14680 90269 14720
rect 90211 14679 90269 14680
rect 90595 14720 90653 14721
rect 90595 14680 90604 14720
rect 90644 14680 90653 14720
rect 90595 14679 90653 14680
rect 91555 14720 91613 14721
rect 91555 14680 91564 14720
rect 91604 14680 91613 14720
rect 91555 14679 91613 14680
rect 91747 14720 91805 14721
rect 91747 14680 91756 14720
rect 91796 14680 91805 14720
rect 91747 14679 91805 14680
rect 92131 14720 92189 14721
rect 92131 14680 92140 14720
rect 92180 14680 92189 14720
rect 92419 14693 92428 14733
rect 92468 14693 92477 14733
rect 92419 14692 92477 14693
rect 92707 14720 92765 14721
rect 92131 14679 92189 14680
rect 92707 14680 92716 14720
rect 92756 14680 92765 14720
rect 92707 14679 92765 14680
rect 93379 14720 93437 14721
rect 93379 14680 93388 14720
rect 93428 14680 93437 14720
rect 93379 14679 93437 14680
rect 93955 14720 94013 14721
rect 93955 14680 93964 14720
rect 94004 14680 94013 14720
rect 93955 14679 94013 14680
rect 94243 14720 94301 14721
rect 94243 14680 94252 14720
rect 94292 14680 94301 14720
rect 94243 14679 94301 14680
rect 94627 14720 94685 14721
rect 94627 14680 94636 14720
rect 94676 14680 94685 14720
rect 94627 14679 94685 14680
rect 95011 14720 95069 14721
rect 95011 14680 95020 14720
rect 95060 14680 95069 14720
rect 95011 14679 95069 14680
rect 95491 14720 95549 14721
rect 95491 14680 95500 14720
rect 95540 14680 95549 14720
rect 95491 14679 95549 14680
rect 95971 14720 96029 14721
rect 95971 14680 95980 14720
rect 96020 14680 96029 14720
rect 95971 14679 96029 14680
rect 96355 14720 96413 14721
rect 96355 14680 96364 14720
rect 96404 14680 96413 14720
rect 96355 14679 96413 14680
rect 97123 14720 97181 14721
rect 97123 14680 97132 14720
rect 97172 14680 97181 14720
rect 97123 14679 97181 14680
rect 97411 14720 97469 14721
rect 97411 14680 97420 14720
rect 97460 14680 97469 14720
rect 97411 14679 97469 14680
rect 97699 14720 97757 14721
rect 97699 14680 97708 14720
rect 97748 14680 97757 14720
rect 97699 14679 97757 14680
rect 98371 14720 98429 14721
rect 98371 14680 98380 14720
rect 98420 14680 98429 14720
rect 98371 14679 98429 14680
rect 651 14552 693 14561
rect 651 14512 652 14552
rect 692 14512 693 14552
rect 651 14503 693 14512
rect 1803 14552 1845 14561
rect 1803 14512 1804 14552
rect 1844 14512 1845 14552
rect 1803 14503 1845 14512
rect 72843 14552 72885 14561
rect 72843 14512 72844 14552
rect 72884 14512 72885 14552
rect 72843 14503 72885 14512
rect 73227 14552 73269 14561
rect 73227 14512 73228 14552
rect 73268 14512 73269 14552
rect 73227 14503 73269 14512
rect 73995 14552 74037 14561
rect 73995 14512 73996 14552
rect 74036 14512 74037 14552
rect 73995 14503 74037 14512
rect 74283 14552 74325 14561
rect 74283 14512 74284 14552
rect 74324 14512 74325 14552
rect 74283 14503 74325 14512
rect 74667 14552 74709 14561
rect 74667 14512 74668 14552
rect 74708 14512 74709 14552
rect 74667 14503 74709 14512
rect 74955 14552 74997 14561
rect 74955 14512 74956 14552
rect 74996 14512 74997 14552
rect 74955 14503 74997 14512
rect 75435 14552 75477 14561
rect 75435 14512 75436 14552
rect 75476 14512 75477 14552
rect 75435 14503 75477 14512
rect 75915 14552 75957 14561
rect 75915 14512 75916 14552
rect 75956 14512 75957 14552
rect 75915 14503 75957 14512
rect 76203 14552 76245 14561
rect 76203 14512 76204 14552
rect 76244 14512 76245 14552
rect 76203 14503 76245 14512
rect 76683 14552 76725 14561
rect 76683 14512 76684 14552
rect 76724 14512 76725 14552
rect 76683 14503 76725 14512
rect 77067 14552 77109 14561
rect 77067 14512 77068 14552
rect 77108 14512 77109 14552
rect 77067 14503 77109 14512
rect 77451 14552 77493 14561
rect 77451 14512 77452 14552
rect 77492 14512 77493 14552
rect 77451 14503 77493 14512
rect 77931 14552 77973 14561
rect 77931 14512 77932 14552
rect 77972 14512 77973 14552
rect 77931 14503 77973 14512
rect 78219 14552 78261 14561
rect 78219 14512 78220 14552
rect 78260 14512 78261 14552
rect 78219 14503 78261 14512
rect 78603 14552 78645 14561
rect 78603 14512 78604 14552
rect 78644 14512 78645 14552
rect 78603 14503 78645 14512
rect 79083 14552 79125 14561
rect 79083 14512 79084 14552
rect 79124 14512 79125 14552
rect 79083 14503 79125 14512
rect 79467 14552 79509 14561
rect 79467 14512 79468 14552
rect 79508 14512 79509 14552
rect 79467 14503 79509 14512
rect 79755 14552 79797 14561
rect 79755 14512 79756 14552
rect 79796 14512 79797 14552
rect 79755 14503 79797 14512
rect 80235 14552 80277 14561
rect 80235 14512 80236 14552
rect 80276 14512 80277 14552
rect 80235 14503 80277 14512
rect 80523 14552 80565 14561
rect 80523 14512 80524 14552
rect 80564 14512 80565 14552
rect 80523 14503 80565 14512
rect 80715 14552 80757 14561
rect 80715 14512 80716 14552
rect 80756 14512 80757 14552
rect 80715 14503 80757 14512
rect 81099 14552 81141 14561
rect 81099 14512 81100 14552
rect 81140 14512 81141 14552
rect 81099 14503 81141 14512
rect 81483 14552 81525 14561
rect 81483 14512 81484 14552
rect 81524 14512 81525 14552
rect 81483 14503 81525 14512
rect 82059 14552 82101 14561
rect 82059 14512 82060 14552
rect 82100 14512 82101 14552
rect 82059 14503 82101 14512
rect 82443 14552 82485 14561
rect 82443 14512 82444 14552
rect 82484 14512 82485 14552
rect 82443 14503 82485 14512
rect 82731 14552 82773 14561
rect 82731 14512 82732 14552
rect 82772 14512 82773 14552
rect 82731 14503 82773 14512
rect 83115 14552 83157 14561
rect 83115 14512 83116 14552
rect 83156 14512 83157 14552
rect 83115 14503 83157 14512
rect 83499 14552 83541 14561
rect 83499 14512 83500 14552
rect 83540 14512 83541 14552
rect 83499 14503 83541 14512
rect 83883 14552 83925 14561
rect 83883 14512 83884 14552
rect 83924 14512 83925 14552
rect 83883 14503 83925 14512
rect 84651 14552 84693 14561
rect 84651 14512 84652 14552
rect 84692 14512 84693 14552
rect 84651 14503 84693 14512
rect 85131 14552 85173 14561
rect 85131 14512 85132 14552
rect 85172 14512 85173 14552
rect 85131 14503 85173 14512
rect 85515 14552 85557 14561
rect 85515 14512 85516 14552
rect 85556 14512 85557 14552
rect 85515 14503 85557 14512
rect 85899 14552 85941 14561
rect 85899 14512 85900 14552
rect 85940 14512 85941 14552
rect 85899 14503 85941 14512
rect 86283 14552 86325 14561
rect 86283 14512 86284 14552
rect 86324 14512 86325 14552
rect 86283 14503 86325 14512
rect 86667 14552 86709 14561
rect 86667 14512 86668 14552
rect 86708 14512 86709 14552
rect 86667 14503 86709 14512
rect 87147 14552 87189 14561
rect 87147 14512 87148 14552
rect 87188 14512 87189 14552
rect 87147 14503 87189 14512
rect 87819 14552 87861 14561
rect 87819 14512 87820 14552
rect 87860 14512 87861 14552
rect 87819 14503 87861 14512
rect 88299 14552 88341 14561
rect 88299 14512 88300 14552
rect 88340 14512 88341 14552
rect 88299 14503 88341 14512
rect 88683 14552 88725 14561
rect 88683 14512 88684 14552
rect 88724 14512 88725 14552
rect 88683 14503 88725 14512
rect 89067 14552 89109 14561
rect 89067 14512 89068 14552
rect 89108 14512 89109 14552
rect 89067 14503 89109 14512
rect 89547 14552 89589 14561
rect 89547 14512 89548 14552
rect 89588 14512 89589 14552
rect 89547 14503 89589 14512
rect 89931 14552 89973 14561
rect 89931 14512 89932 14552
rect 89972 14512 89973 14552
rect 89931 14503 89973 14512
rect 90315 14552 90357 14561
rect 90315 14512 90316 14552
rect 90356 14512 90357 14552
rect 90315 14503 90357 14512
rect 90699 14552 90741 14561
rect 90699 14512 90700 14552
rect 90740 14512 90741 14552
rect 90699 14503 90741 14512
rect 91275 14552 91317 14561
rect 91275 14512 91276 14552
rect 91316 14512 91317 14552
rect 91275 14503 91317 14512
rect 91467 14552 91509 14561
rect 91467 14512 91468 14552
rect 91508 14512 91509 14552
rect 91467 14503 91509 14512
rect 91851 14552 91893 14561
rect 91851 14512 91852 14552
rect 91892 14512 91893 14552
rect 91851 14503 91893 14512
rect 92235 14552 92277 14561
rect 92235 14512 92236 14552
rect 92276 14512 92277 14552
rect 92235 14503 92277 14512
rect 92523 14552 92565 14561
rect 92523 14512 92524 14552
rect 92564 14512 92565 14552
rect 92523 14503 92565 14512
rect 92811 14552 92853 14561
rect 92811 14512 92812 14552
rect 92852 14512 92853 14552
rect 92811 14503 92853 14512
rect 93195 14552 93237 14561
rect 93195 14512 93196 14552
rect 93236 14512 93237 14552
rect 93195 14503 93237 14512
rect 93483 14552 93525 14561
rect 93483 14512 93484 14552
rect 93524 14512 93525 14552
rect 93483 14503 93525 14512
rect 93867 14552 93909 14561
rect 93867 14512 93868 14552
rect 93908 14512 93909 14552
rect 93867 14503 93909 14512
rect 94347 14552 94389 14561
rect 94347 14512 94348 14552
rect 94388 14512 94389 14552
rect 94347 14503 94389 14512
rect 94731 14552 94773 14561
rect 94731 14512 94732 14552
rect 94772 14512 94773 14552
rect 94731 14503 94773 14512
rect 95115 14552 95157 14561
rect 95115 14512 95116 14552
rect 95156 14512 95157 14552
rect 95115 14503 95157 14512
rect 95403 14552 95445 14561
rect 95403 14512 95404 14552
rect 95444 14512 95445 14552
rect 95403 14503 95445 14512
rect 95883 14552 95925 14561
rect 95883 14512 95884 14552
rect 95924 14512 95925 14552
rect 95883 14503 95925 14512
rect 96267 14552 96309 14561
rect 96267 14512 96268 14552
rect 96308 14512 96309 14552
rect 96267 14503 96309 14512
rect 96651 14552 96693 14561
rect 96651 14512 96652 14552
rect 96692 14512 96693 14552
rect 96651 14503 96693 14512
rect 97035 14552 97077 14561
rect 97035 14512 97036 14552
rect 97076 14512 97077 14552
rect 97035 14503 97077 14512
rect 97515 14552 97557 14561
rect 97515 14512 97516 14552
rect 97556 14512 97557 14552
rect 97515 14503 97557 14512
rect 97803 14552 97845 14561
rect 97803 14512 97804 14552
rect 97844 14512 97845 14552
rect 97803 14503 97845 14512
rect 98283 14552 98325 14561
rect 98283 14512 98284 14552
rect 98324 14512 98325 14552
rect 98283 14503 98325 14512
rect 98571 14552 98613 14561
rect 98571 14512 98572 14552
rect 98612 14512 98613 14552
rect 98571 14503 98613 14512
rect 576 14384 99360 14408
rect 576 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 8352 14384
rect 8392 14344 8434 14384
rect 8474 14344 8516 14384
rect 8556 14344 8598 14384
rect 8638 14344 8680 14384
rect 8720 14344 12352 14384
rect 12392 14344 12434 14384
rect 12474 14344 12516 14384
rect 12556 14344 12598 14384
rect 12638 14344 12680 14384
rect 12720 14344 16352 14384
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16720 14344 20352 14384
rect 20392 14344 20434 14384
rect 20474 14344 20516 14384
rect 20556 14344 20598 14384
rect 20638 14344 20680 14384
rect 20720 14344 24352 14384
rect 24392 14344 24434 14384
rect 24474 14344 24516 14384
rect 24556 14344 24598 14384
rect 24638 14344 24680 14384
rect 24720 14344 28352 14384
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28720 14344 32352 14384
rect 32392 14344 32434 14384
rect 32474 14344 32516 14384
rect 32556 14344 32598 14384
rect 32638 14344 32680 14384
rect 32720 14344 36352 14384
rect 36392 14344 36434 14384
rect 36474 14344 36516 14384
rect 36556 14344 36598 14384
rect 36638 14344 36680 14384
rect 36720 14344 40352 14384
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40720 14344 44352 14384
rect 44392 14344 44434 14384
rect 44474 14344 44516 14384
rect 44556 14344 44598 14384
rect 44638 14344 44680 14384
rect 44720 14344 48352 14384
rect 48392 14344 48434 14384
rect 48474 14344 48516 14384
rect 48556 14344 48598 14384
rect 48638 14344 48680 14384
rect 48720 14344 52352 14384
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52720 14344 56352 14384
rect 56392 14344 56434 14384
rect 56474 14344 56516 14384
rect 56556 14344 56598 14384
rect 56638 14344 56680 14384
rect 56720 14344 60352 14384
rect 60392 14344 60434 14384
rect 60474 14344 60516 14384
rect 60556 14344 60598 14384
rect 60638 14344 60680 14384
rect 60720 14344 64352 14384
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64720 14344 68352 14384
rect 68392 14344 68434 14384
rect 68474 14344 68516 14384
rect 68556 14344 68598 14384
rect 68638 14344 68680 14384
rect 68720 14344 99360 14384
rect 576 14320 99360 14344
rect 1035 14216 1077 14225
rect 1035 14176 1036 14216
rect 1076 14176 1077 14216
rect 1035 14167 1077 14176
rect 70627 14048 70685 14049
rect 70627 14008 70636 14048
rect 70676 14008 70685 14048
rect 70627 14007 70685 14008
rect 70819 14048 70877 14049
rect 70819 14008 70828 14048
rect 70868 14008 70877 14048
rect 70819 14007 70877 14008
rect 71299 14048 71357 14049
rect 71299 14008 71308 14048
rect 71348 14008 71357 14048
rect 71299 14007 71357 14008
rect 1219 13964 1277 13965
rect 1219 13924 1228 13964
rect 1268 13924 1277 13964
rect 1219 13923 1277 13924
rect 71403 13880 71445 13889
rect 71403 13840 71404 13880
rect 71444 13840 71445 13880
rect 71403 13831 71445 13840
rect 576 13628 71520 13652
rect 576 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 7112 13628
rect 7152 13588 7194 13628
rect 7234 13588 7276 13628
rect 7316 13588 7358 13628
rect 7398 13588 7440 13628
rect 7480 13588 11112 13628
rect 11152 13588 11194 13628
rect 11234 13588 11276 13628
rect 11316 13588 11358 13628
rect 11398 13588 11440 13628
rect 11480 13588 15112 13628
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15480 13588 19112 13628
rect 19152 13588 19194 13628
rect 19234 13588 19276 13628
rect 19316 13588 19358 13628
rect 19398 13588 19440 13628
rect 19480 13588 23112 13628
rect 23152 13588 23194 13628
rect 23234 13588 23276 13628
rect 23316 13588 23358 13628
rect 23398 13588 23440 13628
rect 23480 13588 27112 13628
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27480 13588 31112 13628
rect 31152 13588 31194 13628
rect 31234 13588 31276 13628
rect 31316 13588 31358 13628
rect 31398 13588 31440 13628
rect 31480 13588 35112 13628
rect 35152 13588 35194 13628
rect 35234 13588 35276 13628
rect 35316 13588 35358 13628
rect 35398 13588 35440 13628
rect 35480 13588 39112 13628
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39480 13588 43112 13628
rect 43152 13588 43194 13628
rect 43234 13588 43276 13628
rect 43316 13588 43358 13628
rect 43398 13588 43440 13628
rect 43480 13588 47112 13628
rect 47152 13588 47194 13628
rect 47234 13588 47276 13628
rect 47316 13588 47358 13628
rect 47398 13588 47440 13628
rect 47480 13588 51112 13628
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51480 13588 55112 13628
rect 55152 13588 55194 13628
rect 55234 13588 55276 13628
rect 55316 13588 55358 13628
rect 55398 13588 55440 13628
rect 55480 13588 59112 13628
rect 59152 13588 59194 13628
rect 59234 13588 59276 13628
rect 59316 13588 59358 13628
rect 59398 13588 59440 13628
rect 59480 13588 63112 13628
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63480 13588 67112 13628
rect 67152 13588 67194 13628
rect 67234 13588 67276 13628
rect 67316 13588 67358 13628
rect 67398 13588 67440 13628
rect 67480 13588 71520 13628
rect 576 13564 71520 13588
rect 70059 13460 70101 13469
rect 70059 13420 70060 13460
rect 70100 13420 70101 13460
rect 70059 13411 70101 13420
rect 70923 13460 70965 13469
rect 70923 13420 70924 13460
rect 70964 13420 70965 13460
rect 70923 13411 70965 13420
rect 71307 13460 71349 13469
rect 71307 13420 71308 13460
rect 71348 13420 71349 13460
rect 71307 13411 71349 13420
rect 1611 13376 1653 13385
rect 1611 13336 1612 13376
rect 1652 13336 1653 13376
rect 1611 13327 1653 13336
rect 835 13292 893 13293
rect 835 13252 844 13292
rect 884 13252 893 13292
rect 835 13251 893 13252
rect 1795 13292 1853 13293
rect 1795 13252 1804 13292
rect 1844 13252 1853 13292
rect 1795 13251 1853 13252
rect 69859 13292 69917 13293
rect 69859 13252 69868 13292
rect 69908 13252 69917 13292
rect 69859 13251 69917 13252
rect 70723 13292 70781 13293
rect 70723 13252 70732 13292
rect 70772 13252 70781 13292
rect 70723 13251 70781 13252
rect 71107 13292 71165 13293
rect 71107 13252 71116 13292
rect 71156 13252 71165 13292
rect 71107 13251 71165 13252
rect 70339 13208 70397 13209
rect 70339 13168 70348 13208
rect 70388 13168 70397 13208
rect 70339 13167 70397 13168
rect 70531 13208 70589 13209
rect 70531 13168 70540 13208
rect 70580 13168 70589 13208
rect 70531 13167 70589 13168
rect 651 13040 693 13049
rect 651 13000 652 13040
rect 692 13000 693 13040
rect 651 12991 693 13000
rect 576 12872 71520 12896
rect 576 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 8352 12872
rect 8392 12832 8434 12872
rect 8474 12832 8516 12872
rect 8556 12832 8598 12872
rect 8638 12832 8680 12872
rect 8720 12832 12352 12872
rect 12392 12832 12434 12872
rect 12474 12832 12516 12872
rect 12556 12832 12598 12872
rect 12638 12832 12680 12872
rect 12720 12832 16352 12872
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16720 12832 20352 12872
rect 20392 12832 20434 12872
rect 20474 12832 20516 12872
rect 20556 12832 20598 12872
rect 20638 12832 20680 12872
rect 20720 12832 24352 12872
rect 24392 12832 24434 12872
rect 24474 12832 24516 12872
rect 24556 12832 24598 12872
rect 24638 12832 24680 12872
rect 24720 12832 28352 12872
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28720 12832 32352 12872
rect 32392 12832 32434 12872
rect 32474 12832 32516 12872
rect 32556 12832 32598 12872
rect 32638 12832 32680 12872
rect 32720 12832 36352 12872
rect 36392 12832 36434 12872
rect 36474 12832 36516 12872
rect 36556 12832 36598 12872
rect 36638 12832 36680 12872
rect 36720 12832 40352 12872
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40720 12832 44352 12872
rect 44392 12832 44434 12872
rect 44474 12832 44516 12872
rect 44556 12832 44598 12872
rect 44638 12832 44680 12872
rect 44720 12832 48352 12872
rect 48392 12832 48434 12872
rect 48474 12832 48516 12872
rect 48556 12832 48598 12872
rect 48638 12832 48680 12872
rect 48720 12832 52352 12872
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52720 12832 56352 12872
rect 56392 12832 56434 12872
rect 56474 12832 56516 12872
rect 56556 12832 56598 12872
rect 56638 12832 56680 12872
rect 56720 12832 60352 12872
rect 60392 12832 60434 12872
rect 60474 12832 60516 12872
rect 60556 12832 60598 12872
rect 60638 12832 60680 12872
rect 60720 12832 64352 12872
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64720 12832 68352 12872
rect 68392 12832 68434 12872
rect 68474 12832 68516 12872
rect 68556 12832 68598 12872
rect 68638 12832 68680 12872
rect 68720 12832 71520 12872
rect 576 12808 71520 12832
rect 70539 12620 70581 12629
rect 70539 12580 70540 12620
rect 70580 12580 70581 12620
rect 70539 12571 70581 12580
rect 70923 12620 70965 12629
rect 70923 12580 70924 12620
rect 70964 12580 70965 12620
rect 70923 12571 70965 12580
rect 71211 12620 71253 12629
rect 71211 12580 71212 12620
rect 71252 12580 71253 12620
rect 71211 12571 71253 12580
rect 70435 12536 70493 12537
rect 70435 12496 70444 12536
rect 70484 12496 70493 12536
rect 70435 12495 70493 12496
rect 70819 12536 70877 12537
rect 70819 12496 70828 12536
rect 70868 12496 70877 12536
rect 70819 12495 70877 12496
rect 71107 12536 71165 12537
rect 71107 12496 71116 12536
rect 71156 12496 71165 12536
rect 71107 12495 71165 12496
rect 835 12452 893 12453
rect 835 12412 844 12452
rect 884 12412 893 12452
rect 835 12411 893 12412
rect 1411 12452 1469 12453
rect 1411 12412 1420 12452
rect 1460 12412 1469 12452
rect 1411 12411 1469 12412
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 651 12319 693 12328
rect 1227 12368 1269 12377
rect 1227 12328 1228 12368
rect 1268 12328 1269 12368
rect 1227 12319 1269 12328
rect 576 12116 71520 12140
rect 576 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 7112 12116
rect 7152 12076 7194 12116
rect 7234 12076 7276 12116
rect 7316 12076 7358 12116
rect 7398 12076 7440 12116
rect 7480 12076 11112 12116
rect 11152 12076 11194 12116
rect 11234 12076 11276 12116
rect 11316 12076 11358 12116
rect 11398 12076 11440 12116
rect 11480 12076 15112 12116
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15480 12076 19112 12116
rect 19152 12076 19194 12116
rect 19234 12076 19276 12116
rect 19316 12076 19358 12116
rect 19398 12076 19440 12116
rect 19480 12076 23112 12116
rect 23152 12076 23194 12116
rect 23234 12076 23276 12116
rect 23316 12076 23358 12116
rect 23398 12076 23440 12116
rect 23480 12076 27112 12116
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27480 12076 31112 12116
rect 31152 12076 31194 12116
rect 31234 12076 31276 12116
rect 31316 12076 31358 12116
rect 31398 12076 31440 12116
rect 31480 12076 35112 12116
rect 35152 12076 35194 12116
rect 35234 12076 35276 12116
rect 35316 12076 35358 12116
rect 35398 12076 35440 12116
rect 35480 12076 39112 12116
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39480 12076 43112 12116
rect 43152 12076 43194 12116
rect 43234 12076 43276 12116
rect 43316 12076 43358 12116
rect 43398 12076 43440 12116
rect 43480 12076 47112 12116
rect 47152 12076 47194 12116
rect 47234 12076 47276 12116
rect 47316 12076 47358 12116
rect 47398 12076 47440 12116
rect 47480 12076 51112 12116
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51480 12076 55112 12116
rect 55152 12076 55194 12116
rect 55234 12076 55276 12116
rect 55316 12076 55358 12116
rect 55398 12076 55440 12116
rect 55480 12076 59112 12116
rect 59152 12076 59194 12116
rect 59234 12076 59276 12116
rect 59316 12076 59358 12116
rect 59398 12076 59440 12116
rect 59480 12076 63112 12116
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63480 12076 67112 12116
rect 67152 12076 67194 12116
rect 67234 12076 67276 12116
rect 67316 12076 67358 12116
rect 67398 12076 67440 12116
rect 67480 12076 71520 12116
rect 576 12052 71520 12076
rect 835 11780 893 11781
rect 835 11740 844 11780
rect 884 11740 893 11780
rect 835 11739 893 11740
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 576 11360 71520 11384
rect 576 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 8352 11360
rect 8392 11320 8434 11360
rect 8474 11320 8516 11360
rect 8556 11320 8598 11360
rect 8638 11320 8680 11360
rect 8720 11320 12352 11360
rect 12392 11320 12434 11360
rect 12474 11320 12516 11360
rect 12556 11320 12598 11360
rect 12638 11320 12680 11360
rect 12720 11320 16352 11360
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16720 11320 20352 11360
rect 20392 11320 20434 11360
rect 20474 11320 20516 11360
rect 20556 11320 20598 11360
rect 20638 11320 20680 11360
rect 20720 11320 24352 11360
rect 24392 11320 24434 11360
rect 24474 11320 24516 11360
rect 24556 11320 24598 11360
rect 24638 11320 24680 11360
rect 24720 11320 28352 11360
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28720 11320 32352 11360
rect 32392 11320 32434 11360
rect 32474 11320 32516 11360
rect 32556 11320 32598 11360
rect 32638 11320 32680 11360
rect 32720 11320 36352 11360
rect 36392 11320 36434 11360
rect 36474 11320 36516 11360
rect 36556 11320 36598 11360
rect 36638 11320 36680 11360
rect 36720 11320 40352 11360
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40720 11320 44352 11360
rect 44392 11320 44434 11360
rect 44474 11320 44516 11360
rect 44556 11320 44598 11360
rect 44638 11320 44680 11360
rect 44720 11320 48352 11360
rect 48392 11320 48434 11360
rect 48474 11320 48516 11360
rect 48556 11320 48598 11360
rect 48638 11320 48680 11360
rect 48720 11320 52352 11360
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52720 11320 56352 11360
rect 56392 11320 56434 11360
rect 56474 11320 56516 11360
rect 56556 11320 56598 11360
rect 56638 11320 56680 11360
rect 56720 11320 60352 11360
rect 60392 11320 60434 11360
rect 60474 11320 60516 11360
rect 60556 11320 60598 11360
rect 60638 11320 60680 11360
rect 60720 11320 64352 11360
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64720 11320 68352 11360
rect 68392 11320 68434 11360
rect 68474 11320 68516 11360
rect 68556 11320 68598 11360
rect 68638 11320 68680 11360
rect 68720 11320 71520 11360
rect 576 11296 71520 11320
rect 1227 11192 1269 11201
rect 1227 11152 1228 11192
rect 1268 11152 1269 11192
rect 1227 11143 1269 11152
rect 835 10940 893 10941
rect 835 10900 844 10940
rect 884 10900 893 10940
rect 835 10899 893 10900
rect 1411 10940 1469 10941
rect 1411 10900 1420 10940
rect 1460 10900 1469 10940
rect 1411 10899 1469 10900
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 576 10604 71520 10628
rect 576 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 7112 10604
rect 7152 10564 7194 10604
rect 7234 10564 7276 10604
rect 7316 10564 7358 10604
rect 7398 10564 7440 10604
rect 7480 10564 11112 10604
rect 11152 10564 11194 10604
rect 11234 10564 11276 10604
rect 11316 10564 11358 10604
rect 11398 10564 11440 10604
rect 11480 10564 15112 10604
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15480 10564 19112 10604
rect 19152 10564 19194 10604
rect 19234 10564 19276 10604
rect 19316 10564 19358 10604
rect 19398 10564 19440 10604
rect 19480 10564 23112 10604
rect 23152 10564 23194 10604
rect 23234 10564 23276 10604
rect 23316 10564 23358 10604
rect 23398 10564 23440 10604
rect 23480 10564 27112 10604
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27480 10564 31112 10604
rect 31152 10564 31194 10604
rect 31234 10564 31276 10604
rect 31316 10564 31358 10604
rect 31398 10564 31440 10604
rect 31480 10564 35112 10604
rect 35152 10564 35194 10604
rect 35234 10564 35276 10604
rect 35316 10564 35358 10604
rect 35398 10564 35440 10604
rect 35480 10564 39112 10604
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39480 10564 43112 10604
rect 43152 10564 43194 10604
rect 43234 10564 43276 10604
rect 43316 10564 43358 10604
rect 43398 10564 43440 10604
rect 43480 10564 47112 10604
rect 47152 10564 47194 10604
rect 47234 10564 47276 10604
rect 47316 10564 47358 10604
rect 47398 10564 47440 10604
rect 47480 10564 51112 10604
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51480 10564 55112 10604
rect 55152 10564 55194 10604
rect 55234 10564 55276 10604
rect 55316 10564 55358 10604
rect 55398 10564 55440 10604
rect 55480 10564 59112 10604
rect 59152 10564 59194 10604
rect 59234 10564 59276 10604
rect 59316 10564 59358 10604
rect 59398 10564 59440 10604
rect 59480 10564 63112 10604
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63480 10564 67112 10604
rect 67152 10564 67194 10604
rect 67234 10564 67276 10604
rect 67316 10564 67358 10604
rect 67398 10564 67440 10604
rect 67480 10564 71520 10604
rect 576 10540 71520 10564
rect 1419 10436 1461 10445
rect 1419 10396 1420 10436
rect 1460 10396 1461 10436
rect 1419 10387 1461 10396
rect 1035 10352 1077 10361
rect 1035 10312 1036 10352
rect 1076 10312 1077 10352
rect 1035 10303 1077 10312
rect 835 10268 893 10269
rect 835 10228 844 10268
rect 884 10228 893 10268
rect 835 10227 893 10228
rect 1219 10268 1277 10269
rect 1219 10228 1228 10268
rect 1268 10228 1277 10268
rect 1219 10227 1277 10228
rect 1603 10268 1661 10269
rect 1603 10228 1612 10268
rect 1652 10228 1661 10268
rect 1603 10227 1661 10228
rect 651 10016 693 10025
rect 651 9976 652 10016
rect 692 9976 693 10016
rect 651 9967 693 9976
rect 576 9848 71520 9872
rect 576 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 8352 9848
rect 8392 9808 8434 9848
rect 8474 9808 8516 9848
rect 8556 9808 8598 9848
rect 8638 9808 8680 9848
rect 8720 9808 12352 9848
rect 12392 9808 12434 9848
rect 12474 9808 12516 9848
rect 12556 9808 12598 9848
rect 12638 9808 12680 9848
rect 12720 9808 16352 9848
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16720 9808 20352 9848
rect 20392 9808 20434 9848
rect 20474 9808 20516 9848
rect 20556 9808 20598 9848
rect 20638 9808 20680 9848
rect 20720 9808 24352 9848
rect 24392 9808 24434 9848
rect 24474 9808 24516 9848
rect 24556 9808 24598 9848
rect 24638 9808 24680 9848
rect 24720 9808 28352 9848
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28720 9808 32352 9848
rect 32392 9808 32434 9848
rect 32474 9808 32516 9848
rect 32556 9808 32598 9848
rect 32638 9808 32680 9848
rect 32720 9808 36352 9848
rect 36392 9808 36434 9848
rect 36474 9808 36516 9848
rect 36556 9808 36598 9848
rect 36638 9808 36680 9848
rect 36720 9808 40352 9848
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40720 9808 44352 9848
rect 44392 9808 44434 9848
rect 44474 9808 44516 9848
rect 44556 9808 44598 9848
rect 44638 9808 44680 9848
rect 44720 9808 48352 9848
rect 48392 9808 48434 9848
rect 48474 9808 48516 9848
rect 48556 9808 48598 9848
rect 48638 9808 48680 9848
rect 48720 9808 52352 9848
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52720 9808 56352 9848
rect 56392 9808 56434 9848
rect 56474 9808 56516 9848
rect 56556 9808 56598 9848
rect 56638 9808 56680 9848
rect 56720 9808 60352 9848
rect 60392 9808 60434 9848
rect 60474 9808 60516 9848
rect 60556 9808 60598 9848
rect 60638 9808 60680 9848
rect 60720 9808 64352 9848
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64720 9808 68352 9848
rect 68392 9808 68434 9848
rect 68474 9808 68516 9848
rect 68556 9808 68598 9848
rect 68638 9808 68680 9848
rect 68720 9808 71520 9848
rect 576 9784 71520 9808
rect 835 9428 893 9429
rect 835 9388 844 9428
rect 884 9388 893 9428
rect 835 9387 893 9388
rect 651 9260 693 9269
rect 651 9220 652 9260
rect 692 9220 693 9260
rect 651 9211 693 9220
rect 576 9092 71520 9116
rect 576 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 7112 9092
rect 7152 9052 7194 9092
rect 7234 9052 7276 9092
rect 7316 9052 7358 9092
rect 7398 9052 7440 9092
rect 7480 9052 11112 9092
rect 11152 9052 11194 9092
rect 11234 9052 11276 9092
rect 11316 9052 11358 9092
rect 11398 9052 11440 9092
rect 11480 9052 15112 9092
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15480 9052 19112 9092
rect 19152 9052 19194 9092
rect 19234 9052 19276 9092
rect 19316 9052 19358 9092
rect 19398 9052 19440 9092
rect 19480 9052 23112 9092
rect 23152 9052 23194 9092
rect 23234 9052 23276 9092
rect 23316 9052 23358 9092
rect 23398 9052 23440 9092
rect 23480 9052 27112 9092
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27480 9052 31112 9092
rect 31152 9052 31194 9092
rect 31234 9052 31276 9092
rect 31316 9052 31358 9092
rect 31398 9052 31440 9092
rect 31480 9052 35112 9092
rect 35152 9052 35194 9092
rect 35234 9052 35276 9092
rect 35316 9052 35358 9092
rect 35398 9052 35440 9092
rect 35480 9052 39112 9092
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39480 9052 43112 9092
rect 43152 9052 43194 9092
rect 43234 9052 43276 9092
rect 43316 9052 43358 9092
rect 43398 9052 43440 9092
rect 43480 9052 47112 9092
rect 47152 9052 47194 9092
rect 47234 9052 47276 9092
rect 47316 9052 47358 9092
rect 47398 9052 47440 9092
rect 47480 9052 51112 9092
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51480 9052 55112 9092
rect 55152 9052 55194 9092
rect 55234 9052 55276 9092
rect 55316 9052 55358 9092
rect 55398 9052 55440 9092
rect 55480 9052 59112 9092
rect 59152 9052 59194 9092
rect 59234 9052 59276 9092
rect 59316 9052 59358 9092
rect 59398 9052 59440 9092
rect 59480 9052 63112 9092
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63480 9052 67112 9092
rect 67152 9052 67194 9092
rect 67234 9052 67276 9092
rect 67316 9052 67358 9092
rect 67398 9052 67440 9092
rect 67480 9052 71520 9092
rect 576 9028 71520 9052
rect 1131 8840 1173 8849
rect 1131 8800 1132 8840
rect 1172 8800 1173 8840
rect 1131 8791 1173 8800
rect 1515 8840 1557 8849
rect 1515 8800 1516 8840
rect 1556 8800 1557 8840
rect 1515 8791 1557 8800
rect 835 8756 893 8757
rect 835 8716 844 8756
rect 884 8716 893 8756
rect 835 8715 893 8716
rect 1315 8756 1373 8757
rect 1315 8716 1324 8756
rect 1364 8716 1373 8756
rect 1315 8715 1373 8716
rect 1699 8756 1757 8757
rect 1699 8716 1708 8756
rect 1748 8716 1757 8756
rect 1699 8715 1757 8716
rect 2083 8756 2141 8757
rect 2083 8716 2092 8756
rect 2132 8716 2141 8756
rect 2083 8715 2141 8716
rect 70915 8672 70973 8673
rect 70915 8632 70924 8672
rect 70964 8632 70973 8672
rect 70915 8631 70973 8632
rect 71107 8672 71165 8673
rect 71107 8632 71116 8672
rect 71156 8632 71165 8672
rect 71107 8631 71165 8632
rect 651 8504 693 8513
rect 651 8464 652 8504
rect 692 8464 693 8504
rect 651 8455 693 8464
rect 1899 8504 1941 8513
rect 1899 8464 1900 8504
rect 1940 8464 1941 8504
rect 1899 8455 1941 8464
rect 576 8336 71520 8360
rect 576 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 8352 8336
rect 8392 8296 8434 8336
rect 8474 8296 8516 8336
rect 8556 8296 8598 8336
rect 8638 8296 8680 8336
rect 8720 8296 12352 8336
rect 12392 8296 12434 8336
rect 12474 8296 12516 8336
rect 12556 8296 12598 8336
rect 12638 8296 12680 8336
rect 12720 8296 16352 8336
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16720 8296 20352 8336
rect 20392 8296 20434 8336
rect 20474 8296 20516 8336
rect 20556 8296 20598 8336
rect 20638 8296 20680 8336
rect 20720 8296 24352 8336
rect 24392 8296 24434 8336
rect 24474 8296 24516 8336
rect 24556 8296 24598 8336
rect 24638 8296 24680 8336
rect 24720 8296 28352 8336
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28720 8296 32352 8336
rect 32392 8296 32434 8336
rect 32474 8296 32516 8336
rect 32556 8296 32598 8336
rect 32638 8296 32680 8336
rect 32720 8296 36352 8336
rect 36392 8296 36434 8336
rect 36474 8296 36516 8336
rect 36556 8296 36598 8336
rect 36638 8296 36680 8336
rect 36720 8296 40352 8336
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40720 8296 44352 8336
rect 44392 8296 44434 8336
rect 44474 8296 44516 8336
rect 44556 8296 44598 8336
rect 44638 8296 44680 8336
rect 44720 8296 48352 8336
rect 48392 8296 48434 8336
rect 48474 8296 48516 8336
rect 48556 8296 48598 8336
rect 48638 8296 48680 8336
rect 48720 8296 52352 8336
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52720 8296 56352 8336
rect 56392 8296 56434 8336
rect 56474 8296 56516 8336
rect 56556 8296 56598 8336
rect 56638 8296 56680 8336
rect 56720 8296 60352 8336
rect 60392 8296 60434 8336
rect 60474 8296 60516 8336
rect 60556 8296 60598 8336
rect 60638 8296 60680 8336
rect 60720 8296 64352 8336
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64720 8296 68352 8336
rect 68392 8296 68434 8336
rect 68474 8296 68516 8336
rect 68556 8296 68598 8336
rect 68638 8296 68680 8336
rect 68720 8296 71520 8336
rect 576 8272 71520 8296
rect 835 7916 893 7917
rect 835 7876 844 7916
rect 884 7876 893 7916
rect 835 7875 893 7876
rect 70819 7916 70877 7917
rect 70819 7876 70828 7916
rect 70868 7876 70877 7916
rect 70819 7875 70877 7876
rect 71203 7916 71261 7917
rect 71203 7876 71212 7916
rect 71252 7876 71261 7916
rect 71203 7875 71261 7876
rect 71019 7832 71061 7841
rect 71019 7792 71020 7832
rect 71060 7792 71061 7832
rect 71019 7783 71061 7792
rect 71403 7832 71445 7841
rect 71403 7792 71404 7832
rect 71444 7792 71445 7832
rect 71403 7783 71445 7792
rect 651 7748 693 7757
rect 651 7708 652 7748
rect 692 7708 693 7748
rect 651 7699 693 7708
rect 576 7580 99360 7604
rect 576 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 7112 7580
rect 7152 7540 7194 7580
rect 7234 7540 7276 7580
rect 7316 7540 7358 7580
rect 7398 7540 7440 7580
rect 7480 7540 11112 7580
rect 11152 7540 11194 7580
rect 11234 7540 11276 7580
rect 11316 7540 11358 7580
rect 11398 7540 11440 7580
rect 11480 7540 15112 7580
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15480 7540 19112 7580
rect 19152 7540 19194 7580
rect 19234 7540 19276 7580
rect 19316 7540 19358 7580
rect 19398 7540 19440 7580
rect 19480 7540 23112 7580
rect 23152 7540 23194 7580
rect 23234 7540 23276 7580
rect 23316 7540 23358 7580
rect 23398 7540 23440 7580
rect 23480 7540 27112 7580
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27480 7540 31112 7580
rect 31152 7540 31194 7580
rect 31234 7540 31276 7580
rect 31316 7540 31358 7580
rect 31398 7540 31440 7580
rect 31480 7540 35112 7580
rect 35152 7540 35194 7580
rect 35234 7540 35276 7580
rect 35316 7540 35358 7580
rect 35398 7540 35440 7580
rect 35480 7540 39112 7580
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39480 7540 43112 7580
rect 43152 7540 43194 7580
rect 43234 7540 43276 7580
rect 43316 7540 43358 7580
rect 43398 7540 43440 7580
rect 43480 7540 47112 7580
rect 47152 7540 47194 7580
rect 47234 7540 47276 7580
rect 47316 7540 47358 7580
rect 47398 7540 47440 7580
rect 47480 7540 51112 7580
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51480 7540 55112 7580
rect 55152 7540 55194 7580
rect 55234 7540 55276 7580
rect 55316 7540 55358 7580
rect 55398 7540 55440 7580
rect 55480 7540 59112 7580
rect 59152 7540 59194 7580
rect 59234 7540 59276 7580
rect 59316 7540 59358 7580
rect 59398 7540 59440 7580
rect 59480 7540 63112 7580
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63480 7540 67112 7580
rect 67152 7540 67194 7580
rect 67234 7540 67276 7580
rect 67316 7540 67358 7580
rect 67398 7540 67440 7580
rect 67480 7540 99360 7580
rect 576 7516 99360 7540
rect 1515 7412 1557 7421
rect 1515 7372 1516 7412
rect 1556 7372 1557 7412
rect 1515 7363 1557 7372
rect 71403 7412 71445 7421
rect 71403 7372 71404 7412
rect 71444 7372 71445 7412
rect 71403 7363 71445 7372
rect 72171 7412 72213 7421
rect 72171 7372 72172 7412
rect 72212 7372 72213 7412
rect 72171 7363 72213 7372
rect 72555 7412 72597 7421
rect 72555 7372 72556 7412
rect 72596 7372 72597 7412
rect 72555 7363 72597 7372
rect 73323 7412 73365 7421
rect 73323 7372 73324 7412
rect 73364 7372 73365 7412
rect 73323 7363 73365 7372
rect 73707 7412 73749 7421
rect 73707 7372 73708 7412
rect 73748 7372 73749 7412
rect 73707 7363 73749 7372
rect 75147 7412 75189 7421
rect 75147 7372 75148 7412
rect 75188 7372 75189 7412
rect 75147 7363 75189 7372
rect 75915 7412 75957 7421
rect 75915 7372 75916 7412
rect 75956 7372 75957 7412
rect 75915 7363 75957 7372
rect 76203 7412 76245 7421
rect 76203 7372 76204 7412
rect 76244 7372 76245 7412
rect 76203 7363 76245 7372
rect 76779 7412 76821 7421
rect 76779 7372 76780 7412
rect 76820 7372 76821 7412
rect 76779 7363 76821 7372
rect 77835 7412 77877 7421
rect 77835 7372 77836 7412
rect 77876 7372 77877 7412
rect 77835 7363 77877 7372
rect 78123 7412 78165 7421
rect 78123 7372 78124 7412
rect 78164 7372 78165 7412
rect 78123 7363 78165 7372
rect 78411 7412 78453 7421
rect 78411 7372 78412 7412
rect 78452 7372 78453 7412
rect 78411 7363 78453 7372
rect 79275 7412 79317 7421
rect 79275 7372 79276 7412
rect 79316 7372 79317 7412
rect 79275 7363 79317 7372
rect 79467 7412 79509 7421
rect 79467 7372 79468 7412
rect 79508 7372 79509 7412
rect 79467 7363 79509 7372
rect 81099 7412 81141 7421
rect 81099 7372 81100 7412
rect 81140 7372 81141 7412
rect 81099 7363 81141 7372
rect 82347 7412 82389 7421
rect 82347 7372 82348 7412
rect 82388 7372 82389 7412
rect 82347 7363 82389 7372
rect 82539 7412 82581 7421
rect 82539 7372 82540 7412
rect 82580 7372 82581 7412
rect 82539 7363 82581 7372
rect 82827 7412 82869 7421
rect 82827 7372 82828 7412
rect 82868 7372 82869 7412
rect 82827 7363 82869 7372
rect 83979 7412 84021 7421
rect 83979 7372 83980 7412
rect 84020 7372 84021 7412
rect 83979 7363 84021 7372
rect 84171 7412 84213 7421
rect 84171 7372 84172 7412
rect 84212 7372 84213 7412
rect 84171 7363 84213 7372
rect 84459 7412 84501 7421
rect 84459 7372 84460 7412
rect 84500 7372 84501 7412
rect 84459 7363 84501 7372
rect 85323 7412 85365 7421
rect 85323 7372 85324 7412
rect 85364 7372 85365 7412
rect 85323 7363 85365 7372
rect 85515 7412 85557 7421
rect 85515 7372 85516 7412
rect 85556 7372 85557 7412
rect 85515 7363 85557 7372
rect 85803 7412 85845 7421
rect 85803 7372 85804 7412
rect 85844 7372 85845 7412
rect 85803 7363 85845 7372
rect 87435 7412 87477 7421
rect 87435 7372 87436 7412
rect 87476 7372 87477 7412
rect 87435 7363 87477 7372
rect 87723 7412 87765 7421
rect 87723 7372 87724 7412
rect 87764 7372 87765 7412
rect 87723 7363 87765 7372
rect 88779 7412 88821 7421
rect 88779 7372 88780 7412
rect 88820 7372 88821 7412
rect 88779 7363 88821 7372
rect 88971 7412 89013 7421
rect 88971 7372 88972 7412
rect 89012 7372 89013 7412
rect 88971 7363 89013 7372
rect 89643 7412 89685 7421
rect 89643 7372 89644 7412
rect 89684 7372 89685 7412
rect 89643 7363 89685 7372
rect 90219 7412 90261 7421
rect 90219 7372 90220 7412
rect 90260 7372 90261 7412
rect 90219 7363 90261 7372
rect 90507 7412 90549 7421
rect 90507 7372 90508 7412
rect 90548 7372 90549 7412
rect 90507 7363 90549 7372
rect 91179 7412 91221 7421
rect 91179 7372 91180 7412
rect 91220 7372 91221 7412
rect 91179 7363 91221 7372
rect 91755 7412 91797 7421
rect 91755 7372 91756 7412
rect 91796 7372 91797 7412
rect 91755 7363 91797 7372
rect 93483 7412 93525 7421
rect 93483 7372 93484 7412
rect 93524 7372 93525 7412
rect 93483 7363 93525 7372
rect 93771 7412 93813 7421
rect 93771 7372 93772 7412
rect 93812 7372 93813 7412
rect 93771 7363 93813 7372
rect 96459 7412 96501 7421
rect 96459 7372 96460 7412
rect 96500 7372 96501 7412
rect 96459 7363 96501 7372
rect 97803 7412 97845 7421
rect 97803 7372 97804 7412
rect 97844 7372 97845 7412
rect 97803 7363 97845 7372
rect 98475 7412 98517 7421
rect 98475 7372 98476 7412
rect 98516 7372 98517 7412
rect 98475 7363 98517 7372
rect 99243 7412 99285 7421
rect 99243 7372 99244 7412
rect 99284 7372 99285 7412
rect 99243 7363 99285 7372
rect 73131 7328 73173 7337
rect 73131 7288 73132 7328
rect 73172 7288 73173 7328
rect 73131 7279 73173 7288
rect 77643 7328 77685 7337
rect 77643 7288 77644 7328
rect 77684 7288 77685 7328
rect 77643 7279 77685 7288
rect 80139 7328 80181 7337
rect 80139 7288 80140 7328
rect 80180 7288 80181 7328
rect 80139 7279 80181 7288
rect 80523 7328 80565 7337
rect 80523 7288 80524 7328
rect 80564 7288 80565 7328
rect 80523 7279 80565 7288
rect 83595 7328 83637 7337
rect 83595 7288 83596 7328
rect 83636 7288 83637 7328
rect 83595 7279 83637 7288
rect 86859 7328 86901 7337
rect 86859 7288 86860 7328
rect 86900 7288 86901 7328
rect 86859 7279 86901 7288
rect 88395 7328 88437 7337
rect 88395 7288 88396 7328
rect 88436 7288 88437 7328
rect 88395 7279 88437 7288
rect 90027 7328 90069 7337
rect 90027 7288 90028 7328
rect 90068 7288 90069 7328
rect 90027 7279 90069 7288
rect 91563 7328 91605 7337
rect 91563 7288 91564 7328
rect 91604 7288 91605 7328
rect 91563 7279 91605 7288
rect 95979 7328 96021 7337
rect 95979 7288 95980 7328
rect 96020 7288 96021 7328
rect 95979 7279 96021 7288
rect 98091 7328 98133 7337
rect 98091 7288 98092 7328
rect 98132 7288 98133 7328
rect 98091 7279 98133 7288
rect 835 7244 893 7245
rect 835 7204 844 7244
rect 884 7204 893 7244
rect 835 7203 893 7204
rect 1699 7244 1757 7245
rect 1699 7204 1708 7244
rect 1748 7204 1757 7244
rect 1699 7203 1757 7204
rect 72355 7244 72413 7245
rect 72355 7204 72364 7244
rect 72404 7204 72413 7244
rect 72355 7203 72413 7204
rect 72931 7244 72989 7245
rect 72931 7204 72940 7244
rect 72980 7204 72989 7244
rect 72931 7203 72989 7204
rect 74275 7244 74333 7245
rect 74275 7204 74284 7244
rect 74324 7204 74333 7244
rect 74275 7203 74333 7204
rect 74659 7244 74717 7245
rect 74659 7204 74668 7244
rect 74708 7204 74717 7244
rect 74659 7203 74717 7204
rect 74859 7244 74901 7253
rect 74859 7204 74860 7244
rect 74900 7204 74901 7244
rect 74859 7195 74901 7204
rect 75523 7244 75581 7245
rect 75523 7204 75532 7244
rect 75572 7204 75581 7244
rect 75523 7203 75581 7204
rect 76491 7244 76533 7253
rect 76491 7204 76492 7244
rect 76532 7204 76533 7244
rect 76491 7195 76533 7204
rect 77347 7244 77405 7245
rect 77347 7204 77356 7244
rect 77396 7204 77405 7244
rect 77347 7203 77405 7204
rect 78787 7244 78845 7245
rect 78787 7204 78796 7244
rect 78836 7204 78845 7244
rect 78787 7203 78845 7204
rect 79747 7244 79805 7245
rect 79747 7204 79756 7244
rect 79796 7204 79805 7244
rect 79747 7203 79805 7204
rect 80323 7244 80381 7245
rect 80323 7204 80332 7244
rect 80372 7204 80381 7244
rect 80323 7203 80381 7204
rect 81571 7244 81629 7245
rect 81571 7204 81580 7244
rect 81620 7204 81629 7244
rect 81571 7203 81629 7204
rect 83203 7244 83261 7245
rect 83203 7204 83212 7244
rect 83252 7204 83261 7244
rect 83203 7203 83261 7204
rect 84835 7244 84893 7245
rect 84835 7204 84844 7244
rect 84884 7204 84893 7244
rect 84835 7203 84893 7204
rect 86275 7244 86333 7245
rect 86275 7204 86284 7244
rect 86324 7204 86333 7244
rect 86275 7203 86333 7204
rect 86659 7244 86717 7245
rect 86659 7204 86668 7244
rect 86708 7204 86717 7244
rect 86659 7203 86717 7204
rect 88195 7244 88253 7245
rect 88195 7204 88204 7244
rect 88244 7204 88253 7244
rect 88195 7203 88253 7204
rect 89251 7244 89309 7245
rect 89251 7204 89260 7244
rect 89300 7204 89309 7244
rect 89251 7203 89309 7204
rect 90787 7244 90845 7245
rect 90787 7204 90796 7244
rect 90836 7204 90845 7244
rect 90787 7203 90845 7204
rect 92323 7244 92381 7245
rect 92323 7204 92332 7244
rect 92372 7204 92381 7244
rect 92323 7203 92381 7204
rect 92707 7244 92765 7245
rect 92707 7204 92716 7244
rect 92756 7204 92765 7244
rect 92707 7203 92765 7204
rect 92907 7244 92949 7253
rect 92907 7204 92908 7244
rect 92948 7204 92949 7244
rect 92907 7195 92949 7204
rect 94243 7244 94301 7245
rect 94243 7204 94252 7244
rect 94292 7204 94301 7244
rect 94243 7203 94301 7204
rect 95203 7244 95261 7245
rect 95203 7204 95212 7244
rect 95252 7204 95261 7244
rect 95203 7203 95261 7204
rect 95595 7244 95637 7253
rect 95595 7204 95596 7244
rect 95636 7204 95637 7244
rect 95595 7195 95637 7204
rect 96171 7244 96213 7253
rect 96171 7204 96172 7244
rect 96212 7204 96213 7244
rect 96171 7195 96213 7204
rect 96835 7244 96893 7245
rect 96835 7204 96844 7244
rect 96884 7204 96893 7244
rect 96835 7203 96893 7204
rect 98659 7244 98717 7245
rect 98659 7204 98668 7244
rect 98708 7204 98717 7244
rect 98659 7203 98717 7204
rect 97315 7173 97373 7174
rect 71299 7160 71357 7161
rect 71299 7120 71308 7160
rect 71348 7120 71357 7160
rect 71299 7119 71357 7120
rect 72067 7160 72125 7161
rect 72067 7120 72076 7160
rect 72116 7120 72125 7160
rect 73603 7160 73661 7161
rect 72067 7119 72125 7120
rect 73432 7149 73474 7158
rect 73432 7109 73433 7149
rect 73473 7109 73474 7149
rect 73603 7120 73612 7160
rect 73652 7120 73661 7160
rect 73603 7119 73661 7120
rect 74947 7160 75005 7161
rect 74947 7120 74956 7160
rect 74996 7120 75005 7160
rect 74947 7119 75005 7120
rect 75235 7160 75293 7161
rect 75235 7120 75244 7160
rect 75284 7120 75293 7160
rect 75235 7119 75293 7120
rect 76003 7160 76061 7161
rect 76003 7120 76012 7160
rect 76052 7120 76061 7160
rect 76003 7119 76061 7120
rect 76291 7160 76349 7161
rect 76291 7120 76300 7160
rect 76340 7120 76349 7160
rect 76291 7119 76349 7120
rect 76579 7160 76637 7161
rect 76579 7120 76588 7160
rect 76628 7120 76637 7160
rect 76579 7119 76637 7120
rect 76867 7160 76925 7161
rect 76867 7120 76876 7160
rect 76916 7120 76925 7160
rect 76867 7119 76925 7120
rect 77539 7160 77597 7161
rect 77539 7120 77548 7160
rect 77588 7120 77597 7160
rect 77539 7119 77597 7120
rect 77923 7160 77981 7161
rect 77923 7120 77932 7160
rect 77972 7120 77981 7160
rect 77923 7119 77981 7120
rect 78211 7160 78269 7161
rect 78211 7120 78220 7160
rect 78260 7120 78269 7160
rect 78211 7119 78269 7120
rect 78499 7160 78557 7161
rect 78499 7120 78508 7160
rect 78548 7120 78557 7160
rect 78499 7119 78557 7120
rect 79171 7160 79229 7161
rect 79171 7120 79180 7160
rect 79220 7120 79229 7160
rect 79171 7119 79229 7120
rect 79555 7160 79613 7161
rect 79555 7120 79564 7160
rect 79604 7120 79613 7160
rect 79555 7119 79613 7120
rect 80611 7160 80669 7161
rect 80611 7120 80620 7160
rect 80660 7120 80669 7160
rect 80611 7119 80669 7120
rect 80803 7160 80861 7161
rect 80803 7120 80812 7160
rect 80852 7120 80861 7160
rect 80803 7119 80861 7120
rect 81187 7160 81245 7161
rect 81187 7120 81196 7160
rect 81236 7120 81245 7160
rect 81187 7119 81245 7120
rect 82051 7160 82109 7161
rect 82051 7120 82060 7160
rect 82100 7120 82109 7160
rect 82051 7119 82109 7120
rect 82243 7160 82301 7161
rect 82243 7120 82252 7160
rect 82292 7120 82301 7160
rect 82243 7119 82301 7120
rect 82627 7160 82685 7161
rect 82627 7120 82636 7160
rect 82676 7120 82685 7160
rect 82627 7119 82685 7120
rect 82915 7160 82973 7161
rect 82915 7120 82924 7160
rect 82964 7120 82973 7160
rect 82915 7119 82973 7120
rect 83683 7160 83741 7161
rect 83683 7120 83692 7160
rect 83732 7120 83741 7160
rect 83683 7119 83741 7120
rect 83875 7160 83933 7161
rect 83875 7120 83884 7160
rect 83924 7120 83933 7160
rect 83875 7119 83933 7120
rect 84259 7160 84317 7161
rect 84259 7120 84268 7160
rect 84308 7120 84317 7160
rect 84259 7119 84317 7120
rect 84547 7160 84605 7161
rect 84547 7120 84556 7160
rect 84596 7120 84605 7160
rect 84547 7119 84605 7120
rect 85219 7160 85277 7161
rect 85219 7120 85228 7160
rect 85268 7120 85277 7160
rect 85219 7119 85277 7120
rect 85603 7160 85661 7161
rect 85603 7120 85612 7160
rect 85652 7120 85661 7160
rect 85603 7119 85661 7120
rect 85891 7160 85949 7161
rect 85891 7120 85900 7160
rect 85940 7120 85949 7160
rect 85891 7119 85949 7120
rect 86947 7160 87005 7161
rect 86947 7120 86956 7160
rect 86996 7120 87005 7160
rect 86947 7119 87005 7120
rect 87139 7160 87197 7161
rect 87139 7120 87148 7160
rect 87188 7120 87197 7160
rect 87139 7119 87197 7120
rect 87523 7160 87581 7161
rect 87523 7120 87532 7160
rect 87572 7120 87581 7160
rect 87523 7119 87581 7120
rect 87811 7160 87869 7161
rect 87811 7120 87820 7160
rect 87860 7120 87869 7160
rect 87811 7119 87869 7120
rect 88483 7160 88541 7161
rect 88483 7120 88492 7160
rect 88532 7120 88541 7160
rect 88483 7119 88541 7120
rect 88675 7160 88733 7161
rect 88675 7120 88684 7160
rect 88724 7120 88733 7160
rect 88675 7119 88733 7120
rect 89059 7160 89117 7161
rect 89059 7120 89068 7160
rect 89108 7120 89117 7160
rect 89059 7119 89117 7120
rect 89731 7160 89789 7161
rect 89731 7120 89740 7160
rect 89780 7120 89789 7160
rect 89731 7119 89789 7120
rect 89923 7160 89981 7161
rect 89923 7120 89932 7160
rect 89972 7120 89981 7160
rect 89923 7119 89981 7120
rect 90307 7160 90365 7161
rect 90307 7120 90316 7160
rect 90356 7120 90365 7160
rect 90307 7119 90365 7120
rect 90595 7160 90653 7161
rect 90595 7120 90604 7160
rect 90644 7120 90653 7160
rect 90595 7119 90653 7120
rect 91267 7160 91325 7161
rect 91267 7120 91276 7160
rect 91316 7120 91325 7160
rect 91267 7119 91325 7120
rect 91459 7160 91517 7161
rect 91459 7120 91468 7160
rect 91508 7120 91517 7160
rect 91459 7119 91517 7120
rect 91843 7160 91901 7161
rect 91843 7120 91852 7160
rect 91892 7120 91901 7160
rect 91843 7119 91901 7120
rect 92995 7160 93053 7161
rect 92995 7120 93004 7160
rect 93044 7120 93053 7160
rect 92995 7119 93053 7120
rect 93187 7160 93245 7161
rect 93187 7120 93196 7160
rect 93236 7120 93245 7160
rect 93187 7119 93245 7120
rect 93571 7160 93629 7161
rect 93571 7120 93580 7160
rect 93620 7120 93629 7160
rect 93571 7119 93629 7120
rect 93859 7160 93917 7161
rect 93859 7120 93868 7160
rect 93908 7120 93917 7160
rect 93859 7119 93917 7120
rect 94531 7160 94589 7161
rect 94531 7120 94540 7160
rect 94580 7120 94589 7160
rect 94531 7119 94589 7120
rect 94723 7160 94781 7161
rect 94723 7120 94732 7160
rect 94772 7120 94781 7160
rect 94723 7119 94781 7120
rect 94827 7160 94869 7169
rect 94827 7120 94828 7160
rect 94868 7120 94869 7160
rect 94827 7111 94869 7120
rect 95683 7160 95741 7161
rect 95683 7120 95692 7160
rect 95732 7120 95741 7160
rect 95683 7119 95741 7120
rect 95875 7160 95933 7161
rect 95875 7120 95884 7160
rect 95924 7120 95933 7160
rect 95875 7119 95933 7120
rect 96259 7160 96317 7161
rect 96259 7120 96268 7160
rect 96308 7120 96317 7160
rect 96259 7119 96317 7120
rect 96547 7160 96605 7161
rect 96547 7120 96556 7160
rect 96596 7120 96605 7160
rect 96547 7119 96605 7120
rect 97227 7160 97269 7169
rect 97227 7120 97228 7160
rect 97268 7120 97269 7160
rect 97315 7133 97324 7173
rect 97364 7133 97373 7173
rect 97315 7132 97373 7133
rect 97507 7160 97565 7161
rect 97227 7111 97269 7120
rect 97507 7120 97516 7160
rect 97556 7120 97565 7160
rect 97507 7119 97565 7120
rect 97891 7160 97949 7161
rect 97891 7120 97900 7160
rect 97940 7120 97949 7160
rect 97891 7119 97949 7120
rect 98179 7160 98237 7161
rect 98179 7120 98188 7160
rect 98228 7120 98237 7160
rect 98179 7119 98237 7120
rect 98947 7160 99005 7161
rect 98947 7120 98956 7160
rect 98996 7120 99005 7160
rect 98947 7119 99005 7120
rect 99139 7160 99197 7161
rect 99139 7120 99148 7160
rect 99188 7120 99197 7160
rect 99139 7119 99197 7120
rect 73432 7100 73474 7109
rect 87243 7076 87285 7085
rect 87243 7036 87244 7076
rect 87284 7036 87285 7076
rect 87243 7027 87285 7036
rect 94443 7076 94485 7085
rect 94443 7036 94444 7076
rect 94484 7036 94485 7076
rect 94443 7027 94485 7036
rect 98859 7076 98901 7085
rect 98859 7036 98860 7076
rect 98900 7036 98901 7076
rect 98859 7027 98901 7036
rect 651 6992 693 7001
rect 651 6952 652 6992
rect 692 6952 693 6992
rect 651 6943 693 6952
rect 74091 6992 74133 7001
rect 74091 6952 74092 6992
rect 74132 6952 74133 6992
rect 74091 6943 74133 6952
rect 74475 6992 74517 7001
rect 74475 6952 74476 6992
rect 74516 6952 74517 6992
rect 74475 6943 74517 6952
rect 75723 6992 75765 7001
rect 75723 6952 75724 6992
rect 75764 6952 75765 6992
rect 75723 6943 75765 6952
rect 77163 6992 77205 7001
rect 77163 6952 77164 6992
rect 77204 6952 77205 6992
rect 77163 6943 77205 6952
rect 78987 6992 79029 7001
rect 78987 6952 78988 6992
rect 79028 6952 79029 6992
rect 78987 6943 79029 6952
rect 79947 6992 79989 7001
rect 79947 6952 79948 6992
rect 79988 6952 79989 6992
rect 79947 6943 79989 6952
rect 80907 6992 80949 7001
rect 80907 6952 80908 6992
rect 80948 6952 80949 6992
rect 80907 6943 80949 6952
rect 81771 6992 81813 7001
rect 81771 6952 81772 6992
rect 81812 6952 81813 6992
rect 81771 6943 81813 6952
rect 81963 6992 82005 7001
rect 81963 6952 81964 6992
rect 82004 6952 82005 6992
rect 81963 6943 82005 6952
rect 83403 6992 83445 7001
rect 83403 6952 83404 6992
rect 83444 6952 83445 6992
rect 83403 6943 83445 6952
rect 85035 6992 85077 7001
rect 85035 6952 85036 6992
rect 85076 6952 85077 6992
rect 85035 6943 85077 6952
rect 86091 6992 86133 7001
rect 86091 6952 86092 6992
rect 86132 6952 86133 6992
rect 86091 6943 86133 6952
rect 86475 6992 86517 7001
rect 86475 6952 86476 6992
rect 86516 6952 86517 6992
rect 86475 6943 86517 6952
rect 88011 6992 88053 7001
rect 88011 6952 88012 6992
rect 88052 6952 88053 6992
rect 88011 6943 88053 6952
rect 89451 6992 89493 7001
rect 89451 6952 89452 6992
rect 89492 6952 89493 6992
rect 89451 6943 89493 6952
rect 90987 6992 91029 7001
rect 90987 6952 90988 6992
rect 91028 6952 91029 6992
rect 90987 6943 91029 6952
rect 92139 6992 92181 7001
rect 92139 6952 92140 6992
rect 92180 6952 92181 6992
rect 92139 6943 92181 6952
rect 92523 6992 92565 7001
rect 92523 6952 92524 6992
rect 92564 6952 92565 6992
rect 92523 6943 92565 6952
rect 93291 6992 93333 7001
rect 93291 6952 93292 6992
rect 93332 6952 93333 6992
rect 93291 6943 93333 6952
rect 94059 6992 94101 7001
rect 94059 6952 94060 6992
rect 94100 6952 94101 6992
rect 94059 6943 94101 6952
rect 95403 6992 95445 7001
rect 95403 6952 95404 6992
rect 95444 6952 95445 6992
rect 95403 6943 95445 6952
rect 97035 6992 97077 7001
rect 97035 6952 97036 6992
rect 97076 6952 97077 6992
rect 97035 6943 97077 6952
rect 97611 6992 97653 7001
rect 97611 6952 97612 6992
rect 97652 6952 97653 6992
rect 97611 6943 97653 6952
rect 576 6824 99360 6848
rect 576 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 8352 6824
rect 8392 6784 8434 6824
rect 8474 6784 8516 6824
rect 8556 6784 8598 6824
rect 8638 6784 8680 6824
rect 8720 6784 12352 6824
rect 12392 6784 12434 6824
rect 12474 6784 12516 6824
rect 12556 6784 12598 6824
rect 12638 6784 12680 6824
rect 12720 6784 16352 6824
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16720 6784 20352 6824
rect 20392 6784 20434 6824
rect 20474 6784 20516 6824
rect 20556 6784 20598 6824
rect 20638 6784 20680 6824
rect 20720 6784 24352 6824
rect 24392 6784 24434 6824
rect 24474 6784 24516 6824
rect 24556 6784 24598 6824
rect 24638 6784 24680 6824
rect 24720 6784 28352 6824
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28720 6784 32352 6824
rect 32392 6784 32434 6824
rect 32474 6784 32516 6824
rect 32556 6784 32598 6824
rect 32638 6784 32680 6824
rect 32720 6784 36352 6824
rect 36392 6784 36434 6824
rect 36474 6784 36516 6824
rect 36556 6784 36598 6824
rect 36638 6784 36680 6824
rect 36720 6784 40352 6824
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40720 6784 44352 6824
rect 44392 6784 44434 6824
rect 44474 6784 44516 6824
rect 44556 6784 44598 6824
rect 44638 6784 44680 6824
rect 44720 6784 48352 6824
rect 48392 6784 48434 6824
rect 48474 6784 48516 6824
rect 48556 6784 48598 6824
rect 48638 6784 48680 6824
rect 48720 6784 52352 6824
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52720 6784 56352 6824
rect 56392 6784 56434 6824
rect 56474 6784 56516 6824
rect 56556 6784 56598 6824
rect 56638 6784 56680 6824
rect 56720 6784 60352 6824
rect 60392 6784 60434 6824
rect 60474 6784 60516 6824
rect 60556 6784 60598 6824
rect 60638 6784 60680 6824
rect 60720 6784 64352 6824
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64720 6784 68352 6824
rect 68392 6784 68434 6824
rect 68474 6784 68516 6824
rect 68556 6784 68598 6824
rect 68638 6784 68680 6824
rect 68720 6784 99360 6824
rect 576 6760 99360 6784
rect 1707 6656 1749 6665
rect 1707 6616 1708 6656
rect 1748 6616 1749 6656
rect 1707 6607 1749 6616
rect 73707 6656 73749 6665
rect 73707 6616 73708 6656
rect 73748 6616 73749 6656
rect 73707 6607 73749 6616
rect 74187 6656 74229 6665
rect 74187 6616 74188 6656
rect 74228 6616 74229 6656
rect 74187 6607 74229 6616
rect 74571 6656 74613 6665
rect 74571 6616 74572 6656
rect 74612 6616 74613 6656
rect 74571 6607 74613 6616
rect 75051 6656 75093 6665
rect 75051 6616 75052 6656
rect 75092 6616 75093 6656
rect 75051 6607 75093 6616
rect 75435 6656 75477 6665
rect 75435 6616 75436 6656
rect 75476 6616 75477 6656
rect 75435 6607 75477 6616
rect 75819 6656 75861 6665
rect 75819 6616 75820 6656
rect 75860 6616 75861 6656
rect 75819 6607 75861 6616
rect 76203 6656 76245 6665
rect 76203 6616 76204 6656
rect 76244 6616 76245 6656
rect 76203 6607 76245 6616
rect 76683 6656 76725 6665
rect 76683 6616 76684 6656
rect 76724 6616 76725 6656
rect 76683 6607 76725 6616
rect 77067 6656 77109 6665
rect 77067 6616 77068 6656
rect 77108 6616 77109 6656
rect 77067 6607 77109 6616
rect 77451 6656 77493 6665
rect 77451 6616 77452 6656
rect 77492 6616 77493 6656
rect 77451 6607 77493 6616
rect 77835 6656 77877 6665
rect 77835 6616 77836 6656
rect 77876 6616 77877 6656
rect 77835 6607 77877 6616
rect 78315 6656 78357 6665
rect 78315 6616 78316 6656
rect 78356 6616 78357 6656
rect 78315 6607 78357 6616
rect 78699 6656 78741 6665
rect 78699 6616 78700 6656
rect 78740 6616 78741 6656
rect 78699 6607 78741 6616
rect 79083 6656 79125 6665
rect 79083 6616 79084 6656
rect 79124 6616 79125 6656
rect 79083 6607 79125 6616
rect 79467 6656 79509 6665
rect 79467 6616 79468 6656
rect 79508 6616 79509 6656
rect 79467 6607 79509 6616
rect 79947 6656 79989 6665
rect 79947 6616 79948 6656
rect 79988 6616 79989 6656
rect 79947 6607 79989 6616
rect 80331 6656 80373 6665
rect 80331 6616 80332 6656
rect 80372 6616 80373 6656
rect 80331 6607 80373 6616
rect 80715 6656 80757 6665
rect 80715 6616 80716 6656
rect 80756 6616 80757 6656
rect 80715 6607 80757 6616
rect 80907 6656 80949 6665
rect 80907 6616 80908 6656
rect 80948 6616 80949 6656
rect 80907 6607 80949 6616
rect 81483 6656 81525 6665
rect 81483 6616 81484 6656
rect 81524 6616 81525 6656
rect 81483 6607 81525 6616
rect 81867 6656 81909 6665
rect 81867 6616 81868 6656
rect 81908 6616 81909 6656
rect 81867 6607 81909 6616
rect 82251 6656 82293 6665
rect 82251 6616 82252 6656
rect 82292 6616 82293 6656
rect 82251 6607 82293 6616
rect 82731 6656 82773 6665
rect 82731 6616 82732 6656
rect 82772 6616 82773 6656
rect 82731 6607 82773 6616
rect 83115 6656 83157 6665
rect 83115 6616 83116 6656
rect 83156 6616 83157 6656
rect 83115 6607 83157 6616
rect 83307 6656 83349 6665
rect 83307 6616 83308 6656
rect 83348 6616 83349 6656
rect 83307 6607 83349 6616
rect 83883 6656 83925 6665
rect 83883 6616 83884 6656
rect 83924 6616 83925 6656
rect 83883 6607 83925 6616
rect 84267 6656 84309 6665
rect 84267 6616 84268 6656
rect 84308 6616 84309 6656
rect 84267 6607 84309 6616
rect 84651 6656 84693 6665
rect 84651 6616 84652 6656
rect 84692 6616 84693 6656
rect 84651 6607 84693 6616
rect 85035 6656 85077 6665
rect 85035 6616 85036 6656
rect 85076 6616 85077 6656
rect 85035 6607 85077 6616
rect 85515 6656 85557 6665
rect 85515 6616 85516 6656
rect 85556 6616 85557 6656
rect 85515 6607 85557 6616
rect 85899 6656 85941 6665
rect 85899 6616 85900 6656
rect 85940 6616 85941 6656
rect 85899 6607 85941 6616
rect 86283 6656 86325 6665
rect 86283 6616 86284 6656
rect 86324 6616 86325 6656
rect 86283 6607 86325 6616
rect 86667 6656 86709 6665
rect 86667 6616 86668 6656
rect 86708 6616 86709 6656
rect 86667 6607 86709 6616
rect 87051 6656 87093 6665
rect 87051 6616 87052 6656
rect 87092 6616 87093 6656
rect 87051 6607 87093 6616
rect 87531 6656 87573 6665
rect 87531 6616 87532 6656
rect 87572 6616 87573 6656
rect 87531 6607 87573 6616
rect 87723 6656 87765 6665
rect 87723 6616 87724 6656
rect 87764 6616 87765 6656
rect 87723 6607 87765 6616
rect 88299 6656 88341 6665
rect 88299 6616 88300 6656
rect 88340 6616 88341 6656
rect 88299 6607 88341 6616
rect 88683 6656 88725 6665
rect 88683 6616 88684 6656
rect 88724 6616 88725 6656
rect 88683 6607 88725 6616
rect 89067 6656 89109 6665
rect 89067 6616 89068 6656
rect 89108 6616 89109 6656
rect 89067 6607 89109 6616
rect 89451 6656 89493 6665
rect 89451 6616 89452 6656
rect 89492 6616 89493 6656
rect 89451 6607 89493 6616
rect 89931 6656 89973 6665
rect 89931 6616 89932 6656
rect 89972 6616 89973 6656
rect 89931 6607 89973 6616
rect 90315 6656 90357 6665
rect 90315 6616 90316 6656
rect 90356 6616 90357 6656
rect 90315 6607 90357 6616
rect 90699 6656 90741 6665
rect 90699 6616 90700 6656
rect 90740 6616 90741 6656
rect 90699 6607 90741 6616
rect 91083 6656 91125 6665
rect 91083 6616 91084 6656
rect 91124 6616 91125 6656
rect 91083 6607 91125 6616
rect 91467 6656 91509 6665
rect 91467 6616 91468 6656
rect 91508 6616 91509 6656
rect 91467 6607 91509 6616
rect 92331 6656 92373 6665
rect 92331 6616 92332 6656
rect 92372 6616 92373 6656
rect 92331 6607 92373 6616
rect 92715 6656 92757 6665
rect 92715 6616 92716 6656
rect 92756 6616 92757 6656
rect 92715 6607 92757 6616
rect 93099 6656 93141 6665
rect 93099 6616 93100 6656
rect 93140 6616 93141 6656
rect 93099 6607 93141 6616
rect 93579 6656 93621 6665
rect 93579 6616 93580 6656
rect 93620 6616 93621 6656
rect 93579 6607 93621 6616
rect 93771 6656 93813 6665
rect 93771 6616 93772 6656
rect 93812 6616 93813 6656
rect 93771 6607 93813 6616
rect 94347 6656 94389 6665
rect 94347 6616 94348 6656
rect 94388 6616 94389 6656
rect 94347 6607 94389 6616
rect 94731 6656 94773 6665
rect 94731 6616 94732 6656
rect 94772 6616 94773 6656
rect 94731 6607 94773 6616
rect 95115 6656 95157 6665
rect 95115 6616 95116 6656
rect 95156 6616 95157 6656
rect 95115 6607 95157 6616
rect 95595 6656 95637 6665
rect 95595 6616 95596 6656
rect 95636 6616 95637 6656
rect 95595 6607 95637 6616
rect 95979 6656 96021 6665
rect 95979 6616 95980 6656
rect 96020 6616 96021 6656
rect 95979 6607 96021 6616
rect 96363 6656 96405 6665
rect 96363 6616 96364 6656
rect 96404 6616 96405 6656
rect 96363 6607 96405 6616
rect 96747 6656 96789 6665
rect 96747 6616 96748 6656
rect 96788 6616 96789 6656
rect 96747 6607 96789 6616
rect 97035 6656 97077 6665
rect 97035 6616 97036 6656
rect 97076 6616 97077 6656
rect 97035 6607 97077 6616
rect 97515 6656 97557 6665
rect 97515 6616 97516 6656
rect 97556 6616 97557 6656
rect 97515 6607 97557 6616
rect 97899 6656 97941 6665
rect 97899 6616 97900 6656
rect 97940 6616 97941 6656
rect 97899 6607 97941 6616
rect 98379 6656 98421 6665
rect 98379 6616 98380 6656
rect 98420 6616 98421 6656
rect 98379 6607 98421 6616
rect 73323 6572 73365 6581
rect 73323 6532 73324 6572
rect 73364 6532 73365 6572
rect 73323 6523 73365 6532
rect 73219 6488 73277 6489
rect 73219 6448 73228 6488
rect 73268 6448 73277 6488
rect 73219 6447 73277 6448
rect 80995 6488 81053 6489
rect 80995 6448 81004 6488
rect 81044 6448 81053 6488
rect 80995 6447 81053 6448
rect 83395 6488 83453 6489
rect 83395 6448 83404 6488
rect 83444 6448 83453 6488
rect 83395 6447 83453 6448
rect 98467 6488 98525 6489
rect 98467 6448 98476 6488
rect 98516 6448 98525 6488
rect 98467 6447 98525 6448
rect 1507 6404 1565 6405
rect 1507 6364 1516 6404
rect 1556 6364 1565 6404
rect 1507 6363 1565 6364
rect 1891 6404 1949 6405
rect 1891 6364 1900 6404
rect 1940 6364 1949 6404
rect 1891 6363 1949 6364
rect 73507 6404 73565 6405
rect 73507 6364 73516 6404
rect 73556 6364 73565 6404
rect 73507 6363 73565 6364
rect 73987 6404 74045 6405
rect 73987 6364 73996 6404
rect 74036 6364 74045 6404
rect 73987 6363 74045 6364
rect 74371 6404 74429 6405
rect 74371 6364 74380 6404
rect 74420 6364 74429 6404
rect 74371 6363 74429 6364
rect 74851 6404 74909 6405
rect 74851 6364 74860 6404
rect 74900 6364 74909 6404
rect 74851 6363 74909 6364
rect 75235 6404 75293 6405
rect 75235 6364 75244 6404
rect 75284 6364 75293 6404
rect 75235 6363 75293 6364
rect 75619 6404 75677 6405
rect 75619 6364 75628 6404
rect 75668 6364 75677 6404
rect 75619 6363 75677 6364
rect 76003 6404 76061 6405
rect 76003 6364 76012 6404
rect 76052 6364 76061 6404
rect 76003 6363 76061 6364
rect 76483 6404 76541 6405
rect 76483 6364 76492 6404
rect 76532 6364 76541 6404
rect 76483 6363 76541 6364
rect 76867 6404 76925 6405
rect 76867 6364 76876 6404
rect 76916 6364 76925 6404
rect 76867 6363 76925 6364
rect 77251 6404 77309 6405
rect 77251 6364 77260 6404
rect 77300 6364 77309 6404
rect 77251 6363 77309 6364
rect 77635 6404 77693 6405
rect 77635 6364 77644 6404
rect 77684 6364 77693 6404
rect 77635 6363 77693 6364
rect 78115 6404 78173 6405
rect 78115 6364 78124 6404
rect 78164 6364 78173 6404
rect 78115 6363 78173 6364
rect 78499 6404 78557 6405
rect 78499 6364 78508 6404
rect 78548 6364 78557 6404
rect 78499 6363 78557 6364
rect 78883 6404 78941 6405
rect 78883 6364 78892 6404
rect 78932 6364 78941 6404
rect 78883 6363 78941 6364
rect 79267 6404 79325 6405
rect 79267 6364 79276 6404
rect 79316 6364 79325 6404
rect 79267 6363 79325 6364
rect 79747 6404 79805 6405
rect 79747 6364 79756 6404
rect 79796 6364 79805 6404
rect 79747 6363 79805 6364
rect 80131 6404 80189 6405
rect 80131 6364 80140 6404
rect 80180 6364 80189 6404
rect 80131 6363 80189 6364
rect 80515 6404 80573 6405
rect 80515 6364 80524 6404
rect 80564 6364 80573 6404
rect 80515 6363 80573 6364
rect 81283 6404 81341 6405
rect 81283 6364 81292 6404
rect 81332 6364 81341 6404
rect 81283 6363 81341 6364
rect 81667 6404 81725 6405
rect 81667 6364 81676 6404
rect 81716 6364 81725 6404
rect 81667 6363 81725 6364
rect 82051 6404 82109 6405
rect 82051 6364 82060 6404
rect 82100 6364 82109 6404
rect 82051 6363 82109 6364
rect 82531 6404 82589 6405
rect 82531 6364 82540 6404
rect 82580 6364 82589 6404
rect 82531 6363 82589 6364
rect 82915 6404 82973 6405
rect 82915 6364 82924 6404
rect 82964 6364 82973 6404
rect 82915 6363 82973 6364
rect 83683 6404 83741 6405
rect 83683 6364 83692 6404
rect 83732 6364 83741 6404
rect 83683 6363 83741 6364
rect 84067 6404 84125 6405
rect 84067 6364 84076 6404
rect 84116 6364 84125 6404
rect 84067 6363 84125 6364
rect 84451 6404 84509 6405
rect 84451 6364 84460 6404
rect 84500 6364 84509 6404
rect 84451 6363 84509 6364
rect 84835 6404 84893 6405
rect 84835 6364 84844 6404
rect 84884 6364 84893 6404
rect 84835 6363 84893 6364
rect 85315 6404 85373 6405
rect 85315 6364 85324 6404
rect 85364 6364 85373 6404
rect 85315 6363 85373 6364
rect 85699 6404 85757 6405
rect 85699 6364 85708 6404
rect 85748 6364 85757 6404
rect 85699 6363 85757 6364
rect 86083 6404 86141 6405
rect 86083 6364 86092 6404
rect 86132 6364 86141 6404
rect 86083 6363 86141 6364
rect 86467 6404 86525 6405
rect 86467 6364 86476 6404
rect 86516 6364 86525 6404
rect 86467 6363 86525 6364
rect 86851 6404 86909 6405
rect 86851 6364 86860 6404
rect 86900 6364 86909 6404
rect 86851 6363 86909 6364
rect 87331 6404 87389 6405
rect 87331 6364 87340 6404
rect 87380 6364 87389 6404
rect 87331 6363 87389 6364
rect 87907 6404 87965 6405
rect 87907 6364 87916 6404
rect 87956 6364 87965 6404
rect 87907 6363 87965 6364
rect 88099 6404 88157 6405
rect 88099 6364 88108 6404
rect 88148 6364 88157 6404
rect 88099 6363 88157 6364
rect 88483 6404 88541 6405
rect 88483 6364 88492 6404
rect 88532 6364 88541 6404
rect 88483 6363 88541 6364
rect 88867 6404 88925 6405
rect 88867 6364 88876 6404
rect 88916 6364 88925 6404
rect 88867 6363 88925 6364
rect 89251 6404 89309 6405
rect 89251 6364 89260 6404
rect 89300 6364 89309 6404
rect 89251 6363 89309 6364
rect 89731 6404 89789 6405
rect 89731 6364 89740 6404
rect 89780 6364 89789 6404
rect 89731 6363 89789 6364
rect 90115 6404 90173 6405
rect 90115 6364 90124 6404
rect 90164 6364 90173 6404
rect 90115 6363 90173 6364
rect 90499 6404 90557 6405
rect 90499 6364 90508 6404
rect 90548 6364 90557 6404
rect 90499 6363 90557 6364
rect 90883 6404 90941 6405
rect 90883 6364 90892 6404
rect 90932 6364 90941 6404
rect 90883 6363 90941 6364
rect 91267 6404 91325 6405
rect 91267 6364 91276 6404
rect 91316 6364 91325 6404
rect 91267 6363 91325 6364
rect 91747 6404 91805 6405
rect 91747 6364 91756 6404
rect 91796 6364 91805 6404
rect 91747 6363 91805 6364
rect 92131 6404 92189 6405
rect 92131 6364 92140 6404
rect 92180 6364 92189 6404
rect 92131 6363 92189 6364
rect 92515 6404 92573 6405
rect 92515 6364 92524 6404
rect 92564 6364 92573 6404
rect 92515 6363 92573 6364
rect 92899 6404 92957 6405
rect 92899 6364 92908 6404
rect 92948 6364 92957 6404
rect 92899 6363 92957 6364
rect 93379 6404 93437 6405
rect 93379 6364 93388 6404
rect 93428 6364 93437 6404
rect 93379 6363 93437 6364
rect 93955 6404 94013 6405
rect 93955 6364 93964 6404
rect 94004 6364 94013 6404
rect 93955 6363 94013 6364
rect 94147 6404 94205 6405
rect 94147 6364 94156 6404
rect 94196 6364 94205 6404
rect 94147 6363 94205 6364
rect 94531 6404 94589 6405
rect 94531 6364 94540 6404
rect 94580 6364 94589 6404
rect 94531 6363 94589 6364
rect 94915 6404 94973 6405
rect 94915 6364 94924 6404
rect 94964 6364 94973 6404
rect 94915 6363 94973 6364
rect 95395 6404 95453 6405
rect 95395 6364 95404 6404
rect 95444 6364 95453 6404
rect 95395 6363 95453 6364
rect 95779 6404 95837 6405
rect 95779 6364 95788 6404
rect 95828 6364 95837 6404
rect 95779 6363 95837 6364
rect 96163 6404 96221 6405
rect 96163 6364 96172 6404
rect 96212 6364 96221 6404
rect 96163 6363 96221 6364
rect 96547 6404 96605 6405
rect 96547 6364 96556 6404
rect 96596 6364 96605 6404
rect 96547 6363 96605 6364
rect 97219 6404 97277 6405
rect 97219 6364 97228 6404
rect 97268 6364 97277 6404
rect 97219 6363 97277 6364
rect 97699 6404 97757 6405
rect 97699 6364 97708 6404
rect 97748 6364 97757 6404
rect 97699 6363 97757 6364
rect 98083 6404 98141 6405
rect 98083 6364 98092 6404
rect 98132 6364 98141 6404
rect 98083 6363 98141 6364
rect 1323 6320 1365 6329
rect 1323 6280 1324 6320
rect 1364 6280 1365 6320
rect 1323 6271 1365 6280
rect 91947 6320 91989 6329
rect 91947 6280 91948 6320
rect 91988 6280 91989 6320
rect 91947 6271 91989 6280
rect 576 6068 99360 6092
rect 576 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 7112 6068
rect 7152 6028 7194 6068
rect 7234 6028 7276 6068
rect 7316 6028 7358 6068
rect 7398 6028 7440 6068
rect 7480 6028 11112 6068
rect 11152 6028 11194 6068
rect 11234 6028 11276 6068
rect 11316 6028 11358 6068
rect 11398 6028 11440 6068
rect 11480 6028 15112 6068
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15480 6028 19112 6068
rect 19152 6028 19194 6068
rect 19234 6028 19276 6068
rect 19316 6028 19358 6068
rect 19398 6028 19440 6068
rect 19480 6028 23112 6068
rect 23152 6028 23194 6068
rect 23234 6028 23276 6068
rect 23316 6028 23358 6068
rect 23398 6028 23440 6068
rect 23480 6028 27112 6068
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27480 6028 31112 6068
rect 31152 6028 31194 6068
rect 31234 6028 31276 6068
rect 31316 6028 31358 6068
rect 31398 6028 31440 6068
rect 31480 6028 35112 6068
rect 35152 6028 35194 6068
rect 35234 6028 35276 6068
rect 35316 6028 35358 6068
rect 35398 6028 35440 6068
rect 35480 6028 39112 6068
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39480 6028 43112 6068
rect 43152 6028 43194 6068
rect 43234 6028 43276 6068
rect 43316 6028 43358 6068
rect 43398 6028 43440 6068
rect 43480 6028 47112 6068
rect 47152 6028 47194 6068
rect 47234 6028 47276 6068
rect 47316 6028 47358 6068
rect 47398 6028 47440 6068
rect 47480 6028 51112 6068
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51480 6028 55112 6068
rect 55152 6028 55194 6068
rect 55234 6028 55276 6068
rect 55316 6028 55358 6068
rect 55398 6028 55440 6068
rect 55480 6028 59112 6068
rect 59152 6028 59194 6068
rect 59234 6028 59276 6068
rect 59316 6028 59358 6068
rect 59398 6028 59440 6068
rect 59480 6028 63112 6068
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63480 6028 67112 6068
rect 67152 6028 67194 6068
rect 67234 6028 67276 6068
rect 67316 6028 67358 6068
rect 67398 6028 67440 6068
rect 67480 6028 99360 6068
rect 576 6004 99360 6028
rect 81099 5900 81141 5909
rect 81099 5860 81100 5900
rect 81140 5860 81141 5900
rect 81099 5851 81141 5860
rect 83499 5900 83541 5909
rect 83499 5860 83500 5900
rect 83540 5860 83541 5900
rect 83499 5851 83541 5860
rect 91179 5900 91221 5909
rect 91179 5860 91180 5900
rect 91220 5860 91221 5900
rect 91179 5851 91221 5860
rect 94059 5900 94101 5909
rect 94059 5860 94060 5900
rect 94100 5860 94101 5900
rect 94059 5851 94101 5860
rect 835 5732 893 5733
rect 835 5692 844 5732
rect 884 5692 893 5732
rect 835 5691 893 5692
rect 80899 5732 80957 5733
rect 80899 5692 80908 5732
rect 80948 5692 80957 5732
rect 80899 5691 80957 5692
rect 83299 5732 83357 5733
rect 83299 5692 83308 5732
rect 83348 5692 83357 5732
rect 83299 5691 83357 5692
rect 91075 5648 91133 5649
rect 91075 5608 91084 5648
rect 91124 5608 91133 5648
rect 91075 5607 91133 5608
rect 93955 5648 94013 5649
rect 93955 5608 93964 5648
rect 94004 5608 94013 5648
rect 93955 5607 94013 5608
rect 651 5480 693 5489
rect 651 5440 652 5480
rect 692 5440 693 5480
rect 651 5431 693 5440
rect 576 5312 99360 5336
rect 576 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 8352 5312
rect 8392 5272 8434 5312
rect 8474 5272 8516 5312
rect 8556 5272 8598 5312
rect 8638 5272 8680 5312
rect 8720 5272 12352 5312
rect 12392 5272 12434 5312
rect 12474 5272 12516 5312
rect 12556 5272 12598 5312
rect 12638 5272 12680 5312
rect 12720 5272 16352 5312
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16720 5272 20352 5312
rect 20392 5272 20434 5312
rect 20474 5272 20516 5312
rect 20556 5272 20598 5312
rect 20638 5272 20680 5312
rect 20720 5272 24352 5312
rect 24392 5272 24434 5312
rect 24474 5272 24516 5312
rect 24556 5272 24598 5312
rect 24638 5272 24680 5312
rect 24720 5272 28352 5312
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28720 5272 32352 5312
rect 32392 5272 32434 5312
rect 32474 5272 32516 5312
rect 32556 5272 32598 5312
rect 32638 5272 32680 5312
rect 32720 5272 36352 5312
rect 36392 5272 36434 5312
rect 36474 5272 36516 5312
rect 36556 5272 36598 5312
rect 36638 5272 36680 5312
rect 36720 5272 40352 5312
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40720 5272 44352 5312
rect 44392 5272 44434 5312
rect 44474 5272 44516 5312
rect 44556 5272 44598 5312
rect 44638 5272 44680 5312
rect 44720 5272 48352 5312
rect 48392 5272 48434 5312
rect 48474 5272 48516 5312
rect 48556 5272 48598 5312
rect 48638 5272 48680 5312
rect 48720 5272 52352 5312
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52720 5272 56352 5312
rect 56392 5272 56434 5312
rect 56474 5272 56516 5312
rect 56556 5272 56598 5312
rect 56638 5272 56680 5312
rect 56720 5272 60352 5312
rect 60392 5272 60434 5312
rect 60474 5272 60516 5312
rect 60556 5272 60598 5312
rect 60638 5272 60680 5312
rect 60720 5272 64352 5312
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64720 5272 68352 5312
rect 68392 5272 68434 5312
rect 68474 5272 68516 5312
rect 68556 5272 68598 5312
rect 68638 5272 68680 5312
rect 68720 5272 72352 5312
rect 72392 5272 72434 5312
rect 72474 5272 72516 5312
rect 72556 5272 72598 5312
rect 72638 5272 72680 5312
rect 72720 5272 76352 5312
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76720 5272 80352 5312
rect 80392 5272 80434 5312
rect 80474 5272 80516 5312
rect 80556 5272 80598 5312
rect 80638 5272 80680 5312
rect 80720 5272 84352 5312
rect 84392 5272 84434 5312
rect 84474 5272 84516 5312
rect 84556 5272 84598 5312
rect 84638 5272 84680 5312
rect 84720 5272 88352 5312
rect 88392 5272 88434 5312
rect 88474 5272 88516 5312
rect 88556 5272 88598 5312
rect 88638 5272 88680 5312
rect 88720 5272 92352 5312
rect 92392 5272 92434 5312
rect 92474 5272 92516 5312
rect 92556 5272 92598 5312
rect 92638 5272 92680 5312
rect 92720 5272 96352 5312
rect 96392 5272 96434 5312
rect 96474 5272 96516 5312
rect 96556 5272 96598 5312
rect 96638 5272 96680 5312
rect 96720 5272 99360 5312
rect 576 5248 99360 5272
rect 1027 4892 1085 4893
rect 1027 4852 1036 4892
rect 1076 4852 1085 4892
rect 1027 4851 1085 4852
rect 1411 4892 1469 4893
rect 1411 4852 1420 4892
rect 1460 4852 1469 4892
rect 1411 4851 1469 4852
rect 1795 4892 1853 4893
rect 1795 4852 1804 4892
rect 1844 4852 1853 4892
rect 1795 4851 1853 4852
rect 2179 4892 2237 4893
rect 2179 4852 2188 4892
rect 2228 4852 2237 4892
rect 2179 4851 2237 4852
rect 843 4724 885 4733
rect 843 4684 844 4724
rect 884 4684 885 4724
rect 843 4675 885 4684
rect 1227 4724 1269 4733
rect 1227 4684 1228 4724
rect 1268 4684 1269 4724
rect 1227 4675 1269 4684
rect 1611 4724 1653 4733
rect 1611 4684 1612 4724
rect 1652 4684 1653 4724
rect 1611 4675 1653 4684
rect 1995 4724 2037 4733
rect 1995 4684 1996 4724
rect 2036 4684 2037 4724
rect 1995 4675 2037 4684
rect 576 4556 99516 4580
rect 576 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 7112 4556
rect 7152 4516 7194 4556
rect 7234 4516 7276 4556
rect 7316 4516 7358 4556
rect 7398 4516 7440 4556
rect 7480 4516 11112 4556
rect 11152 4516 11194 4556
rect 11234 4516 11276 4556
rect 11316 4516 11358 4556
rect 11398 4516 11440 4556
rect 11480 4516 15112 4556
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15480 4516 19112 4556
rect 19152 4516 19194 4556
rect 19234 4516 19276 4556
rect 19316 4516 19358 4556
rect 19398 4516 19440 4556
rect 19480 4516 23112 4556
rect 23152 4516 23194 4556
rect 23234 4516 23276 4556
rect 23316 4516 23358 4556
rect 23398 4516 23440 4556
rect 23480 4516 27112 4556
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27480 4516 31112 4556
rect 31152 4516 31194 4556
rect 31234 4516 31276 4556
rect 31316 4516 31358 4556
rect 31398 4516 31440 4556
rect 31480 4516 35112 4556
rect 35152 4516 35194 4556
rect 35234 4516 35276 4556
rect 35316 4516 35358 4556
rect 35398 4516 35440 4556
rect 35480 4516 39112 4556
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39480 4516 43112 4556
rect 43152 4516 43194 4556
rect 43234 4516 43276 4556
rect 43316 4516 43358 4556
rect 43398 4516 43440 4556
rect 43480 4516 47112 4556
rect 47152 4516 47194 4556
rect 47234 4516 47276 4556
rect 47316 4516 47358 4556
rect 47398 4516 47440 4556
rect 47480 4516 51112 4556
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51480 4516 55112 4556
rect 55152 4516 55194 4556
rect 55234 4516 55276 4556
rect 55316 4516 55358 4556
rect 55398 4516 55440 4556
rect 55480 4516 59112 4556
rect 59152 4516 59194 4556
rect 59234 4516 59276 4556
rect 59316 4516 59358 4556
rect 59398 4516 59440 4556
rect 59480 4516 63112 4556
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63480 4516 67112 4556
rect 67152 4516 67194 4556
rect 67234 4516 67276 4556
rect 67316 4516 67358 4556
rect 67398 4516 67440 4556
rect 67480 4516 71112 4556
rect 71152 4516 71194 4556
rect 71234 4516 71276 4556
rect 71316 4516 71358 4556
rect 71398 4516 71440 4556
rect 71480 4516 75112 4556
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75480 4516 79112 4556
rect 79152 4516 79194 4556
rect 79234 4516 79276 4556
rect 79316 4516 79358 4556
rect 79398 4516 79440 4556
rect 79480 4516 83112 4556
rect 83152 4516 83194 4556
rect 83234 4516 83276 4556
rect 83316 4516 83358 4556
rect 83398 4516 83440 4556
rect 83480 4516 87112 4556
rect 87152 4516 87194 4556
rect 87234 4516 87276 4556
rect 87316 4516 87358 4556
rect 87398 4516 87440 4556
rect 87480 4516 91112 4556
rect 91152 4516 91194 4556
rect 91234 4516 91276 4556
rect 91316 4516 91358 4556
rect 91398 4516 91440 4556
rect 91480 4516 95112 4556
rect 95152 4516 95194 4556
rect 95234 4516 95276 4556
rect 95316 4516 95358 4556
rect 95398 4516 95440 4556
rect 95480 4516 99112 4556
rect 99152 4516 99194 4556
rect 99234 4516 99276 4556
rect 99316 4516 99358 4556
rect 99398 4516 99440 4556
rect 99480 4516 99516 4556
rect 576 4492 99516 4516
rect 651 4388 693 4397
rect 651 4348 652 4388
rect 692 4348 693 4388
rect 651 4339 693 4348
rect 835 4220 893 4221
rect 835 4180 844 4220
rect 884 4180 893 4220
rect 835 4179 893 4180
rect 1219 4220 1277 4221
rect 1219 4180 1228 4220
rect 1268 4180 1277 4220
rect 1219 4179 1277 4180
rect 1035 3968 1077 3977
rect 1035 3928 1036 3968
rect 1076 3928 1077 3968
rect 1035 3919 1077 3928
rect 576 3800 99360 3824
rect 576 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 8352 3800
rect 8392 3760 8434 3800
rect 8474 3760 8516 3800
rect 8556 3760 8598 3800
rect 8638 3760 8680 3800
rect 8720 3760 12352 3800
rect 12392 3760 12434 3800
rect 12474 3760 12516 3800
rect 12556 3760 12598 3800
rect 12638 3760 12680 3800
rect 12720 3760 16352 3800
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16720 3760 20352 3800
rect 20392 3760 20434 3800
rect 20474 3760 20516 3800
rect 20556 3760 20598 3800
rect 20638 3760 20680 3800
rect 20720 3760 24352 3800
rect 24392 3760 24434 3800
rect 24474 3760 24516 3800
rect 24556 3760 24598 3800
rect 24638 3760 24680 3800
rect 24720 3760 28352 3800
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28720 3760 32352 3800
rect 32392 3760 32434 3800
rect 32474 3760 32516 3800
rect 32556 3760 32598 3800
rect 32638 3760 32680 3800
rect 32720 3760 36352 3800
rect 36392 3760 36434 3800
rect 36474 3760 36516 3800
rect 36556 3760 36598 3800
rect 36638 3760 36680 3800
rect 36720 3760 40352 3800
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40720 3760 44352 3800
rect 44392 3760 44434 3800
rect 44474 3760 44516 3800
rect 44556 3760 44598 3800
rect 44638 3760 44680 3800
rect 44720 3760 48352 3800
rect 48392 3760 48434 3800
rect 48474 3760 48516 3800
rect 48556 3760 48598 3800
rect 48638 3760 48680 3800
rect 48720 3760 52352 3800
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52720 3760 56352 3800
rect 56392 3760 56434 3800
rect 56474 3760 56516 3800
rect 56556 3760 56598 3800
rect 56638 3760 56680 3800
rect 56720 3760 60352 3800
rect 60392 3760 60434 3800
rect 60474 3760 60516 3800
rect 60556 3760 60598 3800
rect 60638 3760 60680 3800
rect 60720 3760 64352 3800
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64720 3760 68352 3800
rect 68392 3760 68434 3800
rect 68474 3760 68516 3800
rect 68556 3760 68598 3800
rect 68638 3760 68680 3800
rect 68720 3760 72352 3800
rect 72392 3760 72434 3800
rect 72474 3760 72516 3800
rect 72556 3760 72598 3800
rect 72638 3760 72680 3800
rect 72720 3760 76352 3800
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76720 3760 80352 3800
rect 80392 3760 80434 3800
rect 80474 3760 80516 3800
rect 80556 3760 80598 3800
rect 80638 3760 80680 3800
rect 80720 3760 84352 3800
rect 84392 3760 84434 3800
rect 84474 3760 84516 3800
rect 84556 3760 84598 3800
rect 84638 3760 84680 3800
rect 84720 3760 88352 3800
rect 88392 3760 88434 3800
rect 88474 3760 88516 3800
rect 88556 3760 88598 3800
rect 88638 3760 88680 3800
rect 88720 3760 92352 3800
rect 92392 3760 92434 3800
rect 92474 3760 92516 3800
rect 92556 3760 92598 3800
rect 92638 3760 92680 3800
rect 92720 3760 96352 3800
rect 96392 3760 96434 3800
rect 96474 3760 96516 3800
rect 96556 3760 96598 3800
rect 96638 3760 96680 3800
rect 96720 3760 99360 3800
rect 576 3736 99360 3760
rect 835 3380 893 3381
rect 835 3340 844 3380
rect 884 3340 893 3380
rect 835 3339 893 3340
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 576 3044 99516 3068
rect 576 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 7112 3044
rect 7152 3004 7194 3044
rect 7234 3004 7276 3044
rect 7316 3004 7358 3044
rect 7398 3004 7440 3044
rect 7480 3004 11112 3044
rect 11152 3004 11194 3044
rect 11234 3004 11276 3044
rect 11316 3004 11358 3044
rect 11398 3004 11440 3044
rect 11480 3004 15112 3044
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15480 3004 19112 3044
rect 19152 3004 19194 3044
rect 19234 3004 19276 3044
rect 19316 3004 19358 3044
rect 19398 3004 19440 3044
rect 19480 3004 23112 3044
rect 23152 3004 23194 3044
rect 23234 3004 23276 3044
rect 23316 3004 23358 3044
rect 23398 3004 23440 3044
rect 23480 3004 27112 3044
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27480 3004 31112 3044
rect 31152 3004 31194 3044
rect 31234 3004 31276 3044
rect 31316 3004 31358 3044
rect 31398 3004 31440 3044
rect 31480 3004 35112 3044
rect 35152 3004 35194 3044
rect 35234 3004 35276 3044
rect 35316 3004 35358 3044
rect 35398 3004 35440 3044
rect 35480 3004 39112 3044
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39480 3004 43112 3044
rect 43152 3004 43194 3044
rect 43234 3004 43276 3044
rect 43316 3004 43358 3044
rect 43398 3004 43440 3044
rect 43480 3004 47112 3044
rect 47152 3004 47194 3044
rect 47234 3004 47276 3044
rect 47316 3004 47358 3044
rect 47398 3004 47440 3044
rect 47480 3004 51112 3044
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51480 3004 55112 3044
rect 55152 3004 55194 3044
rect 55234 3004 55276 3044
rect 55316 3004 55358 3044
rect 55398 3004 55440 3044
rect 55480 3004 59112 3044
rect 59152 3004 59194 3044
rect 59234 3004 59276 3044
rect 59316 3004 59358 3044
rect 59398 3004 59440 3044
rect 59480 3004 63112 3044
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63480 3004 67112 3044
rect 67152 3004 67194 3044
rect 67234 3004 67276 3044
rect 67316 3004 67358 3044
rect 67398 3004 67440 3044
rect 67480 3004 71112 3044
rect 71152 3004 71194 3044
rect 71234 3004 71276 3044
rect 71316 3004 71358 3044
rect 71398 3004 71440 3044
rect 71480 3004 75112 3044
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75480 3004 79112 3044
rect 79152 3004 79194 3044
rect 79234 3004 79276 3044
rect 79316 3004 79358 3044
rect 79398 3004 79440 3044
rect 79480 3004 83112 3044
rect 83152 3004 83194 3044
rect 83234 3004 83276 3044
rect 83316 3004 83358 3044
rect 83398 3004 83440 3044
rect 83480 3004 87112 3044
rect 87152 3004 87194 3044
rect 87234 3004 87276 3044
rect 87316 3004 87358 3044
rect 87398 3004 87440 3044
rect 87480 3004 91112 3044
rect 91152 3004 91194 3044
rect 91234 3004 91276 3044
rect 91316 3004 91358 3044
rect 91398 3004 91440 3044
rect 91480 3004 95112 3044
rect 95152 3004 95194 3044
rect 95234 3004 95276 3044
rect 95316 3004 95358 3044
rect 95398 3004 95440 3044
rect 95480 3004 99112 3044
rect 99152 3004 99194 3044
rect 99234 3004 99276 3044
rect 99316 3004 99358 3044
rect 99398 3004 99440 3044
rect 99480 3004 99516 3044
rect 576 2980 99516 3004
rect 835 2708 893 2709
rect 835 2668 844 2708
rect 884 2668 893 2708
rect 835 2667 893 2668
rect 651 2456 693 2465
rect 651 2416 652 2456
rect 692 2416 693 2456
rect 651 2407 693 2416
rect 576 2288 99360 2312
rect 576 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 8352 2288
rect 8392 2248 8434 2288
rect 8474 2248 8516 2288
rect 8556 2248 8598 2288
rect 8638 2248 8680 2288
rect 8720 2248 12352 2288
rect 12392 2248 12434 2288
rect 12474 2248 12516 2288
rect 12556 2248 12598 2288
rect 12638 2248 12680 2288
rect 12720 2248 16352 2288
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16720 2248 20352 2288
rect 20392 2248 20434 2288
rect 20474 2248 20516 2288
rect 20556 2248 20598 2288
rect 20638 2248 20680 2288
rect 20720 2248 24352 2288
rect 24392 2248 24434 2288
rect 24474 2248 24516 2288
rect 24556 2248 24598 2288
rect 24638 2248 24680 2288
rect 24720 2248 28352 2288
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28720 2248 32352 2288
rect 32392 2248 32434 2288
rect 32474 2248 32516 2288
rect 32556 2248 32598 2288
rect 32638 2248 32680 2288
rect 32720 2248 36352 2288
rect 36392 2248 36434 2288
rect 36474 2248 36516 2288
rect 36556 2248 36598 2288
rect 36638 2248 36680 2288
rect 36720 2248 40352 2288
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40720 2248 44352 2288
rect 44392 2248 44434 2288
rect 44474 2248 44516 2288
rect 44556 2248 44598 2288
rect 44638 2248 44680 2288
rect 44720 2248 48352 2288
rect 48392 2248 48434 2288
rect 48474 2248 48516 2288
rect 48556 2248 48598 2288
rect 48638 2248 48680 2288
rect 48720 2248 52352 2288
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52720 2248 56352 2288
rect 56392 2248 56434 2288
rect 56474 2248 56516 2288
rect 56556 2248 56598 2288
rect 56638 2248 56680 2288
rect 56720 2248 60352 2288
rect 60392 2248 60434 2288
rect 60474 2248 60516 2288
rect 60556 2248 60598 2288
rect 60638 2248 60680 2288
rect 60720 2248 64352 2288
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64720 2248 68352 2288
rect 68392 2248 68434 2288
rect 68474 2248 68516 2288
rect 68556 2248 68598 2288
rect 68638 2248 68680 2288
rect 68720 2248 72352 2288
rect 72392 2248 72434 2288
rect 72474 2248 72516 2288
rect 72556 2248 72598 2288
rect 72638 2248 72680 2288
rect 72720 2248 76352 2288
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76720 2248 80352 2288
rect 80392 2248 80434 2288
rect 80474 2248 80516 2288
rect 80556 2248 80598 2288
rect 80638 2248 80680 2288
rect 80720 2248 84352 2288
rect 84392 2248 84434 2288
rect 84474 2248 84516 2288
rect 84556 2248 84598 2288
rect 84638 2248 84680 2288
rect 84720 2248 88352 2288
rect 88392 2248 88434 2288
rect 88474 2248 88516 2288
rect 88556 2248 88598 2288
rect 88638 2248 88680 2288
rect 88720 2248 92352 2288
rect 92392 2248 92434 2288
rect 92474 2248 92516 2288
rect 92556 2248 92598 2288
rect 92638 2248 92680 2288
rect 92720 2248 96352 2288
rect 96392 2248 96434 2288
rect 96474 2248 96516 2288
rect 96556 2248 96598 2288
rect 96638 2248 96680 2288
rect 96720 2248 99360 2288
rect 576 2224 99360 2248
rect 576 1532 99516 1556
rect 576 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 7112 1532
rect 7152 1492 7194 1532
rect 7234 1492 7276 1532
rect 7316 1492 7358 1532
rect 7398 1492 7440 1532
rect 7480 1492 11112 1532
rect 11152 1492 11194 1532
rect 11234 1492 11276 1532
rect 11316 1492 11358 1532
rect 11398 1492 11440 1532
rect 11480 1492 15112 1532
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15480 1492 19112 1532
rect 19152 1492 19194 1532
rect 19234 1492 19276 1532
rect 19316 1492 19358 1532
rect 19398 1492 19440 1532
rect 19480 1492 23112 1532
rect 23152 1492 23194 1532
rect 23234 1492 23276 1532
rect 23316 1492 23358 1532
rect 23398 1492 23440 1532
rect 23480 1492 27112 1532
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27480 1492 31112 1532
rect 31152 1492 31194 1532
rect 31234 1492 31276 1532
rect 31316 1492 31358 1532
rect 31398 1492 31440 1532
rect 31480 1492 35112 1532
rect 35152 1492 35194 1532
rect 35234 1492 35276 1532
rect 35316 1492 35358 1532
rect 35398 1492 35440 1532
rect 35480 1492 39112 1532
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39480 1492 43112 1532
rect 43152 1492 43194 1532
rect 43234 1492 43276 1532
rect 43316 1492 43358 1532
rect 43398 1492 43440 1532
rect 43480 1492 47112 1532
rect 47152 1492 47194 1532
rect 47234 1492 47276 1532
rect 47316 1492 47358 1532
rect 47398 1492 47440 1532
rect 47480 1492 51112 1532
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51480 1492 55112 1532
rect 55152 1492 55194 1532
rect 55234 1492 55276 1532
rect 55316 1492 55358 1532
rect 55398 1492 55440 1532
rect 55480 1492 59112 1532
rect 59152 1492 59194 1532
rect 59234 1492 59276 1532
rect 59316 1492 59358 1532
rect 59398 1492 59440 1532
rect 59480 1492 63112 1532
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63480 1492 67112 1532
rect 67152 1492 67194 1532
rect 67234 1492 67276 1532
rect 67316 1492 67358 1532
rect 67398 1492 67440 1532
rect 67480 1492 71112 1532
rect 71152 1492 71194 1532
rect 71234 1492 71276 1532
rect 71316 1492 71358 1532
rect 71398 1492 71440 1532
rect 71480 1492 75112 1532
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75480 1492 79112 1532
rect 79152 1492 79194 1532
rect 79234 1492 79276 1532
rect 79316 1492 79358 1532
rect 79398 1492 79440 1532
rect 79480 1492 83112 1532
rect 83152 1492 83194 1532
rect 83234 1492 83276 1532
rect 83316 1492 83358 1532
rect 83398 1492 83440 1532
rect 83480 1492 87112 1532
rect 87152 1492 87194 1532
rect 87234 1492 87276 1532
rect 87316 1492 87358 1532
rect 87398 1492 87440 1532
rect 87480 1492 91112 1532
rect 91152 1492 91194 1532
rect 91234 1492 91276 1532
rect 91316 1492 91358 1532
rect 91398 1492 91440 1532
rect 91480 1492 95112 1532
rect 95152 1492 95194 1532
rect 95234 1492 95276 1532
rect 95316 1492 95358 1532
rect 95398 1492 95440 1532
rect 95480 1492 99112 1532
rect 99152 1492 99194 1532
rect 99234 1492 99276 1532
rect 99316 1492 99358 1532
rect 99398 1492 99440 1532
rect 99480 1492 99516 1532
rect 576 1468 99516 1492
rect 576 776 99360 800
rect 576 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 8352 776
rect 8392 736 8434 776
rect 8474 736 8516 776
rect 8556 736 8598 776
rect 8638 736 8680 776
rect 8720 736 12352 776
rect 12392 736 12434 776
rect 12474 736 12516 776
rect 12556 736 12598 776
rect 12638 736 12680 776
rect 12720 736 16352 776
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16720 736 20352 776
rect 20392 736 20434 776
rect 20474 736 20516 776
rect 20556 736 20598 776
rect 20638 736 20680 776
rect 20720 736 24352 776
rect 24392 736 24434 776
rect 24474 736 24516 776
rect 24556 736 24598 776
rect 24638 736 24680 776
rect 24720 736 28352 776
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28720 736 32352 776
rect 32392 736 32434 776
rect 32474 736 32516 776
rect 32556 736 32598 776
rect 32638 736 32680 776
rect 32720 736 36352 776
rect 36392 736 36434 776
rect 36474 736 36516 776
rect 36556 736 36598 776
rect 36638 736 36680 776
rect 36720 736 40352 776
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40720 736 44352 776
rect 44392 736 44434 776
rect 44474 736 44516 776
rect 44556 736 44598 776
rect 44638 736 44680 776
rect 44720 736 48352 776
rect 48392 736 48434 776
rect 48474 736 48516 776
rect 48556 736 48598 776
rect 48638 736 48680 776
rect 48720 736 52352 776
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52720 736 56352 776
rect 56392 736 56434 776
rect 56474 736 56516 776
rect 56556 736 56598 776
rect 56638 736 56680 776
rect 56720 736 60352 776
rect 60392 736 60434 776
rect 60474 736 60516 776
rect 60556 736 60598 776
rect 60638 736 60680 776
rect 60720 736 64352 776
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64720 736 68352 776
rect 68392 736 68434 776
rect 68474 736 68516 776
rect 68556 736 68598 776
rect 68638 736 68680 776
rect 68720 736 72352 776
rect 72392 736 72434 776
rect 72474 736 72516 776
rect 72556 736 72598 776
rect 72638 736 72680 776
rect 72720 736 76352 776
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76720 736 80352 776
rect 80392 736 80434 776
rect 80474 736 80516 776
rect 80556 736 80598 776
rect 80638 736 80680 776
rect 80720 736 84352 776
rect 84392 736 84434 776
rect 84474 736 84516 776
rect 84556 736 84598 776
rect 84638 736 84680 776
rect 84720 736 88352 776
rect 88392 736 88434 776
rect 88474 736 88516 776
rect 88556 736 88598 776
rect 88638 736 88680 776
rect 88720 736 92352 776
rect 92392 736 92434 776
rect 92474 736 92516 776
rect 92556 736 92598 776
rect 92638 736 92680 776
rect 92720 736 96352 776
rect 96392 736 96434 776
rect 96474 736 96516 776
rect 96556 736 96598 776
rect 96638 736 96680 776
rect 96720 736 99360 776
rect 576 712 99360 736
<< via1 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 8352 38536 8392 38576
rect 8434 38536 8474 38576
rect 8516 38536 8556 38576
rect 8598 38536 8638 38576
rect 8680 38536 8720 38576
rect 12352 38536 12392 38576
rect 12434 38536 12474 38576
rect 12516 38536 12556 38576
rect 12598 38536 12638 38576
rect 12680 38536 12720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 20352 38536 20392 38576
rect 20434 38536 20474 38576
rect 20516 38536 20556 38576
rect 20598 38536 20638 38576
rect 20680 38536 20720 38576
rect 24352 38536 24392 38576
rect 24434 38536 24474 38576
rect 24516 38536 24556 38576
rect 24598 38536 24638 38576
rect 24680 38536 24720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 32352 38536 32392 38576
rect 32434 38536 32474 38576
rect 32516 38536 32556 38576
rect 32598 38536 32638 38576
rect 32680 38536 32720 38576
rect 36352 38536 36392 38576
rect 36434 38536 36474 38576
rect 36516 38536 36556 38576
rect 36598 38536 36638 38576
rect 36680 38536 36720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 44352 38536 44392 38576
rect 44434 38536 44474 38576
rect 44516 38536 44556 38576
rect 44598 38536 44638 38576
rect 44680 38536 44720 38576
rect 48352 38536 48392 38576
rect 48434 38536 48474 38576
rect 48516 38536 48556 38576
rect 48598 38536 48638 38576
rect 48680 38536 48720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 56352 38536 56392 38576
rect 56434 38536 56474 38576
rect 56516 38536 56556 38576
rect 56598 38536 56638 38576
rect 56680 38536 56720 38576
rect 60352 38536 60392 38576
rect 60434 38536 60474 38576
rect 60516 38536 60556 38576
rect 60598 38536 60638 38576
rect 60680 38536 60720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 68352 38536 68392 38576
rect 68434 38536 68474 38576
rect 68516 38536 68556 38576
rect 68598 38536 68638 38576
rect 68680 38536 68720 38576
rect 72352 38536 72392 38576
rect 72434 38536 72474 38576
rect 72516 38536 72556 38576
rect 72598 38536 72638 38576
rect 72680 38536 72720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 80352 38536 80392 38576
rect 80434 38536 80474 38576
rect 80516 38536 80556 38576
rect 80598 38536 80638 38576
rect 80680 38536 80720 38576
rect 84352 38536 84392 38576
rect 84434 38536 84474 38576
rect 84516 38536 84556 38576
rect 84598 38536 84638 38576
rect 84680 38536 84720 38576
rect 88352 38536 88392 38576
rect 88434 38536 88474 38576
rect 88516 38536 88556 38576
rect 88598 38536 88638 38576
rect 88680 38536 88720 38576
rect 92352 38536 92392 38576
rect 92434 38536 92474 38576
rect 92516 38536 92556 38576
rect 92598 38536 92638 38576
rect 92680 38536 92720 38576
rect 96352 38536 96392 38576
rect 96434 38536 96474 38576
rect 96516 38536 96556 38576
rect 96598 38536 96638 38576
rect 96680 38536 96720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 7112 37780 7152 37820
rect 7194 37780 7234 37820
rect 7276 37780 7316 37820
rect 7358 37780 7398 37820
rect 7440 37780 7480 37820
rect 11112 37780 11152 37820
rect 11194 37780 11234 37820
rect 11276 37780 11316 37820
rect 11358 37780 11398 37820
rect 11440 37780 11480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 19112 37780 19152 37820
rect 19194 37780 19234 37820
rect 19276 37780 19316 37820
rect 19358 37780 19398 37820
rect 19440 37780 19480 37820
rect 23112 37780 23152 37820
rect 23194 37780 23234 37820
rect 23276 37780 23316 37820
rect 23358 37780 23398 37820
rect 23440 37780 23480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 31112 37780 31152 37820
rect 31194 37780 31234 37820
rect 31276 37780 31316 37820
rect 31358 37780 31398 37820
rect 31440 37780 31480 37820
rect 35112 37780 35152 37820
rect 35194 37780 35234 37820
rect 35276 37780 35316 37820
rect 35358 37780 35398 37820
rect 35440 37780 35480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 43112 37780 43152 37820
rect 43194 37780 43234 37820
rect 43276 37780 43316 37820
rect 43358 37780 43398 37820
rect 43440 37780 43480 37820
rect 47112 37780 47152 37820
rect 47194 37780 47234 37820
rect 47276 37780 47316 37820
rect 47358 37780 47398 37820
rect 47440 37780 47480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 55112 37780 55152 37820
rect 55194 37780 55234 37820
rect 55276 37780 55316 37820
rect 55358 37780 55398 37820
rect 55440 37780 55480 37820
rect 59112 37780 59152 37820
rect 59194 37780 59234 37820
rect 59276 37780 59316 37820
rect 59358 37780 59398 37820
rect 59440 37780 59480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 67112 37780 67152 37820
rect 67194 37780 67234 37820
rect 67276 37780 67316 37820
rect 67358 37780 67398 37820
rect 67440 37780 67480 37820
rect 71112 37780 71152 37820
rect 71194 37780 71234 37820
rect 71276 37780 71316 37820
rect 71358 37780 71398 37820
rect 71440 37780 71480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 79112 37780 79152 37820
rect 79194 37780 79234 37820
rect 79276 37780 79316 37820
rect 79358 37780 79398 37820
rect 79440 37780 79480 37820
rect 83112 37780 83152 37820
rect 83194 37780 83234 37820
rect 83276 37780 83316 37820
rect 83358 37780 83398 37820
rect 83440 37780 83480 37820
rect 87112 37780 87152 37820
rect 87194 37780 87234 37820
rect 87276 37780 87316 37820
rect 87358 37780 87398 37820
rect 87440 37780 87480 37820
rect 91112 37780 91152 37820
rect 91194 37780 91234 37820
rect 91276 37780 91316 37820
rect 91358 37780 91398 37820
rect 91440 37780 91480 37820
rect 95112 37780 95152 37820
rect 95194 37780 95234 37820
rect 95276 37780 95316 37820
rect 95358 37780 95398 37820
rect 95440 37780 95480 37820
rect 99112 37780 99152 37820
rect 99194 37780 99234 37820
rect 99276 37780 99316 37820
rect 99358 37780 99398 37820
rect 99440 37780 99480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 8352 37024 8392 37064
rect 8434 37024 8474 37064
rect 8516 37024 8556 37064
rect 8598 37024 8638 37064
rect 8680 37024 8720 37064
rect 12352 37024 12392 37064
rect 12434 37024 12474 37064
rect 12516 37024 12556 37064
rect 12598 37024 12638 37064
rect 12680 37024 12720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 20352 37024 20392 37064
rect 20434 37024 20474 37064
rect 20516 37024 20556 37064
rect 20598 37024 20638 37064
rect 20680 37024 20720 37064
rect 24352 37024 24392 37064
rect 24434 37024 24474 37064
rect 24516 37024 24556 37064
rect 24598 37024 24638 37064
rect 24680 37024 24720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 32352 37024 32392 37064
rect 32434 37024 32474 37064
rect 32516 37024 32556 37064
rect 32598 37024 32638 37064
rect 32680 37024 32720 37064
rect 36352 37024 36392 37064
rect 36434 37024 36474 37064
rect 36516 37024 36556 37064
rect 36598 37024 36638 37064
rect 36680 37024 36720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 44352 37024 44392 37064
rect 44434 37024 44474 37064
rect 44516 37024 44556 37064
rect 44598 37024 44638 37064
rect 44680 37024 44720 37064
rect 48352 37024 48392 37064
rect 48434 37024 48474 37064
rect 48516 37024 48556 37064
rect 48598 37024 48638 37064
rect 48680 37024 48720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 56352 37024 56392 37064
rect 56434 37024 56474 37064
rect 56516 37024 56556 37064
rect 56598 37024 56638 37064
rect 56680 37024 56720 37064
rect 60352 37024 60392 37064
rect 60434 37024 60474 37064
rect 60516 37024 60556 37064
rect 60598 37024 60638 37064
rect 60680 37024 60720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 68352 37024 68392 37064
rect 68434 37024 68474 37064
rect 68516 37024 68556 37064
rect 68598 37024 68638 37064
rect 68680 37024 68720 37064
rect 72352 37024 72392 37064
rect 72434 37024 72474 37064
rect 72516 37024 72556 37064
rect 72598 37024 72638 37064
rect 72680 37024 72720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 80352 37024 80392 37064
rect 80434 37024 80474 37064
rect 80516 37024 80556 37064
rect 80598 37024 80638 37064
rect 80680 37024 80720 37064
rect 84352 37024 84392 37064
rect 84434 37024 84474 37064
rect 84516 37024 84556 37064
rect 84598 37024 84638 37064
rect 84680 37024 84720 37064
rect 88352 37024 88392 37064
rect 88434 37024 88474 37064
rect 88516 37024 88556 37064
rect 88598 37024 88638 37064
rect 88680 37024 88720 37064
rect 92352 37024 92392 37064
rect 92434 37024 92474 37064
rect 92516 37024 92556 37064
rect 92598 37024 92638 37064
rect 92680 37024 92720 37064
rect 96352 37024 96392 37064
rect 96434 37024 96474 37064
rect 96516 37024 96556 37064
rect 96598 37024 96638 37064
rect 96680 37024 96720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 7112 36268 7152 36308
rect 7194 36268 7234 36308
rect 7276 36268 7316 36308
rect 7358 36268 7398 36308
rect 7440 36268 7480 36308
rect 11112 36268 11152 36308
rect 11194 36268 11234 36308
rect 11276 36268 11316 36308
rect 11358 36268 11398 36308
rect 11440 36268 11480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 19112 36268 19152 36308
rect 19194 36268 19234 36308
rect 19276 36268 19316 36308
rect 19358 36268 19398 36308
rect 19440 36268 19480 36308
rect 23112 36268 23152 36308
rect 23194 36268 23234 36308
rect 23276 36268 23316 36308
rect 23358 36268 23398 36308
rect 23440 36268 23480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 31112 36268 31152 36308
rect 31194 36268 31234 36308
rect 31276 36268 31316 36308
rect 31358 36268 31398 36308
rect 31440 36268 31480 36308
rect 35112 36268 35152 36308
rect 35194 36268 35234 36308
rect 35276 36268 35316 36308
rect 35358 36268 35398 36308
rect 35440 36268 35480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 43112 36268 43152 36308
rect 43194 36268 43234 36308
rect 43276 36268 43316 36308
rect 43358 36268 43398 36308
rect 43440 36268 43480 36308
rect 47112 36268 47152 36308
rect 47194 36268 47234 36308
rect 47276 36268 47316 36308
rect 47358 36268 47398 36308
rect 47440 36268 47480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 55112 36268 55152 36308
rect 55194 36268 55234 36308
rect 55276 36268 55316 36308
rect 55358 36268 55398 36308
rect 55440 36268 55480 36308
rect 59112 36268 59152 36308
rect 59194 36268 59234 36308
rect 59276 36268 59316 36308
rect 59358 36268 59398 36308
rect 59440 36268 59480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 67112 36268 67152 36308
rect 67194 36268 67234 36308
rect 67276 36268 67316 36308
rect 67358 36268 67398 36308
rect 67440 36268 67480 36308
rect 71112 36268 71152 36308
rect 71194 36268 71234 36308
rect 71276 36268 71316 36308
rect 71358 36268 71398 36308
rect 71440 36268 71480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 79112 36268 79152 36308
rect 79194 36268 79234 36308
rect 79276 36268 79316 36308
rect 79358 36268 79398 36308
rect 79440 36268 79480 36308
rect 83112 36268 83152 36308
rect 83194 36268 83234 36308
rect 83276 36268 83316 36308
rect 83358 36268 83398 36308
rect 83440 36268 83480 36308
rect 87112 36268 87152 36308
rect 87194 36268 87234 36308
rect 87276 36268 87316 36308
rect 87358 36268 87398 36308
rect 87440 36268 87480 36308
rect 91112 36268 91152 36308
rect 91194 36268 91234 36308
rect 91276 36268 91316 36308
rect 91358 36268 91398 36308
rect 91440 36268 91480 36308
rect 95112 36268 95152 36308
rect 95194 36268 95234 36308
rect 95276 36268 95316 36308
rect 95358 36268 95398 36308
rect 95440 36268 95480 36308
rect 99112 36268 99152 36308
rect 99194 36268 99234 36308
rect 99276 36268 99316 36308
rect 99358 36268 99398 36308
rect 99440 36268 99480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 8352 35512 8392 35552
rect 8434 35512 8474 35552
rect 8516 35512 8556 35552
rect 8598 35512 8638 35552
rect 8680 35512 8720 35552
rect 12352 35512 12392 35552
rect 12434 35512 12474 35552
rect 12516 35512 12556 35552
rect 12598 35512 12638 35552
rect 12680 35512 12720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 20352 35512 20392 35552
rect 20434 35512 20474 35552
rect 20516 35512 20556 35552
rect 20598 35512 20638 35552
rect 20680 35512 20720 35552
rect 24352 35512 24392 35552
rect 24434 35512 24474 35552
rect 24516 35512 24556 35552
rect 24598 35512 24638 35552
rect 24680 35512 24720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 32352 35512 32392 35552
rect 32434 35512 32474 35552
rect 32516 35512 32556 35552
rect 32598 35512 32638 35552
rect 32680 35512 32720 35552
rect 36352 35512 36392 35552
rect 36434 35512 36474 35552
rect 36516 35512 36556 35552
rect 36598 35512 36638 35552
rect 36680 35512 36720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 44352 35512 44392 35552
rect 44434 35512 44474 35552
rect 44516 35512 44556 35552
rect 44598 35512 44638 35552
rect 44680 35512 44720 35552
rect 48352 35512 48392 35552
rect 48434 35512 48474 35552
rect 48516 35512 48556 35552
rect 48598 35512 48638 35552
rect 48680 35512 48720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 56352 35512 56392 35552
rect 56434 35512 56474 35552
rect 56516 35512 56556 35552
rect 56598 35512 56638 35552
rect 56680 35512 56720 35552
rect 60352 35512 60392 35552
rect 60434 35512 60474 35552
rect 60516 35512 60556 35552
rect 60598 35512 60638 35552
rect 60680 35512 60720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 68352 35512 68392 35552
rect 68434 35512 68474 35552
rect 68516 35512 68556 35552
rect 68598 35512 68638 35552
rect 68680 35512 68720 35552
rect 72352 35512 72392 35552
rect 72434 35512 72474 35552
rect 72516 35512 72556 35552
rect 72598 35512 72638 35552
rect 72680 35512 72720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 80352 35512 80392 35552
rect 80434 35512 80474 35552
rect 80516 35512 80556 35552
rect 80598 35512 80638 35552
rect 80680 35512 80720 35552
rect 84352 35512 84392 35552
rect 84434 35512 84474 35552
rect 84516 35512 84556 35552
rect 84598 35512 84638 35552
rect 84680 35512 84720 35552
rect 88352 35512 88392 35552
rect 88434 35512 88474 35552
rect 88516 35512 88556 35552
rect 88598 35512 88638 35552
rect 88680 35512 88720 35552
rect 92352 35512 92392 35552
rect 92434 35512 92474 35552
rect 92516 35512 92556 35552
rect 92598 35512 92638 35552
rect 92680 35512 92720 35552
rect 96352 35512 96392 35552
rect 96434 35512 96474 35552
rect 96516 35512 96556 35552
rect 96598 35512 96638 35552
rect 96680 35512 96720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 7112 34756 7152 34796
rect 7194 34756 7234 34796
rect 7276 34756 7316 34796
rect 7358 34756 7398 34796
rect 7440 34756 7480 34796
rect 11112 34756 11152 34796
rect 11194 34756 11234 34796
rect 11276 34756 11316 34796
rect 11358 34756 11398 34796
rect 11440 34756 11480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 19112 34756 19152 34796
rect 19194 34756 19234 34796
rect 19276 34756 19316 34796
rect 19358 34756 19398 34796
rect 19440 34756 19480 34796
rect 23112 34756 23152 34796
rect 23194 34756 23234 34796
rect 23276 34756 23316 34796
rect 23358 34756 23398 34796
rect 23440 34756 23480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 31112 34756 31152 34796
rect 31194 34756 31234 34796
rect 31276 34756 31316 34796
rect 31358 34756 31398 34796
rect 31440 34756 31480 34796
rect 35112 34756 35152 34796
rect 35194 34756 35234 34796
rect 35276 34756 35316 34796
rect 35358 34756 35398 34796
rect 35440 34756 35480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 43112 34756 43152 34796
rect 43194 34756 43234 34796
rect 43276 34756 43316 34796
rect 43358 34756 43398 34796
rect 43440 34756 43480 34796
rect 47112 34756 47152 34796
rect 47194 34756 47234 34796
rect 47276 34756 47316 34796
rect 47358 34756 47398 34796
rect 47440 34756 47480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 55112 34756 55152 34796
rect 55194 34756 55234 34796
rect 55276 34756 55316 34796
rect 55358 34756 55398 34796
rect 55440 34756 55480 34796
rect 59112 34756 59152 34796
rect 59194 34756 59234 34796
rect 59276 34756 59316 34796
rect 59358 34756 59398 34796
rect 59440 34756 59480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 67112 34756 67152 34796
rect 67194 34756 67234 34796
rect 67276 34756 67316 34796
rect 67358 34756 67398 34796
rect 67440 34756 67480 34796
rect 71112 34756 71152 34796
rect 71194 34756 71234 34796
rect 71276 34756 71316 34796
rect 71358 34756 71398 34796
rect 71440 34756 71480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 79112 34756 79152 34796
rect 79194 34756 79234 34796
rect 79276 34756 79316 34796
rect 79358 34756 79398 34796
rect 79440 34756 79480 34796
rect 83112 34756 83152 34796
rect 83194 34756 83234 34796
rect 83276 34756 83316 34796
rect 83358 34756 83398 34796
rect 83440 34756 83480 34796
rect 87112 34756 87152 34796
rect 87194 34756 87234 34796
rect 87276 34756 87316 34796
rect 87358 34756 87398 34796
rect 87440 34756 87480 34796
rect 91112 34756 91152 34796
rect 91194 34756 91234 34796
rect 91276 34756 91316 34796
rect 91358 34756 91398 34796
rect 91440 34756 91480 34796
rect 95112 34756 95152 34796
rect 95194 34756 95234 34796
rect 95276 34756 95316 34796
rect 95358 34756 95398 34796
rect 95440 34756 95480 34796
rect 99112 34756 99152 34796
rect 99194 34756 99234 34796
rect 99276 34756 99316 34796
rect 99358 34756 99398 34796
rect 99440 34756 99480 34796
rect 91468 34420 91508 34460
rect 93388 34420 93428 34460
rect 91660 34168 91700 34208
rect 93580 34168 93620 34208
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 8352 34000 8392 34040
rect 8434 34000 8474 34040
rect 8516 34000 8556 34040
rect 8598 34000 8638 34040
rect 8680 34000 8720 34040
rect 12352 34000 12392 34040
rect 12434 34000 12474 34040
rect 12516 34000 12556 34040
rect 12598 34000 12638 34040
rect 12680 34000 12720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 20352 34000 20392 34040
rect 20434 34000 20474 34040
rect 20516 34000 20556 34040
rect 20598 34000 20638 34040
rect 20680 34000 20720 34040
rect 24352 34000 24392 34040
rect 24434 34000 24474 34040
rect 24516 34000 24556 34040
rect 24598 34000 24638 34040
rect 24680 34000 24720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 32352 34000 32392 34040
rect 32434 34000 32474 34040
rect 32516 34000 32556 34040
rect 32598 34000 32638 34040
rect 32680 34000 32720 34040
rect 36352 34000 36392 34040
rect 36434 34000 36474 34040
rect 36516 34000 36556 34040
rect 36598 34000 36638 34040
rect 36680 34000 36720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 44352 34000 44392 34040
rect 44434 34000 44474 34040
rect 44516 34000 44556 34040
rect 44598 34000 44638 34040
rect 44680 34000 44720 34040
rect 48352 34000 48392 34040
rect 48434 34000 48474 34040
rect 48516 34000 48556 34040
rect 48598 34000 48638 34040
rect 48680 34000 48720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 56352 34000 56392 34040
rect 56434 34000 56474 34040
rect 56516 34000 56556 34040
rect 56598 34000 56638 34040
rect 56680 34000 56720 34040
rect 60352 34000 60392 34040
rect 60434 34000 60474 34040
rect 60516 34000 60556 34040
rect 60598 34000 60638 34040
rect 60680 34000 60720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 68352 34000 68392 34040
rect 68434 34000 68474 34040
rect 68516 34000 68556 34040
rect 68598 34000 68638 34040
rect 68680 34000 68720 34040
rect 95500 33832 95540 33872
rect 73228 33580 73268 33620
rect 73612 33580 73652 33620
rect 74092 33580 74132 33620
rect 74476 33580 74516 33620
rect 74860 33580 74900 33620
rect 75340 33580 75380 33620
rect 75820 33580 75860 33620
rect 76204 33580 76244 33620
rect 76588 33580 76628 33620
rect 76972 33580 77012 33620
rect 77452 33580 77492 33620
rect 77836 33580 77876 33620
rect 78220 33580 78260 33620
rect 78604 33580 78644 33620
rect 78988 33580 79028 33620
rect 79372 33580 79412 33620
rect 79756 33580 79796 33620
rect 80332 33580 80372 33620
rect 80908 33580 80948 33620
rect 81100 33580 81140 33620
rect 81676 33580 81716 33620
rect 82060 33580 82100 33620
rect 82444 33580 82484 33620
rect 82828 33580 82868 33620
rect 83212 33580 83252 33620
rect 83596 33580 83636 33620
rect 83980 33580 84020 33620
rect 84364 33580 84404 33620
rect 84748 33580 84788 33620
rect 85132 33580 85172 33620
rect 85516 33580 85556 33620
rect 85900 33580 85940 33620
rect 86284 33580 86324 33620
rect 86668 33580 86708 33620
rect 87052 33580 87092 33620
rect 87436 33580 87476 33620
rect 87820 33580 87860 33620
rect 88204 33580 88244 33620
rect 88588 33580 88628 33620
rect 88972 33580 89012 33620
rect 89356 33580 89396 33620
rect 89740 33580 89780 33620
rect 90124 33580 90164 33620
rect 90508 33580 90548 33620
rect 90892 33580 90932 33620
rect 91276 33580 91316 33620
rect 91660 33580 91700 33620
rect 91852 33580 91892 33620
rect 92236 33580 92276 33620
rect 92620 33580 92660 33620
rect 93196 33580 93236 33620
rect 93580 33580 93620 33620
rect 94060 33580 94100 33620
rect 94252 33580 94292 33620
rect 94636 33580 94676 33620
rect 95308 33580 95348 33620
rect 95692 33580 95732 33620
rect 96076 33580 96116 33620
rect 96460 33580 96500 33620
rect 96844 33580 96884 33620
rect 97228 33580 97268 33620
rect 97612 33580 97652 33620
rect 97996 33580 98036 33620
rect 98380 33580 98420 33620
rect 80524 33496 80564 33536
rect 81292 33496 81332 33536
rect 82252 33496 82292 33536
rect 92812 33496 92852 33536
rect 73420 33412 73460 33452
rect 73804 33412 73844 33452
rect 74284 33412 74324 33452
rect 74668 33412 74708 33452
rect 75052 33412 75092 33452
rect 75532 33412 75572 33452
rect 76012 33412 76052 33452
rect 76396 33412 76436 33452
rect 76780 33412 76820 33452
rect 77164 33412 77204 33452
rect 77644 33412 77684 33452
rect 78028 33412 78068 33452
rect 78412 33412 78452 33452
rect 78796 33412 78836 33452
rect 79180 33412 79220 33452
rect 79564 33412 79604 33452
rect 79948 33412 79988 33452
rect 80716 33412 80756 33452
rect 81484 33412 81524 33452
rect 81868 33412 81908 33452
rect 82636 33412 82676 33452
rect 83020 33412 83060 33452
rect 83404 33412 83444 33452
rect 83788 33412 83828 33452
rect 84172 33412 84212 33452
rect 84556 33412 84596 33452
rect 84940 33412 84980 33452
rect 85324 33412 85364 33452
rect 85708 33412 85748 33452
rect 86092 33412 86132 33452
rect 86476 33412 86516 33452
rect 86860 33412 86900 33452
rect 87244 33412 87284 33452
rect 87628 33412 87668 33452
rect 88012 33412 88052 33452
rect 88396 33412 88436 33452
rect 88780 33412 88820 33452
rect 89164 33412 89204 33452
rect 89548 33412 89588 33452
rect 89932 33412 89972 33452
rect 90316 33412 90356 33452
rect 90700 33412 90740 33452
rect 91084 33412 91124 33452
rect 91468 33412 91508 33452
rect 92044 33412 92084 33452
rect 92428 33412 92468 33452
rect 93004 33412 93044 33452
rect 93388 33412 93428 33452
rect 93868 33412 93908 33452
rect 94444 33412 94484 33452
rect 94828 33412 94868 33452
rect 95116 33412 95156 33452
rect 95884 33412 95924 33452
rect 96268 33412 96308 33452
rect 96652 33412 96692 33452
rect 97036 33412 97076 33452
rect 97420 33412 97460 33452
rect 97804 33412 97844 33452
rect 98188 33412 98228 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 7112 33244 7152 33284
rect 7194 33244 7234 33284
rect 7276 33244 7316 33284
rect 7358 33244 7398 33284
rect 7440 33244 7480 33284
rect 11112 33244 11152 33284
rect 11194 33244 11234 33284
rect 11276 33244 11316 33284
rect 11358 33244 11398 33284
rect 11440 33244 11480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 19112 33244 19152 33284
rect 19194 33244 19234 33284
rect 19276 33244 19316 33284
rect 19358 33244 19398 33284
rect 19440 33244 19480 33284
rect 23112 33244 23152 33284
rect 23194 33244 23234 33284
rect 23276 33244 23316 33284
rect 23358 33244 23398 33284
rect 23440 33244 23480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 31112 33244 31152 33284
rect 31194 33244 31234 33284
rect 31276 33244 31316 33284
rect 31358 33244 31398 33284
rect 31440 33244 31480 33284
rect 35112 33244 35152 33284
rect 35194 33244 35234 33284
rect 35276 33244 35316 33284
rect 35358 33244 35398 33284
rect 35440 33244 35480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 43112 33244 43152 33284
rect 43194 33244 43234 33284
rect 43276 33244 43316 33284
rect 43358 33244 43398 33284
rect 43440 33244 43480 33284
rect 47112 33244 47152 33284
rect 47194 33244 47234 33284
rect 47276 33244 47316 33284
rect 47358 33244 47398 33284
rect 47440 33244 47480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 55112 33244 55152 33284
rect 55194 33244 55234 33284
rect 55276 33244 55316 33284
rect 55358 33244 55398 33284
rect 55440 33244 55480 33284
rect 59112 33244 59152 33284
rect 59194 33244 59234 33284
rect 59276 33244 59316 33284
rect 59358 33244 59398 33284
rect 59440 33244 59480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 67112 33244 67152 33284
rect 67194 33244 67234 33284
rect 67276 33244 67316 33284
rect 67358 33244 67398 33284
rect 67440 33244 67480 33284
rect 74188 33076 74228 33116
rect 77068 33076 77108 33116
rect 78892 33076 78932 33116
rect 86476 33076 86516 33116
rect 90892 33076 90932 33116
rect 92332 33076 92372 33116
rect 94060 33076 94100 33116
rect 74860 32992 74900 33032
rect 76012 32992 76052 33032
rect 83308 32992 83348 33032
rect 84844 32992 84884 33032
rect 88108 32992 88148 33032
rect 92716 32992 92756 33032
rect 94924 32992 94964 33032
rect 96940 32992 96980 33032
rect 72652 32908 72692 32948
rect 74380 32908 74420 32948
rect 74668 32908 74708 32948
rect 75820 32908 75860 32948
rect 77260 32908 77300 32948
rect 78700 32908 78740 32948
rect 79372 32908 79412 32948
rect 80620 32908 80660 32948
rect 82060 32908 82100 32948
rect 83116 32908 83156 32948
rect 83596 32908 83636 32948
rect 84652 32908 84692 32948
rect 86284 32908 86324 32948
rect 86956 32908 86996 32948
rect 87916 32908 87956 32948
rect 88396 32908 88436 32948
rect 88972 32908 89012 32948
rect 90028 32908 90068 32948
rect 90700 32919 90740 32959
rect 91084 32908 91124 32948
rect 92524 32908 92564 32948
rect 93100 32908 93140 32948
rect 93868 32908 93908 32948
rect 95116 32908 95156 32948
rect 96748 32908 96788 32948
rect 98668 32908 98708 32948
rect 71500 32824 71540 32864
rect 71596 32824 71636 32864
rect 72364 32824 72404 32864
rect 73036 32824 73076 32864
rect 73612 32824 73652 32864
rect 73996 32824 74036 32864
rect 75148 32824 75188 32864
rect 75436 32824 75476 32864
rect 76204 32824 76244 32864
rect 76300 32824 76340 32864
rect 76588 32824 76628 32864
rect 76876 32824 76916 32864
rect 77452 32824 77492 32864
rect 77548 32824 77588 32864
rect 77836 32824 77876 32864
rect 78124 32824 78164 32864
rect 78316 32824 78356 32864
rect 78412 32824 78452 32864
rect 79084 32824 79124 32864
rect 79468 32824 79508 32864
rect 79660 32824 79700 32864
rect 79756 32824 79796 32864
rect 80046 32837 80086 32877
rect 80236 32824 80276 32864
rect 81004 32824 81044 32864
rect 81100 32824 81140 32864
rect 81388 32824 81428 32864
rect 81676 32824 81716 32864
rect 82252 32824 82292 32864
rect 82348 32824 82388 32864
rect 82636 32824 82676 32864
rect 82924 32824 82964 32864
rect 83500 32824 83540 32864
rect 83788 32824 83828 32864
rect 83884 32824 83924 32864
rect 84172 32824 84212 32864
rect 84460 32824 84500 32864
rect 85036 32824 85076 32864
rect 85132 32824 85172 32864
rect 85420 32824 85460 32864
rect 85708 32824 85748 32864
rect 85996 32824 86036 32864
rect 86668 32824 86708 32864
rect 87052 32824 87092 32864
rect 87244 32824 87284 32864
rect 87340 32824 87380 32864
rect 87628 32824 87668 32864
rect 88300 32824 88340 32864
rect 88588 32824 88628 32864
rect 88684 32824 88724 32864
rect 89452 32824 89492 32864
rect 89644 32824 89684 32864
rect 89740 32824 89780 32864
rect 89932 32824 89972 32864
rect 90316 32824 90356 32864
rect 91180 32824 91220 32864
rect 91372 32824 91412 32864
rect 91468 32824 91508 32864
rect 91756 32837 91796 32877
rect 92044 32824 92084 32864
rect 92812 32824 92852 32864
rect 93004 32824 93044 32864
rect 93292 32824 93332 32864
rect 93388 32824 93428 32864
rect 93676 32824 93716 32864
rect 94252 32824 94292 32864
rect 94348 32824 94388 32864
rect 94636 32824 94676 32864
rect 94828 32824 94868 32864
rect 95212 32824 95252 32864
rect 95500 32824 95540 32864
rect 95692 32824 95732 32864
rect 95788 32824 95828 32864
rect 96076 32824 96116 32864
rect 96364 32824 96404 32864
rect 97228 32824 97268 32864
rect 97516 32824 97556 32864
rect 97804 32824 97844 32864
rect 98092 32824 98132 32864
rect 98860 32824 98900 32864
rect 99148 32824 99188 32864
rect 85900 32740 85940 32780
rect 93580 32740 93620 32780
rect 94540 32740 94580 32780
rect 95980 32740 96020 32780
rect 72460 32656 72500 32696
rect 72844 32656 72884 32696
rect 73132 32656 73172 32696
rect 73708 32656 73748 32696
rect 73900 32656 73940 32696
rect 75052 32656 75092 32696
rect 75340 32656 75380 32696
rect 76492 32656 76532 32696
rect 76780 32656 76820 32696
rect 77740 32656 77780 32696
rect 78028 32656 78068 32696
rect 79180 32656 79220 32696
rect 79948 32656 79988 32696
rect 80332 32656 80372 32696
rect 80812 32656 80852 32696
rect 81292 32656 81332 32696
rect 81580 32656 81620 32696
rect 81868 32656 81908 32696
rect 82540 32656 82580 32696
rect 82828 32656 82868 32696
rect 84076 32656 84116 32696
rect 84364 32656 84404 32696
rect 85324 32656 85364 32696
rect 85612 32656 85652 32696
rect 86764 32656 86804 32696
rect 87532 32656 87572 32696
rect 89164 32656 89204 32696
rect 89356 32656 89396 32696
rect 90220 32656 90260 32696
rect 91660 32656 91700 32696
rect 91948 32656 91988 32696
rect 95404 32656 95444 32696
rect 96268 32656 96308 32696
rect 97132 32656 97172 32696
rect 97420 32656 97460 32696
rect 97708 32656 97748 32696
rect 97996 32656 98036 32696
rect 98476 32656 98516 32696
rect 98956 32656 98996 32696
rect 99244 32656 99284 32696
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 8352 32488 8392 32528
rect 8434 32488 8474 32528
rect 8516 32488 8556 32528
rect 8598 32488 8638 32528
rect 8680 32488 8720 32528
rect 12352 32488 12392 32528
rect 12434 32488 12474 32528
rect 12516 32488 12556 32528
rect 12598 32488 12638 32528
rect 12680 32488 12720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 20352 32488 20392 32528
rect 20434 32488 20474 32528
rect 20516 32488 20556 32528
rect 20598 32488 20638 32528
rect 20680 32488 20720 32528
rect 24352 32488 24392 32528
rect 24434 32488 24474 32528
rect 24516 32488 24556 32528
rect 24598 32488 24638 32528
rect 24680 32488 24720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 32352 32488 32392 32528
rect 32434 32488 32474 32528
rect 32516 32488 32556 32528
rect 32598 32488 32638 32528
rect 32680 32488 32720 32528
rect 36352 32488 36392 32528
rect 36434 32488 36474 32528
rect 36516 32488 36556 32528
rect 36598 32488 36638 32528
rect 36680 32488 36720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 44352 32488 44392 32528
rect 44434 32488 44474 32528
rect 44516 32488 44556 32528
rect 44598 32488 44638 32528
rect 44680 32488 44720 32528
rect 48352 32488 48392 32528
rect 48434 32488 48474 32528
rect 48516 32488 48556 32528
rect 48598 32488 48638 32528
rect 48680 32488 48720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 56352 32488 56392 32528
rect 56434 32488 56474 32528
rect 56516 32488 56556 32528
rect 56598 32488 56638 32528
rect 56680 32488 56720 32528
rect 60352 32488 60392 32528
rect 60434 32488 60474 32528
rect 60516 32488 60556 32528
rect 60598 32488 60638 32528
rect 60680 32488 60720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 68352 32488 68392 32528
rect 68434 32488 68474 32528
rect 68516 32488 68556 32528
rect 68598 32488 68638 32528
rect 68680 32488 68720 32528
rect 70732 32320 70772 32360
rect 71404 32320 71444 32360
rect 70924 32068 70964 32108
rect 71212 32068 71252 32108
rect 70732 31900 70772 31940
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 7112 31732 7152 31772
rect 7194 31732 7234 31772
rect 7276 31732 7316 31772
rect 7358 31732 7398 31772
rect 7440 31732 7480 31772
rect 11112 31732 11152 31772
rect 11194 31732 11234 31772
rect 11276 31732 11316 31772
rect 11358 31732 11398 31772
rect 11440 31732 11480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 19112 31732 19152 31772
rect 19194 31732 19234 31772
rect 19276 31732 19316 31772
rect 19358 31732 19398 31772
rect 19440 31732 19480 31772
rect 23112 31732 23152 31772
rect 23194 31732 23234 31772
rect 23276 31732 23316 31772
rect 23358 31732 23398 31772
rect 23440 31732 23480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 31112 31732 31152 31772
rect 31194 31732 31234 31772
rect 31276 31732 31316 31772
rect 31358 31732 31398 31772
rect 31440 31732 31480 31772
rect 35112 31732 35152 31772
rect 35194 31732 35234 31772
rect 35276 31732 35316 31772
rect 35358 31732 35398 31772
rect 35440 31732 35480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 43112 31732 43152 31772
rect 43194 31732 43234 31772
rect 43276 31732 43316 31772
rect 43358 31732 43398 31772
rect 43440 31732 43480 31772
rect 47112 31732 47152 31772
rect 47194 31732 47234 31772
rect 47276 31732 47316 31772
rect 47358 31732 47398 31772
rect 47440 31732 47480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 55112 31732 55152 31772
rect 55194 31732 55234 31772
rect 55276 31732 55316 31772
rect 55358 31732 55398 31772
rect 55440 31732 55480 31772
rect 59112 31732 59152 31772
rect 59194 31732 59234 31772
rect 59276 31732 59316 31772
rect 59358 31732 59398 31772
rect 59440 31732 59480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 67112 31732 67152 31772
rect 67194 31732 67234 31772
rect 67276 31732 67316 31772
rect 67358 31732 67398 31772
rect 67440 31732 67480 31772
rect 70828 31564 70868 31604
rect 71116 31480 71156 31520
rect 70636 31396 70676 31436
rect 71020 31312 71060 31352
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 8352 30976 8392 31016
rect 8434 30976 8474 31016
rect 8516 30976 8556 31016
rect 8598 30976 8638 31016
rect 8680 30976 8720 31016
rect 12352 30976 12392 31016
rect 12434 30976 12474 31016
rect 12516 30976 12556 31016
rect 12598 30976 12638 31016
rect 12680 30976 12720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 20352 30976 20392 31016
rect 20434 30976 20474 31016
rect 20516 30976 20556 31016
rect 20598 30976 20638 31016
rect 20680 30976 20720 31016
rect 24352 30976 24392 31016
rect 24434 30976 24474 31016
rect 24516 30976 24556 31016
rect 24598 30976 24638 31016
rect 24680 30976 24720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 32352 30976 32392 31016
rect 32434 30976 32474 31016
rect 32516 30976 32556 31016
rect 32598 30976 32638 31016
rect 32680 30976 32720 31016
rect 36352 30976 36392 31016
rect 36434 30976 36474 31016
rect 36516 30976 36556 31016
rect 36598 30976 36638 31016
rect 36680 30976 36720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 44352 30976 44392 31016
rect 44434 30976 44474 31016
rect 44516 30976 44556 31016
rect 44598 30976 44638 31016
rect 44680 30976 44720 31016
rect 48352 30976 48392 31016
rect 48434 30976 48474 31016
rect 48516 30976 48556 31016
rect 48598 30976 48638 31016
rect 48680 30976 48720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 56352 30976 56392 31016
rect 56434 30976 56474 31016
rect 56516 30976 56556 31016
rect 56598 30976 56638 31016
rect 56680 30976 56720 31016
rect 60352 30976 60392 31016
rect 60434 30976 60474 31016
rect 60516 30976 60556 31016
rect 60598 30976 60638 31016
rect 60680 30976 60720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 68352 30976 68392 31016
rect 68434 30976 68474 31016
rect 68516 30976 68556 31016
rect 68598 30976 68638 31016
rect 68680 30976 68720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 7112 30220 7152 30260
rect 7194 30220 7234 30260
rect 7276 30220 7316 30260
rect 7358 30220 7398 30260
rect 7440 30220 7480 30260
rect 11112 30220 11152 30260
rect 11194 30220 11234 30260
rect 11276 30220 11316 30260
rect 11358 30220 11398 30260
rect 11440 30220 11480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 19112 30220 19152 30260
rect 19194 30220 19234 30260
rect 19276 30220 19316 30260
rect 19358 30220 19398 30260
rect 19440 30220 19480 30260
rect 23112 30220 23152 30260
rect 23194 30220 23234 30260
rect 23276 30220 23316 30260
rect 23358 30220 23398 30260
rect 23440 30220 23480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 31112 30220 31152 30260
rect 31194 30220 31234 30260
rect 31276 30220 31316 30260
rect 31358 30220 31398 30260
rect 31440 30220 31480 30260
rect 35112 30220 35152 30260
rect 35194 30220 35234 30260
rect 35276 30220 35316 30260
rect 35358 30220 35398 30260
rect 35440 30220 35480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 43112 30220 43152 30260
rect 43194 30220 43234 30260
rect 43276 30220 43316 30260
rect 43358 30220 43398 30260
rect 43440 30220 43480 30260
rect 47112 30220 47152 30260
rect 47194 30220 47234 30260
rect 47276 30220 47316 30260
rect 47358 30220 47398 30260
rect 47440 30220 47480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 55112 30220 55152 30260
rect 55194 30220 55234 30260
rect 55276 30220 55316 30260
rect 55358 30220 55398 30260
rect 55440 30220 55480 30260
rect 59112 30220 59152 30260
rect 59194 30220 59234 30260
rect 59276 30220 59316 30260
rect 59358 30220 59398 30260
rect 59440 30220 59480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 67112 30220 67152 30260
rect 67194 30220 67234 30260
rect 67276 30220 67316 30260
rect 67358 30220 67398 30260
rect 67440 30220 67480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 8352 29464 8392 29504
rect 8434 29464 8474 29504
rect 8516 29464 8556 29504
rect 8598 29464 8638 29504
rect 8680 29464 8720 29504
rect 12352 29464 12392 29504
rect 12434 29464 12474 29504
rect 12516 29464 12556 29504
rect 12598 29464 12638 29504
rect 12680 29464 12720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 20352 29464 20392 29504
rect 20434 29464 20474 29504
rect 20516 29464 20556 29504
rect 20598 29464 20638 29504
rect 20680 29464 20720 29504
rect 24352 29464 24392 29504
rect 24434 29464 24474 29504
rect 24516 29464 24556 29504
rect 24598 29464 24638 29504
rect 24680 29464 24720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 32352 29464 32392 29504
rect 32434 29464 32474 29504
rect 32516 29464 32556 29504
rect 32598 29464 32638 29504
rect 32680 29464 32720 29504
rect 36352 29464 36392 29504
rect 36434 29464 36474 29504
rect 36516 29464 36556 29504
rect 36598 29464 36638 29504
rect 36680 29464 36720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 44352 29464 44392 29504
rect 44434 29464 44474 29504
rect 44516 29464 44556 29504
rect 44598 29464 44638 29504
rect 44680 29464 44720 29504
rect 48352 29464 48392 29504
rect 48434 29464 48474 29504
rect 48516 29464 48556 29504
rect 48598 29464 48638 29504
rect 48680 29464 48720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 56352 29464 56392 29504
rect 56434 29464 56474 29504
rect 56516 29464 56556 29504
rect 56598 29464 56638 29504
rect 56680 29464 56720 29504
rect 60352 29464 60392 29504
rect 60434 29464 60474 29504
rect 60516 29464 60556 29504
rect 60598 29464 60638 29504
rect 60680 29464 60720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 68352 29464 68392 29504
rect 68434 29464 68474 29504
rect 68516 29464 68556 29504
rect 68598 29464 68638 29504
rect 68680 29464 68720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 7112 28708 7152 28748
rect 7194 28708 7234 28748
rect 7276 28708 7316 28748
rect 7358 28708 7398 28748
rect 7440 28708 7480 28748
rect 11112 28708 11152 28748
rect 11194 28708 11234 28748
rect 11276 28708 11316 28748
rect 11358 28708 11398 28748
rect 11440 28708 11480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 19112 28708 19152 28748
rect 19194 28708 19234 28748
rect 19276 28708 19316 28748
rect 19358 28708 19398 28748
rect 19440 28708 19480 28748
rect 23112 28708 23152 28748
rect 23194 28708 23234 28748
rect 23276 28708 23316 28748
rect 23358 28708 23398 28748
rect 23440 28708 23480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 31112 28708 31152 28748
rect 31194 28708 31234 28748
rect 31276 28708 31316 28748
rect 31358 28708 31398 28748
rect 31440 28708 31480 28748
rect 35112 28708 35152 28748
rect 35194 28708 35234 28748
rect 35276 28708 35316 28748
rect 35358 28708 35398 28748
rect 35440 28708 35480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 43112 28708 43152 28748
rect 43194 28708 43234 28748
rect 43276 28708 43316 28748
rect 43358 28708 43398 28748
rect 43440 28708 43480 28748
rect 47112 28708 47152 28748
rect 47194 28708 47234 28748
rect 47276 28708 47316 28748
rect 47358 28708 47398 28748
rect 47440 28708 47480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 55112 28708 55152 28748
rect 55194 28708 55234 28748
rect 55276 28708 55316 28748
rect 55358 28708 55398 28748
rect 55440 28708 55480 28748
rect 59112 28708 59152 28748
rect 59194 28708 59234 28748
rect 59276 28708 59316 28748
rect 59358 28708 59398 28748
rect 59440 28708 59480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 67112 28708 67152 28748
rect 67194 28708 67234 28748
rect 67276 28708 67316 28748
rect 67358 28708 67398 28748
rect 67440 28708 67480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 8352 27952 8392 27992
rect 8434 27952 8474 27992
rect 8516 27952 8556 27992
rect 8598 27952 8638 27992
rect 8680 27952 8720 27992
rect 12352 27952 12392 27992
rect 12434 27952 12474 27992
rect 12516 27952 12556 27992
rect 12598 27952 12638 27992
rect 12680 27952 12720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 20352 27952 20392 27992
rect 20434 27952 20474 27992
rect 20516 27952 20556 27992
rect 20598 27952 20638 27992
rect 20680 27952 20720 27992
rect 24352 27952 24392 27992
rect 24434 27952 24474 27992
rect 24516 27952 24556 27992
rect 24598 27952 24638 27992
rect 24680 27952 24720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 32352 27952 32392 27992
rect 32434 27952 32474 27992
rect 32516 27952 32556 27992
rect 32598 27952 32638 27992
rect 32680 27952 32720 27992
rect 36352 27952 36392 27992
rect 36434 27952 36474 27992
rect 36516 27952 36556 27992
rect 36598 27952 36638 27992
rect 36680 27952 36720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 44352 27952 44392 27992
rect 44434 27952 44474 27992
rect 44516 27952 44556 27992
rect 44598 27952 44638 27992
rect 44680 27952 44720 27992
rect 48352 27952 48392 27992
rect 48434 27952 48474 27992
rect 48516 27952 48556 27992
rect 48598 27952 48638 27992
rect 48680 27952 48720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 56352 27952 56392 27992
rect 56434 27952 56474 27992
rect 56516 27952 56556 27992
rect 56598 27952 56638 27992
rect 56680 27952 56720 27992
rect 60352 27952 60392 27992
rect 60434 27952 60474 27992
rect 60516 27952 60556 27992
rect 60598 27952 60638 27992
rect 60680 27952 60720 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 68352 27952 68392 27992
rect 68434 27952 68474 27992
rect 68516 27952 68556 27992
rect 68598 27952 68638 27992
rect 68680 27952 68720 27992
rect 69964 27616 70004 27656
rect 70156 27616 70196 27656
rect 70924 27616 70964 27656
rect 70540 27532 70580 27572
rect 71212 27532 71252 27572
rect 70348 27448 70388 27488
rect 71020 27364 71060 27404
rect 71404 27364 71444 27404
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 7112 27196 7152 27236
rect 7194 27196 7234 27236
rect 7276 27196 7316 27236
rect 7358 27196 7398 27236
rect 7440 27196 7480 27236
rect 11112 27196 11152 27236
rect 11194 27196 11234 27236
rect 11276 27196 11316 27236
rect 11358 27196 11398 27236
rect 11440 27196 11480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 19112 27196 19152 27236
rect 19194 27196 19234 27236
rect 19276 27196 19316 27236
rect 19358 27196 19398 27236
rect 19440 27196 19480 27236
rect 23112 27196 23152 27236
rect 23194 27196 23234 27236
rect 23276 27196 23316 27236
rect 23358 27196 23398 27236
rect 23440 27196 23480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 31112 27196 31152 27236
rect 31194 27196 31234 27236
rect 31276 27196 31316 27236
rect 31358 27196 31398 27236
rect 31440 27196 31480 27236
rect 35112 27196 35152 27236
rect 35194 27196 35234 27236
rect 35276 27196 35316 27236
rect 35358 27196 35398 27236
rect 35440 27196 35480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 43112 27196 43152 27236
rect 43194 27196 43234 27236
rect 43276 27196 43316 27236
rect 43358 27196 43398 27236
rect 43440 27196 43480 27236
rect 47112 27196 47152 27236
rect 47194 27196 47234 27236
rect 47276 27196 47316 27236
rect 47358 27196 47398 27236
rect 47440 27196 47480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 55112 27196 55152 27236
rect 55194 27196 55234 27236
rect 55276 27196 55316 27236
rect 55358 27196 55398 27236
rect 55440 27196 55480 27236
rect 59112 27196 59152 27236
rect 59194 27196 59234 27236
rect 59276 27196 59316 27236
rect 59358 27196 59398 27236
rect 59440 27196 59480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 67112 27196 67152 27236
rect 67194 27196 67234 27236
rect 67276 27196 67316 27236
rect 67358 27196 67398 27236
rect 67440 27196 67480 27236
rect 69772 26860 69812 26900
rect 70348 26860 70388 26900
rect 70732 26860 70772 26900
rect 71116 26860 71156 26900
rect 69964 26608 70004 26648
rect 70540 26608 70580 26648
rect 70924 26608 70964 26648
rect 71308 26608 71348 26648
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 8352 26440 8392 26480
rect 8434 26440 8474 26480
rect 8516 26440 8556 26480
rect 8598 26440 8638 26480
rect 8680 26440 8720 26480
rect 12352 26440 12392 26480
rect 12434 26440 12474 26480
rect 12516 26440 12556 26480
rect 12598 26440 12638 26480
rect 12680 26440 12720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 20352 26440 20392 26480
rect 20434 26440 20474 26480
rect 20516 26440 20556 26480
rect 20598 26440 20638 26480
rect 20680 26440 20720 26480
rect 24352 26440 24392 26480
rect 24434 26440 24474 26480
rect 24516 26440 24556 26480
rect 24598 26440 24638 26480
rect 24680 26440 24720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 32352 26440 32392 26480
rect 32434 26440 32474 26480
rect 32516 26440 32556 26480
rect 32598 26440 32638 26480
rect 32680 26440 32720 26480
rect 36352 26440 36392 26480
rect 36434 26440 36474 26480
rect 36516 26440 36556 26480
rect 36598 26440 36638 26480
rect 36680 26440 36720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 44352 26440 44392 26480
rect 44434 26440 44474 26480
rect 44516 26440 44556 26480
rect 44598 26440 44638 26480
rect 44680 26440 44720 26480
rect 48352 26440 48392 26480
rect 48434 26440 48474 26480
rect 48516 26440 48556 26480
rect 48598 26440 48638 26480
rect 48680 26440 48720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 56352 26440 56392 26480
rect 56434 26440 56474 26480
rect 56516 26440 56556 26480
rect 56598 26440 56638 26480
rect 56680 26440 56720 26480
rect 60352 26440 60392 26480
rect 60434 26440 60474 26480
rect 60516 26440 60556 26480
rect 60598 26440 60638 26480
rect 60680 26440 60720 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 68352 26440 68392 26480
rect 68434 26440 68474 26480
rect 68516 26440 68556 26480
rect 68598 26440 68638 26480
rect 68680 26440 68720 26480
rect 71020 26272 71060 26312
rect 71404 26272 71444 26312
rect 70924 26104 70964 26144
rect 71308 26104 71348 26144
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 7112 25684 7152 25724
rect 7194 25684 7234 25724
rect 7276 25684 7316 25724
rect 7358 25684 7398 25724
rect 7440 25684 7480 25724
rect 11112 25684 11152 25724
rect 11194 25684 11234 25724
rect 11276 25684 11316 25724
rect 11358 25684 11398 25724
rect 11440 25684 11480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 19112 25684 19152 25724
rect 19194 25684 19234 25724
rect 19276 25684 19316 25724
rect 19358 25684 19398 25724
rect 19440 25684 19480 25724
rect 23112 25684 23152 25724
rect 23194 25684 23234 25724
rect 23276 25684 23316 25724
rect 23358 25684 23398 25724
rect 23440 25684 23480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 31112 25684 31152 25724
rect 31194 25684 31234 25724
rect 31276 25684 31316 25724
rect 31358 25684 31398 25724
rect 31440 25684 31480 25724
rect 35112 25684 35152 25724
rect 35194 25684 35234 25724
rect 35276 25684 35316 25724
rect 35358 25684 35398 25724
rect 35440 25684 35480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 43112 25684 43152 25724
rect 43194 25684 43234 25724
rect 43276 25684 43316 25724
rect 43358 25684 43398 25724
rect 43440 25684 43480 25724
rect 47112 25684 47152 25724
rect 47194 25684 47234 25724
rect 47276 25684 47316 25724
rect 47358 25684 47398 25724
rect 47440 25684 47480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 55112 25684 55152 25724
rect 55194 25684 55234 25724
rect 55276 25684 55316 25724
rect 55358 25684 55398 25724
rect 55440 25684 55480 25724
rect 59112 25684 59152 25724
rect 59194 25684 59234 25724
rect 59276 25684 59316 25724
rect 59358 25684 59398 25724
rect 59440 25684 59480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 67112 25684 67152 25724
rect 67194 25684 67234 25724
rect 67276 25684 67316 25724
rect 67358 25684 67398 25724
rect 67440 25684 67480 25724
rect 72748 25516 72788 25556
rect 73132 25516 73172 25556
rect 73516 25516 73556 25556
rect 74092 25516 74132 25556
rect 75724 25516 75764 25556
rect 75916 25516 75956 25556
rect 76204 25516 76244 25556
rect 76876 25516 76916 25556
rect 77164 25516 77204 25556
rect 77932 25516 77972 25556
rect 78220 25516 78260 25556
rect 78508 25516 78548 25556
rect 78796 25516 78836 25556
rect 79180 25516 79220 25556
rect 79564 25516 79604 25556
rect 79756 25516 79796 25556
rect 80140 25516 80180 25556
rect 80332 25516 80372 25556
rect 80812 25516 80852 25556
rect 81196 25516 81236 25556
rect 81580 25516 81620 25556
rect 82060 25516 82100 25556
rect 82348 25516 82388 25556
rect 82732 25516 82772 25556
rect 83116 25516 83156 25556
rect 83980 25516 84020 25556
rect 84268 25516 84308 25556
rect 84556 25516 84596 25556
rect 84844 25516 84884 25556
rect 85228 25516 85268 25556
rect 85612 25516 85652 25556
rect 85996 25516 86036 25556
rect 86380 25516 86420 25556
rect 87532 25516 87572 25556
rect 87820 25516 87860 25556
rect 88108 25516 88148 25556
rect 88396 25516 88436 25556
rect 88780 25516 88820 25556
rect 89164 25516 89204 25556
rect 89932 25516 89972 25556
rect 90220 25516 90260 25556
rect 90508 25516 90548 25556
rect 90796 25516 90836 25556
rect 91180 25516 91220 25556
rect 91564 25516 91604 25556
rect 92044 25516 92084 25556
rect 92812 25516 92852 25556
rect 93196 25516 93236 25556
rect 93580 25516 93620 25556
rect 94060 25516 94100 25556
rect 94348 25516 94388 25556
rect 94828 25516 94868 25556
rect 95212 25516 95252 25556
rect 96076 25516 96116 25556
rect 96364 25516 96404 25556
rect 96844 25516 96884 25556
rect 97228 25516 97268 25556
rect 97420 25516 97460 25556
rect 97708 25516 97748 25556
rect 98092 25516 98132 25556
rect 98380 25516 98420 25556
rect 98764 25516 98804 25556
rect 74668 25432 74708 25472
rect 75244 25432 75284 25472
rect 76492 25432 76532 25472
rect 77740 25432 77780 25472
rect 83788 25432 83828 25472
rect 87340 25432 87380 25472
rect 89740 25432 89780 25472
rect 72940 25348 72980 25388
rect 73324 25348 73364 25388
rect 73900 25348 73940 25388
rect 74476 25348 74516 25388
rect 74860 25348 74900 25388
rect 75052 25348 75092 25388
rect 75532 25348 75572 25388
rect 77548 25348 77588 25388
rect 83596 25348 83636 25388
rect 87148 25348 87188 25388
rect 89548 25348 89588 25388
rect 95692 25348 95732 25388
rect 98572 25348 98612 25388
rect 652 25264 692 25304
rect 844 25264 884 25304
rect 72652 25264 72692 25304
rect 76012 25264 76052 25304
rect 76300 25264 76340 25304
rect 76588 25264 76628 25304
rect 76780 25264 76820 25304
rect 77068 25264 77108 25304
rect 78028 25264 78068 25304
rect 78316 25264 78356 25304
rect 78604 25264 78644 25304
rect 78892 25264 78932 25304
rect 79071 25253 79111 25293
rect 79468 25253 79508 25293
rect 79852 25264 79892 25304
rect 80044 25264 80084 25304
rect 80428 25264 80468 25304
rect 80716 25253 80756 25293
rect 81100 25253 81140 25293
rect 81484 25264 81524 25304
rect 81964 25264 82004 25304
rect 82252 25253 82292 25293
rect 82636 25264 82676 25304
rect 83212 25264 83252 25304
rect 84076 25264 84116 25304
rect 84364 25264 84404 25304
rect 84652 25264 84692 25304
rect 84940 25264 84980 25304
rect 85132 25264 85172 25304
rect 85516 25264 85556 25304
rect 85900 25264 85940 25304
rect 86476 25264 86516 25304
rect 86764 25264 86804 25304
rect 86956 25264 86996 25304
rect 87628 25264 87668 25304
rect 87916 25264 87956 25304
rect 88204 25264 88244 25304
rect 88492 25264 88532 25304
rect 88684 25264 88724 25304
rect 89068 25264 89108 25304
rect 90028 25264 90068 25304
rect 90316 25264 90356 25304
rect 90604 25264 90644 25304
rect 90892 25264 90932 25304
rect 91276 25264 91316 25304
rect 91455 25253 91495 25293
rect 91948 25264 91988 25304
rect 92332 25264 92372 25304
rect 92524 25264 92564 25304
rect 92908 25264 92948 25304
rect 93087 25253 93127 25293
rect 93676 25264 93716 25304
rect 93964 25264 94004 25304
rect 94252 25253 94292 25293
rect 94924 25264 94964 25304
rect 95308 25264 95348 25304
rect 96172 25264 96212 25304
rect 96460 25264 96500 25304
rect 96748 25264 96788 25304
rect 97127 25253 97167 25293
rect 97516 25264 97556 25304
rect 97804 25264 97844 25304
rect 97996 25264 98036 25304
rect 98860 25264 98900 25304
rect 74284 25096 74324 25136
rect 95884 25096 95924 25136
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 8352 24928 8392 24968
rect 8434 24928 8474 24968
rect 8516 24928 8556 24968
rect 8598 24928 8638 24968
rect 8680 24928 8720 24968
rect 12352 24928 12392 24968
rect 12434 24928 12474 24968
rect 12516 24928 12556 24968
rect 12598 24928 12638 24968
rect 12680 24928 12720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 20352 24928 20392 24968
rect 20434 24928 20474 24968
rect 20516 24928 20556 24968
rect 20598 24928 20638 24968
rect 20680 24928 20720 24968
rect 24352 24928 24392 24968
rect 24434 24928 24474 24968
rect 24516 24928 24556 24968
rect 24598 24928 24638 24968
rect 24680 24928 24720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 32352 24928 32392 24968
rect 32434 24928 32474 24968
rect 32516 24928 32556 24968
rect 32598 24928 32638 24968
rect 32680 24928 32720 24968
rect 36352 24928 36392 24968
rect 36434 24928 36474 24968
rect 36516 24928 36556 24968
rect 36598 24928 36638 24968
rect 36680 24928 36720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 44352 24928 44392 24968
rect 44434 24928 44474 24968
rect 44516 24928 44556 24968
rect 44598 24928 44638 24968
rect 44680 24928 44720 24968
rect 48352 24928 48392 24968
rect 48434 24928 48474 24968
rect 48516 24928 48556 24968
rect 48598 24928 48638 24968
rect 48680 24928 48720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 56352 24928 56392 24968
rect 56434 24928 56474 24968
rect 56516 24928 56556 24968
rect 56598 24928 56638 24968
rect 56680 24928 56720 24968
rect 60352 24928 60392 24968
rect 60434 24928 60474 24968
rect 60516 24928 60556 24968
rect 60598 24928 60638 24968
rect 60680 24928 60720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 68352 24928 68392 24968
rect 68434 24928 68474 24968
rect 68516 24928 68556 24968
rect 68598 24928 68638 24968
rect 68680 24928 68720 24968
rect 73324 24760 73364 24800
rect 73516 24760 73556 24800
rect 73996 24760 74036 24800
rect 74860 24760 74900 24800
rect 75436 24760 75476 24800
rect 75628 24760 75668 24800
rect 76204 24760 76244 24800
rect 76588 24760 76628 24800
rect 77068 24760 77108 24800
rect 77452 24760 77492 24800
rect 78028 24760 78068 24800
rect 78412 24760 78452 24800
rect 78796 24760 78836 24800
rect 79180 24760 79220 24800
rect 79564 24760 79604 24800
rect 79948 24760 79988 24800
rect 81196 24760 81236 24800
rect 81580 24760 81620 24800
rect 81964 24760 82004 24800
rect 82348 24760 82388 24800
rect 83116 24760 83156 24800
rect 83500 24760 83540 24800
rect 83884 24760 83924 24800
rect 84460 24760 84500 24800
rect 84844 24760 84884 24800
rect 85516 24760 85556 24800
rect 86284 24760 86324 24800
rect 87148 24760 87188 24800
rect 87532 24760 87572 24800
rect 88300 24760 88340 24800
rect 88684 24760 88724 24800
rect 89452 24760 89492 24800
rect 89932 24760 89972 24800
rect 90316 24760 90356 24800
rect 90700 24760 90740 24800
rect 91180 24760 91220 24800
rect 91852 24760 91892 24800
rect 92140 24760 92180 24800
rect 92908 24760 92948 24800
rect 93292 24760 93332 24800
rect 93964 24760 94004 24800
rect 94348 24760 94388 24800
rect 94732 24760 94772 24800
rect 95116 24760 95156 24800
rect 95596 24760 95636 24800
rect 95980 24760 96020 24800
rect 96172 24760 96212 24800
rect 96556 24760 96596 24800
rect 96940 24760 96980 24800
rect 97324 24760 97364 24800
rect 97708 24760 97748 24800
rect 98092 24760 98132 24800
rect 652 24592 692 24632
rect 844 24592 884 24632
rect 73228 24592 73268 24632
rect 73612 24592 73652 24632
rect 75724 24592 75764 24632
rect 80428 24592 80468 24632
rect 80620 24592 80660 24632
rect 87724 24592 87764 24632
rect 87820 24592 87860 24632
rect 73804 24508 73844 24548
rect 74188 24508 74228 24548
rect 74668 24508 74708 24548
rect 75244 24508 75284 24548
rect 76012 24508 76052 24548
rect 76396 24508 76436 24548
rect 76876 24508 76916 24548
rect 77260 24508 77300 24548
rect 77644 24508 77684 24548
rect 78220 24508 78260 24548
rect 78604 24508 78644 24548
rect 78988 24508 79028 24548
rect 79372 24508 79412 24548
rect 79756 24508 79796 24548
rect 80140 24508 80180 24548
rect 81004 24508 81044 24548
rect 81388 24508 81428 24548
rect 81772 24508 81812 24548
rect 82156 24508 82196 24548
rect 82540 24508 82580 24548
rect 82924 24508 82964 24548
rect 83308 24508 83348 24548
rect 83692 24508 83732 24548
rect 84076 24508 84116 24548
rect 84652 24508 84692 24548
rect 85036 24508 85076 24548
rect 85324 24508 85364 24548
rect 86092 24508 86132 24548
rect 86572 24508 86612 24548
rect 86956 24508 86996 24548
rect 87340 24508 87380 24548
rect 88108 24508 88148 24548
rect 88492 24508 88532 24548
rect 88876 24508 88916 24548
rect 89260 24508 89300 24548
rect 89740 24508 89780 24548
rect 90124 24508 90164 24548
rect 90508 24508 90548 24548
rect 90988 24508 91028 24548
rect 91660 24508 91700 24548
rect 92332 24508 92372 24548
rect 92716 24508 92756 24548
rect 93100 24508 93140 24548
rect 93484 24508 93524 24548
rect 93772 24508 93812 24548
rect 94156 24508 94196 24548
rect 94540 24508 94580 24548
rect 94924 24508 94964 24548
rect 95404 24508 95444 24548
rect 95788 24508 95828 24548
rect 96364 24508 96404 24548
rect 96748 24508 96788 24548
rect 97132 24508 97172 24548
rect 97516 24508 97556 24548
rect 97900 24508 97940 24548
rect 98284 24508 98324 24548
rect 77836 24424 77876 24464
rect 84268 24424 84308 24464
rect 86764 24424 86804 24464
rect 89068 24424 89108 24464
rect 92524 24424 92564 24464
rect 74380 24340 74420 24380
rect 80812 24340 80852 24380
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 7112 24172 7152 24212
rect 7194 24172 7234 24212
rect 7276 24172 7316 24212
rect 7358 24172 7398 24212
rect 7440 24172 7480 24212
rect 11112 24172 11152 24212
rect 11194 24172 11234 24212
rect 11276 24172 11316 24212
rect 11358 24172 11398 24212
rect 11440 24172 11480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 19112 24172 19152 24212
rect 19194 24172 19234 24212
rect 19276 24172 19316 24212
rect 19358 24172 19398 24212
rect 19440 24172 19480 24212
rect 23112 24172 23152 24212
rect 23194 24172 23234 24212
rect 23276 24172 23316 24212
rect 23358 24172 23398 24212
rect 23440 24172 23480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 31112 24172 31152 24212
rect 31194 24172 31234 24212
rect 31276 24172 31316 24212
rect 31358 24172 31398 24212
rect 31440 24172 31480 24212
rect 35112 24172 35152 24212
rect 35194 24172 35234 24212
rect 35276 24172 35316 24212
rect 35358 24172 35398 24212
rect 35440 24172 35480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 43112 24172 43152 24212
rect 43194 24172 43234 24212
rect 43276 24172 43316 24212
rect 43358 24172 43398 24212
rect 43440 24172 43480 24212
rect 47112 24172 47152 24212
rect 47194 24172 47234 24212
rect 47276 24172 47316 24212
rect 47358 24172 47398 24212
rect 47440 24172 47480 24212
rect 51112 24172 51152 24212
rect 51194 24172 51234 24212
rect 51276 24172 51316 24212
rect 51358 24172 51398 24212
rect 51440 24172 51480 24212
rect 55112 24172 55152 24212
rect 55194 24172 55234 24212
rect 55276 24172 55316 24212
rect 55358 24172 55398 24212
rect 55440 24172 55480 24212
rect 59112 24172 59152 24212
rect 59194 24172 59234 24212
rect 59276 24172 59316 24212
rect 59358 24172 59398 24212
rect 59440 24172 59480 24212
rect 63112 24172 63152 24212
rect 63194 24172 63234 24212
rect 63276 24172 63316 24212
rect 63358 24172 63398 24212
rect 63440 24172 63480 24212
rect 67112 24172 67152 24212
rect 67194 24172 67234 24212
rect 67276 24172 67316 24212
rect 67358 24172 67398 24212
rect 67440 24172 67480 24212
rect 71112 24172 71152 24212
rect 71194 24172 71234 24212
rect 71276 24172 71316 24212
rect 71358 24172 71398 24212
rect 71440 24172 71480 24212
rect 75112 24172 75152 24212
rect 75194 24172 75234 24212
rect 75276 24172 75316 24212
rect 75358 24172 75398 24212
rect 75440 24172 75480 24212
rect 79112 24172 79152 24212
rect 79194 24172 79234 24212
rect 79276 24172 79316 24212
rect 79358 24172 79398 24212
rect 79440 24172 79480 24212
rect 83112 24172 83152 24212
rect 83194 24172 83234 24212
rect 83276 24172 83316 24212
rect 83358 24172 83398 24212
rect 83440 24172 83480 24212
rect 87112 24172 87152 24212
rect 87194 24172 87234 24212
rect 87276 24172 87316 24212
rect 87358 24172 87398 24212
rect 87440 24172 87480 24212
rect 91112 24172 91152 24212
rect 91194 24172 91234 24212
rect 91276 24172 91316 24212
rect 91358 24172 91398 24212
rect 91440 24172 91480 24212
rect 95112 24172 95152 24212
rect 95194 24172 95234 24212
rect 95276 24172 95316 24212
rect 95358 24172 95398 24212
rect 95440 24172 95480 24212
rect 99112 24172 99152 24212
rect 99194 24172 99234 24212
rect 99276 24172 99316 24212
rect 99358 24172 99398 24212
rect 99440 24172 99480 24212
rect 81868 24004 81908 24044
rect 80140 23920 80180 23960
rect 82636 23920 82676 23960
rect 85132 23920 85172 23960
rect 85900 23920 85940 23960
rect 86668 23920 86708 23960
rect 87916 23920 87956 23960
rect 89068 23920 89108 23960
rect 91468 23920 91508 23960
rect 92428 23920 92468 23960
rect 93580 23920 93620 23960
rect 80332 23836 80372 23876
rect 81676 23836 81716 23876
rect 82444 23836 82484 23876
rect 84940 23836 84980 23876
rect 85708 23836 85748 23876
rect 86476 23836 86516 23876
rect 87724 23836 87764 23876
rect 88876 23836 88916 23876
rect 91276 23836 91316 23876
rect 93388 23836 93428 23876
rect 652 23752 692 23792
rect 844 23752 884 23792
rect 92332 23752 92372 23792
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 8352 23416 8392 23456
rect 8434 23416 8474 23456
rect 8516 23416 8556 23456
rect 8598 23416 8638 23456
rect 8680 23416 8720 23456
rect 12352 23416 12392 23456
rect 12434 23416 12474 23456
rect 12516 23416 12556 23456
rect 12598 23416 12638 23456
rect 12680 23416 12720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 20352 23416 20392 23456
rect 20434 23416 20474 23456
rect 20516 23416 20556 23456
rect 20598 23416 20638 23456
rect 20680 23416 20720 23456
rect 24352 23416 24392 23456
rect 24434 23416 24474 23456
rect 24516 23416 24556 23456
rect 24598 23416 24638 23456
rect 24680 23416 24720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 32352 23416 32392 23456
rect 32434 23416 32474 23456
rect 32516 23416 32556 23456
rect 32598 23416 32638 23456
rect 32680 23416 32720 23456
rect 36352 23416 36392 23456
rect 36434 23416 36474 23456
rect 36516 23416 36556 23456
rect 36598 23416 36638 23456
rect 36680 23416 36720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 44352 23416 44392 23456
rect 44434 23416 44474 23456
rect 44516 23416 44556 23456
rect 44598 23416 44638 23456
rect 44680 23416 44720 23456
rect 48352 23416 48392 23456
rect 48434 23416 48474 23456
rect 48516 23416 48556 23456
rect 48598 23416 48638 23456
rect 48680 23416 48720 23456
rect 52352 23416 52392 23456
rect 52434 23416 52474 23456
rect 52516 23416 52556 23456
rect 52598 23416 52638 23456
rect 52680 23416 52720 23456
rect 56352 23416 56392 23456
rect 56434 23416 56474 23456
rect 56516 23416 56556 23456
rect 56598 23416 56638 23456
rect 56680 23416 56720 23456
rect 60352 23416 60392 23456
rect 60434 23416 60474 23456
rect 60516 23416 60556 23456
rect 60598 23416 60638 23456
rect 60680 23416 60720 23456
rect 64352 23416 64392 23456
rect 64434 23416 64474 23456
rect 64516 23416 64556 23456
rect 64598 23416 64638 23456
rect 64680 23416 64720 23456
rect 68352 23416 68392 23456
rect 68434 23416 68474 23456
rect 68516 23416 68556 23456
rect 68598 23416 68638 23456
rect 68680 23416 68720 23456
rect 72352 23416 72392 23456
rect 72434 23416 72474 23456
rect 72516 23416 72556 23456
rect 72598 23416 72638 23456
rect 72680 23416 72720 23456
rect 76352 23416 76392 23456
rect 76434 23416 76474 23456
rect 76516 23416 76556 23456
rect 76598 23416 76638 23456
rect 76680 23416 76720 23456
rect 80352 23416 80392 23456
rect 80434 23416 80474 23456
rect 80516 23416 80556 23456
rect 80598 23416 80638 23456
rect 80680 23416 80720 23456
rect 84352 23416 84392 23456
rect 84434 23416 84474 23456
rect 84516 23416 84556 23456
rect 84598 23416 84638 23456
rect 84680 23416 84720 23456
rect 88352 23416 88392 23456
rect 88434 23416 88474 23456
rect 88516 23416 88556 23456
rect 88598 23416 88638 23456
rect 88680 23416 88720 23456
rect 92352 23416 92392 23456
rect 92434 23416 92474 23456
rect 92516 23416 92556 23456
rect 92598 23416 92638 23456
rect 92680 23416 92720 23456
rect 96352 23416 96392 23456
rect 96434 23416 96474 23456
rect 96516 23416 96556 23456
rect 96598 23416 96638 23456
rect 96680 23416 96720 23456
rect 652 23080 692 23120
rect 844 23080 884 23120
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 7112 22660 7152 22700
rect 7194 22660 7234 22700
rect 7276 22660 7316 22700
rect 7358 22660 7398 22700
rect 7440 22660 7480 22700
rect 11112 22660 11152 22700
rect 11194 22660 11234 22700
rect 11276 22660 11316 22700
rect 11358 22660 11398 22700
rect 11440 22660 11480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 19112 22660 19152 22700
rect 19194 22660 19234 22700
rect 19276 22660 19316 22700
rect 19358 22660 19398 22700
rect 19440 22660 19480 22700
rect 23112 22660 23152 22700
rect 23194 22660 23234 22700
rect 23276 22660 23316 22700
rect 23358 22660 23398 22700
rect 23440 22660 23480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 31112 22660 31152 22700
rect 31194 22660 31234 22700
rect 31276 22660 31316 22700
rect 31358 22660 31398 22700
rect 31440 22660 31480 22700
rect 35112 22660 35152 22700
rect 35194 22660 35234 22700
rect 35276 22660 35316 22700
rect 35358 22660 35398 22700
rect 35440 22660 35480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 43112 22660 43152 22700
rect 43194 22660 43234 22700
rect 43276 22660 43316 22700
rect 43358 22660 43398 22700
rect 43440 22660 43480 22700
rect 47112 22660 47152 22700
rect 47194 22660 47234 22700
rect 47276 22660 47316 22700
rect 47358 22660 47398 22700
rect 47440 22660 47480 22700
rect 51112 22660 51152 22700
rect 51194 22660 51234 22700
rect 51276 22660 51316 22700
rect 51358 22660 51398 22700
rect 51440 22660 51480 22700
rect 55112 22660 55152 22700
rect 55194 22660 55234 22700
rect 55276 22660 55316 22700
rect 55358 22660 55398 22700
rect 55440 22660 55480 22700
rect 59112 22660 59152 22700
rect 59194 22660 59234 22700
rect 59276 22660 59316 22700
rect 59358 22660 59398 22700
rect 59440 22660 59480 22700
rect 63112 22660 63152 22700
rect 63194 22660 63234 22700
rect 63276 22660 63316 22700
rect 63358 22660 63398 22700
rect 63440 22660 63480 22700
rect 67112 22660 67152 22700
rect 67194 22660 67234 22700
rect 67276 22660 67316 22700
rect 67358 22660 67398 22700
rect 67440 22660 67480 22700
rect 71112 22660 71152 22700
rect 71194 22660 71234 22700
rect 71276 22660 71316 22700
rect 71358 22660 71398 22700
rect 71440 22660 71480 22700
rect 75112 22660 75152 22700
rect 75194 22660 75234 22700
rect 75276 22660 75316 22700
rect 75358 22660 75398 22700
rect 75440 22660 75480 22700
rect 79112 22660 79152 22700
rect 79194 22660 79234 22700
rect 79276 22660 79316 22700
rect 79358 22660 79398 22700
rect 79440 22660 79480 22700
rect 83112 22660 83152 22700
rect 83194 22660 83234 22700
rect 83276 22660 83316 22700
rect 83358 22660 83398 22700
rect 83440 22660 83480 22700
rect 87112 22660 87152 22700
rect 87194 22660 87234 22700
rect 87276 22660 87316 22700
rect 87358 22660 87398 22700
rect 87440 22660 87480 22700
rect 91112 22660 91152 22700
rect 91194 22660 91234 22700
rect 91276 22660 91316 22700
rect 91358 22660 91398 22700
rect 91440 22660 91480 22700
rect 95112 22660 95152 22700
rect 95194 22660 95234 22700
rect 95276 22660 95316 22700
rect 95358 22660 95398 22700
rect 95440 22660 95480 22700
rect 99112 22660 99152 22700
rect 99194 22660 99234 22700
rect 99276 22660 99316 22700
rect 99358 22660 99398 22700
rect 99440 22660 99480 22700
rect 652 22408 692 22448
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 8352 21904 8392 21944
rect 8434 21904 8474 21944
rect 8516 21904 8556 21944
rect 8598 21904 8638 21944
rect 8680 21904 8720 21944
rect 12352 21904 12392 21944
rect 12434 21904 12474 21944
rect 12516 21904 12556 21944
rect 12598 21904 12638 21944
rect 12680 21904 12720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 20352 21904 20392 21944
rect 20434 21904 20474 21944
rect 20516 21904 20556 21944
rect 20598 21904 20638 21944
rect 20680 21904 20720 21944
rect 24352 21904 24392 21944
rect 24434 21904 24474 21944
rect 24516 21904 24556 21944
rect 24598 21904 24638 21944
rect 24680 21904 24720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 32352 21904 32392 21944
rect 32434 21904 32474 21944
rect 32516 21904 32556 21944
rect 32598 21904 32638 21944
rect 32680 21904 32720 21944
rect 36352 21904 36392 21944
rect 36434 21904 36474 21944
rect 36516 21904 36556 21944
rect 36598 21904 36638 21944
rect 36680 21904 36720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 44352 21904 44392 21944
rect 44434 21904 44474 21944
rect 44516 21904 44556 21944
rect 44598 21904 44638 21944
rect 44680 21904 44720 21944
rect 48352 21904 48392 21944
rect 48434 21904 48474 21944
rect 48516 21904 48556 21944
rect 48598 21904 48638 21944
rect 48680 21904 48720 21944
rect 52352 21904 52392 21944
rect 52434 21904 52474 21944
rect 52516 21904 52556 21944
rect 52598 21904 52638 21944
rect 52680 21904 52720 21944
rect 56352 21904 56392 21944
rect 56434 21904 56474 21944
rect 56516 21904 56556 21944
rect 56598 21904 56638 21944
rect 56680 21904 56720 21944
rect 60352 21904 60392 21944
rect 60434 21904 60474 21944
rect 60516 21904 60556 21944
rect 60598 21904 60638 21944
rect 60680 21904 60720 21944
rect 64352 21904 64392 21944
rect 64434 21904 64474 21944
rect 64516 21904 64556 21944
rect 64598 21904 64638 21944
rect 64680 21904 64720 21944
rect 68352 21904 68392 21944
rect 68434 21904 68474 21944
rect 68516 21904 68556 21944
rect 68598 21904 68638 21944
rect 68680 21904 68720 21944
rect 72352 21904 72392 21944
rect 72434 21904 72474 21944
rect 72516 21904 72556 21944
rect 72598 21904 72638 21944
rect 72680 21904 72720 21944
rect 76352 21904 76392 21944
rect 76434 21904 76474 21944
rect 76516 21904 76556 21944
rect 76598 21904 76638 21944
rect 76680 21904 76720 21944
rect 80352 21904 80392 21944
rect 80434 21904 80474 21944
rect 80516 21904 80556 21944
rect 80598 21904 80638 21944
rect 80680 21904 80720 21944
rect 84352 21904 84392 21944
rect 84434 21904 84474 21944
rect 84516 21904 84556 21944
rect 84598 21904 84638 21944
rect 84680 21904 84720 21944
rect 88352 21904 88392 21944
rect 88434 21904 88474 21944
rect 88516 21904 88556 21944
rect 88598 21904 88638 21944
rect 88680 21904 88720 21944
rect 92352 21904 92392 21944
rect 92434 21904 92474 21944
rect 92516 21904 92556 21944
rect 92598 21904 92638 21944
rect 92680 21904 92720 21944
rect 96352 21904 96392 21944
rect 96434 21904 96474 21944
rect 96516 21904 96556 21944
rect 96598 21904 96638 21944
rect 96680 21904 96720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 7112 21148 7152 21188
rect 7194 21148 7234 21188
rect 7276 21148 7316 21188
rect 7358 21148 7398 21188
rect 7440 21148 7480 21188
rect 11112 21148 11152 21188
rect 11194 21148 11234 21188
rect 11276 21148 11316 21188
rect 11358 21148 11398 21188
rect 11440 21148 11480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 19112 21148 19152 21188
rect 19194 21148 19234 21188
rect 19276 21148 19316 21188
rect 19358 21148 19398 21188
rect 19440 21148 19480 21188
rect 23112 21148 23152 21188
rect 23194 21148 23234 21188
rect 23276 21148 23316 21188
rect 23358 21148 23398 21188
rect 23440 21148 23480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 31112 21148 31152 21188
rect 31194 21148 31234 21188
rect 31276 21148 31316 21188
rect 31358 21148 31398 21188
rect 31440 21148 31480 21188
rect 35112 21148 35152 21188
rect 35194 21148 35234 21188
rect 35276 21148 35316 21188
rect 35358 21148 35398 21188
rect 35440 21148 35480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 43112 21148 43152 21188
rect 43194 21148 43234 21188
rect 43276 21148 43316 21188
rect 43358 21148 43398 21188
rect 43440 21148 43480 21188
rect 47112 21148 47152 21188
rect 47194 21148 47234 21188
rect 47276 21148 47316 21188
rect 47358 21148 47398 21188
rect 47440 21148 47480 21188
rect 51112 21148 51152 21188
rect 51194 21148 51234 21188
rect 51276 21148 51316 21188
rect 51358 21148 51398 21188
rect 51440 21148 51480 21188
rect 55112 21148 55152 21188
rect 55194 21148 55234 21188
rect 55276 21148 55316 21188
rect 55358 21148 55398 21188
rect 55440 21148 55480 21188
rect 59112 21148 59152 21188
rect 59194 21148 59234 21188
rect 59276 21148 59316 21188
rect 59358 21148 59398 21188
rect 59440 21148 59480 21188
rect 63112 21148 63152 21188
rect 63194 21148 63234 21188
rect 63276 21148 63316 21188
rect 63358 21148 63398 21188
rect 63440 21148 63480 21188
rect 67112 21148 67152 21188
rect 67194 21148 67234 21188
rect 67276 21148 67316 21188
rect 67358 21148 67398 21188
rect 67440 21148 67480 21188
rect 71112 21148 71152 21188
rect 71194 21148 71234 21188
rect 71276 21148 71316 21188
rect 71358 21148 71398 21188
rect 71440 21148 71480 21188
rect 75112 21148 75152 21188
rect 75194 21148 75234 21188
rect 75276 21148 75316 21188
rect 75358 21148 75398 21188
rect 75440 21148 75480 21188
rect 79112 21148 79152 21188
rect 79194 21148 79234 21188
rect 79276 21148 79316 21188
rect 79358 21148 79398 21188
rect 79440 21148 79480 21188
rect 83112 21148 83152 21188
rect 83194 21148 83234 21188
rect 83276 21148 83316 21188
rect 83358 21148 83398 21188
rect 83440 21148 83480 21188
rect 87112 21148 87152 21188
rect 87194 21148 87234 21188
rect 87276 21148 87316 21188
rect 87358 21148 87398 21188
rect 87440 21148 87480 21188
rect 91112 21148 91152 21188
rect 91194 21148 91234 21188
rect 91276 21148 91316 21188
rect 91358 21148 91398 21188
rect 91440 21148 91480 21188
rect 95112 21148 95152 21188
rect 95194 21148 95234 21188
rect 95276 21148 95316 21188
rect 95358 21148 95398 21188
rect 95440 21148 95480 21188
rect 99112 21148 99152 21188
rect 99194 21148 99234 21188
rect 99276 21148 99316 21188
rect 99358 21148 99398 21188
rect 99440 21148 99480 21188
rect 652 20896 692 20936
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 8352 20392 8392 20432
rect 8434 20392 8474 20432
rect 8516 20392 8556 20432
rect 8598 20392 8638 20432
rect 8680 20392 8720 20432
rect 12352 20392 12392 20432
rect 12434 20392 12474 20432
rect 12516 20392 12556 20432
rect 12598 20392 12638 20432
rect 12680 20392 12720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 20352 20392 20392 20432
rect 20434 20392 20474 20432
rect 20516 20392 20556 20432
rect 20598 20392 20638 20432
rect 20680 20392 20720 20432
rect 24352 20392 24392 20432
rect 24434 20392 24474 20432
rect 24516 20392 24556 20432
rect 24598 20392 24638 20432
rect 24680 20392 24720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 32352 20392 32392 20432
rect 32434 20392 32474 20432
rect 32516 20392 32556 20432
rect 32598 20392 32638 20432
rect 32680 20392 32720 20432
rect 36352 20392 36392 20432
rect 36434 20392 36474 20432
rect 36516 20392 36556 20432
rect 36598 20392 36638 20432
rect 36680 20392 36720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 44352 20392 44392 20432
rect 44434 20392 44474 20432
rect 44516 20392 44556 20432
rect 44598 20392 44638 20432
rect 44680 20392 44720 20432
rect 48352 20392 48392 20432
rect 48434 20392 48474 20432
rect 48516 20392 48556 20432
rect 48598 20392 48638 20432
rect 48680 20392 48720 20432
rect 52352 20392 52392 20432
rect 52434 20392 52474 20432
rect 52516 20392 52556 20432
rect 52598 20392 52638 20432
rect 52680 20392 52720 20432
rect 56352 20392 56392 20432
rect 56434 20392 56474 20432
rect 56516 20392 56556 20432
rect 56598 20392 56638 20432
rect 56680 20392 56720 20432
rect 60352 20392 60392 20432
rect 60434 20392 60474 20432
rect 60516 20392 60556 20432
rect 60598 20392 60638 20432
rect 60680 20392 60720 20432
rect 64352 20392 64392 20432
rect 64434 20392 64474 20432
rect 64516 20392 64556 20432
rect 64598 20392 64638 20432
rect 64680 20392 64720 20432
rect 68352 20392 68392 20432
rect 68434 20392 68474 20432
rect 68516 20392 68556 20432
rect 68598 20392 68638 20432
rect 68680 20392 68720 20432
rect 72352 20392 72392 20432
rect 72434 20392 72474 20432
rect 72516 20392 72556 20432
rect 72598 20392 72638 20432
rect 72680 20392 72720 20432
rect 76352 20392 76392 20432
rect 76434 20392 76474 20432
rect 76516 20392 76556 20432
rect 76598 20392 76638 20432
rect 76680 20392 76720 20432
rect 80352 20392 80392 20432
rect 80434 20392 80474 20432
rect 80516 20392 80556 20432
rect 80598 20392 80638 20432
rect 80680 20392 80720 20432
rect 84352 20392 84392 20432
rect 84434 20392 84474 20432
rect 84516 20392 84556 20432
rect 84598 20392 84638 20432
rect 84680 20392 84720 20432
rect 88352 20392 88392 20432
rect 88434 20392 88474 20432
rect 88516 20392 88556 20432
rect 88598 20392 88638 20432
rect 88680 20392 88720 20432
rect 92352 20392 92392 20432
rect 92434 20392 92474 20432
rect 92516 20392 92556 20432
rect 92598 20392 92638 20432
rect 92680 20392 92720 20432
rect 96352 20392 96392 20432
rect 96434 20392 96474 20432
rect 96516 20392 96556 20432
rect 96598 20392 96638 20432
rect 96680 20392 96720 20432
rect 652 19888 692 19928
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 7112 19636 7152 19676
rect 7194 19636 7234 19676
rect 7276 19636 7316 19676
rect 7358 19636 7398 19676
rect 7440 19636 7480 19676
rect 11112 19636 11152 19676
rect 11194 19636 11234 19676
rect 11276 19636 11316 19676
rect 11358 19636 11398 19676
rect 11440 19636 11480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 19112 19636 19152 19676
rect 19194 19636 19234 19676
rect 19276 19636 19316 19676
rect 19358 19636 19398 19676
rect 19440 19636 19480 19676
rect 23112 19636 23152 19676
rect 23194 19636 23234 19676
rect 23276 19636 23316 19676
rect 23358 19636 23398 19676
rect 23440 19636 23480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 31112 19636 31152 19676
rect 31194 19636 31234 19676
rect 31276 19636 31316 19676
rect 31358 19636 31398 19676
rect 31440 19636 31480 19676
rect 35112 19636 35152 19676
rect 35194 19636 35234 19676
rect 35276 19636 35316 19676
rect 35358 19636 35398 19676
rect 35440 19636 35480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 43112 19636 43152 19676
rect 43194 19636 43234 19676
rect 43276 19636 43316 19676
rect 43358 19636 43398 19676
rect 43440 19636 43480 19676
rect 47112 19636 47152 19676
rect 47194 19636 47234 19676
rect 47276 19636 47316 19676
rect 47358 19636 47398 19676
rect 47440 19636 47480 19676
rect 51112 19636 51152 19676
rect 51194 19636 51234 19676
rect 51276 19636 51316 19676
rect 51358 19636 51398 19676
rect 51440 19636 51480 19676
rect 55112 19636 55152 19676
rect 55194 19636 55234 19676
rect 55276 19636 55316 19676
rect 55358 19636 55398 19676
rect 55440 19636 55480 19676
rect 59112 19636 59152 19676
rect 59194 19636 59234 19676
rect 59276 19636 59316 19676
rect 59358 19636 59398 19676
rect 59440 19636 59480 19676
rect 63112 19636 63152 19676
rect 63194 19636 63234 19676
rect 63276 19636 63316 19676
rect 63358 19636 63398 19676
rect 63440 19636 63480 19676
rect 67112 19636 67152 19676
rect 67194 19636 67234 19676
rect 67276 19636 67316 19676
rect 67358 19636 67398 19676
rect 67440 19636 67480 19676
rect 71112 19636 71152 19676
rect 71194 19636 71234 19676
rect 71276 19636 71316 19676
rect 71358 19636 71398 19676
rect 71440 19636 71480 19676
rect 75112 19636 75152 19676
rect 75194 19636 75234 19676
rect 75276 19636 75316 19676
rect 75358 19636 75398 19676
rect 75440 19636 75480 19676
rect 79112 19636 79152 19676
rect 79194 19636 79234 19676
rect 79276 19636 79316 19676
rect 79358 19636 79398 19676
rect 79440 19636 79480 19676
rect 83112 19636 83152 19676
rect 83194 19636 83234 19676
rect 83276 19636 83316 19676
rect 83358 19636 83398 19676
rect 83440 19636 83480 19676
rect 87112 19636 87152 19676
rect 87194 19636 87234 19676
rect 87276 19636 87316 19676
rect 87358 19636 87398 19676
rect 87440 19636 87480 19676
rect 91112 19636 91152 19676
rect 91194 19636 91234 19676
rect 91276 19636 91316 19676
rect 91358 19636 91398 19676
rect 91440 19636 91480 19676
rect 95112 19636 95152 19676
rect 95194 19636 95234 19676
rect 95276 19636 95316 19676
rect 95358 19636 95398 19676
rect 95440 19636 95480 19676
rect 99112 19636 99152 19676
rect 99194 19636 99234 19676
rect 99276 19636 99316 19676
rect 99358 19636 99398 19676
rect 99440 19636 99480 19676
rect 652 19384 692 19424
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 8352 18880 8392 18920
rect 8434 18880 8474 18920
rect 8516 18880 8556 18920
rect 8598 18880 8638 18920
rect 8680 18880 8720 18920
rect 12352 18880 12392 18920
rect 12434 18880 12474 18920
rect 12516 18880 12556 18920
rect 12598 18880 12638 18920
rect 12680 18880 12720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 20352 18880 20392 18920
rect 20434 18880 20474 18920
rect 20516 18880 20556 18920
rect 20598 18880 20638 18920
rect 20680 18880 20720 18920
rect 24352 18880 24392 18920
rect 24434 18880 24474 18920
rect 24516 18880 24556 18920
rect 24598 18880 24638 18920
rect 24680 18880 24720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 32352 18880 32392 18920
rect 32434 18880 32474 18920
rect 32516 18880 32556 18920
rect 32598 18880 32638 18920
rect 32680 18880 32720 18920
rect 36352 18880 36392 18920
rect 36434 18880 36474 18920
rect 36516 18880 36556 18920
rect 36598 18880 36638 18920
rect 36680 18880 36720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 44352 18880 44392 18920
rect 44434 18880 44474 18920
rect 44516 18880 44556 18920
rect 44598 18880 44638 18920
rect 44680 18880 44720 18920
rect 48352 18880 48392 18920
rect 48434 18880 48474 18920
rect 48516 18880 48556 18920
rect 48598 18880 48638 18920
rect 48680 18880 48720 18920
rect 52352 18880 52392 18920
rect 52434 18880 52474 18920
rect 52516 18880 52556 18920
rect 52598 18880 52638 18920
rect 52680 18880 52720 18920
rect 56352 18880 56392 18920
rect 56434 18880 56474 18920
rect 56516 18880 56556 18920
rect 56598 18880 56638 18920
rect 56680 18880 56720 18920
rect 60352 18880 60392 18920
rect 60434 18880 60474 18920
rect 60516 18880 60556 18920
rect 60598 18880 60638 18920
rect 60680 18880 60720 18920
rect 64352 18880 64392 18920
rect 64434 18880 64474 18920
rect 64516 18880 64556 18920
rect 64598 18880 64638 18920
rect 64680 18880 64720 18920
rect 68352 18880 68392 18920
rect 68434 18880 68474 18920
rect 68516 18880 68556 18920
rect 68598 18880 68638 18920
rect 68680 18880 68720 18920
rect 72352 18880 72392 18920
rect 72434 18880 72474 18920
rect 72516 18880 72556 18920
rect 72598 18880 72638 18920
rect 72680 18880 72720 18920
rect 76352 18880 76392 18920
rect 76434 18880 76474 18920
rect 76516 18880 76556 18920
rect 76598 18880 76638 18920
rect 76680 18880 76720 18920
rect 80352 18880 80392 18920
rect 80434 18880 80474 18920
rect 80516 18880 80556 18920
rect 80598 18880 80638 18920
rect 80680 18880 80720 18920
rect 84352 18880 84392 18920
rect 84434 18880 84474 18920
rect 84516 18880 84556 18920
rect 84598 18880 84638 18920
rect 84680 18880 84720 18920
rect 88352 18880 88392 18920
rect 88434 18880 88474 18920
rect 88516 18880 88556 18920
rect 88598 18880 88638 18920
rect 88680 18880 88720 18920
rect 92352 18880 92392 18920
rect 92434 18880 92474 18920
rect 92516 18880 92556 18920
rect 92598 18880 92638 18920
rect 92680 18880 92720 18920
rect 96352 18880 96392 18920
rect 96434 18880 96474 18920
rect 96516 18880 96556 18920
rect 96598 18880 96638 18920
rect 96680 18880 96720 18920
rect 652 18376 692 18416
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 7112 18124 7152 18164
rect 7194 18124 7234 18164
rect 7276 18124 7316 18164
rect 7358 18124 7398 18164
rect 7440 18124 7480 18164
rect 11112 18124 11152 18164
rect 11194 18124 11234 18164
rect 11276 18124 11316 18164
rect 11358 18124 11398 18164
rect 11440 18124 11480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 19112 18124 19152 18164
rect 19194 18124 19234 18164
rect 19276 18124 19316 18164
rect 19358 18124 19398 18164
rect 19440 18124 19480 18164
rect 23112 18124 23152 18164
rect 23194 18124 23234 18164
rect 23276 18124 23316 18164
rect 23358 18124 23398 18164
rect 23440 18124 23480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 31112 18124 31152 18164
rect 31194 18124 31234 18164
rect 31276 18124 31316 18164
rect 31358 18124 31398 18164
rect 31440 18124 31480 18164
rect 35112 18124 35152 18164
rect 35194 18124 35234 18164
rect 35276 18124 35316 18164
rect 35358 18124 35398 18164
rect 35440 18124 35480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 43112 18124 43152 18164
rect 43194 18124 43234 18164
rect 43276 18124 43316 18164
rect 43358 18124 43398 18164
rect 43440 18124 43480 18164
rect 47112 18124 47152 18164
rect 47194 18124 47234 18164
rect 47276 18124 47316 18164
rect 47358 18124 47398 18164
rect 47440 18124 47480 18164
rect 51112 18124 51152 18164
rect 51194 18124 51234 18164
rect 51276 18124 51316 18164
rect 51358 18124 51398 18164
rect 51440 18124 51480 18164
rect 55112 18124 55152 18164
rect 55194 18124 55234 18164
rect 55276 18124 55316 18164
rect 55358 18124 55398 18164
rect 55440 18124 55480 18164
rect 59112 18124 59152 18164
rect 59194 18124 59234 18164
rect 59276 18124 59316 18164
rect 59358 18124 59398 18164
rect 59440 18124 59480 18164
rect 63112 18124 63152 18164
rect 63194 18124 63234 18164
rect 63276 18124 63316 18164
rect 63358 18124 63398 18164
rect 63440 18124 63480 18164
rect 67112 18124 67152 18164
rect 67194 18124 67234 18164
rect 67276 18124 67316 18164
rect 67358 18124 67398 18164
rect 67440 18124 67480 18164
rect 71112 18124 71152 18164
rect 71194 18124 71234 18164
rect 71276 18124 71316 18164
rect 71358 18124 71398 18164
rect 71440 18124 71480 18164
rect 75112 18124 75152 18164
rect 75194 18124 75234 18164
rect 75276 18124 75316 18164
rect 75358 18124 75398 18164
rect 75440 18124 75480 18164
rect 79112 18124 79152 18164
rect 79194 18124 79234 18164
rect 79276 18124 79316 18164
rect 79358 18124 79398 18164
rect 79440 18124 79480 18164
rect 83112 18124 83152 18164
rect 83194 18124 83234 18164
rect 83276 18124 83316 18164
rect 83358 18124 83398 18164
rect 83440 18124 83480 18164
rect 87112 18124 87152 18164
rect 87194 18124 87234 18164
rect 87276 18124 87316 18164
rect 87358 18124 87398 18164
rect 87440 18124 87480 18164
rect 91112 18124 91152 18164
rect 91194 18124 91234 18164
rect 91276 18124 91316 18164
rect 91358 18124 91398 18164
rect 91440 18124 91480 18164
rect 95112 18124 95152 18164
rect 95194 18124 95234 18164
rect 95276 18124 95316 18164
rect 95358 18124 95398 18164
rect 95440 18124 95480 18164
rect 99112 18124 99152 18164
rect 99194 18124 99234 18164
rect 99276 18124 99316 18164
rect 99358 18124 99398 18164
rect 99440 18124 99480 18164
rect 652 17872 692 17912
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 8352 17368 8392 17408
rect 8434 17368 8474 17408
rect 8516 17368 8556 17408
rect 8598 17368 8638 17408
rect 8680 17368 8720 17408
rect 12352 17368 12392 17408
rect 12434 17368 12474 17408
rect 12516 17368 12556 17408
rect 12598 17368 12638 17408
rect 12680 17368 12720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 20352 17368 20392 17408
rect 20434 17368 20474 17408
rect 20516 17368 20556 17408
rect 20598 17368 20638 17408
rect 20680 17368 20720 17408
rect 24352 17368 24392 17408
rect 24434 17368 24474 17408
rect 24516 17368 24556 17408
rect 24598 17368 24638 17408
rect 24680 17368 24720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 32352 17368 32392 17408
rect 32434 17368 32474 17408
rect 32516 17368 32556 17408
rect 32598 17368 32638 17408
rect 32680 17368 32720 17408
rect 36352 17368 36392 17408
rect 36434 17368 36474 17408
rect 36516 17368 36556 17408
rect 36598 17368 36638 17408
rect 36680 17368 36720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 44352 17368 44392 17408
rect 44434 17368 44474 17408
rect 44516 17368 44556 17408
rect 44598 17368 44638 17408
rect 44680 17368 44720 17408
rect 48352 17368 48392 17408
rect 48434 17368 48474 17408
rect 48516 17368 48556 17408
rect 48598 17368 48638 17408
rect 48680 17368 48720 17408
rect 52352 17368 52392 17408
rect 52434 17368 52474 17408
rect 52516 17368 52556 17408
rect 52598 17368 52638 17408
rect 52680 17368 52720 17408
rect 56352 17368 56392 17408
rect 56434 17368 56474 17408
rect 56516 17368 56556 17408
rect 56598 17368 56638 17408
rect 56680 17368 56720 17408
rect 60352 17368 60392 17408
rect 60434 17368 60474 17408
rect 60516 17368 60556 17408
rect 60598 17368 60638 17408
rect 60680 17368 60720 17408
rect 64352 17368 64392 17408
rect 64434 17368 64474 17408
rect 64516 17368 64556 17408
rect 64598 17368 64638 17408
rect 64680 17368 64720 17408
rect 68352 17368 68392 17408
rect 68434 17368 68474 17408
rect 68516 17368 68556 17408
rect 68598 17368 68638 17408
rect 68680 17368 68720 17408
rect 72352 17368 72392 17408
rect 72434 17368 72474 17408
rect 72516 17368 72556 17408
rect 72598 17368 72638 17408
rect 72680 17368 72720 17408
rect 76352 17368 76392 17408
rect 76434 17368 76474 17408
rect 76516 17368 76556 17408
rect 76598 17368 76638 17408
rect 76680 17368 76720 17408
rect 80352 17368 80392 17408
rect 80434 17368 80474 17408
rect 80516 17368 80556 17408
rect 80598 17368 80638 17408
rect 80680 17368 80720 17408
rect 84352 17368 84392 17408
rect 84434 17368 84474 17408
rect 84516 17368 84556 17408
rect 84598 17368 84638 17408
rect 84680 17368 84720 17408
rect 88352 17368 88392 17408
rect 88434 17368 88474 17408
rect 88516 17368 88556 17408
rect 88598 17368 88638 17408
rect 88680 17368 88720 17408
rect 92352 17368 92392 17408
rect 92434 17368 92474 17408
rect 92516 17368 92556 17408
rect 92598 17368 92638 17408
rect 92680 17368 92720 17408
rect 96352 17368 96392 17408
rect 96434 17368 96474 17408
rect 96516 17368 96556 17408
rect 96598 17368 96638 17408
rect 96680 17368 96720 17408
rect 86572 17032 86612 17072
rect 86764 17032 86804 17072
rect 80428 16948 80468 16988
rect 86188 16948 86228 16988
rect 652 16864 692 16904
rect 80620 16780 80660 16820
rect 86380 16780 86420 16820
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 7112 16612 7152 16652
rect 7194 16612 7234 16652
rect 7276 16612 7316 16652
rect 7358 16612 7398 16652
rect 7440 16612 7480 16652
rect 11112 16612 11152 16652
rect 11194 16612 11234 16652
rect 11276 16612 11316 16652
rect 11358 16612 11398 16652
rect 11440 16612 11480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 19112 16612 19152 16652
rect 19194 16612 19234 16652
rect 19276 16612 19316 16652
rect 19358 16612 19398 16652
rect 19440 16612 19480 16652
rect 23112 16612 23152 16652
rect 23194 16612 23234 16652
rect 23276 16612 23316 16652
rect 23358 16612 23398 16652
rect 23440 16612 23480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 31112 16612 31152 16652
rect 31194 16612 31234 16652
rect 31276 16612 31316 16652
rect 31358 16612 31398 16652
rect 31440 16612 31480 16652
rect 35112 16612 35152 16652
rect 35194 16612 35234 16652
rect 35276 16612 35316 16652
rect 35358 16612 35398 16652
rect 35440 16612 35480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 43112 16612 43152 16652
rect 43194 16612 43234 16652
rect 43276 16612 43316 16652
rect 43358 16612 43398 16652
rect 43440 16612 43480 16652
rect 47112 16612 47152 16652
rect 47194 16612 47234 16652
rect 47276 16612 47316 16652
rect 47358 16612 47398 16652
rect 47440 16612 47480 16652
rect 51112 16612 51152 16652
rect 51194 16612 51234 16652
rect 51276 16612 51316 16652
rect 51358 16612 51398 16652
rect 51440 16612 51480 16652
rect 55112 16612 55152 16652
rect 55194 16612 55234 16652
rect 55276 16612 55316 16652
rect 55358 16612 55398 16652
rect 55440 16612 55480 16652
rect 59112 16612 59152 16652
rect 59194 16612 59234 16652
rect 59276 16612 59316 16652
rect 59358 16612 59398 16652
rect 59440 16612 59480 16652
rect 63112 16612 63152 16652
rect 63194 16612 63234 16652
rect 63276 16612 63316 16652
rect 63358 16612 63398 16652
rect 63440 16612 63480 16652
rect 67112 16612 67152 16652
rect 67194 16612 67234 16652
rect 67276 16612 67316 16652
rect 67358 16612 67398 16652
rect 67440 16612 67480 16652
rect 71112 16612 71152 16652
rect 71194 16612 71234 16652
rect 71276 16612 71316 16652
rect 71358 16612 71398 16652
rect 71440 16612 71480 16652
rect 75112 16612 75152 16652
rect 75194 16612 75234 16652
rect 75276 16612 75316 16652
rect 75358 16612 75398 16652
rect 75440 16612 75480 16652
rect 79112 16612 79152 16652
rect 79194 16612 79234 16652
rect 79276 16612 79316 16652
rect 79358 16612 79398 16652
rect 79440 16612 79480 16652
rect 83112 16612 83152 16652
rect 83194 16612 83234 16652
rect 83276 16612 83316 16652
rect 83358 16612 83398 16652
rect 83440 16612 83480 16652
rect 87112 16612 87152 16652
rect 87194 16612 87234 16652
rect 87276 16612 87316 16652
rect 87358 16612 87398 16652
rect 87440 16612 87480 16652
rect 91112 16612 91152 16652
rect 91194 16612 91234 16652
rect 91276 16612 91316 16652
rect 91358 16612 91398 16652
rect 91440 16612 91480 16652
rect 95112 16612 95152 16652
rect 95194 16612 95234 16652
rect 95276 16612 95316 16652
rect 95358 16612 95398 16652
rect 95440 16612 95480 16652
rect 99112 16612 99152 16652
rect 99194 16612 99234 16652
rect 99276 16612 99316 16652
rect 99358 16612 99398 16652
rect 99440 16612 99480 16652
rect 652 16360 692 16400
rect 74476 16360 74516 16400
rect 81580 16360 81620 16400
rect 83116 16360 83156 16400
rect 73900 16276 73940 16316
rect 74284 16276 74324 16316
rect 76780 16276 76820 16316
rect 77164 16276 77204 16316
rect 80524 16276 80564 16316
rect 81196 16276 81236 16316
rect 81772 16276 81812 16316
rect 82156 16276 82196 16316
rect 82540 16276 82580 16316
rect 83308 16276 83348 16316
rect 83788 16276 83828 16316
rect 84652 16276 84692 16316
rect 86572 16276 86612 16316
rect 87436 16276 87476 16316
rect 88204 16276 88244 16316
rect 89356 16276 89396 16316
rect 90604 16276 90644 16316
rect 92236 16276 92276 16316
rect 92428 16276 92468 16316
rect 94060 16276 94100 16316
rect 95596 16276 95636 16316
rect 90988 16192 91028 16232
rect 74092 16024 74132 16064
rect 76972 16024 77012 16064
rect 77356 16024 77396 16064
rect 80332 16024 80372 16064
rect 81388 16024 81428 16064
rect 81964 16024 82004 16064
rect 82732 16024 82772 16064
rect 83980 16024 84020 16064
rect 84844 16024 84884 16064
rect 86380 16024 86420 16064
rect 87628 16024 87668 16064
rect 88012 16024 88052 16064
rect 89164 16024 89204 16064
rect 90796 16024 90836 16064
rect 91084 16024 91124 16064
rect 92044 16024 92084 16064
rect 92620 16024 92660 16064
rect 93868 16024 93908 16064
rect 95788 16024 95828 16064
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 8352 15856 8392 15896
rect 8434 15856 8474 15896
rect 8516 15856 8556 15896
rect 8598 15856 8638 15896
rect 8680 15856 8720 15896
rect 12352 15856 12392 15896
rect 12434 15856 12474 15896
rect 12516 15856 12556 15896
rect 12598 15856 12638 15896
rect 12680 15856 12720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 20352 15856 20392 15896
rect 20434 15856 20474 15896
rect 20516 15856 20556 15896
rect 20598 15856 20638 15896
rect 20680 15856 20720 15896
rect 24352 15856 24392 15896
rect 24434 15856 24474 15896
rect 24516 15856 24556 15896
rect 24598 15856 24638 15896
rect 24680 15856 24720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 32352 15856 32392 15896
rect 32434 15856 32474 15896
rect 32516 15856 32556 15896
rect 32598 15856 32638 15896
rect 32680 15856 32720 15896
rect 36352 15856 36392 15896
rect 36434 15856 36474 15896
rect 36516 15856 36556 15896
rect 36598 15856 36638 15896
rect 36680 15856 36720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 44352 15856 44392 15896
rect 44434 15856 44474 15896
rect 44516 15856 44556 15896
rect 44598 15856 44638 15896
rect 44680 15856 44720 15896
rect 48352 15856 48392 15896
rect 48434 15856 48474 15896
rect 48516 15856 48556 15896
rect 48598 15856 48638 15896
rect 48680 15856 48720 15896
rect 52352 15856 52392 15896
rect 52434 15856 52474 15896
rect 52516 15856 52556 15896
rect 52598 15856 52638 15896
rect 52680 15856 52720 15896
rect 56352 15856 56392 15896
rect 56434 15856 56474 15896
rect 56516 15856 56556 15896
rect 56598 15856 56638 15896
rect 56680 15856 56720 15896
rect 60352 15856 60392 15896
rect 60434 15856 60474 15896
rect 60516 15856 60556 15896
rect 60598 15856 60638 15896
rect 60680 15856 60720 15896
rect 64352 15856 64392 15896
rect 64434 15856 64474 15896
rect 64516 15856 64556 15896
rect 64598 15856 64638 15896
rect 64680 15856 64720 15896
rect 68352 15856 68392 15896
rect 68434 15856 68474 15896
rect 68516 15856 68556 15896
rect 68598 15856 68638 15896
rect 68680 15856 68720 15896
rect 72352 15856 72392 15896
rect 72434 15856 72474 15896
rect 72516 15856 72556 15896
rect 72598 15856 72638 15896
rect 72680 15856 72720 15896
rect 76352 15856 76392 15896
rect 76434 15856 76474 15896
rect 76516 15856 76556 15896
rect 76598 15856 76638 15896
rect 76680 15856 76720 15896
rect 80352 15856 80392 15896
rect 80434 15856 80474 15896
rect 80516 15856 80556 15896
rect 80598 15856 80638 15896
rect 80680 15856 80720 15896
rect 84352 15856 84392 15896
rect 84434 15856 84474 15896
rect 84516 15856 84556 15896
rect 84598 15856 84638 15896
rect 84680 15856 84720 15896
rect 88352 15856 88392 15896
rect 88434 15856 88474 15896
rect 88516 15856 88556 15896
rect 88598 15856 88638 15896
rect 88680 15856 88720 15896
rect 92352 15856 92392 15896
rect 92434 15856 92474 15896
rect 92516 15856 92556 15896
rect 92598 15856 92638 15896
rect 92680 15856 92720 15896
rect 96352 15856 96392 15896
rect 96434 15856 96474 15896
rect 96516 15856 96556 15896
rect 96598 15856 96638 15896
rect 96680 15856 96720 15896
rect 81772 15520 81812 15560
rect 83884 15520 83924 15560
rect 87436 15520 87476 15560
rect 98572 15520 98612 15560
rect 844 15436 884 15476
rect 73708 15436 73748 15476
rect 74284 15436 74324 15476
rect 74860 15436 74900 15476
rect 75340 15436 75380 15476
rect 75820 15436 75860 15476
rect 76204 15436 76244 15476
rect 76588 15436 76628 15476
rect 76972 15436 77012 15476
rect 77356 15436 77396 15476
rect 77740 15436 77780 15476
rect 78124 15436 78164 15476
rect 78604 15436 78644 15476
rect 79179 15425 79219 15465
rect 79372 15436 79412 15476
rect 79756 15436 79796 15476
rect 80236 15436 80276 15476
rect 80716 15436 80756 15476
rect 81100 15436 81140 15476
rect 83020 15436 83060 15476
rect 83404 15436 83444 15476
rect 84172 15436 84212 15476
rect 84556 15436 84596 15476
rect 85036 15436 85076 15476
rect 85420 15436 85460 15476
rect 85804 15436 85844 15476
rect 86188 15436 86228 15476
rect 86572 15436 86612 15476
rect 87052 15436 87092 15476
rect 87916 15436 87956 15476
rect 88300 15436 88340 15476
rect 88684 15436 88724 15476
rect 89068 15436 89108 15476
rect 89452 15436 89492 15476
rect 89836 15436 89876 15476
rect 90508 15436 90548 15476
rect 91084 15436 91124 15476
rect 91468 15436 91508 15476
rect 91948 15436 91988 15476
rect 92524 15436 92564 15476
rect 92716 15436 92756 15476
rect 93388 15436 93428 15476
rect 93772 15436 93812 15476
rect 94252 15436 94292 15476
rect 94636 15436 94676 15476
rect 95020 15436 95060 15476
rect 95692 15436 95732 15476
rect 96076 15436 96116 15476
rect 96460 15436 96500 15476
rect 96844 15436 96884 15476
rect 97228 15436 97268 15476
rect 97612 15436 97652 15476
rect 97996 15436 98036 15476
rect 98380 15436 98420 15476
rect 74092 15352 74132 15392
rect 78796 15352 78836 15392
rect 95500 15352 95540 15392
rect 652 15268 692 15308
rect 73900 15268 73940 15308
rect 75052 15268 75092 15308
rect 75532 15268 75572 15308
rect 76012 15268 76052 15308
rect 76396 15268 76436 15308
rect 76780 15268 76820 15308
rect 77164 15268 77204 15308
rect 77548 15268 77588 15308
rect 77932 15268 77972 15308
rect 78316 15268 78356 15308
rect 78988 15268 79028 15308
rect 79564 15268 79604 15308
rect 79948 15268 79988 15308
rect 80428 15268 80468 15308
rect 80908 15268 80948 15308
rect 81292 15268 81332 15308
rect 81868 15268 81908 15308
rect 83212 15268 83252 15308
rect 83596 15268 83636 15308
rect 83980 15268 84020 15308
rect 84364 15268 84404 15308
rect 84748 15268 84788 15308
rect 85228 15268 85268 15308
rect 85612 15268 85652 15308
rect 85996 15268 86036 15308
rect 86380 15268 86420 15308
rect 86764 15268 86804 15308
rect 87244 15268 87284 15308
rect 87532 15268 87572 15308
rect 88108 15268 88148 15308
rect 88492 15268 88532 15308
rect 88876 15268 88916 15308
rect 89260 15268 89300 15308
rect 89644 15268 89684 15308
rect 90028 15268 90068 15308
rect 90700 15268 90740 15308
rect 90892 15268 90932 15308
rect 91660 15268 91700 15308
rect 92140 15268 92180 15308
rect 92332 15268 92372 15308
rect 92908 15268 92948 15308
rect 93580 15268 93620 15308
rect 93964 15268 94004 15308
rect 94444 15268 94484 15308
rect 94828 15268 94868 15308
rect 95212 15268 95252 15308
rect 95884 15268 95924 15308
rect 96268 15268 96308 15308
rect 96652 15268 96692 15308
rect 97036 15268 97076 15308
rect 97420 15268 97460 15308
rect 97804 15268 97844 15308
rect 98188 15268 98228 15308
rect 98668 15268 98708 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 7112 15100 7152 15140
rect 7194 15100 7234 15140
rect 7276 15100 7316 15140
rect 7358 15100 7398 15140
rect 7440 15100 7480 15140
rect 11112 15100 11152 15140
rect 11194 15100 11234 15140
rect 11276 15100 11316 15140
rect 11358 15100 11398 15140
rect 11440 15100 11480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 19112 15100 19152 15140
rect 19194 15100 19234 15140
rect 19276 15100 19316 15140
rect 19358 15100 19398 15140
rect 19440 15100 19480 15140
rect 23112 15100 23152 15140
rect 23194 15100 23234 15140
rect 23276 15100 23316 15140
rect 23358 15100 23398 15140
rect 23440 15100 23480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 31112 15100 31152 15140
rect 31194 15100 31234 15140
rect 31276 15100 31316 15140
rect 31358 15100 31398 15140
rect 31440 15100 31480 15140
rect 35112 15100 35152 15140
rect 35194 15100 35234 15140
rect 35276 15100 35316 15140
rect 35358 15100 35398 15140
rect 35440 15100 35480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 43112 15100 43152 15140
rect 43194 15100 43234 15140
rect 43276 15100 43316 15140
rect 43358 15100 43398 15140
rect 43440 15100 43480 15140
rect 47112 15100 47152 15140
rect 47194 15100 47234 15140
rect 47276 15100 47316 15140
rect 47358 15100 47398 15140
rect 47440 15100 47480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 55112 15100 55152 15140
rect 55194 15100 55234 15140
rect 55276 15100 55316 15140
rect 55358 15100 55398 15140
rect 55440 15100 55480 15140
rect 59112 15100 59152 15140
rect 59194 15100 59234 15140
rect 59276 15100 59316 15140
rect 59358 15100 59398 15140
rect 59440 15100 59480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 67112 15100 67152 15140
rect 67194 15100 67234 15140
rect 67276 15100 67316 15140
rect 67358 15100 67398 15140
rect 67440 15100 67480 15140
rect 1420 14932 1460 14972
rect 73708 14848 73748 14888
rect 844 14764 884 14804
rect 1612 14764 1652 14804
rect 1996 14764 2036 14804
rect 73036 14764 73076 14804
rect 73516 14764 73556 14804
rect 74476 14764 74516 14804
rect 78892 14764 78932 14804
rect 82252 14764 82292 14804
rect 91084 14764 91124 14804
rect 93004 14764 93044 14804
rect 96844 14764 96884 14804
rect 98764 14764 98804 14804
rect 72748 14680 72788 14720
rect 73900 14680 73940 14720
rect 74188 14680 74228 14720
rect 74860 14680 74900 14720
rect 75340 14680 75380 14720
rect 75820 14680 75860 14720
rect 76108 14680 76148 14720
rect 76588 14680 76628 14720
rect 76972 14680 77012 14720
rect 77356 14680 77396 14720
rect 77836 14680 77876 14720
rect 78124 14680 78164 14720
rect 78700 14680 78740 14720
rect 79372 14680 79412 14720
rect 79660 14680 79700 14720
rect 80140 14680 80180 14720
rect 80428 14680 80468 14720
rect 80812 14680 80852 14720
rect 81004 14680 81044 14720
rect 81388 14680 81428 14720
rect 81964 14680 82004 14720
rect 82636 14680 82676 14720
rect 83020 14680 83060 14720
rect 83404 14680 83444 14720
rect 83788 14680 83828 14720
rect 84556 14680 84596 14720
rect 85036 14680 85076 14720
rect 85420 14680 85460 14720
rect 85804 14680 85844 14720
rect 86380 14680 86420 14720
rect 86764 14680 86804 14720
rect 87052 14680 87092 14720
rect 87916 14680 87956 14720
rect 88204 14680 88244 14720
rect 88588 14680 88628 14720
rect 88972 14680 89012 14720
rect 89644 14680 89684 14720
rect 90028 14680 90068 14720
rect 90220 14680 90260 14720
rect 90604 14680 90644 14720
rect 91564 14680 91604 14720
rect 91756 14680 91796 14720
rect 92140 14680 92180 14720
rect 92428 14693 92468 14733
rect 92716 14680 92756 14720
rect 93388 14680 93428 14720
rect 93964 14680 94004 14720
rect 94252 14680 94292 14720
rect 94636 14680 94676 14720
rect 95020 14680 95060 14720
rect 95500 14680 95540 14720
rect 95980 14680 96020 14720
rect 96364 14680 96404 14720
rect 97132 14680 97172 14720
rect 97420 14680 97460 14720
rect 97708 14680 97748 14720
rect 98380 14680 98420 14720
rect 652 14512 692 14552
rect 1804 14512 1844 14552
rect 72844 14512 72884 14552
rect 73228 14512 73268 14552
rect 73996 14512 74036 14552
rect 74284 14512 74324 14552
rect 74668 14512 74708 14552
rect 74956 14512 74996 14552
rect 75436 14512 75476 14552
rect 75916 14512 75956 14552
rect 76204 14512 76244 14552
rect 76684 14512 76724 14552
rect 77068 14512 77108 14552
rect 77452 14512 77492 14552
rect 77932 14512 77972 14552
rect 78220 14512 78260 14552
rect 78604 14512 78644 14552
rect 79084 14512 79124 14552
rect 79468 14512 79508 14552
rect 79756 14512 79796 14552
rect 80236 14512 80276 14552
rect 80524 14512 80564 14552
rect 80716 14512 80756 14552
rect 81100 14512 81140 14552
rect 81484 14512 81524 14552
rect 82060 14512 82100 14552
rect 82444 14512 82484 14552
rect 82732 14512 82772 14552
rect 83116 14512 83156 14552
rect 83500 14512 83540 14552
rect 83884 14512 83924 14552
rect 84652 14512 84692 14552
rect 85132 14512 85172 14552
rect 85516 14512 85556 14552
rect 85900 14512 85940 14552
rect 86284 14512 86324 14552
rect 86668 14512 86708 14552
rect 87148 14512 87188 14552
rect 87820 14512 87860 14552
rect 88300 14512 88340 14552
rect 88684 14512 88724 14552
rect 89068 14512 89108 14552
rect 89548 14512 89588 14552
rect 89932 14512 89972 14552
rect 90316 14512 90356 14552
rect 90700 14512 90740 14552
rect 91276 14512 91316 14552
rect 91468 14512 91508 14552
rect 91852 14512 91892 14552
rect 92236 14512 92276 14552
rect 92524 14512 92564 14552
rect 92812 14512 92852 14552
rect 93196 14512 93236 14552
rect 93484 14512 93524 14552
rect 93868 14512 93908 14552
rect 94348 14512 94388 14552
rect 94732 14512 94772 14552
rect 95116 14512 95156 14552
rect 95404 14512 95444 14552
rect 95884 14512 95924 14552
rect 96268 14512 96308 14552
rect 96652 14512 96692 14552
rect 97036 14512 97076 14552
rect 97516 14512 97556 14552
rect 97804 14512 97844 14552
rect 98284 14512 98324 14552
rect 98572 14512 98612 14552
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 8352 14344 8392 14384
rect 8434 14344 8474 14384
rect 8516 14344 8556 14384
rect 8598 14344 8638 14384
rect 8680 14344 8720 14384
rect 12352 14344 12392 14384
rect 12434 14344 12474 14384
rect 12516 14344 12556 14384
rect 12598 14344 12638 14384
rect 12680 14344 12720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 20352 14344 20392 14384
rect 20434 14344 20474 14384
rect 20516 14344 20556 14384
rect 20598 14344 20638 14384
rect 20680 14344 20720 14384
rect 24352 14344 24392 14384
rect 24434 14344 24474 14384
rect 24516 14344 24556 14384
rect 24598 14344 24638 14384
rect 24680 14344 24720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 32352 14344 32392 14384
rect 32434 14344 32474 14384
rect 32516 14344 32556 14384
rect 32598 14344 32638 14384
rect 32680 14344 32720 14384
rect 36352 14344 36392 14384
rect 36434 14344 36474 14384
rect 36516 14344 36556 14384
rect 36598 14344 36638 14384
rect 36680 14344 36720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 44352 14344 44392 14384
rect 44434 14344 44474 14384
rect 44516 14344 44556 14384
rect 44598 14344 44638 14384
rect 44680 14344 44720 14384
rect 48352 14344 48392 14384
rect 48434 14344 48474 14384
rect 48516 14344 48556 14384
rect 48598 14344 48638 14384
rect 48680 14344 48720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 56352 14344 56392 14384
rect 56434 14344 56474 14384
rect 56516 14344 56556 14384
rect 56598 14344 56638 14384
rect 56680 14344 56720 14384
rect 60352 14344 60392 14384
rect 60434 14344 60474 14384
rect 60516 14344 60556 14384
rect 60598 14344 60638 14384
rect 60680 14344 60720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 68352 14344 68392 14384
rect 68434 14344 68474 14384
rect 68516 14344 68556 14384
rect 68598 14344 68638 14384
rect 68680 14344 68720 14384
rect 1036 14176 1076 14216
rect 70636 14008 70676 14048
rect 70828 14008 70868 14048
rect 71308 14008 71348 14048
rect 1228 13924 1268 13964
rect 71404 13840 71444 13880
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 7112 13588 7152 13628
rect 7194 13588 7234 13628
rect 7276 13588 7316 13628
rect 7358 13588 7398 13628
rect 7440 13588 7480 13628
rect 11112 13588 11152 13628
rect 11194 13588 11234 13628
rect 11276 13588 11316 13628
rect 11358 13588 11398 13628
rect 11440 13588 11480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 19112 13588 19152 13628
rect 19194 13588 19234 13628
rect 19276 13588 19316 13628
rect 19358 13588 19398 13628
rect 19440 13588 19480 13628
rect 23112 13588 23152 13628
rect 23194 13588 23234 13628
rect 23276 13588 23316 13628
rect 23358 13588 23398 13628
rect 23440 13588 23480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 31112 13588 31152 13628
rect 31194 13588 31234 13628
rect 31276 13588 31316 13628
rect 31358 13588 31398 13628
rect 31440 13588 31480 13628
rect 35112 13588 35152 13628
rect 35194 13588 35234 13628
rect 35276 13588 35316 13628
rect 35358 13588 35398 13628
rect 35440 13588 35480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 43112 13588 43152 13628
rect 43194 13588 43234 13628
rect 43276 13588 43316 13628
rect 43358 13588 43398 13628
rect 43440 13588 43480 13628
rect 47112 13588 47152 13628
rect 47194 13588 47234 13628
rect 47276 13588 47316 13628
rect 47358 13588 47398 13628
rect 47440 13588 47480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 55112 13588 55152 13628
rect 55194 13588 55234 13628
rect 55276 13588 55316 13628
rect 55358 13588 55398 13628
rect 55440 13588 55480 13628
rect 59112 13588 59152 13628
rect 59194 13588 59234 13628
rect 59276 13588 59316 13628
rect 59358 13588 59398 13628
rect 59440 13588 59480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 67112 13588 67152 13628
rect 67194 13588 67234 13628
rect 67276 13588 67316 13628
rect 67358 13588 67398 13628
rect 67440 13588 67480 13628
rect 70060 13420 70100 13460
rect 70924 13420 70964 13460
rect 71308 13420 71348 13460
rect 1612 13336 1652 13376
rect 844 13252 884 13292
rect 1804 13252 1844 13292
rect 69868 13252 69908 13292
rect 70732 13252 70772 13292
rect 71116 13252 71156 13292
rect 70348 13168 70388 13208
rect 70540 13168 70580 13208
rect 652 13000 692 13040
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 8352 12832 8392 12872
rect 8434 12832 8474 12872
rect 8516 12832 8556 12872
rect 8598 12832 8638 12872
rect 8680 12832 8720 12872
rect 12352 12832 12392 12872
rect 12434 12832 12474 12872
rect 12516 12832 12556 12872
rect 12598 12832 12638 12872
rect 12680 12832 12720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 20352 12832 20392 12872
rect 20434 12832 20474 12872
rect 20516 12832 20556 12872
rect 20598 12832 20638 12872
rect 20680 12832 20720 12872
rect 24352 12832 24392 12872
rect 24434 12832 24474 12872
rect 24516 12832 24556 12872
rect 24598 12832 24638 12872
rect 24680 12832 24720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 32352 12832 32392 12872
rect 32434 12832 32474 12872
rect 32516 12832 32556 12872
rect 32598 12832 32638 12872
rect 32680 12832 32720 12872
rect 36352 12832 36392 12872
rect 36434 12832 36474 12872
rect 36516 12832 36556 12872
rect 36598 12832 36638 12872
rect 36680 12832 36720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 44352 12832 44392 12872
rect 44434 12832 44474 12872
rect 44516 12832 44556 12872
rect 44598 12832 44638 12872
rect 44680 12832 44720 12872
rect 48352 12832 48392 12872
rect 48434 12832 48474 12872
rect 48516 12832 48556 12872
rect 48598 12832 48638 12872
rect 48680 12832 48720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 56352 12832 56392 12872
rect 56434 12832 56474 12872
rect 56516 12832 56556 12872
rect 56598 12832 56638 12872
rect 56680 12832 56720 12872
rect 60352 12832 60392 12872
rect 60434 12832 60474 12872
rect 60516 12832 60556 12872
rect 60598 12832 60638 12872
rect 60680 12832 60720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 68352 12832 68392 12872
rect 68434 12832 68474 12872
rect 68516 12832 68556 12872
rect 68598 12832 68638 12872
rect 68680 12832 68720 12872
rect 70540 12580 70580 12620
rect 70924 12580 70964 12620
rect 71212 12580 71252 12620
rect 70444 12496 70484 12536
rect 70828 12496 70868 12536
rect 71116 12496 71156 12536
rect 844 12412 884 12452
rect 1420 12412 1460 12452
rect 652 12328 692 12368
rect 1228 12328 1268 12368
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 7112 12076 7152 12116
rect 7194 12076 7234 12116
rect 7276 12076 7316 12116
rect 7358 12076 7398 12116
rect 7440 12076 7480 12116
rect 11112 12076 11152 12116
rect 11194 12076 11234 12116
rect 11276 12076 11316 12116
rect 11358 12076 11398 12116
rect 11440 12076 11480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 19112 12076 19152 12116
rect 19194 12076 19234 12116
rect 19276 12076 19316 12116
rect 19358 12076 19398 12116
rect 19440 12076 19480 12116
rect 23112 12076 23152 12116
rect 23194 12076 23234 12116
rect 23276 12076 23316 12116
rect 23358 12076 23398 12116
rect 23440 12076 23480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 31112 12076 31152 12116
rect 31194 12076 31234 12116
rect 31276 12076 31316 12116
rect 31358 12076 31398 12116
rect 31440 12076 31480 12116
rect 35112 12076 35152 12116
rect 35194 12076 35234 12116
rect 35276 12076 35316 12116
rect 35358 12076 35398 12116
rect 35440 12076 35480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 43112 12076 43152 12116
rect 43194 12076 43234 12116
rect 43276 12076 43316 12116
rect 43358 12076 43398 12116
rect 43440 12076 43480 12116
rect 47112 12076 47152 12116
rect 47194 12076 47234 12116
rect 47276 12076 47316 12116
rect 47358 12076 47398 12116
rect 47440 12076 47480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 55112 12076 55152 12116
rect 55194 12076 55234 12116
rect 55276 12076 55316 12116
rect 55358 12076 55398 12116
rect 55440 12076 55480 12116
rect 59112 12076 59152 12116
rect 59194 12076 59234 12116
rect 59276 12076 59316 12116
rect 59358 12076 59398 12116
rect 59440 12076 59480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 67112 12076 67152 12116
rect 67194 12076 67234 12116
rect 67276 12076 67316 12116
rect 67358 12076 67398 12116
rect 67440 12076 67480 12116
rect 844 11740 884 11780
rect 652 11488 692 11528
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 8352 11320 8392 11360
rect 8434 11320 8474 11360
rect 8516 11320 8556 11360
rect 8598 11320 8638 11360
rect 8680 11320 8720 11360
rect 12352 11320 12392 11360
rect 12434 11320 12474 11360
rect 12516 11320 12556 11360
rect 12598 11320 12638 11360
rect 12680 11320 12720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 20352 11320 20392 11360
rect 20434 11320 20474 11360
rect 20516 11320 20556 11360
rect 20598 11320 20638 11360
rect 20680 11320 20720 11360
rect 24352 11320 24392 11360
rect 24434 11320 24474 11360
rect 24516 11320 24556 11360
rect 24598 11320 24638 11360
rect 24680 11320 24720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 32352 11320 32392 11360
rect 32434 11320 32474 11360
rect 32516 11320 32556 11360
rect 32598 11320 32638 11360
rect 32680 11320 32720 11360
rect 36352 11320 36392 11360
rect 36434 11320 36474 11360
rect 36516 11320 36556 11360
rect 36598 11320 36638 11360
rect 36680 11320 36720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 44352 11320 44392 11360
rect 44434 11320 44474 11360
rect 44516 11320 44556 11360
rect 44598 11320 44638 11360
rect 44680 11320 44720 11360
rect 48352 11320 48392 11360
rect 48434 11320 48474 11360
rect 48516 11320 48556 11360
rect 48598 11320 48638 11360
rect 48680 11320 48720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 56352 11320 56392 11360
rect 56434 11320 56474 11360
rect 56516 11320 56556 11360
rect 56598 11320 56638 11360
rect 56680 11320 56720 11360
rect 60352 11320 60392 11360
rect 60434 11320 60474 11360
rect 60516 11320 60556 11360
rect 60598 11320 60638 11360
rect 60680 11320 60720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 68352 11320 68392 11360
rect 68434 11320 68474 11360
rect 68516 11320 68556 11360
rect 68598 11320 68638 11360
rect 68680 11320 68720 11360
rect 1228 11152 1268 11192
rect 844 10900 884 10940
rect 1420 10900 1460 10940
rect 652 10732 692 10772
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 7112 10564 7152 10604
rect 7194 10564 7234 10604
rect 7276 10564 7316 10604
rect 7358 10564 7398 10604
rect 7440 10564 7480 10604
rect 11112 10564 11152 10604
rect 11194 10564 11234 10604
rect 11276 10564 11316 10604
rect 11358 10564 11398 10604
rect 11440 10564 11480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 19112 10564 19152 10604
rect 19194 10564 19234 10604
rect 19276 10564 19316 10604
rect 19358 10564 19398 10604
rect 19440 10564 19480 10604
rect 23112 10564 23152 10604
rect 23194 10564 23234 10604
rect 23276 10564 23316 10604
rect 23358 10564 23398 10604
rect 23440 10564 23480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 31112 10564 31152 10604
rect 31194 10564 31234 10604
rect 31276 10564 31316 10604
rect 31358 10564 31398 10604
rect 31440 10564 31480 10604
rect 35112 10564 35152 10604
rect 35194 10564 35234 10604
rect 35276 10564 35316 10604
rect 35358 10564 35398 10604
rect 35440 10564 35480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 43112 10564 43152 10604
rect 43194 10564 43234 10604
rect 43276 10564 43316 10604
rect 43358 10564 43398 10604
rect 43440 10564 43480 10604
rect 47112 10564 47152 10604
rect 47194 10564 47234 10604
rect 47276 10564 47316 10604
rect 47358 10564 47398 10604
rect 47440 10564 47480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 55112 10564 55152 10604
rect 55194 10564 55234 10604
rect 55276 10564 55316 10604
rect 55358 10564 55398 10604
rect 55440 10564 55480 10604
rect 59112 10564 59152 10604
rect 59194 10564 59234 10604
rect 59276 10564 59316 10604
rect 59358 10564 59398 10604
rect 59440 10564 59480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 67112 10564 67152 10604
rect 67194 10564 67234 10604
rect 67276 10564 67316 10604
rect 67358 10564 67398 10604
rect 67440 10564 67480 10604
rect 1420 10396 1460 10436
rect 1036 10312 1076 10352
rect 844 10228 884 10268
rect 1228 10228 1268 10268
rect 1612 10228 1652 10268
rect 652 9976 692 10016
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 8352 9808 8392 9848
rect 8434 9808 8474 9848
rect 8516 9808 8556 9848
rect 8598 9808 8638 9848
rect 8680 9808 8720 9848
rect 12352 9808 12392 9848
rect 12434 9808 12474 9848
rect 12516 9808 12556 9848
rect 12598 9808 12638 9848
rect 12680 9808 12720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 20352 9808 20392 9848
rect 20434 9808 20474 9848
rect 20516 9808 20556 9848
rect 20598 9808 20638 9848
rect 20680 9808 20720 9848
rect 24352 9808 24392 9848
rect 24434 9808 24474 9848
rect 24516 9808 24556 9848
rect 24598 9808 24638 9848
rect 24680 9808 24720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 32352 9808 32392 9848
rect 32434 9808 32474 9848
rect 32516 9808 32556 9848
rect 32598 9808 32638 9848
rect 32680 9808 32720 9848
rect 36352 9808 36392 9848
rect 36434 9808 36474 9848
rect 36516 9808 36556 9848
rect 36598 9808 36638 9848
rect 36680 9808 36720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 44352 9808 44392 9848
rect 44434 9808 44474 9848
rect 44516 9808 44556 9848
rect 44598 9808 44638 9848
rect 44680 9808 44720 9848
rect 48352 9808 48392 9848
rect 48434 9808 48474 9848
rect 48516 9808 48556 9848
rect 48598 9808 48638 9848
rect 48680 9808 48720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 56352 9808 56392 9848
rect 56434 9808 56474 9848
rect 56516 9808 56556 9848
rect 56598 9808 56638 9848
rect 56680 9808 56720 9848
rect 60352 9808 60392 9848
rect 60434 9808 60474 9848
rect 60516 9808 60556 9848
rect 60598 9808 60638 9848
rect 60680 9808 60720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 68352 9808 68392 9848
rect 68434 9808 68474 9848
rect 68516 9808 68556 9848
rect 68598 9808 68638 9848
rect 68680 9808 68720 9848
rect 844 9388 884 9428
rect 652 9220 692 9260
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 7112 9052 7152 9092
rect 7194 9052 7234 9092
rect 7276 9052 7316 9092
rect 7358 9052 7398 9092
rect 7440 9052 7480 9092
rect 11112 9052 11152 9092
rect 11194 9052 11234 9092
rect 11276 9052 11316 9092
rect 11358 9052 11398 9092
rect 11440 9052 11480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 19112 9052 19152 9092
rect 19194 9052 19234 9092
rect 19276 9052 19316 9092
rect 19358 9052 19398 9092
rect 19440 9052 19480 9092
rect 23112 9052 23152 9092
rect 23194 9052 23234 9092
rect 23276 9052 23316 9092
rect 23358 9052 23398 9092
rect 23440 9052 23480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 31112 9052 31152 9092
rect 31194 9052 31234 9092
rect 31276 9052 31316 9092
rect 31358 9052 31398 9092
rect 31440 9052 31480 9092
rect 35112 9052 35152 9092
rect 35194 9052 35234 9092
rect 35276 9052 35316 9092
rect 35358 9052 35398 9092
rect 35440 9052 35480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 43112 9052 43152 9092
rect 43194 9052 43234 9092
rect 43276 9052 43316 9092
rect 43358 9052 43398 9092
rect 43440 9052 43480 9092
rect 47112 9052 47152 9092
rect 47194 9052 47234 9092
rect 47276 9052 47316 9092
rect 47358 9052 47398 9092
rect 47440 9052 47480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 55112 9052 55152 9092
rect 55194 9052 55234 9092
rect 55276 9052 55316 9092
rect 55358 9052 55398 9092
rect 55440 9052 55480 9092
rect 59112 9052 59152 9092
rect 59194 9052 59234 9092
rect 59276 9052 59316 9092
rect 59358 9052 59398 9092
rect 59440 9052 59480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 67112 9052 67152 9092
rect 67194 9052 67234 9092
rect 67276 9052 67316 9092
rect 67358 9052 67398 9092
rect 67440 9052 67480 9092
rect 1132 8800 1172 8840
rect 1516 8800 1556 8840
rect 844 8716 884 8756
rect 1324 8716 1364 8756
rect 1708 8716 1748 8756
rect 2092 8716 2132 8756
rect 70924 8632 70964 8672
rect 71116 8632 71156 8672
rect 652 8464 692 8504
rect 1900 8464 1940 8504
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 8352 8296 8392 8336
rect 8434 8296 8474 8336
rect 8516 8296 8556 8336
rect 8598 8296 8638 8336
rect 8680 8296 8720 8336
rect 12352 8296 12392 8336
rect 12434 8296 12474 8336
rect 12516 8296 12556 8336
rect 12598 8296 12638 8336
rect 12680 8296 12720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 20352 8296 20392 8336
rect 20434 8296 20474 8336
rect 20516 8296 20556 8336
rect 20598 8296 20638 8336
rect 20680 8296 20720 8336
rect 24352 8296 24392 8336
rect 24434 8296 24474 8336
rect 24516 8296 24556 8336
rect 24598 8296 24638 8336
rect 24680 8296 24720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 32352 8296 32392 8336
rect 32434 8296 32474 8336
rect 32516 8296 32556 8336
rect 32598 8296 32638 8336
rect 32680 8296 32720 8336
rect 36352 8296 36392 8336
rect 36434 8296 36474 8336
rect 36516 8296 36556 8336
rect 36598 8296 36638 8336
rect 36680 8296 36720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 44352 8296 44392 8336
rect 44434 8296 44474 8336
rect 44516 8296 44556 8336
rect 44598 8296 44638 8336
rect 44680 8296 44720 8336
rect 48352 8296 48392 8336
rect 48434 8296 48474 8336
rect 48516 8296 48556 8336
rect 48598 8296 48638 8336
rect 48680 8296 48720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 56352 8296 56392 8336
rect 56434 8296 56474 8336
rect 56516 8296 56556 8336
rect 56598 8296 56638 8336
rect 56680 8296 56720 8336
rect 60352 8296 60392 8336
rect 60434 8296 60474 8336
rect 60516 8296 60556 8336
rect 60598 8296 60638 8336
rect 60680 8296 60720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 68352 8296 68392 8336
rect 68434 8296 68474 8336
rect 68516 8296 68556 8336
rect 68598 8296 68638 8336
rect 68680 8296 68720 8336
rect 844 7876 884 7916
rect 70828 7876 70868 7916
rect 71212 7876 71252 7916
rect 71020 7792 71060 7832
rect 71404 7792 71444 7832
rect 652 7708 692 7748
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 7112 7540 7152 7580
rect 7194 7540 7234 7580
rect 7276 7540 7316 7580
rect 7358 7540 7398 7580
rect 7440 7540 7480 7580
rect 11112 7540 11152 7580
rect 11194 7540 11234 7580
rect 11276 7540 11316 7580
rect 11358 7540 11398 7580
rect 11440 7540 11480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 19112 7540 19152 7580
rect 19194 7540 19234 7580
rect 19276 7540 19316 7580
rect 19358 7540 19398 7580
rect 19440 7540 19480 7580
rect 23112 7540 23152 7580
rect 23194 7540 23234 7580
rect 23276 7540 23316 7580
rect 23358 7540 23398 7580
rect 23440 7540 23480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 31112 7540 31152 7580
rect 31194 7540 31234 7580
rect 31276 7540 31316 7580
rect 31358 7540 31398 7580
rect 31440 7540 31480 7580
rect 35112 7540 35152 7580
rect 35194 7540 35234 7580
rect 35276 7540 35316 7580
rect 35358 7540 35398 7580
rect 35440 7540 35480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 43112 7540 43152 7580
rect 43194 7540 43234 7580
rect 43276 7540 43316 7580
rect 43358 7540 43398 7580
rect 43440 7540 43480 7580
rect 47112 7540 47152 7580
rect 47194 7540 47234 7580
rect 47276 7540 47316 7580
rect 47358 7540 47398 7580
rect 47440 7540 47480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 55112 7540 55152 7580
rect 55194 7540 55234 7580
rect 55276 7540 55316 7580
rect 55358 7540 55398 7580
rect 55440 7540 55480 7580
rect 59112 7540 59152 7580
rect 59194 7540 59234 7580
rect 59276 7540 59316 7580
rect 59358 7540 59398 7580
rect 59440 7540 59480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 67112 7540 67152 7580
rect 67194 7540 67234 7580
rect 67276 7540 67316 7580
rect 67358 7540 67398 7580
rect 67440 7540 67480 7580
rect 1516 7372 1556 7412
rect 71404 7372 71444 7412
rect 72172 7372 72212 7412
rect 72556 7372 72596 7412
rect 73324 7372 73364 7412
rect 73708 7372 73748 7412
rect 75148 7372 75188 7412
rect 75916 7372 75956 7412
rect 76204 7372 76244 7412
rect 76780 7372 76820 7412
rect 77836 7372 77876 7412
rect 78124 7372 78164 7412
rect 78412 7372 78452 7412
rect 79276 7372 79316 7412
rect 79468 7372 79508 7412
rect 81100 7372 81140 7412
rect 82348 7372 82388 7412
rect 82540 7372 82580 7412
rect 82828 7372 82868 7412
rect 83980 7372 84020 7412
rect 84172 7372 84212 7412
rect 84460 7372 84500 7412
rect 85324 7372 85364 7412
rect 85516 7372 85556 7412
rect 85804 7372 85844 7412
rect 87436 7372 87476 7412
rect 87724 7372 87764 7412
rect 88780 7372 88820 7412
rect 88972 7372 89012 7412
rect 89644 7372 89684 7412
rect 90220 7372 90260 7412
rect 90508 7372 90548 7412
rect 91180 7372 91220 7412
rect 91756 7372 91796 7412
rect 93484 7372 93524 7412
rect 93772 7372 93812 7412
rect 96460 7372 96500 7412
rect 97804 7372 97844 7412
rect 98476 7372 98516 7412
rect 99244 7372 99284 7412
rect 73132 7288 73172 7328
rect 77644 7288 77684 7328
rect 80140 7288 80180 7328
rect 80524 7288 80564 7328
rect 83596 7288 83636 7328
rect 86860 7288 86900 7328
rect 88396 7288 88436 7328
rect 90028 7288 90068 7328
rect 91564 7288 91604 7328
rect 95980 7288 96020 7328
rect 98092 7288 98132 7328
rect 844 7204 884 7244
rect 1708 7204 1748 7244
rect 72364 7204 72404 7244
rect 72940 7204 72980 7244
rect 74284 7204 74324 7244
rect 74668 7204 74708 7244
rect 74860 7204 74900 7244
rect 75532 7204 75572 7244
rect 76492 7204 76532 7244
rect 77356 7204 77396 7244
rect 78796 7204 78836 7244
rect 79756 7204 79796 7244
rect 80332 7204 80372 7244
rect 81580 7204 81620 7244
rect 83212 7204 83252 7244
rect 84844 7204 84884 7244
rect 86284 7204 86324 7244
rect 86668 7204 86708 7244
rect 88204 7204 88244 7244
rect 89260 7204 89300 7244
rect 90796 7204 90836 7244
rect 92332 7204 92372 7244
rect 92716 7204 92756 7244
rect 92908 7204 92948 7244
rect 94252 7204 94292 7244
rect 95212 7204 95252 7244
rect 95596 7204 95636 7244
rect 96172 7204 96212 7244
rect 96844 7204 96884 7244
rect 98668 7204 98708 7244
rect 71308 7120 71348 7160
rect 72076 7120 72116 7160
rect 73433 7109 73473 7149
rect 73612 7120 73652 7160
rect 74956 7120 74996 7160
rect 75244 7120 75284 7160
rect 76012 7120 76052 7160
rect 76300 7120 76340 7160
rect 76588 7120 76628 7160
rect 76876 7120 76916 7160
rect 77548 7120 77588 7160
rect 77932 7120 77972 7160
rect 78220 7120 78260 7160
rect 78508 7120 78548 7160
rect 79180 7120 79220 7160
rect 79564 7120 79604 7160
rect 80620 7120 80660 7160
rect 80812 7120 80852 7160
rect 81196 7120 81236 7160
rect 82060 7120 82100 7160
rect 82252 7120 82292 7160
rect 82636 7120 82676 7160
rect 82924 7120 82964 7160
rect 83692 7120 83732 7160
rect 83884 7120 83924 7160
rect 84268 7120 84308 7160
rect 84556 7120 84596 7160
rect 85228 7120 85268 7160
rect 85612 7120 85652 7160
rect 85900 7120 85940 7160
rect 86956 7120 86996 7160
rect 87148 7120 87188 7160
rect 87532 7120 87572 7160
rect 87820 7120 87860 7160
rect 88492 7120 88532 7160
rect 88684 7120 88724 7160
rect 89068 7120 89108 7160
rect 89740 7120 89780 7160
rect 89932 7120 89972 7160
rect 90316 7120 90356 7160
rect 90604 7120 90644 7160
rect 91276 7120 91316 7160
rect 91468 7120 91508 7160
rect 91852 7120 91892 7160
rect 93004 7120 93044 7160
rect 93196 7120 93236 7160
rect 93580 7120 93620 7160
rect 93868 7120 93908 7160
rect 94540 7120 94580 7160
rect 94732 7120 94772 7160
rect 94828 7120 94868 7160
rect 95692 7120 95732 7160
rect 95884 7120 95924 7160
rect 96268 7120 96308 7160
rect 96556 7120 96596 7160
rect 97228 7120 97268 7160
rect 97324 7133 97364 7173
rect 97516 7120 97556 7160
rect 97900 7120 97940 7160
rect 98188 7120 98228 7160
rect 98956 7120 98996 7160
rect 99148 7120 99188 7160
rect 87244 7036 87284 7076
rect 94444 7036 94484 7076
rect 98860 7036 98900 7076
rect 652 6952 692 6992
rect 74092 6952 74132 6992
rect 74476 6952 74516 6992
rect 75724 6952 75764 6992
rect 77164 6952 77204 6992
rect 78988 6952 79028 6992
rect 79948 6952 79988 6992
rect 80908 6952 80948 6992
rect 81772 6952 81812 6992
rect 81964 6952 82004 6992
rect 83404 6952 83444 6992
rect 85036 6952 85076 6992
rect 86092 6952 86132 6992
rect 86476 6952 86516 6992
rect 88012 6952 88052 6992
rect 89452 6952 89492 6992
rect 90988 6952 91028 6992
rect 92140 6952 92180 6992
rect 92524 6952 92564 6992
rect 93292 6952 93332 6992
rect 94060 6952 94100 6992
rect 95404 6952 95444 6992
rect 97036 6952 97076 6992
rect 97612 6952 97652 6992
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 8352 6784 8392 6824
rect 8434 6784 8474 6824
rect 8516 6784 8556 6824
rect 8598 6784 8638 6824
rect 8680 6784 8720 6824
rect 12352 6784 12392 6824
rect 12434 6784 12474 6824
rect 12516 6784 12556 6824
rect 12598 6784 12638 6824
rect 12680 6784 12720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 20352 6784 20392 6824
rect 20434 6784 20474 6824
rect 20516 6784 20556 6824
rect 20598 6784 20638 6824
rect 20680 6784 20720 6824
rect 24352 6784 24392 6824
rect 24434 6784 24474 6824
rect 24516 6784 24556 6824
rect 24598 6784 24638 6824
rect 24680 6784 24720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 32352 6784 32392 6824
rect 32434 6784 32474 6824
rect 32516 6784 32556 6824
rect 32598 6784 32638 6824
rect 32680 6784 32720 6824
rect 36352 6784 36392 6824
rect 36434 6784 36474 6824
rect 36516 6784 36556 6824
rect 36598 6784 36638 6824
rect 36680 6784 36720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 44352 6784 44392 6824
rect 44434 6784 44474 6824
rect 44516 6784 44556 6824
rect 44598 6784 44638 6824
rect 44680 6784 44720 6824
rect 48352 6784 48392 6824
rect 48434 6784 48474 6824
rect 48516 6784 48556 6824
rect 48598 6784 48638 6824
rect 48680 6784 48720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 56352 6784 56392 6824
rect 56434 6784 56474 6824
rect 56516 6784 56556 6824
rect 56598 6784 56638 6824
rect 56680 6784 56720 6824
rect 60352 6784 60392 6824
rect 60434 6784 60474 6824
rect 60516 6784 60556 6824
rect 60598 6784 60638 6824
rect 60680 6784 60720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 68352 6784 68392 6824
rect 68434 6784 68474 6824
rect 68516 6784 68556 6824
rect 68598 6784 68638 6824
rect 68680 6784 68720 6824
rect 1708 6616 1748 6656
rect 73708 6616 73748 6656
rect 74188 6616 74228 6656
rect 74572 6616 74612 6656
rect 75052 6616 75092 6656
rect 75436 6616 75476 6656
rect 75820 6616 75860 6656
rect 76204 6616 76244 6656
rect 76684 6616 76724 6656
rect 77068 6616 77108 6656
rect 77452 6616 77492 6656
rect 77836 6616 77876 6656
rect 78316 6616 78356 6656
rect 78700 6616 78740 6656
rect 79084 6616 79124 6656
rect 79468 6616 79508 6656
rect 79948 6616 79988 6656
rect 80332 6616 80372 6656
rect 80716 6616 80756 6656
rect 80908 6616 80948 6656
rect 81484 6616 81524 6656
rect 81868 6616 81908 6656
rect 82252 6616 82292 6656
rect 82732 6616 82772 6656
rect 83116 6616 83156 6656
rect 83308 6616 83348 6656
rect 83884 6616 83924 6656
rect 84268 6616 84308 6656
rect 84652 6616 84692 6656
rect 85036 6616 85076 6656
rect 85516 6616 85556 6656
rect 85900 6616 85940 6656
rect 86284 6616 86324 6656
rect 86668 6616 86708 6656
rect 87052 6616 87092 6656
rect 87532 6616 87572 6656
rect 87724 6616 87764 6656
rect 88300 6616 88340 6656
rect 88684 6616 88724 6656
rect 89068 6616 89108 6656
rect 89452 6616 89492 6656
rect 89932 6616 89972 6656
rect 90316 6616 90356 6656
rect 90700 6616 90740 6656
rect 91084 6616 91124 6656
rect 91468 6616 91508 6656
rect 92332 6616 92372 6656
rect 92716 6616 92756 6656
rect 93100 6616 93140 6656
rect 93580 6616 93620 6656
rect 93772 6616 93812 6656
rect 94348 6616 94388 6656
rect 94732 6616 94772 6656
rect 95116 6616 95156 6656
rect 95596 6616 95636 6656
rect 95980 6616 96020 6656
rect 96364 6616 96404 6656
rect 96748 6616 96788 6656
rect 97036 6616 97076 6656
rect 97516 6616 97556 6656
rect 97900 6616 97940 6656
rect 98380 6616 98420 6656
rect 73324 6532 73364 6572
rect 73228 6448 73268 6488
rect 81004 6448 81044 6488
rect 83404 6448 83444 6488
rect 98476 6448 98516 6488
rect 1516 6364 1556 6404
rect 1900 6364 1940 6404
rect 73516 6364 73556 6404
rect 73996 6364 74036 6404
rect 74380 6364 74420 6404
rect 74860 6364 74900 6404
rect 75244 6364 75284 6404
rect 75628 6364 75668 6404
rect 76012 6364 76052 6404
rect 76492 6364 76532 6404
rect 76876 6364 76916 6404
rect 77260 6364 77300 6404
rect 77644 6364 77684 6404
rect 78124 6364 78164 6404
rect 78508 6364 78548 6404
rect 78892 6364 78932 6404
rect 79276 6364 79316 6404
rect 79756 6364 79796 6404
rect 80140 6364 80180 6404
rect 80524 6364 80564 6404
rect 81292 6364 81332 6404
rect 81676 6364 81716 6404
rect 82060 6364 82100 6404
rect 82540 6364 82580 6404
rect 82924 6364 82964 6404
rect 83692 6364 83732 6404
rect 84076 6364 84116 6404
rect 84460 6364 84500 6404
rect 84844 6364 84884 6404
rect 85324 6364 85364 6404
rect 85708 6364 85748 6404
rect 86092 6364 86132 6404
rect 86476 6364 86516 6404
rect 86860 6364 86900 6404
rect 87340 6364 87380 6404
rect 87916 6364 87956 6404
rect 88108 6364 88148 6404
rect 88492 6364 88532 6404
rect 88876 6364 88916 6404
rect 89260 6364 89300 6404
rect 89740 6364 89780 6404
rect 90124 6364 90164 6404
rect 90508 6364 90548 6404
rect 90892 6364 90932 6404
rect 91276 6364 91316 6404
rect 91756 6364 91796 6404
rect 92140 6364 92180 6404
rect 92524 6364 92564 6404
rect 92908 6364 92948 6404
rect 93388 6364 93428 6404
rect 93964 6364 94004 6404
rect 94156 6364 94196 6404
rect 94540 6364 94580 6404
rect 94924 6364 94964 6404
rect 95404 6364 95444 6404
rect 95788 6364 95828 6404
rect 96172 6364 96212 6404
rect 96556 6364 96596 6404
rect 97228 6364 97268 6404
rect 97708 6364 97748 6404
rect 98092 6364 98132 6404
rect 1324 6280 1364 6320
rect 91948 6280 91988 6320
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 7112 6028 7152 6068
rect 7194 6028 7234 6068
rect 7276 6028 7316 6068
rect 7358 6028 7398 6068
rect 7440 6028 7480 6068
rect 11112 6028 11152 6068
rect 11194 6028 11234 6068
rect 11276 6028 11316 6068
rect 11358 6028 11398 6068
rect 11440 6028 11480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 19112 6028 19152 6068
rect 19194 6028 19234 6068
rect 19276 6028 19316 6068
rect 19358 6028 19398 6068
rect 19440 6028 19480 6068
rect 23112 6028 23152 6068
rect 23194 6028 23234 6068
rect 23276 6028 23316 6068
rect 23358 6028 23398 6068
rect 23440 6028 23480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 31112 6028 31152 6068
rect 31194 6028 31234 6068
rect 31276 6028 31316 6068
rect 31358 6028 31398 6068
rect 31440 6028 31480 6068
rect 35112 6028 35152 6068
rect 35194 6028 35234 6068
rect 35276 6028 35316 6068
rect 35358 6028 35398 6068
rect 35440 6028 35480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 43112 6028 43152 6068
rect 43194 6028 43234 6068
rect 43276 6028 43316 6068
rect 43358 6028 43398 6068
rect 43440 6028 43480 6068
rect 47112 6028 47152 6068
rect 47194 6028 47234 6068
rect 47276 6028 47316 6068
rect 47358 6028 47398 6068
rect 47440 6028 47480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 55112 6028 55152 6068
rect 55194 6028 55234 6068
rect 55276 6028 55316 6068
rect 55358 6028 55398 6068
rect 55440 6028 55480 6068
rect 59112 6028 59152 6068
rect 59194 6028 59234 6068
rect 59276 6028 59316 6068
rect 59358 6028 59398 6068
rect 59440 6028 59480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 67112 6028 67152 6068
rect 67194 6028 67234 6068
rect 67276 6028 67316 6068
rect 67358 6028 67398 6068
rect 67440 6028 67480 6068
rect 81100 5860 81140 5900
rect 83500 5860 83540 5900
rect 91180 5860 91220 5900
rect 94060 5860 94100 5900
rect 844 5692 884 5732
rect 80908 5692 80948 5732
rect 83308 5692 83348 5732
rect 91084 5608 91124 5648
rect 93964 5608 94004 5648
rect 652 5440 692 5480
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 8352 5272 8392 5312
rect 8434 5272 8474 5312
rect 8516 5272 8556 5312
rect 8598 5272 8638 5312
rect 8680 5272 8720 5312
rect 12352 5272 12392 5312
rect 12434 5272 12474 5312
rect 12516 5272 12556 5312
rect 12598 5272 12638 5312
rect 12680 5272 12720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 20352 5272 20392 5312
rect 20434 5272 20474 5312
rect 20516 5272 20556 5312
rect 20598 5272 20638 5312
rect 20680 5272 20720 5312
rect 24352 5272 24392 5312
rect 24434 5272 24474 5312
rect 24516 5272 24556 5312
rect 24598 5272 24638 5312
rect 24680 5272 24720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 32352 5272 32392 5312
rect 32434 5272 32474 5312
rect 32516 5272 32556 5312
rect 32598 5272 32638 5312
rect 32680 5272 32720 5312
rect 36352 5272 36392 5312
rect 36434 5272 36474 5312
rect 36516 5272 36556 5312
rect 36598 5272 36638 5312
rect 36680 5272 36720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 44352 5272 44392 5312
rect 44434 5272 44474 5312
rect 44516 5272 44556 5312
rect 44598 5272 44638 5312
rect 44680 5272 44720 5312
rect 48352 5272 48392 5312
rect 48434 5272 48474 5312
rect 48516 5272 48556 5312
rect 48598 5272 48638 5312
rect 48680 5272 48720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 56352 5272 56392 5312
rect 56434 5272 56474 5312
rect 56516 5272 56556 5312
rect 56598 5272 56638 5312
rect 56680 5272 56720 5312
rect 60352 5272 60392 5312
rect 60434 5272 60474 5312
rect 60516 5272 60556 5312
rect 60598 5272 60638 5312
rect 60680 5272 60720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 68352 5272 68392 5312
rect 68434 5272 68474 5312
rect 68516 5272 68556 5312
rect 68598 5272 68638 5312
rect 68680 5272 68720 5312
rect 72352 5272 72392 5312
rect 72434 5272 72474 5312
rect 72516 5272 72556 5312
rect 72598 5272 72638 5312
rect 72680 5272 72720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 80352 5272 80392 5312
rect 80434 5272 80474 5312
rect 80516 5272 80556 5312
rect 80598 5272 80638 5312
rect 80680 5272 80720 5312
rect 84352 5272 84392 5312
rect 84434 5272 84474 5312
rect 84516 5272 84556 5312
rect 84598 5272 84638 5312
rect 84680 5272 84720 5312
rect 88352 5272 88392 5312
rect 88434 5272 88474 5312
rect 88516 5272 88556 5312
rect 88598 5272 88638 5312
rect 88680 5272 88720 5312
rect 92352 5272 92392 5312
rect 92434 5272 92474 5312
rect 92516 5272 92556 5312
rect 92598 5272 92638 5312
rect 92680 5272 92720 5312
rect 96352 5272 96392 5312
rect 96434 5272 96474 5312
rect 96516 5272 96556 5312
rect 96598 5272 96638 5312
rect 96680 5272 96720 5312
rect 1036 4852 1076 4892
rect 1420 4852 1460 4892
rect 1804 4852 1844 4892
rect 2188 4852 2228 4892
rect 844 4684 884 4724
rect 1228 4684 1268 4724
rect 1612 4684 1652 4724
rect 1996 4684 2036 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 7112 4516 7152 4556
rect 7194 4516 7234 4556
rect 7276 4516 7316 4556
rect 7358 4516 7398 4556
rect 7440 4516 7480 4556
rect 11112 4516 11152 4556
rect 11194 4516 11234 4556
rect 11276 4516 11316 4556
rect 11358 4516 11398 4556
rect 11440 4516 11480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 19112 4516 19152 4556
rect 19194 4516 19234 4556
rect 19276 4516 19316 4556
rect 19358 4516 19398 4556
rect 19440 4516 19480 4556
rect 23112 4516 23152 4556
rect 23194 4516 23234 4556
rect 23276 4516 23316 4556
rect 23358 4516 23398 4556
rect 23440 4516 23480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 31112 4516 31152 4556
rect 31194 4516 31234 4556
rect 31276 4516 31316 4556
rect 31358 4516 31398 4556
rect 31440 4516 31480 4556
rect 35112 4516 35152 4556
rect 35194 4516 35234 4556
rect 35276 4516 35316 4556
rect 35358 4516 35398 4556
rect 35440 4516 35480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 43112 4516 43152 4556
rect 43194 4516 43234 4556
rect 43276 4516 43316 4556
rect 43358 4516 43398 4556
rect 43440 4516 43480 4556
rect 47112 4516 47152 4556
rect 47194 4516 47234 4556
rect 47276 4516 47316 4556
rect 47358 4516 47398 4556
rect 47440 4516 47480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 55112 4516 55152 4556
rect 55194 4516 55234 4556
rect 55276 4516 55316 4556
rect 55358 4516 55398 4556
rect 55440 4516 55480 4556
rect 59112 4516 59152 4556
rect 59194 4516 59234 4556
rect 59276 4516 59316 4556
rect 59358 4516 59398 4556
rect 59440 4516 59480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 67112 4516 67152 4556
rect 67194 4516 67234 4556
rect 67276 4516 67316 4556
rect 67358 4516 67398 4556
rect 67440 4516 67480 4556
rect 71112 4516 71152 4556
rect 71194 4516 71234 4556
rect 71276 4516 71316 4556
rect 71358 4516 71398 4556
rect 71440 4516 71480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 79112 4516 79152 4556
rect 79194 4516 79234 4556
rect 79276 4516 79316 4556
rect 79358 4516 79398 4556
rect 79440 4516 79480 4556
rect 83112 4516 83152 4556
rect 83194 4516 83234 4556
rect 83276 4516 83316 4556
rect 83358 4516 83398 4556
rect 83440 4516 83480 4556
rect 87112 4516 87152 4556
rect 87194 4516 87234 4556
rect 87276 4516 87316 4556
rect 87358 4516 87398 4556
rect 87440 4516 87480 4556
rect 91112 4516 91152 4556
rect 91194 4516 91234 4556
rect 91276 4516 91316 4556
rect 91358 4516 91398 4556
rect 91440 4516 91480 4556
rect 95112 4516 95152 4556
rect 95194 4516 95234 4556
rect 95276 4516 95316 4556
rect 95358 4516 95398 4556
rect 95440 4516 95480 4556
rect 99112 4516 99152 4556
rect 99194 4516 99234 4556
rect 99276 4516 99316 4556
rect 99358 4516 99398 4556
rect 99440 4516 99480 4556
rect 652 4348 692 4388
rect 844 4180 884 4220
rect 1228 4180 1268 4220
rect 1036 3928 1076 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 8352 3760 8392 3800
rect 8434 3760 8474 3800
rect 8516 3760 8556 3800
rect 8598 3760 8638 3800
rect 8680 3760 8720 3800
rect 12352 3760 12392 3800
rect 12434 3760 12474 3800
rect 12516 3760 12556 3800
rect 12598 3760 12638 3800
rect 12680 3760 12720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 20352 3760 20392 3800
rect 20434 3760 20474 3800
rect 20516 3760 20556 3800
rect 20598 3760 20638 3800
rect 20680 3760 20720 3800
rect 24352 3760 24392 3800
rect 24434 3760 24474 3800
rect 24516 3760 24556 3800
rect 24598 3760 24638 3800
rect 24680 3760 24720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 32352 3760 32392 3800
rect 32434 3760 32474 3800
rect 32516 3760 32556 3800
rect 32598 3760 32638 3800
rect 32680 3760 32720 3800
rect 36352 3760 36392 3800
rect 36434 3760 36474 3800
rect 36516 3760 36556 3800
rect 36598 3760 36638 3800
rect 36680 3760 36720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 44352 3760 44392 3800
rect 44434 3760 44474 3800
rect 44516 3760 44556 3800
rect 44598 3760 44638 3800
rect 44680 3760 44720 3800
rect 48352 3760 48392 3800
rect 48434 3760 48474 3800
rect 48516 3760 48556 3800
rect 48598 3760 48638 3800
rect 48680 3760 48720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 56352 3760 56392 3800
rect 56434 3760 56474 3800
rect 56516 3760 56556 3800
rect 56598 3760 56638 3800
rect 56680 3760 56720 3800
rect 60352 3760 60392 3800
rect 60434 3760 60474 3800
rect 60516 3760 60556 3800
rect 60598 3760 60638 3800
rect 60680 3760 60720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 68352 3760 68392 3800
rect 68434 3760 68474 3800
rect 68516 3760 68556 3800
rect 68598 3760 68638 3800
rect 68680 3760 68720 3800
rect 72352 3760 72392 3800
rect 72434 3760 72474 3800
rect 72516 3760 72556 3800
rect 72598 3760 72638 3800
rect 72680 3760 72720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 80352 3760 80392 3800
rect 80434 3760 80474 3800
rect 80516 3760 80556 3800
rect 80598 3760 80638 3800
rect 80680 3760 80720 3800
rect 84352 3760 84392 3800
rect 84434 3760 84474 3800
rect 84516 3760 84556 3800
rect 84598 3760 84638 3800
rect 84680 3760 84720 3800
rect 88352 3760 88392 3800
rect 88434 3760 88474 3800
rect 88516 3760 88556 3800
rect 88598 3760 88638 3800
rect 88680 3760 88720 3800
rect 92352 3760 92392 3800
rect 92434 3760 92474 3800
rect 92516 3760 92556 3800
rect 92598 3760 92638 3800
rect 92680 3760 92720 3800
rect 96352 3760 96392 3800
rect 96434 3760 96474 3800
rect 96516 3760 96556 3800
rect 96598 3760 96638 3800
rect 96680 3760 96720 3800
rect 844 3340 884 3380
rect 652 3172 692 3212
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 7112 3004 7152 3044
rect 7194 3004 7234 3044
rect 7276 3004 7316 3044
rect 7358 3004 7398 3044
rect 7440 3004 7480 3044
rect 11112 3004 11152 3044
rect 11194 3004 11234 3044
rect 11276 3004 11316 3044
rect 11358 3004 11398 3044
rect 11440 3004 11480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 19112 3004 19152 3044
rect 19194 3004 19234 3044
rect 19276 3004 19316 3044
rect 19358 3004 19398 3044
rect 19440 3004 19480 3044
rect 23112 3004 23152 3044
rect 23194 3004 23234 3044
rect 23276 3004 23316 3044
rect 23358 3004 23398 3044
rect 23440 3004 23480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 31112 3004 31152 3044
rect 31194 3004 31234 3044
rect 31276 3004 31316 3044
rect 31358 3004 31398 3044
rect 31440 3004 31480 3044
rect 35112 3004 35152 3044
rect 35194 3004 35234 3044
rect 35276 3004 35316 3044
rect 35358 3004 35398 3044
rect 35440 3004 35480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 43112 3004 43152 3044
rect 43194 3004 43234 3044
rect 43276 3004 43316 3044
rect 43358 3004 43398 3044
rect 43440 3004 43480 3044
rect 47112 3004 47152 3044
rect 47194 3004 47234 3044
rect 47276 3004 47316 3044
rect 47358 3004 47398 3044
rect 47440 3004 47480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 55112 3004 55152 3044
rect 55194 3004 55234 3044
rect 55276 3004 55316 3044
rect 55358 3004 55398 3044
rect 55440 3004 55480 3044
rect 59112 3004 59152 3044
rect 59194 3004 59234 3044
rect 59276 3004 59316 3044
rect 59358 3004 59398 3044
rect 59440 3004 59480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 67112 3004 67152 3044
rect 67194 3004 67234 3044
rect 67276 3004 67316 3044
rect 67358 3004 67398 3044
rect 67440 3004 67480 3044
rect 71112 3004 71152 3044
rect 71194 3004 71234 3044
rect 71276 3004 71316 3044
rect 71358 3004 71398 3044
rect 71440 3004 71480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 79112 3004 79152 3044
rect 79194 3004 79234 3044
rect 79276 3004 79316 3044
rect 79358 3004 79398 3044
rect 79440 3004 79480 3044
rect 83112 3004 83152 3044
rect 83194 3004 83234 3044
rect 83276 3004 83316 3044
rect 83358 3004 83398 3044
rect 83440 3004 83480 3044
rect 87112 3004 87152 3044
rect 87194 3004 87234 3044
rect 87276 3004 87316 3044
rect 87358 3004 87398 3044
rect 87440 3004 87480 3044
rect 91112 3004 91152 3044
rect 91194 3004 91234 3044
rect 91276 3004 91316 3044
rect 91358 3004 91398 3044
rect 91440 3004 91480 3044
rect 95112 3004 95152 3044
rect 95194 3004 95234 3044
rect 95276 3004 95316 3044
rect 95358 3004 95398 3044
rect 95440 3004 95480 3044
rect 99112 3004 99152 3044
rect 99194 3004 99234 3044
rect 99276 3004 99316 3044
rect 99358 3004 99398 3044
rect 99440 3004 99480 3044
rect 844 2668 884 2708
rect 652 2416 692 2456
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 8352 2248 8392 2288
rect 8434 2248 8474 2288
rect 8516 2248 8556 2288
rect 8598 2248 8638 2288
rect 8680 2248 8720 2288
rect 12352 2248 12392 2288
rect 12434 2248 12474 2288
rect 12516 2248 12556 2288
rect 12598 2248 12638 2288
rect 12680 2248 12720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 20352 2248 20392 2288
rect 20434 2248 20474 2288
rect 20516 2248 20556 2288
rect 20598 2248 20638 2288
rect 20680 2248 20720 2288
rect 24352 2248 24392 2288
rect 24434 2248 24474 2288
rect 24516 2248 24556 2288
rect 24598 2248 24638 2288
rect 24680 2248 24720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 32352 2248 32392 2288
rect 32434 2248 32474 2288
rect 32516 2248 32556 2288
rect 32598 2248 32638 2288
rect 32680 2248 32720 2288
rect 36352 2248 36392 2288
rect 36434 2248 36474 2288
rect 36516 2248 36556 2288
rect 36598 2248 36638 2288
rect 36680 2248 36720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 44352 2248 44392 2288
rect 44434 2248 44474 2288
rect 44516 2248 44556 2288
rect 44598 2248 44638 2288
rect 44680 2248 44720 2288
rect 48352 2248 48392 2288
rect 48434 2248 48474 2288
rect 48516 2248 48556 2288
rect 48598 2248 48638 2288
rect 48680 2248 48720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 56352 2248 56392 2288
rect 56434 2248 56474 2288
rect 56516 2248 56556 2288
rect 56598 2248 56638 2288
rect 56680 2248 56720 2288
rect 60352 2248 60392 2288
rect 60434 2248 60474 2288
rect 60516 2248 60556 2288
rect 60598 2248 60638 2288
rect 60680 2248 60720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 68352 2248 68392 2288
rect 68434 2248 68474 2288
rect 68516 2248 68556 2288
rect 68598 2248 68638 2288
rect 68680 2248 68720 2288
rect 72352 2248 72392 2288
rect 72434 2248 72474 2288
rect 72516 2248 72556 2288
rect 72598 2248 72638 2288
rect 72680 2248 72720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 80352 2248 80392 2288
rect 80434 2248 80474 2288
rect 80516 2248 80556 2288
rect 80598 2248 80638 2288
rect 80680 2248 80720 2288
rect 84352 2248 84392 2288
rect 84434 2248 84474 2288
rect 84516 2248 84556 2288
rect 84598 2248 84638 2288
rect 84680 2248 84720 2288
rect 88352 2248 88392 2288
rect 88434 2248 88474 2288
rect 88516 2248 88556 2288
rect 88598 2248 88638 2288
rect 88680 2248 88720 2288
rect 92352 2248 92392 2288
rect 92434 2248 92474 2288
rect 92516 2248 92556 2288
rect 92598 2248 92638 2288
rect 92680 2248 92720 2288
rect 96352 2248 96392 2288
rect 96434 2248 96474 2288
rect 96516 2248 96556 2288
rect 96598 2248 96638 2288
rect 96680 2248 96720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 7112 1492 7152 1532
rect 7194 1492 7234 1532
rect 7276 1492 7316 1532
rect 7358 1492 7398 1532
rect 7440 1492 7480 1532
rect 11112 1492 11152 1532
rect 11194 1492 11234 1532
rect 11276 1492 11316 1532
rect 11358 1492 11398 1532
rect 11440 1492 11480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 19112 1492 19152 1532
rect 19194 1492 19234 1532
rect 19276 1492 19316 1532
rect 19358 1492 19398 1532
rect 19440 1492 19480 1532
rect 23112 1492 23152 1532
rect 23194 1492 23234 1532
rect 23276 1492 23316 1532
rect 23358 1492 23398 1532
rect 23440 1492 23480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 31112 1492 31152 1532
rect 31194 1492 31234 1532
rect 31276 1492 31316 1532
rect 31358 1492 31398 1532
rect 31440 1492 31480 1532
rect 35112 1492 35152 1532
rect 35194 1492 35234 1532
rect 35276 1492 35316 1532
rect 35358 1492 35398 1532
rect 35440 1492 35480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 43112 1492 43152 1532
rect 43194 1492 43234 1532
rect 43276 1492 43316 1532
rect 43358 1492 43398 1532
rect 43440 1492 43480 1532
rect 47112 1492 47152 1532
rect 47194 1492 47234 1532
rect 47276 1492 47316 1532
rect 47358 1492 47398 1532
rect 47440 1492 47480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 55112 1492 55152 1532
rect 55194 1492 55234 1532
rect 55276 1492 55316 1532
rect 55358 1492 55398 1532
rect 55440 1492 55480 1532
rect 59112 1492 59152 1532
rect 59194 1492 59234 1532
rect 59276 1492 59316 1532
rect 59358 1492 59398 1532
rect 59440 1492 59480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 67112 1492 67152 1532
rect 67194 1492 67234 1532
rect 67276 1492 67316 1532
rect 67358 1492 67398 1532
rect 67440 1492 67480 1532
rect 71112 1492 71152 1532
rect 71194 1492 71234 1532
rect 71276 1492 71316 1532
rect 71358 1492 71398 1532
rect 71440 1492 71480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 79112 1492 79152 1532
rect 79194 1492 79234 1532
rect 79276 1492 79316 1532
rect 79358 1492 79398 1532
rect 79440 1492 79480 1532
rect 83112 1492 83152 1532
rect 83194 1492 83234 1532
rect 83276 1492 83316 1532
rect 83358 1492 83398 1532
rect 83440 1492 83480 1532
rect 87112 1492 87152 1532
rect 87194 1492 87234 1532
rect 87276 1492 87316 1532
rect 87358 1492 87398 1532
rect 87440 1492 87480 1532
rect 91112 1492 91152 1532
rect 91194 1492 91234 1532
rect 91276 1492 91316 1532
rect 91358 1492 91398 1532
rect 91440 1492 91480 1532
rect 95112 1492 95152 1532
rect 95194 1492 95234 1532
rect 95276 1492 95316 1532
rect 95358 1492 95398 1532
rect 95440 1492 95480 1532
rect 99112 1492 99152 1532
rect 99194 1492 99234 1532
rect 99276 1492 99316 1532
rect 99358 1492 99398 1532
rect 99440 1492 99480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 8352 736 8392 776
rect 8434 736 8474 776
rect 8516 736 8556 776
rect 8598 736 8638 776
rect 8680 736 8720 776
rect 12352 736 12392 776
rect 12434 736 12474 776
rect 12516 736 12556 776
rect 12598 736 12638 776
rect 12680 736 12720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 20352 736 20392 776
rect 20434 736 20474 776
rect 20516 736 20556 776
rect 20598 736 20638 776
rect 20680 736 20720 776
rect 24352 736 24392 776
rect 24434 736 24474 776
rect 24516 736 24556 776
rect 24598 736 24638 776
rect 24680 736 24720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 32352 736 32392 776
rect 32434 736 32474 776
rect 32516 736 32556 776
rect 32598 736 32638 776
rect 32680 736 32720 776
rect 36352 736 36392 776
rect 36434 736 36474 776
rect 36516 736 36556 776
rect 36598 736 36638 776
rect 36680 736 36720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 44352 736 44392 776
rect 44434 736 44474 776
rect 44516 736 44556 776
rect 44598 736 44638 776
rect 44680 736 44720 776
rect 48352 736 48392 776
rect 48434 736 48474 776
rect 48516 736 48556 776
rect 48598 736 48638 776
rect 48680 736 48720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 56352 736 56392 776
rect 56434 736 56474 776
rect 56516 736 56556 776
rect 56598 736 56638 776
rect 56680 736 56720 776
rect 60352 736 60392 776
rect 60434 736 60474 776
rect 60516 736 60556 776
rect 60598 736 60638 776
rect 60680 736 60720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 68352 736 68392 776
rect 68434 736 68474 776
rect 68516 736 68556 776
rect 68598 736 68638 776
rect 68680 736 68720 776
rect 72352 736 72392 776
rect 72434 736 72474 776
rect 72516 736 72556 776
rect 72598 736 72638 776
rect 72680 736 72720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
rect 80352 736 80392 776
rect 80434 736 80474 776
rect 80516 736 80556 776
rect 80598 736 80638 776
rect 80680 736 80720 776
rect 84352 736 84392 776
rect 84434 736 84474 776
rect 84516 736 84556 776
rect 84598 736 84638 776
rect 84680 736 84720 776
rect 88352 736 88392 776
rect 88434 736 88474 776
rect 88516 736 88556 776
rect 88598 736 88638 776
rect 88680 736 88720 776
rect 92352 736 92392 776
rect 92434 736 92474 776
rect 92516 736 92556 776
rect 92598 736 92638 776
rect 92680 736 92720 776
rect 96352 736 96392 776
rect 96434 736 96474 776
rect 96516 736 96556 776
rect 96598 736 96638 776
rect 96680 736 96720 776
<< metal2 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 8352 38576 8720 38585
rect 8392 38536 8434 38576
rect 8474 38536 8516 38576
rect 8556 38536 8598 38576
rect 8638 38536 8680 38576
rect 8352 38527 8720 38536
rect 12352 38576 12720 38585
rect 12392 38536 12434 38576
rect 12474 38536 12516 38576
rect 12556 38536 12598 38576
rect 12638 38536 12680 38576
rect 12352 38527 12720 38536
rect 16352 38576 16720 38585
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16352 38527 16720 38536
rect 20352 38576 20720 38585
rect 20392 38536 20434 38576
rect 20474 38536 20516 38576
rect 20556 38536 20598 38576
rect 20638 38536 20680 38576
rect 20352 38527 20720 38536
rect 24352 38576 24720 38585
rect 24392 38536 24434 38576
rect 24474 38536 24516 38576
rect 24556 38536 24598 38576
rect 24638 38536 24680 38576
rect 24352 38527 24720 38536
rect 28352 38576 28720 38585
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28352 38527 28720 38536
rect 32352 38576 32720 38585
rect 32392 38536 32434 38576
rect 32474 38536 32516 38576
rect 32556 38536 32598 38576
rect 32638 38536 32680 38576
rect 32352 38527 32720 38536
rect 36352 38576 36720 38585
rect 36392 38536 36434 38576
rect 36474 38536 36516 38576
rect 36556 38536 36598 38576
rect 36638 38536 36680 38576
rect 36352 38527 36720 38536
rect 40352 38576 40720 38585
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40352 38527 40720 38536
rect 44352 38576 44720 38585
rect 44392 38536 44434 38576
rect 44474 38536 44516 38576
rect 44556 38536 44598 38576
rect 44638 38536 44680 38576
rect 44352 38527 44720 38536
rect 48352 38576 48720 38585
rect 48392 38536 48434 38576
rect 48474 38536 48516 38576
rect 48556 38536 48598 38576
rect 48638 38536 48680 38576
rect 48352 38527 48720 38536
rect 52352 38576 52720 38585
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52352 38527 52720 38536
rect 56352 38576 56720 38585
rect 56392 38536 56434 38576
rect 56474 38536 56516 38576
rect 56556 38536 56598 38576
rect 56638 38536 56680 38576
rect 56352 38527 56720 38536
rect 60352 38576 60720 38585
rect 60392 38536 60434 38576
rect 60474 38536 60516 38576
rect 60556 38536 60598 38576
rect 60638 38536 60680 38576
rect 60352 38527 60720 38536
rect 64352 38576 64720 38585
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64352 38527 64720 38536
rect 68352 38576 68720 38585
rect 68392 38536 68434 38576
rect 68474 38536 68516 38576
rect 68556 38536 68598 38576
rect 68638 38536 68680 38576
rect 68352 38527 68720 38536
rect 72352 38576 72720 38585
rect 72392 38536 72434 38576
rect 72474 38536 72516 38576
rect 72556 38536 72598 38576
rect 72638 38536 72680 38576
rect 72352 38527 72720 38536
rect 76352 38576 76720 38585
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76352 38527 76720 38536
rect 80352 38576 80720 38585
rect 80392 38536 80434 38576
rect 80474 38536 80516 38576
rect 80556 38536 80598 38576
rect 80638 38536 80680 38576
rect 80352 38527 80720 38536
rect 84352 38576 84720 38585
rect 84392 38536 84434 38576
rect 84474 38536 84516 38576
rect 84556 38536 84598 38576
rect 84638 38536 84680 38576
rect 84352 38527 84720 38536
rect 88352 38576 88720 38585
rect 88392 38536 88434 38576
rect 88474 38536 88516 38576
rect 88556 38536 88598 38576
rect 88638 38536 88680 38576
rect 88352 38527 88720 38536
rect 92352 38576 92720 38585
rect 92392 38536 92434 38576
rect 92474 38536 92516 38576
rect 92556 38536 92598 38576
rect 92638 38536 92680 38576
rect 92352 38527 92720 38536
rect 96352 38576 96720 38585
rect 96392 38536 96434 38576
rect 96474 38536 96516 38576
rect 96556 38536 96598 38576
rect 96638 38536 96680 38576
rect 96352 38527 96720 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 7112 37820 7480 37829
rect 7152 37780 7194 37820
rect 7234 37780 7276 37820
rect 7316 37780 7358 37820
rect 7398 37780 7440 37820
rect 7112 37771 7480 37780
rect 11112 37820 11480 37829
rect 11152 37780 11194 37820
rect 11234 37780 11276 37820
rect 11316 37780 11358 37820
rect 11398 37780 11440 37820
rect 11112 37771 11480 37780
rect 15112 37820 15480 37829
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15112 37771 15480 37780
rect 19112 37820 19480 37829
rect 19152 37780 19194 37820
rect 19234 37780 19276 37820
rect 19316 37780 19358 37820
rect 19398 37780 19440 37820
rect 19112 37771 19480 37780
rect 23112 37820 23480 37829
rect 23152 37780 23194 37820
rect 23234 37780 23276 37820
rect 23316 37780 23358 37820
rect 23398 37780 23440 37820
rect 23112 37771 23480 37780
rect 27112 37820 27480 37829
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27112 37771 27480 37780
rect 31112 37820 31480 37829
rect 31152 37780 31194 37820
rect 31234 37780 31276 37820
rect 31316 37780 31358 37820
rect 31398 37780 31440 37820
rect 31112 37771 31480 37780
rect 35112 37820 35480 37829
rect 35152 37780 35194 37820
rect 35234 37780 35276 37820
rect 35316 37780 35358 37820
rect 35398 37780 35440 37820
rect 35112 37771 35480 37780
rect 39112 37820 39480 37829
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39112 37771 39480 37780
rect 43112 37820 43480 37829
rect 43152 37780 43194 37820
rect 43234 37780 43276 37820
rect 43316 37780 43358 37820
rect 43398 37780 43440 37820
rect 43112 37771 43480 37780
rect 47112 37820 47480 37829
rect 47152 37780 47194 37820
rect 47234 37780 47276 37820
rect 47316 37780 47358 37820
rect 47398 37780 47440 37820
rect 47112 37771 47480 37780
rect 51112 37820 51480 37829
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51112 37771 51480 37780
rect 55112 37820 55480 37829
rect 55152 37780 55194 37820
rect 55234 37780 55276 37820
rect 55316 37780 55358 37820
rect 55398 37780 55440 37820
rect 55112 37771 55480 37780
rect 59112 37820 59480 37829
rect 59152 37780 59194 37820
rect 59234 37780 59276 37820
rect 59316 37780 59358 37820
rect 59398 37780 59440 37820
rect 59112 37771 59480 37780
rect 63112 37820 63480 37829
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63112 37771 63480 37780
rect 67112 37820 67480 37829
rect 67152 37780 67194 37820
rect 67234 37780 67276 37820
rect 67316 37780 67358 37820
rect 67398 37780 67440 37820
rect 67112 37771 67480 37780
rect 71112 37820 71480 37829
rect 71152 37780 71194 37820
rect 71234 37780 71276 37820
rect 71316 37780 71358 37820
rect 71398 37780 71440 37820
rect 71112 37771 71480 37780
rect 75112 37820 75480 37829
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75112 37771 75480 37780
rect 79112 37820 79480 37829
rect 79152 37780 79194 37820
rect 79234 37780 79276 37820
rect 79316 37780 79358 37820
rect 79398 37780 79440 37820
rect 79112 37771 79480 37780
rect 83112 37820 83480 37829
rect 83152 37780 83194 37820
rect 83234 37780 83276 37820
rect 83316 37780 83358 37820
rect 83398 37780 83440 37820
rect 83112 37771 83480 37780
rect 87112 37820 87480 37829
rect 87152 37780 87194 37820
rect 87234 37780 87276 37820
rect 87316 37780 87358 37820
rect 87398 37780 87440 37820
rect 87112 37771 87480 37780
rect 91112 37820 91480 37829
rect 91152 37780 91194 37820
rect 91234 37780 91276 37820
rect 91316 37780 91358 37820
rect 91398 37780 91440 37820
rect 91112 37771 91480 37780
rect 95112 37820 95480 37829
rect 95152 37780 95194 37820
rect 95234 37780 95276 37820
rect 95316 37780 95358 37820
rect 95398 37780 95440 37820
rect 95112 37771 95480 37780
rect 99112 37820 99480 37829
rect 99152 37780 99194 37820
rect 99234 37780 99276 37820
rect 99316 37780 99358 37820
rect 99398 37780 99440 37820
rect 99112 37771 99480 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 8352 37064 8720 37073
rect 8392 37024 8434 37064
rect 8474 37024 8516 37064
rect 8556 37024 8598 37064
rect 8638 37024 8680 37064
rect 8352 37015 8720 37024
rect 12352 37064 12720 37073
rect 12392 37024 12434 37064
rect 12474 37024 12516 37064
rect 12556 37024 12598 37064
rect 12638 37024 12680 37064
rect 12352 37015 12720 37024
rect 16352 37064 16720 37073
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16352 37015 16720 37024
rect 20352 37064 20720 37073
rect 20392 37024 20434 37064
rect 20474 37024 20516 37064
rect 20556 37024 20598 37064
rect 20638 37024 20680 37064
rect 20352 37015 20720 37024
rect 24352 37064 24720 37073
rect 24392 37024 24434 37064
rect 24474 37024 24516 37064
rect 24556 37024 24598 37064
rect 24638 37024 24680 37064
rect 24352 37015 24720 37024
rect 28352 37064 28720 37073
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28352 37015 28720 37024
rect 32352 37064 32720 37073
rect 32392 37024 32434 37064
rect 32474 37024 32516 37064
rect 32556 37024 32598 37064
rect 32638 37024 32680 37064
rect 32352 37015 32720 37024
rect 36352 37064 36720 37073
rect 36392 37024 36434 37064
rect 36474 37024 36516 37064
rect 36556 37024 36598 37064
rect 36638 37024 36680 37064
rect 36352 37015 36720 37024
rect 40352 37064 40720 37073
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40352 37015 40720 37024
rect 44352 37064 44720 37073
rect 44392 37024 44434 37064
rect 44474 37024 44516 37064
rect 44556 37024 44598 37064
rect 44638 37024 44680 37064
rect 44352 37015 44720 37024
rect 48352 37064 48720 37073
rect 48392 37024 48434 37064
rect 48474 37024 48516 37064
rect 48556 37024 48598 37064
rect 48638 37024 48680 37064
rect 48352 37015 48720 37024
rect 52352 37064 52720 37073
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52352 37015 52720 37024
rect 56352 37064 56720 37073
rect 56392 37024 56434 37064
rect 56474 37024 56516 37064
rect 56556 37024 56598 37064
rect 56638 37024 56680 37064
rect 56352 37015 56720 37024
rect 60352 37064 60720 37073
rect 60392 37024 60434 37064
rect 60474 37024 60516 37064
rect 60556 37024 60598 37064
rect 60638 37024 60680 37064
rect 60352 37015 60720 37024
rect 64352 37064 64720 37073
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64352 37015 64720 37024
rect 68352 37064 68720 37073
rect 68392 37024 68434 37064
rect 68474 37024 68516 37064
rect 68556 37024 68598 37064
rect 68638 37024 68680 37064
rect 68352 37015 68720 37024
rect 72352 37064 72720 37073
rect 72392 37024 72434 37064
rect 72474 37024 72516 37064
rect 72556 37024 72598 37064
rect 72638 37024 72680 37064
rect 72352 37015 72720 37024
rect 76352 37064 76720 37073
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76352 37015 76720 37024
rect 80352 37064 80720 37073
rect 80392 37024 80434 37064
rect 80474 37024 80516 37064
rect 80556 37024 80598 37064
rect 80638 37024 80680 37064
rect 80352 37015 80720 37024
rect 84352 37064 84720 37073
rect 84392 37024 84434 37064
rect 84474 37024 84516 37064
rect 84556 37024 84598 37064
rect 84638 37024 84680 37064
rect 84352 37015 84720 37024
rect 88352 37064 88720 37073
rect 88392 37024 88434 37064
rect 88474 37024 88516 37064
rect 88556 37024 88598 37064
rect 88638 37024 88680 37064
rect 88352 37015 88720 37024
rect 92352 37064 92720 37073
rect 92392 37024 92434 37064
rect 92474 37024 92516 37064
rect 92556 37024 92598 37064
rect 92638 37024 92680 37064
rect 92352 37015 92720 37024
rect 96352 37064 96720 37073
rect 96392 37024 96434 37064
rect 96474 37024 96516 37064
rect 96556 37024 96598 37064
rect 96638 37024 96680 37064
rect 96352 37015 96720 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 7112 36308 7480 36317
rect 7152 36268 7194 36308
rect 7234 36268 7276 36308
rect 7316 36268 7358 36308
rect 7398 36268 7440 36308
rect 7112 36259 7480 36268
rect 11112 36308 11480 36317
rect 11152 36268 11194 36308
rect 11234 36268 11276 36308
rect 11316 36268 11358 36308
rect 11398 36268 11440 36308
rect 11112 36259 11480 36268
rect 15112 36308 15480 36317
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15112 36259 15480 36268
rect 19112 36308 19480 36317
rect 19152 36268 19194 36308
rect 19234 36268 19276 36308
rect 19316 36268 19358 36308
rect 19398 36268 19440 36308
rect 19112 36259 19480 36268
rect 23112 36308 23480 36317
rect 23152 36268 23194 36308
rect 23234 36268 23276 36308
rect 23316 36268 23358 36308
rect 23398 36268 23440 36308
rect 23112 36259 23480 36268
rect 27112 36308 27480 36317
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27112 36259 27480 36268
rect 31112 36308 31480 36317
rect 31152 36268 31194 36308
rect 31234 36268 31276 36308
rect 31316 36268 31358 36308
rect 31398 36268 31440 36308
rect 31112 36259 31480 36268
rect 35112 36308 35480 36317
rect 35152 36268 35194 36308
rect 35234 36268 35276 36308
rect 35316 36268 35358 36308
rect 35398 36268 35440 36308
rect 35112 36259 35480 36268
rect 39112 36308 39480 36317
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39112 36259 39480 36268
rect 43112 36308 43480 36317
rect 43152 36268 43194 36308
rect 43234 36268 43276 36308
rect 43316 36268 43358 36308
rect 43398 36268 43440 36308
rect 43112 36259 43480 36268
rect 47112 36308 47480 36317
rect 47152 36268 47194 36308
rect 47234 36268 47276 36308
rect 47316 36268 47358 36308
rect 47398 36268 47440 36308
rect 47112 36259 47480 36268
rect 51112 36308 51480 36317
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51112 36259 51480 36268
rect 55112 36308 55480 36317
rect 55152 36268 55194 36308
rect 55234 36268 55276 36308
rect 55316 36268 55358 36308
rect 55398 36268 55440 36308
rect 55112 36259 55480 36268
rect 59112 36308 59480 36317
rect 59152 36268 59194 36308
rect 59234 36268 59276 36308
rect 59316 36268 59358 36308
rect 59398 36268 59440 36308
rect 59112 36259 59480 36268
rect 63112 36308 63480 36317
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63112 36259 63480 36268
rect 67112 36308 67480 36317
rect 67152 36268 67194 36308
rect 67234 36268 67276 36308
rect 67316 36268 67358 36308
rect 67398 36268 67440 36308
rect 67112 36259 67480 36268
rect 71112 36308 71480 36317
rect 71152 36268 71194 36308
rect 71234 36268 71276 36308
rect 71316 36268 71358 36308
rect 71398 36268 71440 36308
rect 71112 36259 71480 36268
rect 75112 36308 75480 36317
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75112 36259 75480 36268
rect 79112 36308 79480 36317
rect 79152 36268 79194 36308
rect 79234 36268 79276 36308
rect 79316 36268 79358 36308
rect 79398 36268 79440 36308
rect 79112 36259 79480 36268
rect 83112 36308 83480 36317
rect 83152 36268 83194 36308
rect 83234 36268 83276 36308
rect 83316 36268 83358 36308
rect 83398 36268 83440 36308
rect 83112 36259 83480 36268
rect 87112 36308 87480 36317
rect 87152 36268 87194 36308
rect 87234 36268 87276 36308
rect 87316 36268 87358 36308
rect 87398 36268 87440 36308
rect 87112 36259 87480 36268
rect 91112 36308 91480 36317
rect 91152 36268 91194 36308
rect 91234 36268 91276 36308
rect 91316 36268 91358 36308
rect 91398 36268 91440 36308
rect 91112 36259 91480 36268
rect 95112 36308 95480 36317
rect 95152 36268 95194 36308
rect 95234 36268 95276 36308
rect 95316 36268 95358 36308
rect 95398 36268 95440 36308
rect 95112 36259 95480 36268
rect 99112 36308 99480 36317
rect 99152 36268 99194 36308
rect 99234 36268 99276 36308
rect 99316 36268 99358 36308
rect 99398 36268 99440 36308
rect 99112 36259 99480 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 8352 35552 8720 35561
rect 8392 35512 8434 35552
rect 8474 35512 8516 35552
rect 8556 35512 8598 35552
rect 8638 35512 8680 35552
rect 8352 35503 8720 35512
rect 12352 35552 12720 35561
rect 12392 35512 12434 35552
rect 12474 35512 12516 35552
rect 12556 35512 12598 35552
rect 12638 35512 12680 35552
rect 12352 35503 12720 35512
rect 16352 35552 16720 35561
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16352 35503 16720 35512
rect 20352 35552 20720 35561
rect 20392 35512 20434 35552
rect 20474 35512 20516 35552
rect 20556 35512 20598 35552
rect 20638 35512 20680 35552
rect 20352 35503 20720 35512
rect 24352 35552 24720 35561
rect 24392 35512 24434 35552
rect 24474 35512 24516 35552
rect 24556 35512 24598 35552
rect 24638 35512 24680 35552
rect 24352 35503 24720 35512
rect 28352 35552 28720 35561
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28352 35503 28720 35512
rect 32352 35552 32720 35561
rect 32392 35512 32434 35552
rect 32474 35512 32516 35552
rect 32556 35512 32598 35552
rect 32638 35512 32680 35552
rect 32352 35503 32720 35512
rect 36352 35552 36720 35561
rect 36392 35512 36434 35552
rect 36474 35512 36516 35552
rect 36556 35512 36598 35552
rect 36638 35512 36680 35552
rect 36352 35503 36720 35512
rect 40352 35552 40720 35561
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40352 35503 40720 35512
rect 44352 35552 44720 35561
rect 44392 35512 44434 35552
rect 44474 35512 44516 35552
rect 44556 35512 44598 35552
rect 44638 35512 44680 35552
rect 44352 35503 44720 35512
rect 48352 35552 48720 35561
rect 48392 35512 48434 35552
rect 48474 35512 48516 35552
rect 48556 35512 48598 35552
rect 48638 35512 48680 35552
rect 48352 35503 48720 35512
rect 52352 35552 52720 35561
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52352 35503 52720 35512
rect 56352 35552 56720 35561
rect 56392 35512 56434 35552
rect 56474 35512 56516 35552
rect 56556 35512 56598 35552
rect 56638 35512 56680 35552
rect 56352 35503 56720 35512
rect 60352 35552 60720 35561
rect 60392 35512 60434 35552
rect 60474 35512 60516 35552
rect 60556 35512 60598 35552
rect 60638 35512 60680 35552
rect 60352 35503 60720 35512
rect 64352 35552 64720 35561
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64352 35503 64720 35512
rect 68352 35552 68720 35561
rect 68392 35512 68434 35552
rect 68474 35512 68516 35552
rect 68556 35512 68598 35552
rect 68638 35512 68680 35552
rect 68352 35503 68720 35512
rect 72352 35552 72720 35561
rect 72392 35512 72434 35552
rect 72474 35512 72516 35552
rect 72556 35512 72598 35552
rect 72638 35512 72680 35552
rect 72352 35503 72720 35512
rect 76352 35552 76720 35561
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76352 35503 76720 35512
rect 80352 35552 80720 35561
rect 80392 35512 80434 35552
rect 80474 35512 80516 35552
rect 80556 35512 80598 35552
rect 80638 35512 80680 35552
rect 80352 35503 80720 35512
rect 84352 35552 84720 35561
rect 84392 35512 84434 35552
rect 84474 35512 84516 35552
rect 84556 35512 84598 35552
rect 84638 35512 84680 35552
rect 84352 35503 84720 35512
rect 88352 35552 88720 35561
rect 88392 35512 88434 35552
rect 88474 35512 88516 35552
rect 88556 35512 88598 35552
rect 88638 35512 88680 35552
rect 88352 35503 88720 35512
rect 92352 35552 92720 35561
rect 92392 35512 92434 35552
rect 92474 35512 92516 35552
rect 92556 35512 92598 35552
rect 92638 35512 92680 35552
rect 92352 35503 92720 35512
rect 96352 35552 96720 35561
rect 96392 35512 96434 35552
rect 96474 35512 96516 35552
rect 96556 35512 96598 35552
rect 96638 35512 96680 35552
rect 96352 35503 96720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 7112 34796 7480 34805
rect 7152 34756 7194 34796
rect 7234 34756 7276 34796
rect 7316 34756 7358 34796
rect 7398 34756 7440 34796
rect 7112 34747 7480 34756
rect 11112 34796 11480 34805
rect 11152 34756 11194 34796
rect 11234 34756 11276 34796
rect 11316 34756 11358 34796
rect 11398 34756 11440 34796
rect 11112 34747 11480 34756
rect 15112 34796 15480 34805
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15112 34747 15480 34756
rect 19112 34796 19480 34805
rect 19152 34756 19194 34796
rect 19234 34756 19276 34796
rect 19316 34756 19358 34796
rect 19398 34756 19440 34796
rect 19112 34747 19480 34756
rect 23112 34796 23480 34805
rect 23152 34756 23194 34796
rect 23234 34756 23276 34796
rect 23316 34756 23358 34796
rect 23398 34756 23440 34796
rect 23112 34747 23480 34756
rect 27112 34796 27480 34805
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27112 34747 27480 34756
rect 31112 34796 31480 34805
rect 31152 34756 31194 34796
rect 31234 34756 31276 34796
rect 31316 34756 31358 34796
rect 31398 34756 31440 34796
rect 31112 34747 31480 34756
rect 35112 34796 35480 34805
rect 35152 34756 35194 34796
rect 35234 34756 35276 34796
rect 35316 34756 35358 34796
rect 35398 34756 35440 34796
rect 35112 34747 35480 34756
rect 39112 34796 39480 34805
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39112 34747 39480 34756
rect 43112 34796 43480 34805
rect 43152 34756 43194 34796
rect 43234 34756 43276 34796
rect 43316 34756 43358 34796
rect 43398 34756 43440 34796
rect 43112 34747 43480 34756
rect 47112 34796 47480 34805
rect 47152 34756 47194 34796
rect 47234 34756 47276 34796
rect 47316 34756 47358 34796
rect 47398 34756 47440 34796
rect 47112 34747 47480 34756
rect 51112 34796 51480 34805
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51112 34747 51480 34756
rect 55112 34796 55480 34805
rect 55152 34756 55194 34796
rect 55234 34756 55276 34796
rect 55316 34756 55358 34796
rect 55398 34756 55440 34796
rect 55112 34747 55480 34756
rect 59112 34796 59480 34805
rect 59152 34756 59194 34796
rect 59234 34756 59276 34796
rect 59316 34756 59358 34796
rect 59398 34756 59440 34796
rect 59112 34747 59480 34756
rect 63112 34796 63480 34805
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63112 34747 63480 34756
rect 67112 34796 67480 34805
rect 67152 34756 67194 34796
rect 67234 34756 67276 34796
rect 67316 34756 67358 34796
rect 67398 34756 67440 34796
rect 67112 34747 67480 34756
rect 71112 34796 71480 34805
rect 71152 34756 71194 34796
rect 71234 34756 71276 34796
rect 71316 34756 71358 34796
rect 71398 34756 71440 34796
rect 71112 34747 71480 34756
rect 75112 34796 75480 34805
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75112 34747 75480 34756
rect 79112 34796 79480 34805
rect 79152 34756 79194 34796
rect 79234 34756 79276 34796
rect 79316 34756 79358 34796
rect 79398 34756 79440 34796
rect 79112 34747 79480 34756
rect 83112 34796 83480 34805
rect 83152 34756 83194 34796
rect 83234 34756 83276 34796
rect 83316 34756 83358 34796
rect 83398 34756 83440 34796
rect 83112 34747 83480 34756
rect 87112 34796 87480 34805
rect 87152 34756 87194 34796
rect 87234 34756 87276 34796
rect 87316 34756 87358 34796
rect 87398 34756 87440 34796
rect 87112 34747 87480 34756
rect 91112 34796 91480 34805
rect 91152 34756 91194 34796
rect 91234 34756 91276 34796
rect 91316 34756 91358 34796
rect 91398 34756 91440 34796
rect 91112 34747 91480 34756
rect 95112 34796 95480 34805
rect 95152 34756 95194 34796
rect 95234 34756 95276 34796
rect 95316 34756 95358 34796
rect 95398 34756 95440 34796
rect 95112 34747 95480 34756
rect 99112 34796 99480 34805
rect 99152 34756 99194 34796
rect 99234 34756 99276 34796
rect 99316 34756 99358 34796
rect 99398 34756 99440 34796
rect 99112 34747 99480 34756
rect 91468 34460 91508 34469
rect 91276 34420 91468 34460
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 8352 34040 8720 34049
rect 8392 34000 8434 34040
rect 8474 34000 8516 34040
rect 8556 34000 8598 34040
rect 8638 34000 8680 34040
rect 8352 33991 8720 34000
rect 12352 34040 12720 34049
rect 12392 34000 12434 34040
rect 12474 34000 12516 34040
rect 12556 34000 12598 34040
rect 12638 34000 12680 34040
rect 12352 33991 12720 34000
rect 16352 34040 16720 34049
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16352 33991 16720 34000
rect 20352 34040 20720 34049
rect 20392 34000 20434 34040
rect 20474 34000 20516 34040
rect 20556 34000 20598 34040
rect 20638 34000 20680 34040
rect 20352 33991 20720 34000
rect 24352 34040 24720 34049
rect 24392 34000 24434 34040
rect 24474 34000 24516 34040
rect 24556 34000 24598 34040
rect 24638 34000 24680 34040
rect 24352 33991 24720 34000
rect 28352 34040 28720 34049
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28352 33991 28720 34000
rect 32352 34040 32720 34049
rect 32392 34000 32434 34040
rect 32474 34000 32516 34040
rect 32556 34000 32598 34040
rect 32638 34000 32680 34040
rect 32352 33991 32720 34000
rect 36352 34040 36720 34049
rect 36392 34000 36434 34040
rect 36474 34000 36516 34040
rect 36556 34000 36598 34040
rect 36638 34000 36680 34040
rect 36352 33991 36720 34000
rect 40352 34040 40720 34049
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40352 33991 40720 34000
rect 44352 34040 44720 34049
rect 44392 34000 44434 34040
rect 44474 34000 44516 34040
rect 44556 34000 44598 34040
rect 44638 34000 44680 34040
rect 44352 33991 44720 34000
rect 48352 34040 48720 34049
rect 48392 34000 48434 34040
rect 48474 34000 48516 34040
rect 48556 34000 48598 34040
rect 48638 34000 48680 34040
rect 48352 33991 48720 34000
rect 52352 34040 52720 34049
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52352 33991 52720 34000
rect 56352 34040 56720 34049
rect 56392 34000 56434 34040
rect 56474 34000 56516 34040
rect 56556 34000 56598 34040
rect 56638 34000 56680 34040
rect 56352 33991 56720 34000
rect 60352 34040 60720 34049
rect 60392 34000 60434 34040
rect 60474 34000 60516 34040
rect 60556 34000 60598 34040
rect 60638 34000 60680 34040
rect 60352 33991 60720 34000
rect 64352 34040 64720 34049
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64352 33991 64720 34000
rect 68352 34040 68720 34049
rect 68392 34000 68434 34040
rect 68474 34000 68516 34040
rect 68556 34000 68598 34040
rect 68638 34000 68680 34040
rect 68352 33991 68720 34000
rect 91276 33797 91316 34420
rect 91468 34411 91508 34420
rect 93388 34460 93428 34469
rect 91660 34208 91700 34217
rect 91564 34168 91660 34208
rect 91275 33788 91317 33797
rect 91275 33748 91276 33788
rect 91316 33748 91317 33788
rect 91275 33739 91317 33748
rect 73228 33620 73268 33629
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 7112 33284 7480 33293
rect 7152 33244 7194 33284
rect 7234 33244 7276 33284
rect 7316 33244 7358 33284
rect 7398 33244 7440 33284
rect 7112 33235 7480 33244
rect 11112 33284 11480 33293
rect 11152 33244 11194 33284
rect 11234 33244 11276 33284
rect 11316 33244 11358 33284
rect 11398 33244 11440 33284
rect 11112 33235 11480 33244
rect 15112 33284 15480 33293
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15112 33235 15480 33244
rect 19112 33284 19480 33293
rect 19152 33244 19194 33284
rect 19234 33244 19276 33284
rect 19316 33244 19358 33284
rect 19398 33244 19440 33284
rect 19112 33235 19480 33244
rect 23112 33284 23480 33293
rect 23152 33244 23194 33284
rect 23234 33244 23276 33284
rect 23316 33244 23358 33284
rect 23398 33244 23440 33284
rect 23112 33235 23480 33244
rect 27112 33284 27480 33293
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27112 33235 27480 33244
rect 31112 33284 31480 33293
rect 31152 33244 31194 33284
rect 31234 33244 31276 33284
rect 31316 33244 31358 33284
rect 31398 33244 31440 33284
rect 31112 33235 31480 33244
rect 35112 33284 35480 33293
rect 35152 33244 35194 33284
rect 35234 33244 35276 33284
rect 35316 33244 35358 33284
rect 35398 33244 35440 33284
rect 35112 33235 35480 33244
rect 39112 33284 39480 33293
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39112 33235 39480 33244
rect 43112 33284 43480 33293
rect 43152 33244 43194 33284
rect 43234 33244 43276 33284
rect 43316 33244 43358 33284
rect 43398 33244 43440 33284
rect 43112 33235 43480 33244
rect 47112 33284 47480 33293
rect 47152 33244 47194 33284
rect 47234 33244 47276 33284
rect 47316 33244 47358 33284
rect 47398 33244 47440 33284
rect 47112 33235 47480 33244
rect 51112 33284 51480 33293
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51112 33235 51480 33244
rect 55112 33284 55480 33293
rect 55152 33244 55194 33284
rect 55234 33244 55276 33284
rect 55316 33244 55358 33284
rect 55398 33244 55440 33284
rect 55112 33235 55480 33244
rect 59112 33284 59480 33293
rect 59152 33244 59194 33284
rect 59234 33244 59276 33284
rect 59316 33244 59358 33284
rect 59398 33244 59440 33284
rect 59112 33235 59480 33244
rect 63112 33284 63480 33293
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63112 33235 63480 33244
rect 67112 33284 67480 33293
rect 67152 33244 67194 33284
rect 67234 33244 67276 33284
rect 67316 33244 67358 33284
rect 67398 33244 67440 33284
rect 67112 33235 67480 33244
rect 71787 33284 71829 33293
rect 71787 33244 71788 33284
rect 71828 33244 71829 33284
rect 71787 33235 71829 33244
rect 70731 32948 70773 32957
rect 70731 32908 70732 32948
rect 70772 32908 70773 32948
rect 70731 32899 70773 32908
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 8352 32528 8720 32537
rect 8392 32488 8434 32528
rect 8474 32488 8516 32528
rect 8556 32488 8598 32528
rect 8638 32488 8680 32528
rect 8352 32479 8720 32488
rect 12352 32528 12720 32537
rect 12392 32488 12434 32528
rect 12474 32488 12516 32528
rect 12556 32488 12598 32528
rect 12638 32488 12680 32528
rect 12352 32479 12720 32488
rect 16352 32528 16720 32537
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16352 32479 16720 32488
rect 20352 32528 20720 32537
rect 20392 32488 20434 32528
rect 20474 32488 20516 32528
rect 20556 32488 20598 32528
rect 20638 32488 20680 32528
rect 20352 32479 20720 32488
rect 24352 32528 24720 32537
rect 24392 32488 24434 32528
rect 24474 32488 24516 32528
rect 24556 32488 24598 32528
rect 24638 32488 24680 32528
rect 24352 32479 24720 32488
rect 28352 32528 28720 32537
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28352 32479 28720 32488
rect 32352 32528 32720 32537
rect 32392 32488 32434 32528
rect 32474 32488 32516 32528
rect 32556 32488 32598 32528
rect 32638 32488 32680 32528
rect 32352 32479 32720 32488
rect 36352 32528 36720 32537
rect 36392 32488 36434 32528
rect 36474 32488 36516 32528
rect 36556 32488 36598 32528
rect 36638 32488 36680 32528
rect 36352 32479 36720 32488
rect 40352 32528 40720 32537
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40352 32479 40720 32488
rect 44352 32528 44720 32537
rect 44392 32488 44434 32528
rect 44474 32488 44516 32528
rect 44556 32488 44598 32528
rect 44638 32488 44680 32528
rect 44352 32479 44720 32488
rect 48352 32528 48720 32537
rect 48392 32488 48434 32528
rect 48474 32488 48516 32528
rect 48556 32488 48598 32528
rect 48638 32488 48680 32528
rect 48352 32479 48720 32488
rect 52352 32528 52720 32537
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52352 32479 52720 32488
rect 56352 32528 56720 32537
rect 56392 32488 56434 32528
rect 56474 32488 56516 32528
rect 56556 32488 56598 32528
rect 56638 32488 56680 32528
rect 56352 32479 56720 32488
rect 60352 32528 60720 32537
rect 60392 32488 60434 32528
rect 60474 32488 60516 32528
rect 60556 32488 60598 32528
rect 60638 32488 60680 32528
rect 60352 32479 60720 32488
rect 64352 32528 64720 32537
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64352 32479 64720 32488
rect 68352 32528 68720 32537
rect 68392 32488 68434 32528
rect 68474 32488 68516 32528
rect 68556 32488 68598 32528
rect 68638 32488 68680 32528
rect 68352 32479 68720 32488
rect 70732 32360 70772 32899
rect 71596 32873 71636 32958
rect 71500 32864 71540 32873
rect 71500 32780 71540 32824
rect 71595 32864 71637 32873
rect 71595 32824 71596 32864
rect 71636 32824 71637 32864
rect 71595 32815 71637 32824
rect 70732 32311 70772 32320
rect 71212 32740 71540 32780
rect 70827 32192 70869 32201
rect 70827 32152 70828 32192
rect 70868 32152 70869 32192
rect 70827 32143 70869 32152
rect 70539 32108 70581 32117
rect 70539 32068 70540 32108
rect 70580 32068 70581 32108
rect 70539 32059 70581 32068
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 7112 31772 7480 31781
rect 7152 31732 7194 31772
rect 7234 31732 7276 31772
rect 7316 31732 7358 31772
rect 7398 31732 7440 31772
rect 7112 31723 7480 31732
rect 11112 31772 11480 31781
rect 11152 31732 11194 31772
rect 11234 31732 11276 31772
rect 11316 31732 11358 31772
rect 11398 31732 11440 31772
rect 11112 31723 11480 31732
rect 15112 31772 15480 31781
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15112 31723 15480 31732
rect 19112 31772 19480 31781
rect 19152 31732 19194 31772
rect 19234 31732 19276 31772
rect 19316 31732 19358 31772
rect 19398 31732 19440 31772
rect 19112 31723 19480 31732
rect 23112 31772 23480 31781
rect 23152 31732 23194 31772
rect 23234 31732 23276 31772
rect 23316 31732 23358 31772
rect 23398 31732 23440 31772
rect 23112 31723 23480 31732
rect 27112 31772 27480 31781
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27112 31723 27480 31732
rect 31112 31772 31480 31781
rect 31152 31732 31194 31772
rect 31234 31732 31276 31772
rect 31316 31732 31358 31772
rect 31398 31732 31440 31772
rect 31112 31723 31480 31732
rect 35112 31772 35480 31781
rect 35152 31732 35194 31772
rect 35234 31732 35276 31772
rect 35316 31732 35358 31772
rect 35398 31732 35440 31772
rect 35112 31723 35480 31732
rect 39112 31772 39480 31781
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39112 31723 39480 31732
rect 43112 31772 43480 31781
rect 43152 31732 43194 31772
rect 43234 31732 43276 31772
rect 43316 31732 43358 31772
rect 43398 31732 43440 31772
rect 43112 31723 43480 31732
rect 47112 31772 47480 31781
rect 47152 31732 47194 31772
rect 47234 31732 47276 31772
rect 47316 31732 47358 31772
rect 47398 31732 47440 31772
rect 47112 31723 47480 31732
rect 51112 31772 51480 31781
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51112 31723 51480 31732
rect 55112 31772 55480 31781
rect 55152 31732 55194 31772
rect 55234 31732 55276 31772
rect 55316 31732 55358 31772
rect 55398 31732 55440 31772
rect 55112 31723 55480 31732
rect 59112 31772 59480 31781
rect 59152 31732 59194 31772
rect 59234 31732 59276 31772
rect 59316 31732 59358 31772
rect 59398 31732 59440 31772
rect 59112 31723 59480 31732
rect 63112 31772 63480 31781
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63112 31723 63480 31732
rect 67112 31772 67480 31781
rect 67152 31732 67194 31772
rect 67234 31732 67276 31772
rect 67316 31732 67358 31772
rect 67398 31732 67440 31772
rect 67112 31723 67480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 8352 31016 8720 31025
rect 8392 30976 8434 31016
rect 8474 30976 8516 31016
rect 8556 30976 8598 31016
rect 8638 30976 8680 31016
rect 8352 30967 8720 30976
rect 12352 31016 12720 31025
rect 12392 30976 12434 31016
rect 12474 30976 12516 31016
rect 12556 30976 12598 31016
rect 12638 30976 12680 31016
rect 12352 30967 12720 30976
rect 16352 31016 16720 31025
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16352 30967 16720 30976
rect 20352 31016 20720 31025
rect 20392 30976 20434 31016
rect 20474 30976 20516 31016
rect 20556 30976 20598 31016
rect 20638 30976 20680 31016
rect 20352 30967 20720 30976
rect 24352 31016 24720 31025
rect 24392 30976 24434 31016
rect 24474 30976 24516 31016
rect 24556 30976 24598 31016
rect 24638 30976 24680 31016
rect 24352 30967 24720 30976
rect 28352 31016 28720 31025
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28352 30967 28720 30976
rect 32352 31016 32720 31025
rect 32392 30976 32434 31016
rect 32474 30976 32516 31016
rect 32556 30976 32598 31016
rect 32638 30976 32680 31016
rect 32352 30967 32720 30976
rect 36352 31016 36720 31025
rect 36392 30976 36434 31016
rect 36474 30976 36516 31016
rect 36556 30976 36598 31016
rect 36638 30976 36680 31016
rect 36352 30967 36720 30976
rect 40352 31016 40720 31025
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40352 30967 40720 30976
rect 44352 31016 44720 31025
rect 44392 30976 44434 31016
rect 44474 30976 44516 31016
rect 44556 30976 44598 31016
rect 44638 30976 44680 31016
rect 44352 30967 44720 30976
rect 48352 31016 48720 31025
rect 48392 30976 48434 31016
rect 48474 30976 48516 31016
rect 48556 30976 48598 31016
rect 48638 30976 48680 31016
rect 48352 30967 48720 30976
rect 52352 31016 52720 31025
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52352 30967 52720 30976
rect 56352 31016 56720 31025
rect 56392 30976 56434 31016
rect 56474 30976 56516 31016
rect 56556 30976 56598 31016
rect 56638 30976 56680 31016
rect 56352 30967 56720 30976
rect 60352 31016 60720 31025
rect 60392 30976 60434 31016
rect 60474 30976 60516 31016
rect 60556 30976 60598 31016
rect 60638 30976 60680 31016
rect 60352 30967 60720 30976
rect 64352 31016 64720 31025
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64352 30967 64720 30976
rect 68352 31016 68720 31025
rect 68392 30976 68434 31016
rect 68474 30976 68516 31016
rect 68556 30976 68598 31016
rect 68638 30976 68680 31016
rect 68352 30967 68720 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 7112 30260 7480 30269
rect 7152 30220 7194 30260
rect 7234 30220 7276 30260
rect 7316 30220 7358 30260
rect 7398 30220 7440 30260
rect 7112 30211 7480 30220
rect 11112 30260 11480 30269
rect 11152 30220 11194 30260
rect 11234 30220 11276 30260
rect 11316 30220 11358 30260
rect 11398 30220 11440 30260
rect 11112 30211 11480 30220
rect 15112 30260 15480 30269
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15112 30211 15480 30220
rect 19112 30260 19480 30269
rect 19152 30220 19194 30260
rect 19234 30220 19276 30260
rect 19316 30220 19358 30260
rect 19398 30220 19440 30260
rect 19112 30211 19480 30220
rect 23112 30260 23480 30269
rect 23152 30220 23194 30260
rect 23234 30220 23276 30260
rect 23316 30220 23358 30260
rect 23398 30220 23440 30260
rect 23112 30211 23480 30220
rect 27112 30260 27480 30269
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27112 30211 27480 30220
rect 31112 30260 31480 30269
rect 31152 30220 31194 30260
rect 31234 30220 31276 30260
rect 31316 30220 31358 30260
rect 31398 30220 31440 30260
rect 31112 30211 31480 30220
rect 35112 30260 35480 30269
rect 35152 30220 35194 30260
rect 35234 30220 35276 30260
rect 35316 30220 35358 30260
rect 35398 30220 35440 30260
rect 35112 30211 35480 30220
rect 39112 30260 39480 30269
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39112 30211 39480 30220
rect 43112 30260 43480 30269
rect 43152 30220 43194 30260
rect 43234 30220 43276 30260
rect 43316 30220 43358 30260
rect 43398 30220 43440 30260
rect 43112 30211 43480 30220
rect 47112 30260 47480 30269
rect 47152 30220 47194 30260
rect 47234 30220 47276 30260
rect 47316 30220 47358 30260
rect 47398 30220 47440 30260
rect 47112 30211 47480 30220
rect 51112 30260 51480 30269
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51112 30211 51480 30220
rect 55112 30260 55480 30269
rect 55152 30220 55194 30260
rect 55234 30220 55276 30260
rect 55316 30220 55358 30260
rect 55398 30220 55440 30260
rect 55112 30211 55480 30220
rect 59112 30260 59480 30269
rect 59152 30220 59194 30260
rect 59234 30220 59276 30260
rect 59316 30220 59358 30260
rect 59398 30220 59440 30260
rect 59112 30211 59480 30220
rect 63112 30260 63480 30269
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63112 30211 63480 30220
rect 67112 30260 67480 30269
rect 67152 30220 67194 30260
rect 67234 30220 67276 30260
rect 67316 30220 67358 30260
rect 67398 30220 67440 30260
rect 67112 30211 67480 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 8352 29504 8720 29513
rect 8392 29464 8434 29504
rect 8474 29464 8516 29504
rect 8556 29464 8598 29504
rect 8638 29464 8680 29504
rect 8352 29455 8720 29464
rect 12352 29504 12720 29513
rect 12392 29464 12434 29504
rect 12474 29464 12516 29504
rect 12556 29464 12598 29504
rect 12638 29464 12680 29504
rect 12352 29455 12720 29464
rect 16352 29504 16720 29513
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16352 29455 16720 29464
rect 20352 29504 20720 29513
rect 20392 29464 20434 29504
rect 20474 29464 20516 29504
rect 20556 29464 20598 29504
rect 20638 29464 20680 29504
rect 20352 29455 20720 29464
rect 24352 29504 24720 29513
rect 24392 29464 24434 29504
rect 24474 29464 24516 29504
rect 24556 29464 24598 29504
rect 24638 29464 24680 29504
rect 24352 29455 24720 29464
rect 28352 29504 28720 29513
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28352 29455 28720 29464
rect 32352 29504 32720 29513
rect 32392 29464 32434 29504
rect 32474 29464 32516 29504
rect 32556 29464 32598 29504
rect 32638 29464 32680 29504
rect 32352 29455 32720 29464
rect 36352 29504 36720 29513
rect 36392 29464 36434 29504
rect 36474 29464 36516 29504
rect 36556 29464 36598 29504
rect 36638 29464 36680 29504
rect 36352 29455 36720 29464
rect 40352 29504 40720 29513
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40352 29455 40720 29464
rect 44352 29504 44720 29513
rect 44392 29464 44434 29504
rect 44474 29464 44516 29504
rect 44556 29464 44598 29504
rect 44638 29464 44680 29504
rect 44352 29455 44720 29464
rect 48352 29504 48720 29513
rect 48392 29464 48434 29504
rect 48474 29464 48516 29504
rect 48556 29464 48598 29504
rect 48638 29464 48680 29504
rect 48352 29455 48720 29464
rect 52352 29504 52720 29513
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52352 29455 52720 29464
rect 56352 29504 56720 29513
rect 56392 29464 56434 29504
rect 56474 29464 56516 29504
rect 56556 29464 56598 29504
rect 56638 29464 56680 29504
rect 56352 29455 56720 29464
rect 60352 29504 60720 29513
rect 60392 29464 60434 29504
rect 60474 29464 60516 29504
rect 60556 29464 60598 29504
rect 60638 29464 60680 29504
rect 60352 29455 60720 29464
rect 64352 29504 64720 29513
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64352 29455 64720 29464
rect 68352 29504 68720 29513
rect 68392 29464 68434 29504
rect 68474 29464 68516 29504
rect 68556 29464 68598 29504
rect 68638 29464 68680 29504
rect 68352 29455 68720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 7112 28748 7480 28757
rect 7152 28708 7194 28748
rect 7234 28708 7276 28748
rect 7316 28708 7358 28748
rect 7398 28708 7440 28748
rect 7112 28699 7480 28708
rect 11112 28748 11480 28757
rect 11152 28708 11194 28748
rect 11234 28708 11276 28748
rect 11316 28708 11358 28748
rect 11398 28708 11440 28748
rect 11112 28699 11480 28708
rect 15112 28748 15480 28757
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15112 28699 15480 28708
rect 19112 28748 19480 28757
rect 19152 28708 19194 28748
rect 19234 28708 19276 28748
rect 19316 28708 19358 28748
rect 19398 28708 19440 28748
rect 19112 28699 19480 28708
rect 23112 28748 23480 28757
rect 23152 28708 23194 28748
rect 23234 28708 23276 28748
rect 23316 28708 23358 28748
rect 23398 28708 23440 28748
rect 23112 28699 23480 28708
rect 27112 28748 27480 28757
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27112 28699 27480 28708
rect 31112 28748 31480 28757
rect 31152 28708 31194 28748
rect 31234 28708 31276 28748
rect 31316 28708 31358 28748
rect 31398 28708 31440 28748
rect 31112 28699 31480 28708
rect 35112 28748 35480 28757
rect 35152 28708 35194 28748
rect 35234 28708 35276 28748
rect 35316 28708 35358 28748
rect 35398 28708 35440 28748
rect 35112 28699 35480 28708
rect 39112 28748 39480 28757
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39112 28699 39480 28708
rect 43112 28748 43480 28757
rect 43152 28708 43194 28748
rect 43234 28708 43276 28748
rect 43316 28708 43358 28748
rect 43398 28708 43440 28748
rect 43112 28699 43480 28708
rect 47112 28748 47480 28757
rect 47152 28708 47194 28748
rect 47234 28708 47276 28748
rect 47316 28708 47358 28748
rect 47398 28708 47440 28748
rect 47112 28699 47480 28708
rect 51112 28748 51480 28757
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51112 28699 51480 28708
rect 55112 28748 55480 28757
rect 55152 28708 55194 28748
rect 55234 28708 55276 28748
rect 55316 28708 55358 28748
rect 55398 28708 55440 28748
rect 55112 28699 55480 28708
rect 59112 28748 59480 28757
rect 59152 28708 59194 28748
rect 59234 28708 59276 28748
rect 59316 28708 59358 28748
rect 59398 28708 59440 28748
rect 59112 28699 59480 28708
rect 63112 28748 63480 28757
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63112 28699 63480 28708
rect 67112 28748 67480 28757
rect 67152 28708 67194 28748
rect 67234 28708 67276 28748
rect 67316 28708 67358 28748
rect 67398 28708 67440 28748
rect 67112 28699 67480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 8352 27992 8720 28001
rect 8392 27952 8434 27992
rect 8474 27952 8516 27992
rect 8556 27952 8598 27992
rect 8638 27952 8680 27992
rect 8352 27943 8720 27952
rect 12352 27992 12720 28001
rect 12392 27952 12434 27992
rect 12474 27952 12516 27992
rect 12556 27952 12598 27992
rect 12638 27952 12680 27992
rect 12352 27943 12720 27952
rect 16352 27992 16720 28001
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16352 27943 16720 27952
rect 20352 27992 20720 28001
rect 20392 27952 20434 27992
rect 20474 27952 20516 27992
rect 20556 27952 20598 27992
rect 20638 27952 20680 27992
rect 20352 27943 20720 27952
rect 24352 27992 24720 28001
rect 24392 27952 24434 27992
rect 24474 27952 24516 27992
rect 24556 27952 24598 27992
rect 24638 27952 24680 27992
rect 24352 27943 24720 27952
rect 28352 27992 28720 28001
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28352 27943 28720 27952
rect 32352 27992 32720 28001
rect 32392 27952 32434 27992
rect 32474 27952 32516 27992
rect 32556 27952 32598 27992
rect 32638 27952 32680 27992
rect 32352 27943 32720 27952
rect 36352 27992 36720 28001
rect 36392 27952 36434 27992
rect 36474 27952 36516 27992
rect 36556 27952 36598 27992
rect 36638 27952 36680 27992
rect 36352 27943 36720 27952
rect 40352 27992 40720 28001
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40352 27943 40720 27952
rect 44352 27992 44720 28001
rect 44392 27952 44434 27992
rect 44474 27952 44516 27992
rect 44556 27952 44598 27992
rect 44638 27952 44680 27992
rect 44352 27943 44720 27952
rect 48352 27992 48720 28001
rect 48392 27952 48434 27992
rect 48474 27952 48516 27992
rect 48556 27952 48598 27992
rect 48638 27952 48680 27992
rect 48352 27943 48720 27952
rect 52352 27992 52720 28001
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52352 27943 52720 27952
rect 56352 27992 56720 28001
rect 56392 27952 56434 27992
rect 56474 27952 56516 27992
rect 56556 27952 56598 27992
rect 56638 27952 56680 27992
rect 56352 27943 56720 27952
rect 60352 27992 60720 28001
rect 60392 27952 60434 27992
rect 60474 27952 60516 27992
rect 60556 27952 60598 27992
rect 60638 27952 60680 27992
rect 60352 27943 60720 27952
rect 64352 27992 64720 28001
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64352 27943 64720 27952
rect 68352 27992 68720 28001
rect 68392 27952 68434 27992
rect 68474 27952 68516 27992
rect 68556 27952 68598 27992
rect 68638 27952 68680 27992
rect 68352 27943 68720 27952
rect 70540 27740 70580 32059
rect 70732 31940 70772 31949
rect 70636 31900 70732 31940
rect 70636 31436 70676 31900
rect 70732 31891 70772 31900
rect 70828 31604 70868 32143
rect 70923 32108 70965 32117
rect 70923 32068 70924 32108
rect 70964 32068 70965 32108
rect 70923 32059 70965 32068
rect 71115 32108 71157 32117
rect 71115 32068 71116 32108
rect 71156 32068 71157 32108
rect 71115 32059 71157 32068
rect 71212 32108 71252 32740
rect 71403 32360 71445 32369
rect 71403 32320 71404 32360
rect 71444 32320 71445 32360
rect 71403 32311 71445 32320
rect 71404 32226 71444 32311
rect 70924 31974 70964 32059
rect 70828 31555 70868 31564
rect 71116 31520 71156 32059
rect 71116 31471 71156 31480
rect 70676 31396 71060 31436
rect 70636 31387 70676 31396
rect 71020 31352 71060 31396
rect 71020 31303 71060 31312
rect 70348 27700 70676 27740
rect 69963 27656 70005 27665
rect 69963 27616 69964 27656
rect 70004 27616 70005 27656
rect 69963 27607 70005 27616
rect 70156 27656 70196 27665
rect 70348 27656 70388 27700
rect 70196 27616 70388 27656
rect 70156 27607 70196 27616
rect 69964 27522 70004 27607
rect 70348 27488 70388 27616
rect 70540 27572 70580 27581
rect 70348 27439 70388 27448
rect 70444 27532 70540 27572
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 7112 27236 7480 27245
rect 7152 27196 7194 27236
rect 7234 27196 7276 27236
rect 7316 27196 7358 27236
rect 7398 27196 7440 27236
rect 7112 27187 7480 27196
rect 11112 27236 11480 27245
rect 11152 27196 11194 27236
rect 11234 27196 11276 27236
rect 11316 27196 11358 27236
rect 11398 27196 11440 27236
rect 11112 27187 11480 27196
rect 15112 27236 15480 27245
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15112 27187 15480 27196
rect 19112 27236 19480 27245
rect 19152 27196 19194 27236
rect 19234 27196 19276 27236
rect 19316 27196 19358 27236
rect 19398 27196 19440 27236
rect 19112 27187 19480 27196
rect 23112 27236 23480 27245
rect 23152 27196 23194 27236
rect 23234 27196 23276 27236
rect 23316 27196 23358 27236
rect 23398 27196 23440 27236
rect 23112 27187 23480 27196
rect 27112 27236 27480 27245
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27112 27187 27480 27196
rect 31112 27236 31480 27245
rect 31152 27196 31194 27236
rect 31234 27196 31276 27236
rect 31316 27196 31358 27236
rect 31398 27196 31440 27236
rect 31112 27187 31480 27196
rect 35112 27236 35480 27245
rect 35152 27196 35194 27236
rect 35234 27196 35276 27236
rect 35316 27196 35358 27236
rect 35398 27196 35440 27236
rect 35112 27187 35480 27196
rect 39112 27236 39480 27245
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39112 27187 39480 27196
rect 43112 27236 43480 27245
rect 43152 27196 43194 27236
rect 43234 27196 43276 27236
rect 43316 27196 43358 27236
rect 43398 27196 43440 27236
rect 43112 27187 43480 27196
rect 47112 27236 47480 27245
rect 47152 27196 47194 27236
rect 47234 27196 47276 27236
rect 47316 27196 47358 27236
rect 47398 27196 47440 27236
rect 47112 27187 47480 27196
rect 51112 27236 51480 27245
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51112 27187 51480 27196
rect 55112 27236 55480 27245
rect 55152 27196 55194 27236
rect 55234 27196 55276 27236
rect 55316 27196 55358 27236
rect 55398 27196 55440 27236
rect 55112 27187 55480 27196
rect 59112 27236 59480 27245
rect 59152 27196 59194 27236
rect 59234 27196 59276 27236
rect 59316 27196 59358 27236
rect 59398 27196 59440 27236
rect 59112 27187 59480 27196
rect 63112 27236 63480 27245
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63112 27187 63480 27196
rect 67112 27236 67480 27245
rect 67152 27196 67194 27236
rect 67234 27196 67276 27236
rect 67316 27196 67358 27236
rect 67398 27196 67440 27236
rect 67112 27187 67480 27196
rect 69772 26900 69812 26911
rect 69772 26825 69812 26860
rect 70348 26900 70388 26911
rect 70348 26825 70388 26860
rect 69771 26816 69813 26825
rect 69771 26776 69772 26816
rect 69812 26776 69813 26816
rect 69771 26767 69813 26776
rect 70347 26816 70389 26825
rect 70347 26776 70348 26816
rect 70388 26776 70389 26816
rect 70347 26767 70389 26776
rect 69963 26732 70005 26741
rect 69963 26692 69964 26732
rect 70004 26692 70005 26732
rect 69963 26683 70005 26692
rect 69964 26648 70004 26683
rect 69964 26597 70004 26608
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 8352 26480 8720 26489
rect 8392 26440 8434 26480
rect 8474 26440 8516 26480
rect 8556 26440 8598 26480
rect 8638 26440 8680 26480
rect 8352 26431 8720 26440
rect 12352 26480 12720 26489
rect 12392 26440 12434 26480
rect 12474 26440 12516 26480
rect 12556 26440 12598 26480
rect 12638 26440 12680 26480
rect 12352 26431 12720 26440
rect 16352 26480 16720 26489
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16352 26431 16720 26440
rect 20352 26480 20720 26489
rect 20392 26440 20434 26480
rect 20474 26440 20516 26480
rect 20556 26440 20598 26480
rect 20638 26440 20680 26480
rect 20352 26431 20720 26440
rect 24352 26480 24720 26489
rect 24392 26440 24434 26480
rect 24474 26440 24516 26480
rect 24556 26440 24598 26480
rect 24638 26440 24680 26480
rect 24352 26431 24720 26440
rect 28352 26480 28720 26489
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28352 26431 28720 26440
rect 32352 26480 32720 26489
rect 32392 26440 32434 26480
rect 32474 26440 32516 26480
rect 32556 26440 32598 26480
rect 32638 26440 32680 26480
rect 32352 26431 32720 26440
rect 36352 26480 36720 26489
rect 36392 26440 36434 26480
rect 36474 26440 36516 26480
rect 36556 26440 36598 26480
rect 36638 26440 36680 26480
rect 36352 26431 36720 26440
rect 40352 26480 40720 26489
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40352 26431 40720 26440
rect 44352 26480 44720 26489
rect 44392 26440 44434 26480
rect 44474 26440 44516 26480
rect 44556 26440 44598 26480
rect 44638 26440 44680 26480
rect 44352 26431 44720 26440
rect 48352 26480 48720 26489
rect 48392 26440 48434 26480
rect 48474 26440 48516 26480
rect 48556 26440 48598 26480
rect 48638 26440 48680 26480
rect 48352 26431 48720 26440
rect 52352 26480 52720 26489
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52352 26431 52720 26440
rect 56352 26480 56720 26489
rect 56392 26440 56434 26480
rect 56474 26440 56516 26480
rect 56556 26440 56598 26480
rect 56638 26440 56680 26480
rect 56352 26431 56720 26440
rect 60352 26480 60720 26489
rect 60392 26440 60434 26480
rect 60474 26440 60516 26480
rect 60556 26440 60598 26480
rect 60638 26440 60680 26480
rect 60352 26431 60720 26440
rect 64352 26480 64720 26489
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64352 26431 64720 26440
rect 68352 26480 68720 26489
rect 68392 26440 68434 26480
rect 68474 26440 68516 26480
rect 68556 26440 68598 26480
rect 68638 26440 68680 26480
rect 68352 26431 68720 26440
rect 70444 26321 70484 27532
rect 70540 27523 70580 27532
rect 70540 26648 70580 26657
rect 70540 26405 70580 26608
rect 70539 26396 70581 26405
rect 70539 26356 70540 26396
rect 70580 26356 70581 26396
rect 70539 26347 70581 26356
rect 69291 26312 69333 26321
rect 69291 26272 69292 26312
rect 69332 26272 69333 26312
rect 69291 26263 69333 26272
rect 70443 26312 70485 26321
rect 70443 26272 70444 26312
rect 70484 26272 70485 26312
rect 70443 26263 70485 26272
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 7112 25724 7480 25733
rect 7152 25684 7194 25724
rect 7234 25684 7276 25724
rect 7316 25684 7358 25724
rect 7398 25684 7440 25724
rect 7112 25675 7480 25684
rect 11112 25724 11480 25733
rect 11152 25684 11194 25724
rect 11234 25684 11276 25724
rect 11316 25684 11358 25724
rect 11398 25684 11440 25724
rect 11112 25675 11480 25684
rect 15112 25724 15480 25733
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15112 25675 15480 25684
rect 19112 25724 19480 25733
rect 19152 25684 19194 25724
rect 19234 25684 19276 25724
rect 19316 25684 19358 25724
rect 19398 25684 19440 25724
rect 19112 25675 19480 25684
rect 23112 25724 23480 25733
rect 23152 25684 23194 25724
rect 23234 25684 23276 25724
rect 23316 25684 23358 25724
rect 23398 25684 23440 25724
rect 23112 25675 23480 25684
rect 27112 25724 27480 25733
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27112 25675 27480 25684
rect 31112 25724 31480 25733
rect 31152 25684 31194 25724
rect 31234 25684 31276 25724
rect 31316 25684 31358 25724
rect 31398 25684 31440 25724
rect 31112 25675 31480 25684
rect 35112 25724 35480 25733
rect 35152 25684 35194 25724
rect 35234 25684 35276 25724
rect 35316 25684 35358 25724
rect 35398 25684 35440 25724
rect 35112 25675 35480 25684
rect 39112 25724 39480 25733
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39112 25675 39480 25684
rect 43112 25724 43480 25733
rect 43152 25684 43194 25724
rect 43234 25684 43276 25724
rect 43316 25684 43358 25724
rect 43398 25684 43440 25724
rect 43112 25675 43480 25684
rect 47112 25724 47480 25733
rect 47152 25684 47194 25724
rect 47234 25684 47276 25724
rect 47316 25684 47358 25724
rect 47398 25684 47440 25724
rect 47112 25675 47480 25684
rect 51112 25724 51480 25733
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51112 25675 51480 25684
rect 55112 25724 55480 25733
rect 55152 25684 55194 25724
rect 55234 25684 55276 25724
rect 55316 25684 55358 25724
rect 55398 25684 55440 25724
rect 55112 25675 55480 25684
rect 59112 25724 59480 25733
rect 59152 25684 59194 25724
rect 59234 25684 59276 25724
rect 59316 25684 59358 25724
rect 59398 25684 59440 25724
rect 59112 25675 59480 25684
rect 63112 25724 63480 25733
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63112 25675 63480 25684
rect 67112 25724 67480 25733
rect 67152 25684 67194 25724
rect 67234 25684 67276 25724
rect 67316 25684 67358 25724
rect 67398 25684 67440 25724
rect 67112 25675 67480 25684
rect 652 25304 692 25313
rect 652 24977 692 25264
rect 843 25304 885 25313
rect 843 25264 844 25304
rect 884 25264 885 25304
rect 843 25255 885 25264
rect 844 25170 884 25255
rect 651 24968 693 24977
rect 651 24928 652 24968
rect 692 24928 693 24968
rect 651 24919 693 24928
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 8352 24968 8720 24977
rect 8392 24928 8434 24968
rect 8474 24928 8516 24968
rect 8556 24928 8598 24968
rect 8638 24928 8680 24968
rect 8352 24919 8720 24928
rect 12352 24968 12720 24977
rect 12392 24928 12434 24968
rect 12474 24928 12516 24968
rect 12556 24928 12598 24968
rect 12638 24928 12680 24968
rect 12352 24919 12720 24928
rect 16352 24968 16720 24977
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16352 24919 16720 24928
rect 20352 24968 20720 24977
rect 20392 24928 20434 24968
rect 20474 24928 20516 24968
rect 20556 24928 20598 24968
rect 20638 24928 20680 24968
rect 20352 24919 20720 24928
rect 24352 24968 24720 24977
rect 24392 24928 24434 24968
rect 24474 24928 24516 24968
rect 24556 24928 24598 24968
rect 24638 24928 24680 24968
rect 24352 24919 24720 24928
rect 28352 24968 28720 24977
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28352 24919 28720 24928
rect 32352 24968 32720 24977
rect 32392 24928 32434 24968
rect 32474 24928 32516 24968
rect 32556 24928 32598 24968
rect 32638 24928 32680 24968
rect 32352 24919 32720 24928
rect 36352 24968 36720 24977
rect 36392 24928 36434 24968
rect 36474 24928 36516 24968
rect 36556 24928 36598 24968
rect 36638 24928 36680 24968
rect 36352 24919 36720 24928
rect 40352 24968 40720 24977
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40352 24919 40720 24928
rect 44352 24968 44720 24977
rect 44392 24928 44434 24968
rect 44474 24928 44516 24968
rect 44556 24928 44598 24968
rect 44638 24928 44680 24968
rect 44352 24919 44720 24928
rect 48352 24968 48720 24977
rect 48392 24928 48434 24968
rect 48474 24928 48516 24968
rect 48556 24928 48598 24968
rect 48638 24928 48680 24968
rect 48352 24919 48720 24928
rect 52352 24968 52720 24977
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52352 24919 52720 24928
rect 56352 24968 56720 24977
rect 56392 24928 56434 24968
rect 56474 24928 56516 24968
rect 56556 24928 56598 24968
rect 56638 24928 56680 24968
rect 56352 24919 56720 24928
rect 60352 24968 60720 24977
rect 60392 24928 60434 24968
rect 60474 24928 60516 24968
rect 60556 24928 60598 24968
rect 60638 24928 60680 24968
rect 60352 24919 60720 24928
rect 64352 24968 64720 24977
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64352 24919 64720 24928
rect 68352 24968 68720 24977
rect 68392 24928 68434 24968
rect 68474 24928 68516 24968
rect 68556 24928 68598 24968
rect 68638 24928 68680 24968
rect 68352 24919 68720 24928
rect 652 24632 692 24641
rect 652 24137 692 24592
rect 843 24632 885 24641
rect 843 24592 844 24632
rect 884 24592 885 24632
rect 843 24583 885 24592
rect 844 24498 884 24583
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 7112 24212 7480 24221
rect 7152 24172 7194 24212
rect 7234 24172 7276 24212
rect 7316 24172 7358 24212
rect 7398 24172 7440 24212
rect 7112 24163 7480 24172
rect 11112 24212 11480 24221
rect 11152 24172 11194 24212
rect 11234 24172 11276 24212
rect 11316 24172 11358 24212
rect 11398 24172 11440 24212
rect 11112 24163 11480 24172
rect 15112 24212 15480 24221
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15112 24163 15480 24172
rect 19112 24212 19480 24221
rect 19152 24172 19194 24212
rect 19234 24172 19276 24212
rect 19316 24172 19358 24212
rect 19398 24172 19440 24212
rect 19112 24163 19480 24172
rect 23112 24212 23480 24221
rect 23152 24172 23194 24212
rect 23234 24172 23276 24212
rect 23316 24172 23358 24212
rect 23398 24172 23440 24212
rect 23112 24163 23480 24172
rect 27112 24212 27480 24221
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27112 24163 27480 24172
rect 31112 24212 31480 24221
rect 31152 24172 31194 24212
rect 31234 24172 31276 24212
rect 31316 24172 31358 24212
rect 31398 24172 31440 24212
rect 31112 24163 31480 24172
rect 35112 24212 35480 24221
rect 35152 24172 35194 24212
rect 35234 24172 35276 24212
rect 35316 24172 35358 24212
rect 35398 24172 35440 24212
rect 35112 24163 35480 24172
rect 39112 24212 39480 24221
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39112 24163 39480 24172
rect 43112 24212 43480 24221
rect 43152 24172 43194 24212
rect 43234 24172 43276 24212
rect 43316 24172 43358 24212
rect 43398 24172 43440 24212
rect 43112 24163 43480 24172
rect 47112 24212 47480 24221
rect 47152 24172 47194 24212
rect 47234 24172 47276 24212
rect 47316 24172 47358 24212
rect 47398 24172 47440 24212
rect 47112 24163 47480 24172
rect 51112 24212 51480 24221
rect 51152 24172 51194 24212
rect 51234 24172 51276 24212
rect 51316 24172 51358 24212
rect 51398 24172 51440 24212
rect 51112 24163 51480 24172
rect 55112 24212 55480 24221
rect 55152 24172 55194 24212
rect 55234 24172 55276 24212
rect 55316 24172 55358 24212
rect 55398 24172 55440 24212
rect 55112 24163 55480 24172
rect 59112 24212 59480 24221
rect 59152 24172 59194 24212
rect 59234 24172 59276 24212
rect 59316 24172 59358 24212
rect 59398 24172 59440 24212
rect 59112 24163 59480 24172
rect 63112 24212 63480 24221
rect 63152 24172 63194 24212
rect 63234 24172 63276 24212
rect 63316 24172 63358 24212
rect 63398 24172 63440 24212
rect 63112 24163 63480 24172
rect 67112 24212 67480 24221
rect 67152 24172 67194 24212
rect 67234 24172 67276 24212
rect 67316 24172 67358 24212
rect 67398 24172 67440 24212
rect 67112 24163 67480 24172
rect 651 24128 693 24137
rect 651 24088 652 24128
rect 692 24088 693 24128
rect 651 24079 693 24088
rect 652 23792 692 23801
rect 652 23297 692 23752
rect 843 23792 885 23801
rect 843 23752 844 23792
rect 884 23752 885 23792
rect 843 23743 885 23752
rect 2091 23792 2133 23801
rect 2091 23752 2092 23792
rect 2132 23752 2133 23792
rect 2091 23743 2133 23752
rect 844 23658 884 23743
rect 2092 23297 2132 23743
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 8352 23456 8720 23465
rect 8392 23416 8434 23456
rect 8474 23416 8516 23456
rect 8556 23416 8598 23456
rect 8638 23416 8680 23456
rect 8352 23407 8720 23416
rect 12352 23456 12720 23465
rect 12392 23416 12434 23456
rect 12474 23416 12516 23456
rect 12556 23416 12598 23456
rect 12638 23416 12680 23456
rect 12352 23407 12720 23416
rect 16352 23456 16720 23465
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16352 23407 16720 23416
rect 20352 23456 20720 23465
rect 20392 23416 20434 23456
rect 20474 23416 20516 23456
rect 20556 23416 20598 23456
rect 20638 23416 20680 23456
rect 20352 23407 20720 23416
rect 24352 23456 24720 23465
rect 24392 23416 24434 23456
rect 24474 23416 24516 23456
rect 24556 23416 24598 23456
rect 24638 23416 24680 23456
rect 24352 23407 24720 23416
rect 28352 23456 28720 23465
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28352 23407 28720 23416
rect 32352 23456 32720 23465
rect 32392 23416 32434 23456
rect 32474 23416 32516 23456
rect 32556 23416 32598 23456
rect 32638 23416 32680 23456
rect 32352 23407 32720 23416
rect 36352 23456 36720 23465
rect 36392 23416 36434 23456
rect 36474 23416 36516 23456
rect 36556 23416 36598 23456
rect 36638 23416 36680 23456
rect 36352 23407 36720 23416
rect 40352 23456 40720 23465
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40352 23407 40720 23416
rect 44352 23456 44720 23465
rect 44392 23416 44434 23456
rect 44474 23416 44516 23456
rect 44556 23416 44598 23456
rect 44638 23416 44680 23456
rect 44352 23407 44720 23416
rect 48352 23456 48720 23465
rect 48392 23416 48434 23456
rect 48474 23416 48516 23456
rect 48556 23416 48598 23456
rect 48638 23416 48680 23456
rect 48352 23407 48720 23416
rect 52352 23456 52720 23465
rect 52392 23416 52434 23456
rect 52474 23416 52516 23456
rect 52556 23416 52598 23456
rect 52638 23416 52680 23456
rect 52352 23407 52720 23416
rect 56352 23456 56720 23465
rect 56392 23416 56434 23456
rect 56474 23416 56516 23456
rect 56556 23416 56598 23456
rect 56638 23416 56680 23456
rect 56352 23407 56720 23416
rect 60352 23456 60720 23465
rect 60392 23416 60434 23456
rect 60474 23416 60516 23456
rect 60556 23416 60598 23456
rect 60638 23416 60680 23456
rect 60352 23407 60720 23416
rect 64352 23456 64720 23465
rect 64392 23416 64434 23456
rect 64474 23416 64516 23456
rect 64556 23416 64598 23456
rect 64638 23416 64680 23456
rect 64352 23407 64720 23416
rect 68352 23456 68720 23465
rect 68392 23416 68434 23456
rect 68474 23416 68516 23456
rect 68556 23416 68598 23456
rect 68638 23416 68680 23456
rect 68352 23407 68720 23416
rect 69292 23297 69332 26263
rect 70444 25397 70484 26263
rect 70636 26153 70676 27700
rect 70923 27656 70965 27665
rect 70923 27616 70924 27656
rect 70964 27616 71156 27656
rect 70923 27607 70965 27616
rect 70924 27522 70964 27607
rect 71020 27404 71060 27413
rect 70732 26900 70772 26911
rect 70732 26825 70772 26860
rect 70731 26816 70773 26825
rect 70731 26776 70732 26816
rect 70772 26776 70773 26816
rect 70731 26767 70773 26776
rect 70924 26648 70964 26657
rect 70828 26608 70924 26648
rect 70828 26237 70868 26608
rect 70924 26599 70964 26608
rect 71020 26480 71060 27364
rect 71116 26900 71156 27616
rect 71116 26825 71156 26860
rect 71212 27572 71252 32068
rect 71115 26816 71157 26825
rect 71115 26776 71116 26816
rect 71156 26776 71157 26816
rect 71115 26767 71157 26776
rect 71020 26440 71156 26480
rect 71019 26312 71061 26321
rect 71019 26272 71020 26312
rect 71060 26272 71061 26312
rect 71019 26263 71061 26272
rect 70827 26228 70869 26237
rect 70827 26188 70828 26228
rect 70868 26188 70869 26228
rect 70827 26179 70869 26188
rect 71020 26178 71060 26263
rect 71116 26153 71156 26440
rect 70635 26144 70677 26153
rect 70635 26104 70636 26144
rect 70676 26104 70677 26144
rect 70635 26095 70677 26104
rect 70923 26144 70965 26153
rect 70923 26104 70924 26144
rect 70964 26104 70965 26144
rect 70923 26095 70965 26104
rect 71115 26144 71157 26153
rect 71115 26104 71116 26144
rect 71156 26104 71157 26144
rect 71212 26144 71252 27532
rect 71404 27404 71444 27413
rect 71308 26648 71348 26659
rect 71404 26657 71444 27364
rect 71308 26573 71348 26608
rect 71403 26648 71445 26657
rect 71403 26608 71404 26648
rect 71444 26608 71445 26648
rect 71403 26599 71445 26608
rect 71307 26564 71349 26573
rect 71307 26524 71308 26564
rect 71348 26524 71349 26564
rect 71307 26515 71349 26524
rect 71403 26480 71445 26489
rect 71403 26440 71404 26480
rect 71444 26440 71445 26480
rect 71403 26431 71445 26440
rect 71404 26312 71444 26431
rect 71404 26263 71444 26272
rect 71308 26144 71348 26153
rect 71212 26104 71308 26144
rect 71115 26095 71157 26104
rect 70443 25388 70485 25397
rect 70443 25348 70444 25388
rect 70484 25348 70485 25388
rect 70443 25339 70485 25348
rect 70924 25313 70964 26095
rect 71308 25985 71348 26104
rect 71307 25976 71349 25985
rect 71307 25936 71308 25976
rect 71348 25936 71349 25976
rect 71307 25927 71349 25936
rect 70923 25304 70965 25313
rect 70923 25264 70924 25304
rect 70964 25264 70965 25304
rect 70923 25255 70965 25264
rect 71308 25229 71348 25927
rect 71307 25220 71349 25229
rect 71307 25180 71308 25220
rect 71348 25180 71349 25220
rect 71307 25171 71349 25180
rect 71788 24725 71828 33235
rect 73228 32957 73268 33580
rect 73612 33620 73652 33629
rect 73420 33452 73460 33461
rect 72363 32948 72405 32957
rect 72363 32908 72364 32948
rect 72404 32908 72405 32948
rect 72363 32899 72405 32908
rect 72651 32948 72693 32957
rect 72651 32908 72652 32948
rect 72692 32908 72693 32948
rect 72651 32899 72693 32908
rect 73035 32948 73077 32957
rect 73035 32908 73036 32948
rect 73076 32908 73077 32948
rect 73035 32899 73077 32908
rect 73227 32948 73269 32957
rect 73227 32908 73228 32948
rect 73268 32908 73269 32948
rect 73227 32899 73269 32908
rect 72267 32864 72309 32873
rect 72267 32824 72268 32864
rect 72308 32824 72309 32864
rect 72267 32815 72309 32824
rect 72364 32864 72404 32899
rect 72268 32192 72308 32815
rect 72364 32813 72404 32824
rect 72652 32814 72692 32899
rect 73036 32864 73076 32899
rect 73036 32813 73076 32824
rect 72460 32696 72500 32705
rect 72460 32537 72500 32656
rect 72844 32696 72884 32705
rect 72459 32528 72501 32537
rect 72459 32488 72460 32528
rect 72500 32488 72501 32528
rect 72459 32479 72501 32488
rect 72844 32369 72884 32656
rect 73132 32696 73172 32705
rect 73172 32656 73364 32696
rect 73132 32647 73172 32656
rect 73131 32528 73173 32537
rect 73131 32488 73132 32528
rect 73172 32488 73173 32528
rect 73131 32479 73173 32488
rect 72414 32360 72456 32369
rect 72414 32320 72415 32360
rect 72455 32320 72456 32360
rect 72414 32311 72456 32320
rect 72843 32360 72885 32369
rect 72843 32320 72844 32360
rect 72884 32320 72885 32360
rect 72843 32311 72885 32320
rect 72268 32152 72345 32192
rect 72305 31920 72345 32152
rect 72415 31920 72455 32311
rect 72814 32192 72856 32201
rect 72814 32152 72815 32192
rect 72855 32152 72856 32192
rect 72814 32143 72856 32152
rect 72704 32108 72746 32117
rect 72704 32068 72705 32108
rect 72745 32068 72746 32108
rect 72704 32059 72746 32068
rect 72705 31920 72745 32059
rect 72815 31920 72855 32143
rect 73132 32108 73172 32479
rect 73214 32360 73256 32369
rect 73214 32320 73215 32360
rect 73255 32320 73256 32360
rect 73214 32311 73256 32320
rect 73105 32068 73172 32108
rect 73105 31920 73145 32068
rect 73215 31920 73255 32311
rect 73324 32108 73364 32656
rect 73420 32192 73460 33412
rect 73612 32873 73652 33580
rect 74092 33620 74132 33648
rect 74187 33620 74229 33629
rect 74132 33580 74188 33620
rect 74228 33580 74229 33620
rect 74092 33571 74132 33580
rect 74187 33571 74229 33580
rect 74475 33620 74517 33629
rect 74475 33580 74476 33620
rect 74516 33580 74517 33620
rect 74475 33571 74517 33580
rect 74859 33620 74901 33629
rect 74859 33580 74860 33620
rect 74900 33580 74901 33620
rect 74859 33571 74901 33580
rect 75339 33620 75381 33629
rect 75819 33620 75861 33629
rect 75339 33580 75340 33620
rect 75380 33580 75476 33620
rect 75339 33571 75381 33580
rect 73804 33452 73844 33461
rect 73844 33412 74132 33452
rect 73804 33403 73844 33412
rect 73996 32873 74036 32958
rect 73611 32864 73653 32873
rect 73611 32824 73612 32864
rect 73652 32824 73653 32864
rect 73611 32815 73653 32824
rect 73995 32864 74037 32873
rect 73995 32824 73996 32864
rect 74036 32824 74037 32864
rect 73995 32815 74037 32824
rect 73708 32696 73748 32705
rect 73899 32696 73941 32705
rect 73748 32656 73844 32696
rect 73708 32647 73748 32656
rect 73420 32152 73655 32192
rect 73324 32068 73545 32108
rect 73505 31920 73545 32068
rect 73615 31920 73655 32152
rect 73804 32108 73844 32656
rect 73899 32656 73900 32696
rect 73940 32656 73941 32696
rect 73899 32647 73941 32656
rect 73900 32562 73940 32647
rect 74092 32108 74132 33412
rect 74188 33116 74228 33571
rect 74476 33486 74516 33571
rect 74860 33486 74900 33571
rect 75340 33486 75380 33571
rect 74188 32873 74228 33076
rect 74284 33452 74324 33461
rect 74187 32864 74229 32873
rect 74187 32824 74188 32864
rect 74228 32824 74229 32864
rect 74187 32815 74229 32824
rect 74187 32696 74229 32705
rect 74187 32656 74188 32696
rect 74228 32656 74229 32696
rect 74187 32647 74229 32656
rect 73804 32068 73945 32108
rect 73905 31920 73945 32068
rect 74015 32068 74132 32108
rect 74188 32108 74228 32647
rect 74284 32192 74324 33412
rect 74668 33452 74708 33461
rect 75052 33452 75092 33461
rect 74708 33412 74804 33452
rect 74668 33403 74708 33412
rect 74667 33284 74709 33293
rect 74667 33244 74668 33284
rect 74708 33244 74709 33284
rect 74667 33235 74709 33244
rect 74379 32948 74421 32957
rect 74379 32908 74380 32948
rect 74420 32908 74421 32948
rect 74379 32899 74421 32908
rect 74668 32948 74708 33235
rect 74668 32899 74708 32908
rect 74380 32814 74420 32899
rect 74667 32696 74709 32705
rect 74667 32656 74668 32696
rect 74708 32656 74709 32696
rect 74667 32647 74709 32656
rect 74284 32152 74455 32192
rect 74188 32068 74345 32108
rect 74015 31920 74055 32068
rect 74305 31920 74345 32068
rect 74415 31920 74455 32152
rect 74668 32108 74708 32647
rect 74764 32192 74804 33412
rect 75092 33412 75284 33452
rect 75052 33403 75092 33412
rect 74860 33032 74900 33043
rect 74860 32957 74900 32992
rect 74859 32948 74901 32957
rect 74859 32908 74860 32948
rect 74900 32908 74901 32948
rect 74859 32899 74901 32908
rect 75147 32948 75189 32957
rect 75147 32908 75148 32948
rect 75188 32908 75189 32948
rect 75147 32899 75189 32908
rect 75148 32864 75188 32899
rect 75148 32813 75188 32824
rect 75051 32696 75093 32705
rect 75051 32656 75052 32696
rect 75092 32656 75093 32696
rect 75051 32647 75093 32656
rect 75052 32562 75092 32647
rect 74764 32152 74855 32192
rect 74668 32068 74745 32108
rect 74705 31920 74745 32068
rect 74815 31920 74855 32152
rect 75104 32108 75146 32117
rect 75244 32108 75284 33412
rect 75436 33209 75476 33580
rect 75819 33580 75820 33620
rect 75860 33580 75861 33620
rect 75819 33571 75861 33580
rect 76203 33620 76245 33629
rect 76588 33620 76628 33629
rect 76203 33580 76204 33620
rect 76244 33580 76245 33620
rect 76203 33571 76245 33580
rect 76300 33580 76588 33620
rect 75820 33486 75860 33571
rect 75532 33452 75572 33461
rect 75435 33200 75477 33209
rect 75435 33160 75436 33200
rect 75476 33160 75477 33200
rect 75435 33151 75477 33160
rect 75436 32864 75476 33151
rect 75436 32815 75476 32824
rect 75340 32696 75380 32705
rect 75340 32117 75380 32656
rect 75435 32696 75477 32705
rect 75435 32656 75436 32696
rect 75476 32656 75477 32696
rect 75435 32647 75477 32656
rect 75436 32192 75476 32647
rect 75532 32276 75572 33412
rect 76012 33452 76052 33461
rect 76052 33412 76148 33452
rect 76012 33403 76052 33412
rect 76011 33032 76053 33041
rect 76011 32992 76012 33032
rect 76052 32992 76053 33032
rect 76011 32983 76053 32992
rect 75819 32948 75861 32957
rect 75819 32908 75820 32948
rect 75860 32908 75861 32948
rect 75819 32899 75861 32908
rect 75820 32814 75860 32899
rect 76012 32898 76052 32983
rect 75904 32276 75946 32285
rect 75532 32236 75655 32276
rect 75436 32152 75545 32192
rect 75104 32068 75105 32108
rect 75145 32068 75146 32108
rect 75104 32059 75146 32068
rect 75215 32068 75284 32108
rect 75339 32108 75381 32117
rect 75339 32068 75340 32108
rect 75380 32068 75381 32108
rect 75105 31920 75145 32059
rect 75215 31920 75255 32068
rect 75339 32059 75381 32068
rect 75505 31920 75545 32152
rect 75615 31920 75655 32236
rect 75904 32236 75905 32276
rect 75945 32236 75946 32276
rect 75904 32227 75946 32236
rect 75905 31920 75945 32227
rect 76108 32108 76148 33412
rect 76204 33125 76244 33571
rect 76300 33209 76340 33580
rect 76588 33571 76628 33580
rect 76972 33620 77012 33648
rect 77067 33620 77109 33629
rect 77012 33580 77068 33620
rect 77108 33580 77109 33620
rect 76972 33571 77012 33580
rect 77067 33571 77109 33580
rect 77451 33620 77493 33629
rect 77451 33580 77452 33620
rect 77492 33580 77493 33620
rect 77451 33571 77493 33580
rect 77835 33620 77877 33629
rect 77835 33580 77836 33620
rect 77876 33580 77877 33620
rect 77835 33571 77877 33580
rect 78220 33620 78260 33629
rect 76396 33452 76436 33461
rect 76780 33452 76820 33461
rect 76299 33200 76341 33209
rect 76299 33160 76300 33200
rect 76340 33160 76341 33200
rect 76299 33151 76341 33160
rect 76203 33116 76245 33125
rect 76203 33076 76204 33116
rect 76244 33076 76245 33116
rect 76203 33067 76245 33076
rect 76204 32873 76244 32958
rect 76203 32864 76245 32873
rect 76203 32824 76204 32864
rect 76244 32824 76245 32864
rect 76203 32815 76245 32824
rect 76300 32864 76340 33151
rect 76300 32815 76340 32824
rect 76299 32696 76341 32705
rect 76299 32656 76300 32696
rect 76340 32656 76341 32696
rect 76299 32647 76341 32656
rect 76015 32068 76148 32108
rect 76300 32108 76340 32647
rect 76396 32192 76436 33412
rect 76684 33412 76780 33452
rect 76587 33032 76629 33041
rect 76587 32992 76588 33032
rect 76628 32992 76629 33032
rect 76587 32983 76629 32992
rect 76588 32873 76628 32983
rect 76587 32864 76629 32873
rect 76587 32824 76588 32864
rect 76628 32824 76629 32864
rect 76587 32815 76629 32824
rect 76492 32696 76532 32705
rect 76492 32285 76532 32656
rect 76684 32444 76724 33412
rect 76780 33403 76820 33412
rect 77068 33116 77108 33571
rect 77452 33486 77492 33571
rect 77068 33067 77108 33076
rect 77164 33452 77204 33461
rect 76875 33032 76917 33041
rect 76875 32992 76876 33032
rect 76916 32992 76917 33032
rect 76875 32983 76917 32992
rect 76876 32873 76916 32983
rect 76875 32864 76917 32873
rect 76875 32824 76876 32864
rect 76916 32824 76917 32864
rect 76875 32815 76917 32824
rect 76971 32780 77013 32789
rect 76971 32740 76972 32780
rect 77012 32740 77013 32780
rect 76971 32731 77013 32740
rect 76779 32696 76821 32705
rect 76779 32656 76780 32696
rect 76820 32656 76821 32696
rect 76779 32647 76821 32656
rect 76780 32562 76820 32647
rect 76684 32404 76820 32444
rect 76780 32360 76820 32404
rect 76780 32320 76855 32360
rect 76491 32276 76533 32285
rect 76491 32236 76492 32276
rect 76532 32236 76533 32276
rect 76491 32227 76533 32236
rect 76396 32152 76455 32192
rect 76300 32068 76345 32108
rect 76015 31920 76055 32068
rect 76305 31920 76345 32068
rect 76415 31920 76455 32152
rect 76704 32108 76746 32117
rect 76704 32068 76705 32108
rect 76745 32068 76746 32108
rect 76704 32059 76746 32068
rect 76705 31920 76745 32059
rect 76815 31920 76855 32320
rect 76972 32117 77012 32731
rect 77067 32192 77109 32201
rect 77164 32192 77204 33412
rect 77644 33452 77684 33461
rect 77451 33032 77493 33041
rect 77451 32992 77452 33032
rect 77492 32992 77493 33032
rect 77451 32983 77493 32992
rect 77259 32948 77301 32957
rect 77259 32908 77260 32948
rect 77300 32908 77301 32948
rect 77259 32899 77301 32908
rect 77260 32814 77300 32899
rect 77452 32864 77492 32983
rect 77548 32873 77588 32958
rect 77452 32815 77492 32824
rect 77547 32864 77589 32873
rect 77547 32824 77548 32864
rect 77588 32824 77589 32864
rect 77547 32815 77589 32824
rect 77504 32360 77546 32369
rect 77504 32320 77505 32360
rect 77545 32320 77546 32360
rect 77504 32311 77546 32320
rect 77067 32152 77068 32192
rect 77108 32152 77116 32192
rect 77164 32152 77255 32192
rect 77067 32143 77116 32152
rect 76971 32108 77013 32117
rect 76971 32068 76972 32108
rect 77012 32068 77013 32108
rect 77076 32108 77116 32143
rect 77076 32068 77145 32108
rect 76971 32059 77013 32068
rect 77105 31920 77145 32068
rect 77215 31920 77255 32152
rect 77505 31920 77545 32311
rect 77644 32108 77684 33412
rect 77836 33041 77876 33571
rect 78028 33452 78068 33461
rect 77932 33412 78028 33452
rect 77835 33032 77877 33041
rect 77835 32992 77836 33032
rect 77876 32992 77877 33032
rect 77835 32983 77877 32992
rect 77836 32864 77876 32983
rect 77836 32815 77876 32824
rect 77740 32696 77780 32705
rect 77740 32201 77780 32656
rect 77835 32696 77877 32705
rect 77835 32656 77836 32696
rect 77876 32656 77877 32696
rect 77835 32647 77877 32656
rect 77739 32192 77781 32201
rect 77739 32152 77740 32192
rect 77780 32152 77781 32192
rect 77836 32192 77876 32647
rect 77932 32276 77972 33412
rect 78028 33403 78068 33412
rect 78123 33032 78165 33041
rect 78220 33032 78260 33580
rect 78603 33620 78645 33629
rect 78603 33580 78604 33620
rect 78644 33580 78645 33620
rect 78603 33571 78645 33580
rect 78987 33620 79029 33629
rect 78987 33580 78988 33620
rect 79028 33580 79029 33620
rect 78987 33571 79029 33580
rect 79371 33620 79413 33629
rect 79755 33620 79797 33629
rect 79371 33580 79372 33620
rect 79412 33580 79508 33620
rect 79371 33571 79413 33580
rect 78604 33486 78644 33571
rect 78412 33452 78452 33461
rect 78796 33452 78836 33461
rect 78452 33412 78548 33452
rect 78412 33403 78452 33412
rect 78123 32992 78124 33032
rect 78164 32992 78260 33032
rect 78411 33032 78453 33041
rect 78411 32992 78412 33032
rect 78452 32992 78453 33032
rect 78123 32983 78165 32992
rect 78411 32983 78453 32992
rect 78124 32864 78164 32983
rect 78316 32873 78356 32958
rect 78124 32815 78164 32824
rect 78315 32864 78357 32873
rect 78315 32824 78316 32864
rect 78356 32824 78357 32864
rect 78315 32815 78357 32824
rect 78412 32864 78452 32983
rect 78412 32815 78452 32824
rect 78028 32696 78068 32705
rect 78028 32453 78068 32656
rect 78027 32444 78069 32453
rect 78027 32404 78028 32444
rect 78068 32404 78069 32444
rect 78027 32395 78069 32404
rect 78304 32276 78346 32285
rect 77932 32236 78055 32276
rect 77836 32152 77945 32192
rect 77739 32143 77781 32152
rect 77615 32068 77684 32108
rect 77615 31920 77655 32068
rect 77905 31920 77945 32152
rect 78015 31920 78055 32236
rect 78304 32236 78305 32276
rect 78345 32236 78346 32276
rect 78304 32227 78346 32236
rect 78305 31920 78345 32227
rect 78508 32108 78548 33412
rect 78700 32957 78740 33042
rect 78699 32948 78741 32957
rect 78699 32908 78700 32948
rect 78740 32908 78741 32948
rect 78699 32899 78741 32908
rect 78699 32780 78741 32789
rect 78699 32740 78700 32780
rect 78740 32740 78741 32780
rect 78699 32731 78741 32740
rect 78700 32192 78740 32731
rect 78796 32192 78836 33412
rect 78892 33116 78932 33125
rect 78988 33116 79028 33571
rect 79372 33486 79412 33571
rect 79180 33452 79220 33461
rect 79220 33412 79316 33452
rect 79180 33403 79220 33412
rect 78932 33076 79028 33116
rect 78892 33067 78932 33076
rect 79083 33032 79125 33041
rect 79083 32992 79084 33032
rect 79124 32992 79125 33032
rect 79083 32983 79125 32992
rect 78987 32864 79029 32873
rect 78987 32824 78988 32864
rect 79028 32824 79029 32864
rect 78987 32815 79029 32824
rect 79084 32864 79124 32983
rect 79084 32815 79124 32824
rect 78988 32192 79028 32815
rect 79180 32696 79220 32705
rect 79180 32285 79220 32656
rect 79179 32276 79221 32285
rect 79179 32236 79180 32276
rect 79220 32236 79221 32276
rect 79179 32227 79221 32236
rect 78700 32152 78745 32192
rect 78796 32152 78855 32192
rect 78988 32152 79145 32192
rect 78415 32068 78548 32108
rect 78415 31920 78455 32068
rect 78705 31920 78745 32152
rect 78815 31920 78855 32152
rect 79105 31920 79145 32152
rect 79276 32108 79316 33412
rect 79371 32948 79413 32957
rect 79371 32908 79372 32948
rect 79412 32908 79413 32948
rect 79371 32899 79413 32908
rect 79372 32814 79412 32899
rect 79468 32864 79508 33580
rect 79755 33580 79756 33620
rect 79796 33580 79797 33620
rect 79755 33571 79797 33580
rect 80331 33620 80373 33629
rect 80331 33580 80332 33620
rect 80372 33580 80373 33620
rect 80331 33571 80373 33580
rect 80908 33620 80948 33631
rect 79468 32815 79508 32824
rect 79564 33452 79604 33461
rect 79467 32696 79509 32705
rect 79467 32656 79468 32696
rect 79508 32656 79509 32696
rect 79467 32647 79509 32656
rect 79215 32068 79316 32108
rect 79468 32108 79508 32647
rect 79564 32192 79604 33412
rect 79660 32873 79700 32958
rect 79756 32957 79796 33571
rect 80332 33486 80372 33571
rect 80908 33545 80948 33580
rect 81100 33620 81140 33629
rect 80523 33536 80565 33545
rect 80523 33496 80524 33536
rect 80564 33496 80565 33536
rect 80523 33487 80565 33496
rect 80907 33536 80949 33545
rect 80907 33496 80908 33536
rect 80948 33496 80949 33536
rect 80907 33487 80949 33496
rect 79948 33452 79988 33461
rect 79852 33412 79948 33452
rect 79755 32948 79797 32957
rect 79755 32908 79756 32948
rect 79796 32908 79797 32948
rect 79755 32899 79797 32908
rect 79659 32864 79701 32873
rect 79659 32824 79660 32864
rect 79700 32824 79701 32864
rect 79659 32815 79701 32824
rect 79756 32864 79796 32899
rect 79756 32814 79796 32824
rect 79755 32360 79797 32369
rect 79755 32320 79756 32360
rect 79796 32320 79797 32360
rect 79755 32311 79797 32320
rect 79564 32152 79655 32192
rect 79468 32068 79545 32108
rect 79215 31920 79255 32068
rect 79505 31920 79545 32068
rect 79615 31920 79655 32152
rect 79756 32108 79796 32311
rect 79852 32192 79892 33412
rect 79948 33403 79988 33412
rect 80044 32957 80084 32970
rect 80236 32957 80276 32959
rect 80043 32948 80085 32957
rect 80235 32948 80277 32957
rect 80043 32908 80044 32948
rect 80084 32908 80086 32948
rect 80043 32899 80086 32908
rect 80235 32908 80236 32948
rect 80276 32908 80277 32948
rect 80524 32948 80564 33487
rect 80716 33452 80756 33461
rect 80620 32957 80660 33042
rect 80619 32948 80661 32957
rect 80524 32908 80620 32948
rect 80660 32908 80661 32948
rect 80235 32899 80277 32908
rect 80619 32899 80661 32908
rect 80046 32877 80086 32899
rect 80046 32828 80086 32837
rect 80236 32864 80276 32899
rect 80236 32815 80276 32824
rect 80716 32780 80756 33412
rect 81100 33293 81140 33580
rect 81291 33620 81333 33629
rect 81291 33580 81292 33620
rect 81332 33580 81333 33620
rect 81291 33571 81333 33580
rect 81676 33620 81716 33631
rect 81292 33536 81332 33571
rect 81676 33545 81716 33580
rect 82060 33620 82100 33631
rect 82444 33629 82484 33714
rect 82060 33545 82100 33580
rect 82443 33620 82485 33629
rect 82443 33580 82444 33620
rect 82484 33580 82485 33620
rect 82443 33571 82485 33580
rect 82828 33620 82868 33631
rect 82828 33545 82868 33580
rect 83115 33620 83157 33629
rect 83115 33580 83116 33620
rect 83156 33580 83157 33620
rect 83115 33571 83157 33580
rect 83212 33620 83252 33631
rect 87436 33629 87476 33714
rect 87820 33629 87860 33714
rect 88588 33629 88628 33714
rect 88972 33629 89012 33714
rect 90124 33629 90164 33714
rect 90508 33629 90548 33714
rect 81292 33485 81332 33496
rect 81675 33536 81717 33545
rect 81675 33496 81676 33536
rect 81716 33496 81717 33536
rect 81675 33487 81717 33496
rect 82059 33536 82101 33545
rect 82251 33536 82293 33545
rect 82059 33496 82060 33536
rect 82100 33496 82101 33536
rect 82059 33487 82101 33496
rect 82156 33496 82252 33536
rect 82292 33496 82293 33536
rect 81484 33452 81524 33461
rect 81388 33412 81484 33452
rect 81099 33284 81141 33293
rect 81099 33244 81100 33284
rect 81140 33244 81141 33284
rect 81099 33235 81141 33244
rect 81388 33116 81428 33412
rect 81484 33403 81524 33412
rect 81196 33076 81428 33116
rect 81004 32873 81044 32958
rect 81100 32957 81140 32959
rect 81099 32948 81141 32957
rect 81099 32908 81100 32948
rect 81140 32908 81141 32948
rect 81099 32899 81141 32908
rect 81003 32864 81045 32873
rect 81003 32824 81004 32864
rect 81044 32824 81045 32864
rect 81003 32815 81045 32824
rect 81100 32864 81140 32899
rect 81100 32815 81140 32824
rect 80428 32740 80756 32780
rect 79947 32696 79989 32705
rect 79947 32656 79948 32696
rect 79988 32656 79989 32696
rect 79947 32647 79989 32656
rect 80235 32696 80277 32705
rect 80235 32656 80236 32696
rect 80276 32656 80277 32696
rect 80235 32647 80277 32656
rect 80332 32696 80372 32705
rect 79948 32562 79988 32647
rect 80236 32192 80276 32647
rect 80332 32369 80372 32656
rect 80331 32360 80373 32369
rect 80331 32320 80332 32360
rect 80372 32320 80373 32360
rect 80331 32311 80373 32320
rect 79852 32152 80055 32192
rect 80236 32152 80345 32192
rect 79756 32068 79945 32108
rect 79905 31920 79945 32068
rect 80015 31920 80055 32152
rect 80305 31920 80345 32152
rect 80428 32108 80468 32740
rect 80812 32696 80852 32705
rect 80704 32360 80746 32369
rect 80704 32320 80705 32360
rect 80745 32320 80746 32360
rect 80704 32311 80746 32320
rect 80415 32068 80468 32108
rect 80415 31920 80455 32068
rect 80705 31920 80745 32311
rect 80812 32108 80852 32656
rect 81104 32276 81146 32285
rect 81104 32236 81105 32276
rect 81145 32236 81146 32276
rect 81104 32227 81146 32236
rect 80812 32068 80855 32108
rect 80815 31920 80855 32068
rect 81105 31920 81145 32227
rect 81196 32192 81236 33076
rect 81387 32948 81429 32957
rect 81387 32908 81388 32948
rect 81428 32908 81429 32948
rect 81387 32899 81429 32908
rect 81388 32864 81428 32899
rect 81388 32813 81428 32824
rect 81676 32864 81716 33487
rect 81868 33452 81908 33461
rect 81676 32815 81716 32824
rect 81772 33412 81868 33452
rect 81483 32780 81525 32789
rect 81483 32740 81484 32780
rect 81524 32740 81525 32780
rect 81483 32731 81525 32740
rect 81292 32696 81332 32705
rect 81292 32369 81332 32656
rect 81291 32360 81333 32369
rect 81291 32320 81292 32360
rect 81332 32320 81333 32360
rect 81291 32311 81333 32320
rect 81196 32152 81255 32192
rect 81215 31920 81255 32152
rect 81484 32108 81524 32731
rect 81580 32696 81620 32705
rect 81580 32285 81620 32656
rect 81579 32276 81621 32285
rect 81579 32236 81580 32276
rect 81620 32236 81621 32276
rect 81579 32227 81621 32236
rect 81772 32108 81812 33412
rect 81868 33403 81908 33412
rect 82060 32948 82100 32957
rect 82156 32948 82196 33496
rect 82251 33487 82293 33496
rect 82827 33536 82869 33545
rect 82827 33496 82828 33536
rect 82868 33496 82869 33536
rect 82827 33487 82869 33496
rect 82252 33402 82292 33487
rect 82636 33452 82676 33461
rect 82444 33412 82636 33452
rect 82100 32908 82196 32948
rect 82251 32948 82293 32957
rect 82251 32908 82252 32948
rect 82292 32908 82293 32948
rect 82060 32899 82100 32908
rect 82251 32899 82293 32908
rect 82252 32864 82292 32899
rect 82348 32873 82388 32958
rect 82252 32813 82292 32824
rect 82347 32864 82389 32873
rect 82347 32824 82348 32864
rect 82388 32824 82389 32864
rect 82347 32815 82389 32824
rect 81868 32696 81908 32705
rect 81868 32276 81908 32656
rect 82304 32360 82346 32369
rect 82304 32320 82305 32360
rect 82345 32320 82346 32360
rect 82304 32311 82346 32320
rect 81868 32236 82055 32276
rect 81484 32068 81545 32108
rect 81505 31920 81545 32068
rect 81615 32068 81812 32108
rect 81904 32108 81946 32117
rect 81904 32068 81905 32108
rect 81945 32068 81946 32108
rect 81615 31920 81655 32068
rect 81904 32059 81946 32068
rect 81905 31920 81945 32059
rect 82015 31920 82055 32236
rect 82305 31920 82345 32311
rect 82444 32108 82484 33412
rect 82636 33403 82676 33412
rect 82636 32864 82676 32873
rect 82828 32864 82868 33487
rect 83020 33452 83060 33461
rect 82924 32864 82964 32873
rect 82676 32824 82924 32864
rect 82636 32815 82676 32824
rect 82924 32815 82964 32824
rect 82540 32696 82580 32705
rect 82540 32117 82580 32656
rect 82635 32696 82677 32705
rect 82635 32656 82636 32696
rect 82676 32656 82677 32696
rect 82635 32647 82677 32656
rect 82828 32696 82868 32705
rect 82636 32192 82676 32647
rect 82828 32369 82868 32656
rect 82827 32360 82869 32369
rect 82827 32320 82828 32360
rect 82868 32320 82869 32360
rect 82827 32311 82869 32320
rect 83020 32192 83060 33412
rect 83116 33209 83156 33571
rect 83212 33545 83252 33580
rect 83596 33620 83636 33629
rect 83980 33620 84020 33629
rect 83211 33536 83253 33545
rect 83211 33496 83212 33536
rect 83252 33496 83253 33536
rect 83211 33487 83253 33496
rect 83499 33536 83541 33545
rect 83499 33496 83500 33536
rect 83540 33496 83541 33536
rect 83499 33487 83541 33496
rect 83404 33452 83444 33461
rect 83115 33200 83157 33209
rect 83115 33160 83116 33200
rect 83156 33160 83157 33200
rect 83115 33151 83157 33160
rect 83116 32948 83156 33151
rect 83307 33032 83349 33041
rect 83307 32992 83308 33032
rect 83348 32992 83349 33032
rect 83307 32983 83349 32992
rect 83116 32899 83156 32908
rect 83308 32898 83348 32983
rect 83115 32780 83157 32789
rect 83115 32740 83116 32780
rect 83156 32740 83157 32780
rect 83115 32731 83157 32740
rect 82636 32152 82745 32192
rect 82415 32068 82484 32108
rect 82539 32108 82581 32117
rect 82539 32068 82540 32108
rect 82580 32068 82581 32108
rect 82415 31920 82455 32068
rect 82539 32059 82581 32068
rect 82705 31920 82745 32152
rect 82815 32152 83060 32192
rect 82815 31920 82855 32152
rect 83116 32108 83156 32731
rect 83404 32108 83444 33412
rect 83500 32864 83540 33487
rect 83596 33125 83636 33580
rect 83884 33580 83980 33620
rect 83788 33452 83828 33461
rect 83692 33412 83788 33452
rect 83595 33116 83637 33125
rect 83595 33076 83596 33116
rect 83636 33076 83637 33116
rect 83595 33067 83637 33076
rect 83595 32948 83637 32957
rect 83595 32908 83596 32948
rect 83636 32908 83637 32948
rect 83595 32899 83637 32908
rect 83500 32815 83540 32824
rect 83596 32814 83636 32899
rect 83504 32360 83546 32369
rect 83504 32320 83505 32360
rect 83545 32320 83546 32360
rect 83504 32311 83546 32320
rect 83105 32068 83156 32108
rect 83215 32068 83444 32108
rect 83105 31920 83145 32068
rect 83215 31920 83255 32068
rect 83505 31920 83545 32311
rect 83692 32108 83732 33412
rect 83788 33403 83828 33412
rect 83884 33041 83924 33580
rect 83980 33571 84020 33580
rect 84364 33620 84404 33629
rect 84172 33452 84212 33461
rect 83980 33412 84172 33452
rect 83883 33032 83925 33041
rect 83883 32992 83884 33032
rect 83924 32992 83925 33032
rect 83883 32983 83925 32992
rect 83788 32873 83828 32958
rect 83787 32864 83829 32873
rect 83787 32824 83788 32864
rect 83828 32824 83829 32864
rect 83787 32815 83829 32824
rect 83884 32864 83924 32983
rect 83884 32815 83924 32824
rect 83883 32696 83925 32705
rect 83883 32656 83884 32696
rect 83924 32656 83925 32696
rect 83883 32647 83925 32656
rect 83615 32068 83732 32108
rect 83884 32108 83924 32647
rect 83980 32192 84020 33412
rect 84172 33403 84212 33412
rect 84171 33032 84213 33041
rect 84171 32992 84172 33032
rect 84212 32992 84213 33032
rect 84364 33032 84404 33580
rect 84748 33620 84788 33629
rect 84556 33452 84596 33461
rect 84459 33032 84501 33041
rect 84364 32992 84460 33032
rect 84500 32992 84501 33032
rect 84171 32983 84213 32992
rect 84459 32983 84501 32992
rect 84172 32864 84212 32983
rect 84172 32815 84212 32824
rect 84460 32864 84500 32983
rect 84460 32815 84500 32824
rect 84267 32780 84309 32789
rect 84267 32740 84268 32780
rect 84308 32740 84309 32780
rect 84267 32731 84309 32740
rect 84076 32696 84116 32705
rect 84076 32369 84116 32656
rect 84075 32360 84117 32369
rect 84075 32320 84076 32360
rect 84116 32320 84117 32360
rect 84268 32360 84308 32731
rect 84363 32696 84405 32705
rect 84363 32656 84364 32696
rect 84404 32656 84405 32696
rect 84363 32647 84405 32656
rect 84364 32562 84404 32647
rect 84268 32320 84345 32360
rect 84075 32311 84117 32320
rect 83980 32152 84055 32192
rect 83884 32068 83945 32108
rect 83615 31920 83655 32068
rect 83905 31920 83945 32068
rect 84015 31920 84055 32152
rect 84305 31920 84345 32320
rect 84556 32108 84596 33412
rect 84651 33200 84693 33209
rect 84651 33160 84652 33200
rect 84692 33160 84693 33200
rect 84651 33151 84693 33160
rect 84652 32948 84692 33151
rect 84748 33041 84788 33580
rect 85132 33620 85172 33629
rect 85516 33620 85556 33629
rect 84940 33452 84980 33461
rect 84747 33032 84789 33041
rect 84747 32992 84748 33032
rect 84788 32992 84789 33032
rect 84747 32983 84789 32992
rect 84844 33032 84884 33043
rect 84844 32957 84884 32992
rect 84652 32899 84692 32908
rect 84843 32948 84885 32957
rect 84843 32908 84844 32948
rect 84884 32908 84885 32948
rect 84843 32899 84885 32908
rect 84940 32780 84980 33412
rect 85132 33125 85172 33580
rect 85420 33580 85516 33620
rect 85324 33452 85364 33461
rect 85228 33412 85324 33452
rect 85131 33116 85173 33125
rect 85131 33076 85132 33116
rect 85172 33076 85173 33116
rect 85131 33067 85173 33076
rect 85035 33032 85077 33041
rect 85035 32992 85036 33032
rect 85076 32992 85077 33032
rect 85035 32983 85077 32992
rect 85036 32864 85076 32983
rect 85132 32873 85172 32958
rect 85036 32815 85076 32824
rect 85131 32864 85173 32873
rect 85131 32824 85132 32864
rect 85172 32824 85173 32864
rect 85131 32815 85173 32824
rect 84844 32740 84980 32780
rect 84415 32068 84596 32108
rect 84704 32108 84746 32117
rect 84844 32108 84884 32740
rect 85104 32360 85146 32369
rect 85104 32320 85105 32360
rect 85145 32320 85146 32360
rect 85104 32311 85146 32320
rect 84704 32068 84705 32108
rect 84745 32068 84746 32108
rect 84415 31920 84455 32068
rect 84704 32059 84746 32068
rect 84815 32068 84884 32108
rect 84705 31920 84745 32059
rect 84815 31920 84855 32068
rect 85105 31920 85145 32311
rect 85228 32108 85268 33412
rect 85324 33403 85364 33412
rect 85420 32873 85460 33580
rect 85516 33571 85556 33580
rect 85899 33620 85941 33629
rect 85899 33580 85900 33620
rect 85940 33580 85941 33620
rect 85899 33571 85941 33580
rect 86283 33620 86325 33629
rect 86283 33580 86284 33620
rect 86324 33580 86325 33620
rect 86283 33571 86325 33580
rect 86667 33620 86709 33629
rect 86667 33580 86668 33620
rect 86708 33580 86709 33620
rect 86667 33571 86709 33580
rect 87052 33620 87092 33629
rect 87435 33620 87477 33629
rect 85708 33452 85748 33461
rect 85516 33412 85708 33452
rect 85419 32864 85461 32873
rect 85419 32824 85420 32864
rect 85460 32824 85461 32864
rect 85419 32815 85461 32824
rect 85324 32696 85364 32705
rect 85324 32117 85364 32656
rect 85419 32696 85461 32705
rect 85419 32656 85420 32696
rect 85460 32656 85461 32696
rect 85419 32647 85461 32656
rect 85215 32068 85268 32108
rect 85323 32108 85365 32117
rect 85323 32068 85324 32108
rect 85364 32068 85365 32108
rect 85420 32108 85460 32647
rect 85516 32192 85556 33412
rect 85708 33403 85748 33412
rect 85900 33041 85940 33571
rect 86284 33486 86324 33571
rect 86668 33486 86708 33571
rect 87052 33461 87092 33580
rect 87340 33580 87436 33620
rect 87476 33580 87477 33620
rect 86092 33452 86132 33461
rect 86476 33452 86516 33461
rect 85899 33032 85941 33041
rect 85899 32992 85900 33032
rect 85940 32992 85941 33032
rect 85899 32983 85941 32992
rect 85708 32873 85748 32958
rect 85996 32873 86036 32958
rect 85707 32864 85749 32873
rect 85707 32824 85708 32864
rect 85748 32824 85749 32864
rect 85707 32815 85749 32824
rect 85995 32864 86037 32873
rect 85995 32824 85996 32864
rect 86036 32824 86037 32864
rect 85995 32815 86037 32824
rect 85899 32780 85941 32789
rect 85899 32740 85900 32780
rect 85940 32740 85941 32780
rect 85899 32731 85941 32740
rect 85612 32696 85652 32705
rect 85612 32369 85652 32656
rect 85900 32646 85940 32731
rect 85611 32360 85653 32369
rect 85611 32320 85612 32360
rect 85652 32320 85653 32360
rect 85611 32311 85653 32320
rect 85904 32360 85946 32369
rect 85904 32320 85905 32360
rect 85945 32320 85946 32360
rect 85904 32311 85946 32320
rect 85516 32152 85655 32192
rect 85420 32068 85545 32108
rect 85215 31920 85255 32068
rect 85323 32059 85365 32068
rect 85505 31920 85545 32068
rect 85615 31920 85655 32152
rect 85905 31920 85945 32311
rect 86092 32108 86132 33412
rect 86380 33412 86476 33452
rect 86283 33284 86325 33293
rect 86283 33244 86284 33284
rect 86324 33244 86325 33284
rect 86283 33235 86325 33244
rect 86284 32948 86324 33235
rect 86284 32899 86324 32908
rect 86283 32780 86325 32789
rect 86283 32740 86284 32780
rect 86324 32740 86325 32780
rect 86283 32731 86325 32740
rect 86284 32192 86324 32731
rect 86380 32276 86420 33412
rect 86476 33403 86516 33412
rect 86860 33452 86900 33461
rect 86860 33293 86900 33412
rect 87051 33452 87093 33461
rect 87051 33412 87052 33452
rect 87092 33412 87093 33452
rect 87051 33403 87093 33412
rect 87244 33452 87284 33461
rect 86859 33284 86901 33293
rect 86859 33244 86860 33284
rect 86900 33244 86901 33284
rect 86859 33235 86901 33244
rect 86475 33200 86517 33209
rect 86475 33160 86476 33200
rect 86516 33160 86517 33200
rect 86475 33151 86517 33160
rect 87051 33200 87093 33209
rect 87051 33160 87052 33200
rect 87092 33160 87093 33200
rect 87051 33151 87093 33160
rect 86476 33116 86516 33151
rect 86476 33065 86516 33076
rect 86859 33116 86901 33125
rect 86859 33076 86860 33116
rect 86900 33076 86901 33116
rect 86859 33067 86901 33076
rect 86667 33032 86709 33041
rect 86667 32992 86668 33032
rect 86708 32992 86709 33032
rect 86667 32983 86709 32992
rect 86668 32864 86708 32983
rect 86668 32815 86708 32824
rect 86667 32696 86709 32705
rect 86667 32656 86668 32696
rect 86708 32656 86709 32696
rect 86667 32647 86709 32656
rect 86764 32696 86804 32705
rect 86380 32236 86455 32276
rect 86284 32152 86345 32192
rect 86015 32068 86132 32108
rect 86015 31920 86055 32068
rect 86305 31920 86345 32152
rect 86415 31920 86455 32236
rect 86668 32192 86708 32647
rect 86764 32369 86804 32656
rect 86763 32360 86805 32369
rect 86763 32320 86764 32360
rect 86804 32320 86805 32360
rect 86763 32311 86805 32320
rect 86668 32152 86745 32192
rect 86705 31920 86745 32152
rect 86860 32108 86900 33067
rect 86955 32948 86997 32957
rect 86955 32908 86956 32948
rect 86996 32908 86997 32948
rect 86955 32899 86997 32908
rect 86956 32814 86996 32899
rect 87052 32864 87092 33151
rect 87244 33125 87284 33412
rect 87340 33209 87380 33580
rect 87435 33571 87477 33580
rect 87819 33620 87861 33629
rect 87819 33580 87820 33620
rect 87860 33580 87861 33620
rect 87819 33571 87861 33580
rect 88204 33620 88244 33629
rect 87628 33452 87668 33461
rect 88012 33452 88052 33461
rect 87436 33412 87628 33452
rect 87339 33200 87381 33209
rect 87339 33160 87340 33200
rect 87380 33160 87381 33200
rect 87339 33151 87381 33160
rect 87243 33116 87285 33125
rect 87243 33076 87244 33116
rect 87284 33076 87285 33116
rect 87243 33067 87285 33076
rect 87244 32873 87284 32958
rect 87052 32815 87092 32824
rect 87243 32864 87285 32873
rect 87243 32824 87244 32864
rect 87284 32824 87285 32864
rect 87243 32815 87285 32824
rect 87340 32864 87380 33151
rect 87340 32815 87380 32824
rect 87104 32360 87146 32369
rect 87104 32320 87105 32360
rect 87145 32320 87146 32360
rect 87104 32311 87146 32320
rect 86815 32068 86900 32108
rect 86815 31920 86855 32068
rect 87105 31920 87145 32311
rect 87436 32192 87476 33412
rect 87628 33403 87668 33412
rect 87724 33412 88012 33452
rect 87627 33200 87669 33209
rect 87627 33160 87628 33200
rect 87668 33160 87669 33200
rect 87627 33151 87669 33160
rect 87628 32864 87668 33151
rect 87628 32815 87668 32824
rect 87532 32696 87572 32705
rect 87532 32369 87572 32656
rect 87627 32696 87669 32705
rect 87627 32656 87628 32696
rect 87668 32656 87669 32696
rect 87627 32647 87669 32656
rect 87531 32360 87573 32369
rect 87531 32320 87532 32360
rect 87572 32320 87573 32360
rect 87531 32311 87573 32320
rect 87628 32192 87668 32647
rect 87215 32152 87476 32192
rect 87532 32152 87668 32192
rect 87215 31920 87255 32152
rect 87532 32108 87572 32152
rect 87724 32108 87764 33412
rect 88012 33403 88052 33412
rect 87915 33284 87957 33293
rect 87915 33244 87916 33284
rect 87956 33244 87957 33284
rect 87915 33235 87957 33244
rect 87916 32948 87956 33235
rect 88204 33200 88244 33580
rect 88587 33620 88629 33629
rect 88587 33580 88588 33620
rect 88628 33580 88629 33620
rect 88587 33571 88629 33580
rect 88971 33620 89013 33629
rect 88971 33580 88972 33620
rect 89012 33580 89013 33620
rect 88971 33571 89013 33580
rect 89355 33620 89397 33629
rect 89547 33620 89589 33629
rect 89355 33580 89356 33620
rect 89396 33580 89492 33620
rect 89355 33571 89397 33580
rect 89356 33486 89396 33571
rect 88396 33452 88436 33461
rect 88780 33452 88820 33461
rect 89164 33452 89204 33461
rect 88299 33200 88341 33209
rect 88204 33160 88300 33200
rect 88340 33160 88341 33200
rect 88299 33151 88341 33160
rect 88011 33116 88053 33125
rect 88011 33076 88012 33116
rect 88052 33076 88053 33116
rect 88011 33067 88053 33076
rect 87916 32899 87956 32908
rect 87915 32780 87957 32789
rect 87915 32740 87916 32780
rect 87956 32740 87957 32780
rect 87915 32731 87957 32740
rect 87916 32108 87956 32731
rect 88012 32192 88052 33067
rect 88107 33032 88149 33041
rect 88107 32992 88108 33032
rect 88148 32992 88149 33032
rect 88107 32983 88149 32992
rect 88108 32898 88148 32983
rect 88300 32864 88340 33151
rect 88396 33125 88436 33412
rect 88492 33412 88780 33452
rect 88395 33116 88437 33125
rect 88395 33076 88396 33116
rect 88436 33076 88437 33116
rect 88395 33067 88437 33076
rect 88395 32948 88437 32957
rect 88395 32908 88396 32948
rect 88436 32908 88437 32948
rect 88395 32899 88437 32908
rect 88300 32815 88340 32824
rect 88396 32814 88436 32899
rect 88012 32152 88055 32192
rect 87505 32068 87572 32108
rect 87615 32068 87764 32108
rect 87905 32068 87956 32108
rect 87505 31920 87545 32068
rect 87615 31920 87655 32068
rect 87905 31920 87945 32068
rect 88015 31920 88055 32152
rect 88304 32108 88346 32117
rect 88492 32108 88532 33412
rect 88780 33403 88820 33412
rect 88876 33412 89164 33452
rect 88683 33032 88725 33041
rect 88683 32992 88684 33032
rect 88724 32992 88725 33032
rect 88683 32983 88725 32992
rect 88588 32873 88628 32958
rect 88587 32864 88629 32873
rect 88587 32824 88588 32864
rect 88628 32824 88629 32864
rect 88587 32815 88629 32824
rect 88684 32864 88724 32983
rect 88684 32815 88724 32824
rect 88779 32864 88821 32873
rect 88779 32824 88780 32864
rect 88820 32824 88821 32864
rect 88779 32815 88821 32824
rect 88780 32192 88820 32815
rect 88304 32068 88305 32108
rect 88345 32068 88346 32108
rect 88304 32059 88346 32068
rect 88415 32068 88532 32108
rect 88705 32152 88820 32192
rect 88305 31920 88345 32059
rect 88415 31920 88455 32068
rect 88705 31920 88745 32152
rect 88876 32108 88916 33412
rect 89164 33403 89204 33412
rect 88971 33284 89013 33293
rect 88971 33244 88972 33284
rect 89012 33244 89013 33284
rect 88971 33235 89013 33244
rect 88972 32948 89012 33235
rect 89452 33041 89492 33580
rect 89547 33580 89548 33620
rect 89588 33580 89589 33620
rect 89547 33571 89589 33580
rect 89740 33620 89780 33629
rect 89548 33452 89588 33571
rect 89548 33293 89588 33412
rect 89547 33284 89589 33293
rect 89547 33244 89548 33284
rect 89588 33244 89589 33284
rect 89547 33235 89589 33244
rect 89740 33209 89780 33580
rect 90123 33620 90165 33629
rect 90123 33580 90124 33620
rect 90164 33580 90165 33620
rect 90123 33571 90165 33580
rect 90507 33620 90549 33629
rect 90507 33580 90508 33620
rect 90548 33580 90549 33620
rect 90507 33571 90549 33580
rect 90891 33620 90933 33629
rect 90891 33580 90892 33620
rect 90932 33580 90933 33620
rect 90891 33571 90933 33580
rect 91179 33620 91221 33629
rect 91179 33580 91180 33620
rect 91220 33580 91221 33620
rect 91179 33571 91221 33580
rect 91276 33620 91316 33739
rect 91276 33571 91316 33580
rect 90892 33486 90932 33571
rect 89932 33452 89972 33461
rect 90316 33452 90356 33461
rect 90700 33452 90740 33461
rect 91084 33452 91124 33461
rect 89836 33412 89932 33452
rect 89739 33200 89781 33209
rect 89739 33160 89740 33200
rect 89780 33160 89781 33200
rect 89739 33151 89781 33160
rect 89451 33032 89493 33041
rect 89451 32992 89452 33032
rect 89492 32992 89493 33032
rect 89451 32983 89493 32992
rect 89739 33032 89781 33041
rect 89739 32992 89740 33032
rect 89780 32992 89781 33032
rect 89739 32983 89781 32992
rect 88972 32899 89012 32908
rect 89067 32948 89109 32957
rect 89067 32908 89068 32948
rect 89108 32908 89109 32948
rect 89067 32899 89109 32908
rect 89068 32192 89108 32899
rect 89452 32864 89492 32983
rect 89644 32873 89684 32958
rect 89452 32815 89492 32824
rect 89643 32864 89685 32873
rect 89643 32824 89644 32864
rect 89684 32824 89685 32864
rect 89643 32815 89685 32824
rect 89740 32864 89780 32983
rect 89740 32815 89780 32824
rect 89164 32696 89204 32705
rect 89164 32276 89204 32656
rect 89356 32696 89396 32705
rect 89164 32236 89255 32276
rect 89068 32152 89145 32192
rect 88815 32068 88916 32108
rect 88815 31920 88855 32068
rect 89105 31920 89145 32152
rect 89215 31920 89255 32236
rect 89356 32117 89396 32656
rect 89836 32192 89876 33412
rect 89932 33403 89972 33412
rect 90124 33412 90316 33452
rect 89931 33032 89973 33041
rect 89931 32992 89932 33032
rect 89972 32992 89973 33032
rect 89931 32983 89973 32992
rect 89932 32864 89972 32983
rect 90027 32948 90069 32957
rect 90027 32908 90028 32948
rect 90068 32908 90069 32948
rect 90027 32899 90069 32908
rect 89932 32815 89972 32824
rect 90028 32814 90068 32899
rect 89931 32696 89973 32705
rect 89931 32656 89932 32696
rect 89972 32656 89973 32696
rect 89931 32647 89973 32656
rect 89615 32152 89876 32192
rect 89355 32108 89397 32117
rect 89355 32068 89356 32108
rect 89396 32068 89397 32108
rect 89355 32059 89397 32068
rect 89504 32108 89546 32117
rect 89504 32068 89505 32108
rect 89545 32068 89546 32108
rect 89504 32059 89546 32068
rect 89505 31920 89545 32059
rect 89615 31920 89655 32152
rect 89932 32108 89972 32647
rect 90124 32108 90164 33412
rect 90316 33403 90356 33412
rect 90508 33412 90700 33452
rect 90315 33284 90357 33293
rect 90315 33244 90316 33284
rect 90356 33244 90357 33284
rect 90315 33235 90357 33244
rect 90316 32864 90356 33235
rect 90316 32815 90356 32824
rect 90411 32864 90453 32873
rect 90411 32824 90412 32864
rect 90452 32824 90453 32864
rect 90411 32815 90453 32824
rect 90220 32696 90260 32705
rect 90220 32117 90260 32656
rect 90412 32192 90452 32815
rect 90305 32152 90452 32192
rect 89905 32068 89972 32108
rect 90015 32068 90164 32108
rect 90219 32108 90261 32117
rect 90219 32068 90220 32108
rect 90260 32068 90261 32108
rect 89905 31920 89945 32068
rect 90015 31920 90055 32068
rect 90219 32059 90261 32068
rect 90305 31920 90345 32152
rect 90508 32108 90548 33412
rect 90700 33403 90740 33412
rect 90988 33412 91084 33452
rect 90699 33200 90741 33209
rect 90699 33160 90700 33200
rect 90740 33160 90741 33200
rect 90699 33151 90741 33160
rect 90700 32959 90740 33151
rect 90891 33116 90933 33125
rect 90891 33076 90892 33116
rect 90932 33076 90933 33116
rect 90891 33067 90933 33076
rect 90892 32982 90932 33067
rect 90700 32910 90740 32919
rect 90795 32696 90837 32705
rect 90795 32656 90796 32696
rect 90836 32656 90837 32696
rect 90795 32647 90837 32656
rect 90796 32444 90836 32647
rect 90415 32068 90548 32108
rect 90705 32404 90836 32444
rect 90415 31920 90455 32068
rect 90705 31920 90745 32404
rect 90988 32360 91028 33412
rect 91084 33403 91124 33412
rect 91180 33041 91220 33571
rect 91468 33452 91508 33461
rect 91276 33412 91468 33452
rect 91179 33032 91221 33041
rect 91179 32992 91180 33032
rect 91220 32992 91221 33032
rect 91179 32983 91221 32992
rect 91083 32948 91125 32957
rect 91083 32908 91084 32948
rect 91124 32908 91125 32948
rect 91083 32899 91125 32908
rect 91084 32814 91124 32899
rect 91180 32864 91220 32983
rect 91180 32815 91220 32824
rect 91276 32360 91316 33412
rect 91468 33403 91508 33412
rect 91467 33032 91509 33041
rect 91467 32992 91468 33032
rect 91508 32992 91509 33032
rect 91467 32983 91509 32992
rect 91371 32864 91413 32873
rect 91371 32824 91372 32864
rect 91412 32824 91413 32864
rect 91371 32815 91413 32824
rect 91468 32864 91508 32983
rect 91468 32815 91508 32824
rect 91372 32730 91412 32815
rect 91467 32612 91509 32621
rect 91467 32572 91468 32612
rect 91508 32572 91509 32612
rect 91467 32563 91509 32572
rect 90815 32320 91028 32360
rect 91215 32320 91316 32360
rect 90815 31920 90855 32320
rect 91104 32276 91146 32285
rect 91104 32236 91105 32276
rect 91145 32236 91146 32276
rect 91104 32227 91146 32236
rect 91105 31920 91145 32227
rect 91215 31920 91255 32320
rect 91468 32108 91508 32563
rect 91564 32360 91604 34168
rect 91660 34159 91700 34168
rect 91659 33788 91701 33797
rect 91659 33748 91660 33788
rect 91700 33748 91701 33788
rect 91659 33739 91701 33748
rect 91660 33620 91700 33739
rect 93196 33629 93236 33714
rect 93388 33629 93428 34420
rect 93580 34208 93620 34217
rect 93484 34168 93580 34208
rect 91851 33620 91893 33629
rect 91700 33580 91796 33620
rect 91660 33571 91700 33580
rect 91756 33125 91796 33580
rect 91851 33580 91852 33620
rect 91892 33580 91893 33620
rect 91851 33571 91893 33580
rect 92236 33620 92276 33629
rect 92620 33620 92660 33629
rect 92276 33580 92372 33620
rect 92236 33571 92276 33580
rect 91852 33486 91892 33571
rect 92044 33452 92084 33461
rect 92084 33412 92180 33452
rect 92044 33403 92084 33412
rect 91755 33116 91797 33125
rect 91755 33076 91756 33116
rect 91796 33076 92084 33116
rect 91755 33067 91797 33076
rect 91756 32877 91796 33067
rect 91851 32948 91893 32957
rect 91851 32908 91852 32948
rect 91892 32908 91893 32948
rect 91851 32899 91893 32908
rect 91756 32828 91796 32837
rect 91852 32780 91892 32899
rect 92044 32864 92084 33076
rect 92044 32815 92084 32824
rect 91756 32740 91892 32780
rect 91659 32696 91701 32705
rect 91659 32656 91660 32696
rect 91700 32656 91701 32696
rect 91659 32647 91701 32656
rect 91660 32562 91700 32647
rect 91564 32320 91655 32360
rect 91468 32068 91545 32108
rect 91505 31920 91545 32068
rect 91615 31920 91655 32320
rect 91756 32108 91796 32740
rect 91948 32696 91988 32705
rect 91852 32656 91948 32696
rect 91852 32285 91892 32656
rect 91948 32647 91988 32656
rect 92140 32360 92180 33412
rect 92332 33209 92372 33580
rect 92523 33536 92565 33545
rect 92523 33496 92524 33536
rect 92564 33496 92565 33536
rect 92523 33487 92565 33496
rect 92428 33452 92468 33461
rect 92331 33200 92373 33209
rect 92331 33160 92332 33200
rect 92372 33160 92373 33200
rect 92331 33151 92373 33160
rect 92332 33116 92372 33151
rect 92332 33065 92372 33076
rect 92331 32864 92373 32873
rect 92331 32824 92332 32864
rect 92372 32824 92373 32864
rect 92331 32815 92373 32824
rect 92015 32320 92180 32360
rect 91851 32276 91893 32285
rect 91851 32236 91852 32276
rect 91892 32236 91893 32276
rect 91851 32227 91893 32236
rect 91756 32068 91945 32108
rect 91905 31920 91945 32068
rect 92015 31920 92055 32320
rect 92332 32192 92372 32815
rect 92428 32360 92468 33412
rect 92524 32948 92564 33487
rect 92620 33461 92660 33580
rect 93195 33620 93237 33629
rect 93195 33580 93196 33620
rect 93236 33580 93237 33620
rect 93195 33571 93237 33580
rect 93387 33620 93429 33629
rect 93387 33580 93388 33620
rect 93428 33580 93429 33620
rect 93387 33571 93429 33580
rect 92811 33536 92853 33545
rect 92811 33496 92812 33536
rect 92852 33496 92853 33536
rect 92811 33487 92853 33496
rect 92619 33452 92661 33461
rect 92619 33412 92620 33452
rect 92660 33412 92661 33452
rect 92619 33403 92661 33412
rect 92812 33402 92852 33487
rect 93004 33452 93044 33461
rect 93388 33452 93428 33461
rect 92908 33412 93004 33452
rect 92811 33116 92853 33125
rect 92811 33076 92812 33116
rect 92852 33076 92853 33116
rect 92811 33067 92853 33076
rect 92715 33032 92757 33041
rect 92715 32992 92716 33032
rect 92756 32992 92757 33032
rect 92715 32983 92757 32992
rect 92524 32899 92564 32908
rect 92716 32898 92756 32983
rect 92812 32864 92852 33067
rect 92812 32815 92852 32824
rect 92619 32780 92661 32789
rect 92619 32740 92620 32780
rect 92660 32740 92661 32780
rect 92619 32731 92661 32740
rect 92305 32152 92372 32192
rect 92415 32320 92468 32360
rect 92305 31920 92345 32152
rect 92415 31920 92455 32320
rect 92620 32108 92660 32731
rect 92908 32360 92948 33412
rect 93004 33403 93044 33412
rect 93196 33412 93388 33452
rect 93003 33116 93045 33125
rect 93003 33076 93004 33116
rect 93044 33076 93045 33116
rect 93003 33067 93045 33076
rect 93004 32864 93044 33067
rect 93099 32948 93141 32957
rect 93099 32908 93100 32948
rect 93140 32908 93141 32948
rect 93099 32899 93141 32908
rect 93004 32815 93044 32824
rect 93100 32814 93140 32899
rect 93003 32696 93045 32705
rect 93003 32656 93004 32696
rect 93044 32656 93045 32696
rect 93003 32647 93045 32656
rect 92815 32320 92948 32360
rect 92620 32068 92745 32108
rect 92705 31920 92745 32068
rect 92815 31920 92855 32320
rect 93004 32108 93044 32647
rect 93196 32360 93236 33412
rect 93388 33403 93428 33412
rect 93387 33200 93429 33209
rect 93387 33160 93388 33200
rect 93428 33160 93429 33200
rect 93387 33151 93429 33160
rect 93291 32864 93333 32873
rect 93291 32824 93292 32864
rect 93332 32824 93333 32864
rect 93291 32815 93333 32824
rect 93388 32864 93428 33151
rect 93388 32815 93428 32824
rect 93292 32730 93332 32815
rect 93484 32360 93524 34168
rect 93580 34159 93620 34168
rect 95500 33872 95540 33883
rect 95500 33797 95540 33832
rect 95499 33788 95541 33797
rect 95499 33748 95500 33788
rect 95540 33748 95541 33788
rect 95499 33739 95541 33748
rect 95307 33704 95349 33713
rect 95307 33664 95308 33704
rect 95348 33664 95349 33704
rect 95307 33655 95349 33664
rect 93579 33620 93621 33629
rect 93579 33580 93580 33620
rect 93620 33580 93621 33620
rect 93579 33571 93621 33580
rect 94060 33620 94100 33629
rect 94251 33620 94293 33629
rect 94100 33580 94252 33620
rect 94292 33580 94293 33620
rect 93580 33200 93620 33571
rect 93771 33536 93813 33545
rect 93771 33496 93772 33536
rect 93812 33496 93813 33536
rect 93771 33487 93813 33496
rect 93675 33200 93717 33209
rect 93580 33160 93676 33200
rect 93716 33160 93717 33200
rect 93772 33200 93812 33487
rect 93868 33452 93908 33461
rect 93908 33412 94004 33452
rect 93868 33403 93908 33412
rect 93772 33160 93908 33200
rect 93675 33151 93717 33160
rect 93676 32864 93716 33151
rect 93771 33032 93813 33041
rect 93771 32992 93772 33032
rect 93812 32992 93813 33032
rect 93771 32983 93813 32992
rect 93676 32815 93716 32824
rect 93579 32780 93621 32789
rect 93579 32740 93580 32780
rect 93620 32740 93621 32780
rect 93579 32731 93621 32740
rect 93580 32646 93620 32731
rect 93196 32320 93255 32360
rect 93484 32320 93655 32360
rect 93004 32068 93145 32108
rect 93105 31920 93145 32068
rect 93215 31920 93255 32320
rect 93504 32108 93546 32117
rect 93504 32068 93505 32108
rect 93545 32068 93546 32108
rect 93504 32059 93546 32068
rect 93505 31920 93545 32059
rect 93615 31920 93655 32320
rect 93772 32117 93812 32983
rect 93868 32948 93908 33160
rect 93868 32899 93908 32908
rect 93867 32780 93909 32789
rect 93867 32740 93868 32780
rect 93908 32740 93909 32780
rect 93867 32731 93909 32740
rect 93771 32108 93813 32117
rect 93771 32068 93772 32108
rect 93812 32068 93813 32108
rect 93868 32108 93908 32731
rect 93964 32360 94004 33412
rect 94060 33116 94100 33580
rect 94251 33571 94293 33580
rect 94635 33620 94677 33629
rect 94635 33580 94636 33620
rect 94676 33580 94677 33620
rect 94635 33571 94677 33580
rect 95308 33620 95348 33655
rect 95692 33629 95732 33714
rect 96075 33704 96117 33713
rect 96075 33664 96076 33704
rect 96116 33664 96117 33704
rect 96075 33655 96117 33664
rect 96459 33704 96501 33713
rect 96459 33664 96460 33704
rect 96500 33664 96501 33704
rect 96459 33655 96501 33664
rect 94252 33486 94292 33571
rect 94444 33452 94484 33461
rect 94347 33200 94389 33209
rect 94347 33160 94348 33200
rect 94388 33160 94389 33200
rect 94347 33151 94389 33160
rect 94060 33067 94100 33076
rect 94155 32948 94197 32957
rect 94155 32908 94156 32948
rect 94196 32908 94197 32948
rect 94155 32899 94197 32908
rect 93964 32320 94055 32360
rect 93868 32068 93945 32108
rect 93771 32059 93813 32068
rect 93905 31920 93945 32068
rect 94015 31920 94055 32320
rect 94156 32108 94196 32899
rect 94251 32864 94293 32873
rect 94251 32824 94252 32864
rect 94292 32824 94293 32864
rect 94251 32815 94293 32824
rect 94348 32864 94388 33151
rect 94348 32815 94388 32824
rect 94252 32730 94292 32815
rect 94444 32360 94484 33412
rect 94636 33125 94676 33571
rect 95308 33569 95348 33580
rect 95691 33620 95733 33629
rect 95691 33580 95692 33620
rect 95732 33580 95733 33620
rect 95691 33571 95733 33580
rect 96076 33620 96116 33655
rect 94828 33452 94868 33461
rect 94732 33412 94828 33452
rect 94635 33116 94677 33125
rect 94635 33076 94636 33116
rect 94676 33076 94677 33116
rect 94635 33067 94677 33076
rect 94636 32864 94676 33067
rect 94636 32815 94676 32824
rect 94539 32780 94581 32789
rect 94539 32740 94540 32780
rect 94580 32740 94581 32780
rect 94539 32731 94581 32740
rect 94540 32646 94580 32731
rect 94415 32320 94484 32360
rect 94732 32360 94772 33412
rect 94828 33403 94868 33412
rect 95116 33452 95156 33461
rect 95884 33452 95924 33461
rect 95156 33412 95348 33452
rect 95116 33403 95156 33412
rect 94827 33200 94869 33209
rect 94827 33160 94828 33200
rect 94868 33160 94869 33200
rect 94827 33151 94869 33160
rect 94828 32864 94868 33151
rect 95211 33116 95253 33125
rect 95211 33076 95212 33116
rect 95252 33076 95253 33116
rect 95211 33067 95253 33076
rect 94923 33032 94965 33041
rect 94923 32992 94924 33032
rect 94964 32992 94965 33032
rect 94923 32983 94965 32992
rect 94924 32898 94964 32983
rect 95115 32948 95157 32957
rect 95115 32908 95116 32948
rect 95156 32908 95157 32948
rect 95115 32899 95157 32908
rect 94828 32815 94868 32824
rect 95019 32864 95061 32873
rect 95019 32824 95020 32864
rect 95060 32824 95061 32864
rect 95019 32815 95061 32824
rect 94732 32320 94855 32360
rect 94156 32068 94345 32108
rect 94305 31920 94345 32068
rect 94415 31920 94455 32320
rect 94704 32108 94746 32117
rect 94704 32068 94705 32108
rect 94745 32068 94746 32108
rect 94704 32059 94746 32068
rect 94705 31920 94745 32059
rect 94815 31920 94855 32320
rect 95020 32108 95060 32815
rect 95116 32814 95156 32899
rect 95212 32864 95252 33067
rect 95212 32815 95252 32824
rect 95308 32360 95348 33412
rect 95596 33412 95884 33452
rect 95499 33116 95541 33125
rect 95499 33076 95500 33116
rect 95540 33076 95541 33116
rect 95499 33067 95541 33076
rect 95500 32864 95540 33067
rect 95500 32815 95540 32824
rect 95215 32320 95348 32360
rect 95404 32696 95444 32705
rect 95020 32068 95145 32108
rect 95105 31920 95145 32068
rect 95215 31920 95255 32320
rect 95404 32117 95444 32656
rect 95499 32696 95541 32705
rect 95499 32656 95500 32696
rect 95540 32656 95541 32696
rect 95499 32647 95541 32656
rect 95403 32108 95445 32117
rect 95403 32068 95404 32108
rect 95444 32068 95445 32108
rect 95500 32108 95540 32647
rect 95596 32360 95636 33412
rect 95884 33403 95924 33412
rect 95691 33116 95733 33125
rect 95691 33076 95692 33116
rect 95732 33076 95733 33116
rect 95691 33067 95733 33076
rect 95692 32864 95732 33067
rect 96076 32873 96116 33580
rect 96460 33620 96500 33655
rect 96460 33569 96500 33580
rect 96747 33620 96789 33629
rect 96747 33580 96748 33620
rect 96788 33580 96789 33620
rect 96747 33571 96789 33580
rect 96844 33620 96884 33629
rect 96939 33620 96981 33629
rect 97228 33620 97268 33629
rect 97612 33620 97652 33629
rect 96884 33580 96940 33620
rect 96980 33580 96981 33620
rect 96844 33571 96884 33580
rect 96939 33571 96981 33580
rect 97132 33580 97228 33620
rect 96268 33452 96308 33461
rect 96652 33452 96692 33461
rect 96172 33412 96268 33452
rect 95692 32815 95732 32824
rect 95787 32864 95829 32873
rect 95787 32824 95788 32864
rect 95828 32824 95829 32864
rect 95787 32815 95829 32824
rect 96075 32864 96117 32873
rect 96075 32824 96076 32864
rect 96116 32824 96117 32864
rect 96075 32815 96117 32824
rect 95788 32730 95828 32815
rect 95979 32780 96021 32789
rect 95979 32740 95980 32780
rect 96020 32740 96021 32780
rect 95979 32731 96021 32740
rect 95980 32646 96020 32731
rect 96076 32730 96116 32815
rect 95596 32320 95655 32360
rect 95500 32068 95545 32108
rect 95403 32059 95445 32068
rect 95505 31920 95545 32068
rect 95615 31920 95655 32320
rect 95904 32276 95946 32285
rect 95904 32236 95905 32276
rect 95945 32236 95946 32276
rect 95904 32227 95946 32236
rect 95905 31920 95945 32227
rect 96172 32192 96212 33412
rect 96268 33403 96308 33412
rect 96460 33412 96652 33452
rect 96363 32864 96405 32873
rect 96363 32824 96364 32864
rect 96404 32824 96405 32864
rect 96363 32815 96405 32824
rect 96364 32730 96404 32815
rect 96268 32696 96308 32705
rect 96268 32285 96308 32656
rect 96460 32360 96500 33412
rect 96652 33403 96692 33412
rect 96748 32948 96788 33571
rect 97036 33452 97076 33461
rect 96748 32899 96788 32908
rect 96940 33032 96980 33041
rect 96940 32873 96980 32992
rect 96939 32864 96981 32873
rect 96939 32824 96940 32864
rect 96980 32824 96981 32864
rect 96939 32815 96981 32824
rect 97036 32444 97076 33412
rect 97132 32873 97172 33580
rect 97228 33571 97268 33580
rect 97516 33580 97612 33620
rect 97227 33452 97269 33461
rect 97420 33452 97460 33461
rect 97227 33412 97228 33452
rect 97268 33412 97269 33452
rect 97227 33403 97269 33412
rect 97324 33412 97420 33452
rect 97131 32864 97173 32873
rect 97131 32824 97132 32864
rect 97172 32824 97173 32864
rect 97131 32815 97173 32824
rect 97228 32864 97268 33403
rect 97228 32815 97268 32824
rect 96844 32404 97076 32444
rect 97132 32696 97172 32705
rect 96844 32360 96884 32404
rect 96415 32320 96500 32360
rect 96815 32320 96884 32360
rect 96267 32276 96309 32285
rect 96267 32236 96268 32276
rect 96308 32236 96309 32276
rect 96267 32227 96309 32236
rect 96015 32152 96212 32192
rect 96015 31920 96055 32152
rect 96304 32108 96346 32117
rect 96304 32068 96305 32108
rect 96345 32068 96346 32108
rect 96304 32059 96346 32068
rect 96305 31920 96345 32059
rect 96415 31920 96455 32320
rect 96704 32192 96746 32201
rect 96704 32152 96705 32192
rect 96745 32152 96746 32192
rect 96704 32143 96746 32152
rect 96705 31920 96745 32143
rect 96815 31920 96855 32320
rect 97132 32285 97172 32656
rect 97324 32360 97364 33412
rect 97420 33403 97460 33412
rect 97516 32873 97556 33580
rect 97612 33571 97652 33580
rect 97996 33620 98036 33629
rect 97804 33452 97844 33461
rect 97612 33412 97804 33452
rect 97515 32864 97557 32873
rect 97515 32824 97516 32864
rect 97556 32824 97557 32864
rect 97515 32815 97557 32824
rect 97215 32320 97364 32360
rect 97420 32696 97460 32705
rect 97131 32276 97173 32285
rect 97131 32236 97132 32276
rect 97172 32236 97173 32276
rect 97131 32227 97173 32236
rect 97104 32108 97146 32117
rect 97104 32068 97105 32108
rect 97145 32068 97146 32108
rect 97104 32059 97146 32068
rect 97105 31920 97145 32059
rect 97215 31920 97255 32320
rect 97420 32201 97460 32656
rect 97515 32696 97557 32705
rect 97515 32656 97516 32696
rect 97556 32656 97557 32696
rect 97515 32647 97557 32656
rect 97419 32192 97461 32201
rect 97419 32152 97420 32192
rect 97460 32152 97461 32192
rect 97419 32143 97461 32152
rect 97516 32108 97556 32647
rect 97612 32360 97652 33412
rect 97804 33403 97844 33412
rect 97803 32864 97845 32873
rect 97803 32824 97804 32864
rect 97844 32824 97845 32864
rect 97996 32864 98036 33580
rect 98379 33620 98421 33629
rect 98379 33580 98380 33620
rect 98420 33580 98421 33620
rect 98379 33571 98421 33580
rect 98380 33486 98420 33571
rect 98188 33452 98228 33461
rect 98091 32864 98133 32873
rect 97996 32824 98092 32864
rect 98132 32824 98133 32864
rect 97803 32815 97845 32824
rect 98091 32815 98133 32824
rect 97804 32730 97844 32815
rect 98092 32730 98132 32815
rect 97708 32696 97748 32705
rect 97612 32320 97655 32360
rect 97505 32068 97556 32108
rect 97505 31920 97545 32068
rect 97615 31920 97655 32320
rect 97708 32117 97748 32656
rect 97995 32696 98037 32705
rect 97995 32656 97996 32696
rect 98036 32656 98037 32696
rect 97995 32647 98037 32656
rect 97996 32562 98036 32647
rect 98188 32360 98228 33412
rect 98668 32948 98708 32957
rect 98668 32864 98708 32908
rect 98860 32864 98900 32873
rect 98668 32824 98860 32864
rect 98015 32320 98228 32360
rect 98476 32696 98516 32705
rect 97707 32108 97749 32117
rect 97707 32068 97708 32108
rect 97748 32068 97749 32108
rect 97707 32059 97749 32068
rect 97904 32108 97946 32117
rect 97904 32068 97905 32108
rect 97945 32068 97946 32108
rect 97904 32059 97946 32068
rect 97905 31920 97945 32059
rect 98015 31920 98055 32320
rect 98304 32192 98346 32201
rect 98476 32192 98516 32656
rect 98304 32152 98305 32192
rect 98345 32152 98346 32192
rect 98304 32143 98346 32152
rect 98390 32152 98516 32192
rect 98305 31920 98345 32143
rect 98390 32108 98430 32152
rect 98390 32068 98455 32108
rect 98415 31920 98455 32068
rect 71883 26732 71925 26741
rect 71883 26692 71884 26732
rect 71924 26692 71925 26732
rect 71883 26683 71925 26692
rect 71884 26069 71924 26683
rect 72305 26657 72345 26796
rect 72304 26648 72346 26657
rect 72304 26608 72305 26648
rect 72345 26608 72346 26648
rect 72304 26599 72346 26608
rect 72415 26489 72455 26796
rect 72705 26573 72745 26796
rect 72704 26564 72746 26573
rect 72704 26524 72705 26564
rect 72745 26524 72746 26564
rect 72815 26564 72855 26796
rect 72815 26524 72884 26564
rect 72704 26515 72746 26524
rect 72414 26480 72456 26489
rect 72414 26440 72415 26480
rect 72455 26440 72456 26480
rect 72414 26431 72456 26440
rect 72844 26321 72884 26524
rect 73105 26489 73145 26796
rect 73104 26480 73146 26489
rect 73104 26440 73105 26480
rect 73145 26440 73146 26480
rect 73104 26431 73146 26440
rect 73215 26396 73255 26796
rect 73505 26480 73545 26796
rect 73615 26648 73655 26796
rect 73420 26440 73545 26480
rect 73612 26608 73655 26648
rect 73215 26356 73268 26396
rect 72843 26312 72885 26321
rect 72843 26272 72844 26312
rect 72884 26272 72885 26312
rect 72843 26263 72885 26272
rect 71883 26060 71925 26069
rect 71883 26020 71884 26060
rect 71924 26020 71925 26060
rect 71883 26011 71925 26020
rect 73131 25724 73173 25733
rect 73131 25684 73132 25724
rect 73172 25684 73173 25724
rect 73131 25675 73173 25684
rect 72747 25556 72789 25565
rect 72747 25516 72748 25556
rect 72788 25516 72789 25556
rect 72747 25507 72789 25516
rect 73132 25556 73172 25675
rect 73228 25565 73268 26356
rect 73420 26237 73460 26440
rect 73419 26228 73461 26237
rect 73419 26188 73420 26228
rect 73460 26188 73461 26228
rect 73419 26179 73461 26188
rect 73612 26153 73652 26608
rect 73905 26396 73945 26796
rect 74015 26480 74055 26796
rect 73708 26356 73945 26396
rect 73996 26440 74055 26480
rect 73611 26144 73653 26153
rect 73611 26104 73612 26144
rect 73652 26104 73653 26144
rect 73611 26095 73653 26104
rect 73132 25507 73172 25516
rect 73227 25556 73269 25565
rect 73227 25516 73228 25556
rect 73268 25516 73269 25556
rect 73227 25507 73269 25516
rect 73516 25556 73556 25565
rect 73708 25556 73748 26356
rect 73803 25724 73845 25733
rect 73803 25684 73804 25724
rect 73844 25684 73845 25724
rect 73803 25675 73845 25684
rect 73556 25516 73748 25556
rect 73516 25507 73556 25516
rect 72748 25422 72788 25507
rect 72939 25388 72981 25397
rect 72939 25348 72940 25388
rect 72980 25348 72981 25388
rect 72939 25339 72981 25348
rect 73324 25388 73364 25399
rect 72651 25304 72693 25313
rect 72651 25264 72652 25304
rect 72692 25264 72693 25304
rect 72651 25255 72693 25264
rect 72652 25170 72692 25255
rect 72940 25254 72980 25339
rect 73324 25313 73364 25348
rect 73323 25304 73365 25313
rect 73323 25264 73324 25304
rect 73364 25264 73365 25304
rect 73323 25255 73365 25264
rect 73323 24968 73365 24977
rect 73323 24928 73324 24968
rect 73364 24928 73365 24968
rect 73323 24919 73365 24928
rect 73324 24800 73364 24919
rect 73324 24751 73364 24760
rect 73515 24800 73557 24809
rect 73515 24760 73516 24800
rect 73556 24760 73557 24800
rect 73515 24751 73557 24760
rect 71787 24716 71829 24725
rect 71787 24676 71788 24716
rect 71828 24676 71829 24716
rect 71787 24667 71829 24676
rect 73516 24666 73556 24751
rect 71019 24632 71061 24641
rect 71019 24592 71020 24632
rect 71060 24592 71061 24632
rect 71019 24583 71061 24592
rect 73227 24632 73269 24641
rect 73227 24592 73228 24632
rect 73268 24592 73269 24632
rect 73227 24583 73269 24592
rect 73612 24632 73652 24643
rect 651 23288 693 23297
rect 651 23248 652 23288
rect 692 23248 693 23288
rect 651 23239 693 23248
rect 2091 23288 2133 23297
rect 2091 23248 2092 23288
rect 2132 23248 2133 23288
rect 2091 23239 2133 23248
rect 69291 23288 69333 23297
rect 69291 23248 69292 23288
rect 69332 23248 69333 23288
rect 69291 23239 69333 23248
rect 652 23120 692 23129
rect 556 23080 652 23120
rect 556 22457 596 23080
rect 652 23071 692 23080
rect 843 23120 885 23129
rect 843 23080 844 23120
rect 884 23080 885 23120
rect 843 23071 885 23080
rect 1995 23120 2037 23129
rect 1995 23080 1996 23120
rect 2036 23080 2037 23120
rect 1995 23071 2037 23080
rect 844 22986 884 23071
rect 555 22448 597 22457
rect 555 22408 556 22448
rect 596 22408 597 22448
rect 555 22399 597 22408
rect 652 22448 692 22457
rect 652 21617 692 22408
rect 651 21608 693 21617
rect 651 21568 652 21608
rect 692 21568 693 21608
rect 651 21559 693 21568
rect 652 20936 692 20945
rect 652 20777 692 20896
rect 651 20768 693 20777
rect 651 20728 652 20768
rect 692 20728 693 20768
rect 651 20719 693 20728
rect 651 19928 693 19937
rect 651 19888 652 19928
rect 692 19888 693 19928
rect 651 19879 693 19888
rect 652 19794 692 19879
rect 652 19424 692 19433
rect 652 19097 692 19384
rect 651 19088 693 19097
rect 651 19048 652 19088
rect 692 19048 693 19088
rect 651 19039 693 19048
rect 652 18416 692 18425
rect 652 18257 692 18376
rect 651 18248 693 18257
rect 651 18208 652 18248
rect 692 18208 693 18248
rect 651 18199 693 18208
rect 652 17912 692 17921
rect 652 17417 692 17872
rect 651 17408 693 17417
rect 651 17368 652 17408
rect 692 17368 693 17408
rect 651 17359 693 17368
rect 652 16904 692 16913
rect 652 16577 692 16864
rect 651 16568 693 16577
rect 651 16528 652 16568
rect 692 16528 693 16568
rect 651 16519 693 16528
rect 652 16400 692 16409
rect 652 15737 692 16360
rect 651 15728 693 15737
rect 651 15688 652 15728
rect 692 15688 693 15728
rect 651 15679 693 15688
rect 844 15476 884 15485
rect 652 15308 692 15317
rect 652 14897 692 15268
rect 844 14981 884 15436
rect 843 14972 885 14981
rect 843 14932 844 14972
rect 884 14932 885 14972
rect 843 14923 885 14932
rect 1419 14972 1461 14981
rect 1419 14932 1420 14972
rect 1460 14932 1461 14972
rect 1419 14923 1461 14932
rect 651 14888 693 14897
rect 651 14848 652 14888
rect 692 14848 693 14888
rect 651 14839 693 14848
rect 1420 14838 1460 14923
rect 1996 14813 2036 23071
rect 844 14804 884 14813
rect 1612 14804 1652 14813
rect 884 14764 1076 14804
rect 844 14755 884 14764
rect 652 14552 692 14561
rect 652 14057 692 14512
rect 1036 14216 1076 14764
rect 1612 14552 1652 14764
rect 1995 14804 2037 14813
rect 1995 14764 1996 14804
rect 2036 14764 2037 14804
rect 1995 14755 2037 14764
rect 1996 14669 2036 14755
rect 1804 14552 1844 14561
rect 1612 14512 1804 14552
rect 1036 14167 1076 14176
rect 651 14048 693 14057
rect 651 14008 652 14048
rect 692 14008 693 14048
rect 651 13999 693 14008
rect 1804 13973 1844 14512
rect 1227 13964 1269 13973
rect 1227 13924 1228 13964
rect 1268 13924 1269 13964
rect 1227 13915 1269 13924
rect 1803 13964 1845 13973
rect 1803 13924 1804 13964
rect 1844 13924 1845 13964
rect 1803 13915 1845 13924
rect 1228 13830 1268 13915
rect 843 13376 885 13385
rect 843 13336 844 13376
rect 884 13336 885 13376
rect 843 13327 885 13336
rect 1611 13376 1653 13385
rect 1611 13336 1612 13376
rect 1652 13336 1653 13376
rect 1611 13327 1653 13336
rect 844 13292 884 13327
rect 844 13241 884 13252
rect 1612 13242 1652 13327
rect 1804 13292 1844 13915
rect 651 13208 693 13217
rect 651 13168 652 13208
rect 692 13168 693 13208
rect 651 13159 693 13168
rect 652 13040 692 13159
rect 652 12991 692 13000
rect 844 12452 884 12461
rect 651 12368 693 12377
rect 651 12328 652 12368
rect 692 12328 693 12368
rect 844 12368 884 12412
rect 1420 12452 1460 12461
rect 1804 12452 1844 13252
rect 1460 12412 1844 12452
rect 1228 12368 1268 12377
rect 844 12328 1228 12368
rect 651 12319 693 12328
rect 1228 12319 1268 12328
rect 652 12234 692 12319
rect 844 11780 884 11789
rect 884 11740 1268 11780
rect 844 11731 884 11740
rect 651 11528 693 11537
rect 651 11488 652 11528
rect 692 11488 693 11528
rect 651 11479 693 11488
rect 652 11394 692 11479
rect 1228 11192 1268 11740
rect 1228 11143 1268 11152
rect 844 10940 884 10949
rect 1420 10940 1460 12412
rect 651 10772 693 10781
rect 651 10732 652 10772
rect 692 10732 693 10772
rect 651 10723 693 10732
rect 652 10638 692 10723
rect 844 10529 884 10900
rect 1324 10900 1420 10940
rect 843 10520 885 10529
rect 843 10480 844 10520
rect 884 10480 885 10520
rect 843 10471 885 10480
rect 1036 10352 1076 10361
rect 844 10312 1036 10352
rect 844 10268 884 10312
rect 1036 10303 1076 10312
rect 844 10219 884 10228
rect 1227 10268 1269 10277
rect 1324 10268 1364 10900
rect 1420 10891 1460 10900
rect 1419 10520 1461 10529
rect 1419 10480 1420 10520
rect 1460 10480 1461 10520
rect 1419 10471 1461 10480
rect 1420 10436 1460 10471
rect 1420 10385 1460 10396
rect 1227 10228 1228 10268
rect 1268 10228 1364 10268
rect 1611 10268 1653 10277
rect 1611 10228 1612 10268
rect 1652 10228 1748 10268
rect 1227 10219 1269 10228
rect 1611 10219 1653 10228
rect 1228 10134 1268 10219
rect 1612 10134 1652 10219
rect 652 10016 692 10025
rect 652 9857 692 9976
rect 651 9848 693 9857
rect 651 9808 652 9848
rect 692 9808 693 9848
rect 651 9799 693 9808
rect 844 9428 884 9437
rect 748 9388 844 9428
rect 652 9260 692 9269
rect 652 9017 692 9220
rect 651 9008 693 9017
rect 651 8968 652 9008
rect 692 8968 693 9008
rect 651 8959 693 8968
rect 748 8849 788 9388
rect 844 9379 884 9388
rect 747 8840 789 8849
rect 1132 8840 1172 8849
rect 747 8800 748 8840
rect 788 8800 789 8840
rect 747 8791 789 8800
rect 844 8800 1132 8840
rect 844 8756 884 8800
rect 1132 8791 1172 8800
rect 1515 8840 1557 8849
rect 1515 8800 1516 8840
rect 1556 8800 1557 8840
rect 1515 8791 1557 8800
rect 844 8707 884 8716
rect 1324 8756 1364 8765
rect 652 8504 692 8513
rect 1324 8504 1364 8716
rect 1516 8706 1556 8791
rect 1708 8756 1748 10228
rect 1708 8707 1748 8716
rect 2092 8756 2132 23239
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 7112 22700 7480 22709
rect 7152 22660 7194 22700
rect 7234 22660 7276 22700
rect 7316 22660 7358 22700
rect 7398 22660 7440 22700
rect 7112 22651 7480 22660
rect 11112 22700 11480 22709
rect 11152 22660 11194 22700
rect 11234 22660 11276 22700
rect 11316 22660 11358 22700
rect 11398 22660 11440 22700
rect 11112 22651 11480 22660
rect 15112 22700 15480 22709
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15112 22651 15480 22660
rect 19112 22700 19480 22709
rect 19152 22660 19194 22700
rect 19234 22660 19276 22700
rect 19316 22660 19358 22700
rect 19398 22660 19440 22700
rect 19112 22651 19480 22660
rect 23112 22700 23480 22709
rect 23152 22660 23194 22700
rect 23234 22660 23276 22700
rect 23316 22660 23358 22700
rect 23398 22660 23440 22700
rect 23112 22651 23480 22660
rect 27112 22700 27480 22709
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27112 22651 27480 22660
rect 31112 22700 31480 22709
rect 31152 22660 31194 22700
rect 31234 22660 31276 22700
rect 31316 22660 31358 22700
rect 31398 22660 31440 22700
rect 31112 22651 31480 22660
rect 35112 22700 35480 22709
rect 35152 22660 35194 22700
rect 35234 22660 35276 22700
rect 35316 22660 35358 22700
rect 35398 22660 35440 22700
rect 35112 22651 35480 22660
rect 39112 22700 39480 22709
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39112 22651 39480 22660
rect 43112 22700 43480 22709
rect 43152 22660 43194 22700
rect 43234 22660 43276 22700
rect 43316 22660 43358 22700
rect 43398 22660 43440 22700
rect 43112 22651 43480 22660
rect 47112 22700 47480 22709
rect 47152 22660 47194 22700
rect 47234 22660 47276 22700
rect 47316 22660 47358 22700
rect 47398 22660 47440 22700
rect 47112 22651 47480 22660
rect 51112 22700 51480 22709
rect 51152 22660 51194 22700
rect 51234 22660 51276 22700
rect 51316 22660 51358 22700
rect 51398 22660 51440 22700
rect 51112 22651 51480 22660
rect 55112 22700 55480 22709
rect 55152 22660 55194 22700
rect 55234 22660 55276 22700
rect 55316 22660 55358 22700
rect 55398 22660 55440 22700
rect 55112 22651 55480 22660
rect 59112 22700 59480 22709
rect 59152 22660 59194 22700
rect 59234 22660 59276 22700
rect 59316 22660 59358 22700
rect 59398 22660 59440 22700
rect 59112 22651 59480 22660
rect 63112 22700 63480 22709
rect 63152 22660 63194 22700
rect 63234 22660 63276 22700
rect 63316 22660 63358 22700
rect 63398 22660 63440 22700
rect 63112 22651 63480 22660
rect 67112 22700 67480 22709
rect 67152 22660 67194 22700
rect 67234 22660 67276 22700
rect 67316 22660 67358 22700
rect 67398 22660 67440 22700
rect 67112 22651 67480 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 8352 21944 8720 21953
rect 8392 21904 8434 21944
rect 8474 21904 8516 21944
rect 8556 21904 8598 21944
rect 8638 21904 8680 21944
rect 8352 21895 8720 21904
rect 12352 21944 12720 21953
rect 12392 21904 12434 21944
rect 12474 21904 12516 21944
rect 12556 21904 12598 21944
rect 12638 21904 12680 21944
rect 12352 21895 12720 21904
rect 16352 21944 16720 21953
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16352 21895 16720 21904
rect 20352 21944 20720 21953
rect 20392 21904 20434 21944
rect 20474 21904 20516 21944
rect 20556 21904 20598 21944
rect 20638 21904 20680 21944
rect 20352 21895 20720 21904
rect 24352 21944 24720 21953
rect 24392 21904 24434 21944
rect 24474 21904 24516 21944
rect 24556 21904 24598 21944
rect 24638 21904 24680 21944
rect 24352 21895 24720 21904
rect 28352 21944 28720 21953
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28352 21895 28720 21904
rect 32352 21944 32720 21953
rect 32392 21904 32434 21944
rect 32474 21904 32516 21944
rect 32556 21904 32598 21944
rect 32638 21904 32680 21944
rect 32352 21895 32720 21904
rect 36352 21944 36720 21953
rect 36392 21904 36434 21944
rect 36474 21904 36516 21944
rect 36556 21904 36598 21944
rect 36638 21904 36680 21944
rect 36352 21895 36720 21904
rect 40352 21944 40720 21953
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40352 21895 40720 21904
rect 44352 21944 44720 21953
rect 44392 21904 44434 21944
rect 44474 21904 44516 21944
rect 44556 21904 44598 21944
rect 44638 21904 44680 21944
rect 44352 21895 44720 21904
rect 48352 21944 48720 21953
rect 48392 21904 48434 21944
rect 48474 21904 48516 21944
rect 48556 21904 48598 21944
rect 48638 21904 48680 21944
rect 48352 21895 48720 21904
rect 52352 21944 52720 21953
rect 52392 21904 52434 21944
rect 52474 21904 52516 21944
rect 52556 21904 52598 21944
rect 52638 21904 52680 21944
rect 52352 21895 52720 21904
rect 56352 21944 56720 21953
rect 56392 21904 56434 21944
rect 56474 21904 56516 21944
rect 56556 21904 56598 21944
rect 56638 21904 56680 21944
rect 56352 21895 56720 21904
rect 60352 21944 60720 21953
rect 60392 21904 60434 21944
rect 60474 21904 60516 21944
rect 60556 21904 60598 21944
rect 60638 21904 60680 21944
rect 60352 21895 60720 21904
rect 64352 21944 64720 21953
rect 64392 21904 64434 21944
rect 64474 21904 64516 21944
rect 64556 21904 64598 21944
rect 64638 21904 64680 21944
rect 64352 21895 64720 21904
rect 68352 21944 68720 21953
rect 68392 21904 68434 21944
rect 68474 21904 68516 21944
rect 68556 21904 68598 21944
rect 68638 21904 68680 21944
rect 68352 21895 68720 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 7112 21188 7480 21197
rect 7152 21148 7194 21188
rect 7234 21148 7276 21188
rect 7316 21148 7358 21188
rect 7398 21148 7440 21188
rect 7112 21139 7480 21148
rect 11112 21188 11480 21197
rect 11152 21148 11194 21188
rect 11234 21148 11276 21188
rect 11316 21148 11358 21188
rect 11398 21148 11440 21188
rect 11112 21139 11480 21148
rect 15112 21188 15480 21197
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15112 21139 15480 21148
rect 19112 21188 19480 21197
rect 19152 21148 19194 21188
rect 19234 21148 19276 21188
rect 19316 21148 19358 21188
rect 19398 21148 19440 21188
rect 19112 21139 19480 21148
rect 23112 21188 23480 21197
rect 23152 21148 23194 21188
rect 23234 21148 23276 21188
rect 23316 21148 23358 21188
rect 23398 21148 23440 21188
rect 23112 21139 23480 21148
rect 27112 21188 27480 21197
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27112 21139 27480 21148
rect 31112 21188 31480 21197
rect 31152 21148 31194 21188
rect 31234 21148 31276 21188
rect 31316 21148 31358 21188
rect 31398 21148 31440 21188
rect 31112 21139 31480 21148
rect 35112 21188 35480 21197
rect 35152 21148 35194 21188
rect 35234 21148 35276 21188
rect 35316 21148 35358 21188
rect 35398 21148 35440 21188
rect 35112 21139 35480 21148
rect 39112 21188 39480 21197
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39112 21139 39480 21148
rect 43112 21188 43480 21197
rect 43152 21148 43194 21188
rect 43234 21148 43276 21188
rect 43316 21148 43358 21188
rect 43398 21148 43440 21188
rect 43112 21139 43480 21148
rect 47112 21188 47480 21197
rect 47152 21148 47194 21188
rect 47234 21148 47276 21188
rect 47316 21148 47358 21188
rect 47398 21148 47440 21188
rect 47112 21139 47480 21148
rect 51112 21188 51480 21197
rect 51152 21148 51194 21188
rect 51234 21148 51276 21188
rect 51316 21148 51358 21188
rect 51398 21148 51440 21188
rect 51112 21139 51480 21148
rect 55112 21188 55480 21197
rect 55152 21148 55194 21188
rect 55234 21148 55276 21188
rect 55316 21148 55358 21188
rect 55398 21148 55440 21188
rect 55112 21139 55480 21148
rect 59112 21188 59480 21197
rect 59152 21148 59194 21188
rect 59234 21148 59276 21188
rect 59316 21148 59358 21188
rect 59398 21148 59440 21188
rect 59112 21139 59480 21148
rect 63112 21188 63480 21197
rect 63152 21148 63194 21188
rect 63234 21148 63276 21188
rect 63316 21148 63358 21188
rect 63398 21148 63440 21188
rect 63112 21139 63480 21148
rect 67112 21188 67480 21197
rect 67152 21148 67194 21188
rect 67234 21148 67276 21188
rect 67316 21148 67358 21188
rect 67398 21148 67440 21188
rect 67112 21139 67480 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 8352 20432 8720 20441
rect 8392 20392 8434 20432
rect 8474 20392 8516 20432
rect 8556 20392 8598 20432
rect 8638 20392 8680 20432
rect 8352 20383 8720 20392
rect 12352 20432 12720 20441
rect 12392 20392 12434 20432
rect 12474 20392 12516 20432
rect 12556 20392 12598 20432
rect 12638 20392 12680 20432
rect 12352 20383 12720 20392
rect 16352 20432 16720 20441
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16352 20383 16720 20392
rect 20352 20432 20720 20441
rect 20392 20392 20434 20432
rect 20474 20392 20516 20432
rect 20556 20392 20598 20432
rect 20638 20392 20680 20432
rect 20352 20383 20720 20392
rect 24352 20432 24720 20441
rect 24392 20392 24434 20432
rect 24474 20392 24516 20432
rect 24556 20392 24598 20432
rect 24638 20392 24680 20432
rect 24352 20383 24720 20392
rect 28352 20432 28720 20441
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28352 20383 28720 20392
rect 32352 20432 32720 20441
rect 32392 20392 32434 20432
rect 32474 20392 32516 20432
rect 32556 20392 32598 20432
rect 32638 20392 32680 20432
rect 32352 20383 32720 20392
rect 36352 20432 36720 20441
rect 36392 20392 36434 20432
rect 36474 20392 36516 20432
rect 36556 20392 36598 20432
rect 36638 20392 36680 20432
rect 36352 20383 36720 20392
rect 40352 20432 40720 20441
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40352 20383 40720 20392
rect 44352 20432 44720 20441
rect 44392 20392 44434 20432
rect 44474 20392 44516 20432
rect 44556 20392 44598 20432
rect 44638 20392 44680 20432
rect 44352 20383 44720 20392
rect 48352 20432 48720 20441
rect 48392 20392 48434 20432
rect 48474 20392 48516 20432
rect 48556 20392 48598 20432
rect 48638 20392 48680 20432
rect 48352 20383 48720 20392
rect 52352 20432 52720 20441
rect 52392 20392 52434 20432
rect 52474 20392 52516 20432
rect 52556 20392 52598 20432
rect 52638 20392 52680 20432
rect 52352 20383 52720 20392
rect 56352 20432 56720 20441
rect 56392 20392 56434 20432
rect 56474 20392 56516 20432
rect 56556 20392 56598 20432
rect 56638 20392 56680 20432
rect 56352 20383 56720 20392
rect 60352 20432 60720 20441
rect 60392 20392 60434 20432
rect 60474 20392 60516 20432
rect 60556 20392 60598 20432
rect 60638 20392 60680 20432
rect 60352 20383 60720 20392
rect 64352 20432 64720 20441
rect 64392 20392 64434 20432
rect 64474 20392 64516 20432
rect 64556 20392 64598 20432
rect 64638 20392 64680 20432
rect 64352 20383 64720 20392
rect 68352 20432 68720 20441
rect 68392 20392 68434 20432
rect 68474 20392 68516 20432
rect 68556 20392 68598 20432
rect 68638 20392 68680 20432
rect 68352 20383 68720 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 7112 19676 7480 19685
rect 7152 19636 7194 19676
rect 7234 19636 7276 19676
rect 7316 19636 7358 19676
rect 7398 19636 7440 19676
rect 7112 19627 7480 19636
rect 11112 19676 11480 19685
rect 11152 19636 11194 19676
rect 11234 19636 11276 19676
rect 11316 19636 11358 19676
rect 11398 19636 11440 19676
rect 11112 19627 11480 19636
rect 15112 19676 15480 19685
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15112 19627 15480 19636
rect 19112 19676 19480 19685
rect 19152 19636 19194 19676
rect 19234 19636 19276 19676
rect 19316 19636 19358 19676
rect 19398 19636 19440 19676
rect 19112 19627 19480 19636
rect 23112 19676 23480 19685
rect 23152 19636 23194 19676
rect 23234 19636 23276 19676
rect 23316 19636 23358 19676
rect 23398 19636 23440 19676
rect 23112 19627 23480 19636
rect 27112 19676 27480 19685
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27112 19627 27480 19636
rect 31112 19676 31480 19685
rect 31152 19636 31194 19676
rect 31234 19636 31276 19676
rect 31316 19636 31358 19676
rect 31398 19636 31440 19676
rect 31112 19627 31480 19636
rect 35112 19676 35480 19685
rect 35152 19636 35194 19676
rect 35234 19636 35276 19676
rect 35316 19636 35358 19676
rect 35398 19636 35440 19676
rect 35112 19627 35480 19636
rect 39112 19676 39480 19685
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39112 19627 39480 19636
rect 43112 19676 43480 19685
rect 43152 19636 43194 19676
rect 43234 19636 43276 19676
rect 43316 19636 43358 19676
rect 43398 19636 43440 19676
rect 43112 19627 43480 19636
rect 47112 19676 47480 19685
rect 47152 19636 47194 19676
rect 47234 19636 47276 19676
rect 47316 19636 47358 19676
rect 47398 19636 47440 19676
rect 47112 19627 47480 19636
rect 51112 19676 51480 19685
rect 51152 19636 51194 19676
rect 51234 19636 51276 19676
rect 51316 19636 51358 19676
rect 51398 19636 51440 19676
rect 51112 19627 51480 19636
rect 55112 19676 55480 19685
rect 55152 19636 55194 19676
rect 55234 19636 55276 19676
rect 55316 19636 55358 19676
rect 55398 19636 55440 19676
rect 55112 19627 55480 19636
rect 59112 19676 59480 19685
rect 59152 19636 59194 19676
rect 59234 19636 59276 19676
rect 59316 19636 59358 19676
rect 59398 19636 59440 19676
rect 59112 19627 59480 19636
rect 63112 19676 63480 19685
rect 63152 19636 63194 19676
rect 63234 19636 63276 19676
rect 63316 19636 63358 19676
rect 63398 19636 63440 19676
rect 63112 19627 63480 19636
rect 67112 19676 67480 19685
rect 67152 19636 67194 19676
rect 67234 19636 67276 19676
rect 67316 19636 67358 19676
rect 67398 19636 67440 19676
rect 67112 19627 67480 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 8352 18920 8720 18929
rect 8392 18880 8434 18920
rect 8474 18880 8516 18920
rect 8556 18880 8598 18920
rect 8638 18880 8680 18920
rect 8352 18871 8720 18880
rect 12352 18920 12720 18929
rect 12392 18880 12434 18920
rect 12474 18880 12516 18920
rect 12556 18880 12598 18920
rect 12638 18880 12680 18920
rect 12352 18871 12720 18880
rect 16352 18920 16720 18929
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16352 18871 16720 18880
rect 20352 18920 20720 18929
rect 20392 18880 20434 18920
rect 20474 18880 20516 18920
rect 20556 18880 20598 18920
rect 20638 18880 20680 18920
rect 20352 18871 20720 18880
rect 24352 18920 24720 18929
rect 24392 18880 24434 18920
rect 24474 18880 24516 18920
rect 24556 18880 24598 18920
rect 24638 18880 24680 18920
rect 24352 18871 24720 18880
rect 28352 18920 28720 18929
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28352 18871 28720 18880
rect 32352 18920 32720 18929
rect 32392 18880 32434 18920
rect 32474 18880 32516 18920
rect 32556 18880 32598 18920
rect 32638 18880 32680 18920
rect 32352 18871 32720 18880
rect 36352 18920 36720 18929
rect 36392 18880 36434 18920
rect 36474 18880 36516 18920
rect 36556 18880 36598 18920
rect 36638 18880 36680 18920
rect 36352 18871 36720 18880
rect 40352 18920 40720 18929
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40352 18871 40720 18880
rect 44352 18920 44720 18929
rect 44392 18880 44434 18920
rect 44474 18880 44516 18920
rect 44556 18880 44598 18920
rect 44638 18880 44680 18920
rect 44352 18871 44720 18880
rect 48352 18920 48720 18929
rect 48392 18880 48434 18920
rect 48474 18880 48516 18920
rect 48556 18880 48598 18920
rect 48638 18880 48680 18920
rect 48352 18871 48720 18880
rect 52352 18920 52720 18929
rect 52392 18880 52434 18920
rect 52474 18880 52516 18920
rect 52556 18880 52598 18920
rect 52638 18880 52680 18920
rect 52352 18871 52720 18880
rect 56352 18920 56720 18929
rect 56392 18880 56434 18920
rect 56474 18880 56516 18920
rect 56556 18880 56598 18920
rect 56638 18880 56680 18920
rect 56352 18871 56720 18880
rect 60352 18920 60720 18929
rect 60392 18880 60434 18920
rect 60474 18880 60516 18920
rect 60556 18880 60598 18920
rect 60638 18880 60680 18920
rect 60352 18871 60720 18880
rect 64352 18920 64720 18929
rect 64392 18880 64434 18920
rect 64474 18880 64516 18920
rect 64556 18880 64598 18920
rect 64638 18880 64680 18920
rect 64352 18871 64720 18880
rect 68352 18920 68720 18929
rect 68392 18880 68434 18920
rect 68474 18880 68516 18920
rect 68556 18880 68598 18920
rect 68638 18880 68680 18920
rect 68352 18871 68720 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 7112 18164 7480 18173
rect 7152 18124 7194 18164
rect 7234 18124 7276 18164
rect 7316 18124 7358 18164
rect 7398 18124 7440 18164
rect 7112 18115 7480 18124
rect 11112 18164 11480 18173
rect 11152 18124 11194 18164
rect 11234 18124 11276 18164
rect 11316 18124 11358 18164
rect 11398 18124 11440 18164
rect 11112 18115 11480 18124
rect 15112 18164 15480 18173
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15112 18115 15480 18124
rect 19112 18164 19480 18173
rect 19152 18124 19194 18164
rect 19234 18124 19276 18164
rect 19316 18124 19358 18164
rect 19398 18124 19440 18164
rect 19112 18115 19480 18124
rect 23112 18164 23480 18173
rect 23152 18124 23194 18164
rect 23234 18124 23276 18164
rect 23316 18124 23358 18164
rect 23398 18124 23440 18164
rect 23112 18115 23480 18124
rect 27112 18164 27480 18173
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27112 18115 27480 18124
rect 31112 18164 31480 18173
rect 31152 18124 31194 18164
rect 31234 18124 31276 18164
rect 31316 18124 31358 18164
rect 31398 18124 31440 18164
rect 31112 18115 31480 18124
rect 35112 18164 35480 18173
rect 35152 18124 35194 18164
rect 35234 18124 35276 18164
rect 35316 18124 35358 18164
rect 35398 18124 35440 18164
rect 35112 18115 35480 18124
rect 39112 18164 39480 18173
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39112 18115 39480 18124
rect 43112 18164 43480 18173
rect 43152 18124 43194 18164
rect 43234 18124 43276 18164
rect 43316 18124 43358 18164
rect 43398 18124 43440 18164
rect 43112 18115 43480 18124
rect 47112 18164 47480 18173
rect 47152 18124 47194 18164
rect 47234 18124 47276 18164
rect 47316 18124 47358 18164
rect 47398 18124 47440 18164
rect 47112 18115 47480 18124
rect 51112 18164 51480 18173
rect 51152 18124 51194 18164
rect 51234 18124 51276 18164
rect 51316 18124 51358 18164
rect 51398 18124 51440 18164
rect 51112 18115 51480 18124
rect 55112 18164 55480 18173
rect 55152 18124 55194 18164
rect 55234 18124 55276 18164
rect 55316 18124 55358 18164
rect 55398 18124 55440 18164
rect 55112 18115 55480 18124
rect 59112 18164 59480 18173
rect 59152 18124 59194 18164
rect 59234 18124 59276 18164
rect 59316 18124 59358 18164
rect 59398 18124 59440 18164
rect 59112 18115 59480 18124
rect 63112 18164 63480 18173
rect 63152 18124 63194 18164
rect 63234 18124 63276 18164
rect 63316 18124 63358 18164
rect 63398 18124 63440 18164
rect 63112 18115 63480 18124
rect 67112 18164 67480 18173
rect 67152 18124 67194 18164
rect 67234 18124 67276 18164
rect 67316 18124 67358 18164
rect 67398 18124 67440 18164
rect 67112 18115 67480 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 8352 17408 8720 17417
rect 8392 17368 8434 17408
rect 8474 17368 8516 17408
rect 8556 17368 8598 17408
rect 8638 17368 8680 17408
rect 8352 17359 8720 17368
rect 12352 17408 12720 17417
rect 12392 17368 12434 17408
rect 12474 17368 12516 17408
rect 12556 17368 12598 17408
rect 12638 17368 12680 17408
rect 12352 17359 12720 17368
rect 16352 17408 16720 17417
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16352 17359 16720 17368
rect 20352 17408 20720 17417
rect 20392 17368 20434 17408
rect 20474 17368 20516 17408
rect 20556 17368 20598 17408
rect 20638 17368 20680 17408
rect 20352 17359 20720 17368
rect 24352 17408 24720 17417
rect 24392 17368 24434 17408
rect 24474 17368 24516 17408
rect 24556 17368 24598 17408
rect 24638 17368 24680 17408
rect 24352 17359 24720 17368
rect 28352 17408 28720 17417
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28352 17359 28720 17368
rect 32352 17408 32720 17417
rect 32392 17368 32434 17408
rect 32474 17368 32516 17408
rect 32556 17368 32598 17408
rect 32638 17368 32680 17408
rect 32352 17359 32720 17368
rect 36352 17408 36720 17417
rect 36392 17368 36434 17408
rect 36474 17368 36516 17408
rect 36556 17368 36598 17408
rect 36638 17368 36680 17408
rect 36352 17359 36720 17368
rect 40352 17408 40720 17417
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40352 17359 40720 17368
rect 44352 17408 44720 17417
rect 44392 17368 44434 17408
rect 44474 17368 44516 17408
rect 44556 17368 44598 17408
rect 44638 17368 44680 17408
rect 44352 17359 44720 17368
rect 48352 17408 48720 17417
rect 48392 17368 48434 17408
rect 48474 17368 48516 17408
rect 48556 17368 48598 17408
rect 48638 17368 48680 17408
rect 48352 17359 48720 17368
rect 52352 17408 52720 17417
rect 52392 17368 52434 17408
rect 52474 17368 52516 17408
rect 52556 17368 52598 17408
rect 52638 17368 52680 17408
rect 52352 17359 52720 17368
rect 56352 17408 56720 17417
rect 56392 17368 56434 17408
rect 56474 17368 56516 17408
rect 56556 17368 56598 17408
rect 56638 17368 56680 17408
rect 56352 17359 56720 17368
rect 60352 17408 60720 17417
rect 60392 17368 60434 17408
rect 60474 17368 60516 17408
rect 60556 17368 60598 17408
rect 60638 17368 60680 17408
rect 60352 17359 60720 17368
rect 64352 17408 64720 17417
rect 64392 17368 64434 17408
rect 64474 17368 64516 17408
rect 64556 17368 64598 17408
rect 64638 17368 64680 17408
rect 64352 17359 64720 17368
rect 68352 17408 68720 17417
rect 68392 17368 68434 17408
rect 68474 17368 68516 17408
rect 68556 17368 68598 17408
rect 68638 17368 68680 17408
rect 68352 17359 68720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 7112 16652 7480 16661
rect 7152 16612 7194 16652
rect 7234 16612 7276 16652
rect 7316 16612 7358 16652
rect 7398 16612 7440 16652
rect 7112 16603 7480 16612
rect 11112 16652 11480 16661
rect 11152 16612 11194 16652
rect 11234 16612 11276 16652
rect 11316 16612 11358 16652
rect 11398 16612 11440 16652
rect 11112 16603 11480 16612
rect 15112 16652 15480 16661
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15112 16603 15480 16612
rect 19112 16652 19480 16661
rect 19152 16612 19194 16652
rect 19234 16612 19276 16652
rect 19316 16612 19358 16652
rect 19398 16612 19440 16652
rect 19112 16603 19480 16612
rect 23112 16652 23480 16661
rect 23152 16612 23194 16652
rect 23234 16612 23276 16652
rect 23316 16612 23358 16652
rect 23398 16612 23440 16652
rect 23112 16603 23480 16612
rect 27112 16652 27480 16661
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27112 16603 27480 16612
rect 31112 16652 31480 16661
rect 31152 16612 31194 16652
rect 31234 16612 31276 16652
rect 31316 16612 31358 16652
rect 31398 16612 31440 16652
rect 31112 16603 31480 16612
rect 35112 16652 35480 16661
rect 35152 16612 35194 16652
rect 35234 16612 35276 16652
rect 35316 16612 35358 16652
rect 35398 16612 35440 16652
rect 35112 16603 35480 16612
rect 39112 16652 39480 16661
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39112 16603 39480 16612
rect 43112 16652 43480 16661
rect 43152 16612 43194 16652
rect 43234 16612 43276 16652
rect 43316 16612 43358 16652
rect 43398 16612 43440 16652
rect 43112 16603 43480 16612
rect 47112 16652 47480 16661
rect 47152 16612 47194 16652
rect 47234 16612 47276 16652
rect 47316 16612 47358 16652
rect 47398 16612 47440 16652
rect 47112 16603 47480 16612
rect 51112 16652 51480 16661
rect 51152 16612 51194 16652
rect 51234 16612 51276 16652
rect 51316 16612 51358 16652
rect 51398 16612 51440 16652
rect 51112 16603 51480 16612
rect 55112 16652 55480 16661
rect 55152 16612 55194 16652
rect 55234 16612 55276 16652
rect 55316 16612 55358 16652
rect 55398 16612 55440 16652
rect 55112 16603 55480 16612
rect 59112 16652 59480 16661
rect 59152 16612 59194 16652
rect 59234 16612 59276 16652
rect 59316 16612 59358 16652
rect 59398 16612 59440 16652
rect 59112 16603 59480 16612
rect 63112 16652 63480 16661
rect 63152 16612 63194 16652
rect 63234 16612 63276 16652
rect 63316 16612 63358 16652
rect 63398 16612 63440 16652
rect 63112 16603 63480 16612
rect 67112 16652 67480 16661
rect 67152 16612 67194 16652
rect 67234 16612 67276 16652
rect 67316 16612 67358 16652
rect 67398 16612 67440 16652
rect 67112 16603 67480 16612
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 8352 15896 8720 15905
rect 8392 15856 8434 15896
rect 8474 15856 8516 15896
rect 8556 15856 8598 15896
rect 8638 15856 8680 15896
rect 8352 15847 8720 15856
rect 12352 15896 12720 15905
rect 12392 15856 12434 15896
rect 12474 15856 12516 15896
rect 12556 15856 12598 15896
rect 12638 15856 12680 15896
rect 12352 15847 12720 15856
rect 16352 15896 16720 15905
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16352 15847 16720 15856
rect 20352 15896 20720 15905
rect 20392 15856 20434 15896
rect 20474 15856 20516 15896
rect 20556 15856 20598 15896
rect 20638 15856 20680 15896
rect 20352 15847 20720 15856
rect 24352 15896 24720 15905
rect 24392 15856 24434 15896
rect 24474 15856 24516 15896
rect 24556 15856 24598 15896
rect 24638 15856 24680 15896
rect 24352 15847 24720 15856
rect 28352 15896 28720 15905
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28352 15847 28720 15856
rect 32352 15896 32720 15905
rect 32392 15856 32434 15896
rect 32474 15856 32516 15896
rect 32556 15856 32598 15896
rect 32638 15856 32680 15896
rect 32352 15847 32720 15856
rect 36352 15896 36720 15905
rect 36392 15856 36434 15896
rect 36474 15856 36516 15896
rect 36556 15856 36598 15896
rect 36638 15856 36680 15896
rect 36352 15847 36720 15856
rect 40352 15896 40720 15905
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40352 15847 40720 15856
rect 44352 15896 44720 15905
rect 44392 15856 44434 15896
rect 44474 15856 44516 15896
rect 44556 15856 44598 15896
rect 44638 15856 44680 15896
rect 44352 15847 44720 15856
rect 48352 15896 48720 15905
rect 48392 15856 48434 15896
rect 48474 15856 48516 15896
rect 48556 15856 48598 15896
rect 48638 15856 48680 15896
rect 48352 15847 48720 15856
rect 52352 15896 52720 15905
rect 52392 15856 52434 15896
rect 52474 15856 52516 15896
rect 52556 15856 52598 15896
rect 52638 15856 52680 15896
rect 52352 15847 52720 15856
rect 56352 15896 56720 15905
rect 56392 15856 56434 15896
rect 56474 15856 56516 15896
rect 56556 15856 56598 15896
rect 56638 15856 56680 15896
rect 56352 15847 56720 15856
rect 60352 15896 60720 15905
rect 60392 15856 60434 15896
rect 60474 15856 60516 15896
rect 60556 15856 60598 15896
rect 60638 15856 60680 15896
rect 60352 15847 60720 15856
rect 64352 15896 64720 15905
rect 64392 15856 64434 15896
rect 64474 15856 64516 15896
rect 64556 15856 64598 15896
rect 64638 15856 64680 15896
rect 64352 15847 64720 15856
rect 68352 15896 68720 15905
rect 68392 15856 68434 15896
rect 68474 15856 68516 15896
rect 68556 15856 68598 15896
rect 68638 15856 68680 15896
rect 68352 15847 68720 15856
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 7112 15140 7480 15149
rect 7152 15100 7194 15140
rect 7234 15100 7276 15140
rect 7316 15100 7358 15140
rect 7398 15100 7440 15140
rect 7112 15091 7480 15100
rect 11112 15140 11480 15149
rect 11152 15100 11194 15140
rect 11234 15100 11276 15140
rect 11316 15100 11358 15140
rect 11398 15100 11440 15140
rect 11112 15091 11480 15100
rect 15112 15140 15480 15149
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15112 15091 15480 15100
rect 19112 15140 19480 15149
rect 19152 15100 19194 15140
rect 19234 15100 19276 15140
rect 19316 15100 19358 15140
rect 19398 15100 19440 15140
rect 19112 15091 19480 15100
rect 23112 15140 23480 15149
rect 23152 15100 23194 15140
rect 23234 15100 23276 15140
rect 23316 15100 23358 15140
rect 23398 15100 23440 15140
rect 23112 15091 23480 15100
rect 27112 15140 27480 15149
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27112 15091 27480 15100
rect 31112 15140 31480 15149
rect 31152 15100 31194 15140
rect 31234 15100 31276 15140
rect 31316 15100 31358 15140
rect 31398 15100 31440 15140
rect 31112 15091 31480 15100
rect 35112 15140 35480 15149
rect 35152 15100 35194 15140
rect 35234 15100 35276 15140
rect 35316 15100 35358 15140
rect 35398 15100 35440 15140
rect 35112 15091 35480 15100
rect 39112 15140 39480 15149
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39112 15091 39480 15100
rect 43112 15140 43480 15149
rect 43152 15100 43194 15140
rect 43234 15100 43276 15140
rect 43316 15100 43358 15140
rect 43398 15100 43440 15140
rect 43112 15091 43480 15100
rect 47112 15140 47480 15149
rect 47152 15100 47194 15140
rect 47234 15100 47276 15140
rect 47316 15100 47358 15140
rect 47398 15100 47440 15140
rect 47112 15091 47480 15100
rect 51112 15140 51480 15149
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51112 15091 51480 15100
rect 55112 15140 55480 15149
rect 55152 15100 55194 15140
rect 55234 15100 55276 15140
rect 55316 15100 55358 15140
rect 55398 15100 55440 15140
rect 55112 15091 55480 15100
rect 59112 15140 59480 15149
rect 59152 15100 59194 15140
rect 59234 15100 59276 15140
rect 59316 15100 59358 15140
rect 59398 15100 59440 15140
rect 59112 15091 59480 15100
rect 63112 15140 63480 15149
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63112 15091 63480 15100
rect 67112 15140 67480 15149
rect 67152 15100 67194 15140
rect 67234 15100 67276 15140
rect 67316 15100 67358 15140
rect 67398 15100 67440 15140
rect 71020 15140 71060 24583
rect 73228 24498 73268 24583
rect 73612 24557 73652 24592
rect 73611 24548 73653 24557
rect 73611 24508 73612 24548
rect 73652 24508 73653 24548
rect 73611 24499 73653 24508
rect 73804 24548 73844 25675
rect 73900 25388 73940 25397
rect 73900 25145 73940 25348
rect 73899 25136 73941 25145
rect 73899 25096 73900 25136
rect 73940 25096 73941 25136
rect 73899 25087 73941 25096
rect 73996 24977 74036 26440
rect 74305 26396 74345 26796
rect 74092 26356 74345 26396
rect 74092 25556 74132 26356
rect 74415 26312 74455 26796
rect 74705 26396 74745 26796
rect 74092 25507 74132 25516
rect 74380 26272 74455 26312
rect 74668 26356 74745 26396
rect 74815 26396 74855 26796
rect 75105 26396 75145 26796
rect 75215 26489 75255 26796
rect 75214 26480 75256 26489
rect 75214 26440 75215 26480
rect 75255 26440 75256 26480
rect 75214 26431 75256 26440
rect 75505 26396 75545 26796
rect 74815 26356 74900 26396
rect 74283 25136 74325 25145
rect 74283 25096 74284 25136
rect 74324 25096 74325 25136
rect 74283 25087 74325 25096
rect 73995 24968 74037 24977
rect 73995 24928 73996 24968
rect 74036 24928 74037 24968
rect 73995 24919 74037 24928
rect 73996 24800 74036 24811
rect 73996 24725 74036 24760
rect 73995 24716 74037 24725
rect 73995 24676 73996 24716
rect 74036 24676 74037 24716
rect 73995 24667 74037 24676
rect 74187 24716 74229 24725
rect 74187 24676 74188 24716
rect 74228 24676 74229 24716
rect 74187 24667 74229 24676
rect 73804 24499 73844 24508
rect 74188 24548 74228 24667
rect 74284 24557 74324 25087
rect 74380 24809 74420 26272
rect 74668 26069 74708 26356
rect 74667 26060 74709 26069
rect 74667 26020 74668 26060
rect 74708 26020 74709 26060
rect 74667 26011 74709 26020
rect 74860 25565 74900 26356
rect 74956 26356 75145 26396
rect 75436 26356 75545 26396
rect 75615 26396 75655 26796
rect 75905 26396 75945 26796
rect 76015 26396 76055 26796
rect 76203 26480 76245 26489
rect 76203 26440 76204 26480
rect 76244 26440 76245 26480
rect 76203 26431 76245 26440
rect 75615 26356 75668 26396
rect 74859 25556 74901 25565
rect 74859 25516 74860 25556
rect 74900 25516 74901 25556
rect 74859 25507 74901 25516
rect 74668 25472 74708 25483
rect 74668 25397 74708 25432
rect 74475 25388 74517 25397
rect 74475 25348 74476 25388
rect 74516 25348 74517 25388
rect 74475 25339 74517 25348
rect 74667 25388 74709 25397
rect 74860 25388 74900 25397
rect 74667 25348 74668 25388
rect 74708 25348 74709 25388
rect 74667 25339 74709 25348
rect 74764 25348 74860 25388
rect 74476 25254 74516 25339
rect 74379 24800 74421 24809
rect 74379 24760 74380 24800
rect 74420 24760 74421 24800
rect 74379 24751 74421 24760
rect 74188 24499 74228 24508
rect 74283 24548 74325 24557
rect 74283 24508 74284 24548
rect 74324 24508 74325 24548
rect 74283 24499 74325 24508
rect 74667 24548 74709 24557
rect 74667 24508 74668 24548
rect 74708 24508 74709 24548
rect 74667 24499 74709 24508
rect 74668 24414 74708 24499
rect 74764 24389 74804 25348
rect 74860 25339 74900 25348
rect 74860 24800 74900 24809
rect 74956 24800 74996 26356
rect 75243 25472 75285 25481
rect 75243 25432 75244 25472
rect 75284 25432 75285 25472
rect 75243 25423 75285 25432
rect 75051 25388 75093 25397
rect 75051 25348 75052 25388
rect 75092 25348 75093 25388
rect 75051 25339 75093 25348
rect 75052 25254 75092 25339
rect 75244 25338 75284 25423
rect 74900 24760 74996 24800
rect 75436 24800 75476 26356
rect 75531 25472 75573 25481
rect 75531 25432 75532 25472
rect 75572 25432 75573 25472
rect 75531 25423 75573 25432
rect 75532 25388 75572 25423
rect 75532 25313 75572 25348
rect 75531 25304 75573 25313
rect 75531 25264 75532 25304
rect 75572 25264 75573 25304
rect 75531 25255 75573 25264
rect 75532 25224 75572 25255
rect 74860 24751 74900 24760
rect 75436 24751 75476 24760
rect 75628 24800 75668 26356
rect 75724 26356 75945 26396
rect 76012 26356 76055 26396
rect 75724 25556 75764 26356
rect 75724 25507 75764 25516
rect 75915 25556 75957 25565
rect 75915 25516 75916 25556
rect 75956 25516 75957 25556
rect 75915 25507 75957 25516
rect 75916 25422 75956 25507
rect 76012 25481 76052 26356
rect 76204 25556 76244 26431
rect 76305 26396 76345 26796
rect 76415 26480 76455 26796
rect 76705 26480 76745 26796
rect 76415 26440 76532 26480
rect 76305 26356 76436 26396
rect 76204 25507 76244 25516
rect 76011 25472 76053 25481
rect 76011 25432 76012 25472
rect 76052 25432 76053 25472
rect 76011 25423 76053 25432
rect 76011 25304 76053 25313
rect 76011 25264 76012 25304
rect 76052 25264 76053 25304
rect 76011 25255 76053 25264
rect 76299 25304 76341 25313
rect 76299 25264 76300 25304
rect 76340 25264 76341 25304
rect 76299 25255 76341 25264
rect 76012 25170 76052 25255
rect 76300 25170 76340 25255
rect 75628 24751 75668 24760
rect 76204 24800 76244 24809
rect 76396 24800 76436 26356
rect 76492 25649 76532 26440
rect 76684 26440 76745 26480
rect 76491 25640 76533 25649
rect 76491 25600 76492 25640
rect 76532 25600 76533 25640
rect 76491 25591 76533 25600
rect 76491 25472 76533 25481
rect 76491 25432 76492 25472
rect 76532 25432 76533 25472
rect 76491 25423 76533 25432
rect 76492 25338 76532 25423
rect 76587 25304 76629 25313
rect 76587 25264 76588 25304
rect 76628 25264 76629 25304
rect 76587 25255 76629 25264
rect 76588 25170 76628 25255
rect 76244 24760 76436 24800
rect 76588 24800 76628 24809
rect 76684 24800 76724 26440
rect 76815 26396 76855 26796
rect 77105 26396 77145 26796
rect 77215 26489 77255 26796
rect 77214 26480 77256 26489
rect 77214 26440 77215 26480
rect 77255 26440 77256 26480
rect 77214 26431 77256 26440
rect 77505 26396 77545 26796
rect 76780 26356 76855 26396
rect 76972 26356 77145 26396
rect 77452 26356 77545 26396
rect 77615 26396 77655 26796
rect 77905 26480 77945 26796
rect 77836 26440 77945 26480
rect 77615 26356 77684 26396
rect 76780 25565 76820 26356
rect 76875 25640 76917 25649
rect 76875 25600 76876 25640
rect 76916 25600 76917 25640
rect 76875 25591 76917 25600
rect 76779 25556 76821 25565
rect 76779 25516 76780 25556
rect 76820 25516 76821 25556
rect 76779 25507 76821 25516
rect 76876 25556 76916 25591
rect 76876 25505 76916 25516
rect 76779 25304 76821 25313
rect 76779 25264 76780 25304
rect 76820 25264 76821 25304
rect 76779 25255 76821 25264
rect 76780 25170 76820 25255
rect 76875 24968 76917 24977
rect 76875 24928 76876 24968
rect 76916 24928 76917 24968
rect 76875 24919 76917 24928
rect 76628 24760 76724 24800
rect 76204 24751 76244 24760
rect 76588 24751 76628 24760
rect 75723 24716 75765 24725
rect 75723 24676 75724 24716
rect 75764 24676 75765 24716
rect 75723 24667 75765 24676
rect 75724 24632 75764 24667
rect 75724 24581 75764 24592
rect 76876 24557 76916 24919
rect 76972 24800 77012 26356
rect 77163 25556 77205 25565
rect 77163 25516 77164 25556
rect 77204 25516 77205 25556
rect 77163 25507 77205 25516
rect 77164 25422 77204 25507
rect 77068 25304 77108 25313
rect 77068 24977 77108 25264
rect 77067 24968 77109 24977
rect 77067 24928 77068 24968
rect 77108 24928 77109 24968
rect 77067 24919 77109 24928
rect 77068 24800 77108 24809
rect 76972 24760 77068 24800
rect 77068 24751 77108 24760
rect 77452 24800 77492 26356
rect 77644 25565 77684 26356
rect 77643 25556 77685 25565
rect 77643 25516 77644 25556
rect 77684 25516 77685 25556
rect 77643 25507 77685 25516
rect 77740 25472 77780 25481
rect 77547 25388 77589 25397
rect 77547 25348 77548 25388
rect 77588 25348 77589 25388
rect 77547 25339 77589 25348
rect 77452 24751 77492 24760
rect 75243 24548 75285 24557
rect 75243 24508 75244 24548
rect 75284 24508 75285 24548
rect 75243 24499 75285 24508
rect 76011 24548 76053 24557
rect 76011 24508 76012 24548
rect 76052 24508 76053 24548
rect 76011 24499 76053 24508
rect 76395 24548 76437 24557
rect 76395 24508 76396 24548
rect 76436 24508 76437 24548
rect 76395 24499 76437 24508
rect 76875 24548 76917 24557
rect 76875 24508 76876 24548
rect 76916 24508 76917 24548
rect 76875 24499 76917 24508
rect 77259 24548 77301 24557
rect 77259 24508 77260 24548
rect 77300 24508 77301 24548
rect 77548 24548 77588 25339
rect 77740 25313 77780 25432
rect 77739 25304 77781 25313
rect 77739 25264 77740 25304
rect 77780 25264 77781 25304
rect 77739 25255 77781 25264
rect 77836 25220 77876 26440
rect 78015 26396 78055 26796
rect 78305 26396 78345 26796
rect 78415 26648 78455 26796
rect 78415 26608 78644 26648
rect 78507 26480 78549 26489
rect 78507 26440 78508 26480
rect 78548 26440 78549 26480
rect 78507 26431 78549 26440
rect 78015 26356 78260 26396
rect 78305 26356 78452 26396
rect 77931 25556 77973 25565
rect 77931 25516 77932 25556
rect 77972 25516 77973 25556
rect 77931 25507 77973 25516
rect 78220 25556 78260 26356
rect 78220 25507 78260 25516
rect 77932 25422 77972 25507
rect 78027 25304 78069 25313
rect 78027 25264 78028 25304
rect 78068 25264 78069 25304
rect 78027 25255 78069 25264
rect 78315 25304 78357 25313
rect 78315 25264 78316 25304
rect 78356 25264 78357 25304
rect 78315 25255 78357 25264
rect 77836 25180 77972 25220
rect 77932 24800 77972 25180
rect 78028 25170 78068 25255
rect 78316 25170 78356 25255
rect 78028 24800 78068 24809
rect 77932 24760 78028 24800
rect 78028 24751 78068 24760
rect 78412 24800 78452 26356
rect 78508 25556 78548 26431
rect 78604 25565 78644 26608
rect 78705 26396 78745 26796
rect 78815 26396 78855 26796
rect 79105 26480 79145 26796
rect 78700 26356 78745 26396
rect 78796 26356 78855 26396
rect 79084 26440 79145 26480
rect 78508 25507 78548 25516
rect 78603 25556 78645 25565
rect 78603 25516 78604 25556
rect 78644 25516 78645 25556
rect 78603 25507 78645 25516
rect 78412 24751 78452 24760
rect 78604 25304 78644 25313
rect 78604 24557 78644 25264
rect 78700 24800 78740 26356
rect 78796 25556 78836 26356
rect 78796 25507 78836 25516
rect 79084 25388 79124 26440
rect 79215 26396 79255 26796
rect 79505 26480 79545 26796
rect 79180 26356 79255 26396
rect 79468 26440 79545 26480
rect 79180 25556 79220 26356
rect 79180 25507 79220 25516
rect 79468 25388 79508 26440
rect 79615 26396 79655 26796
rect 79564 26356 79655 26396
rect 79905 26396 79945 26796
rect 80015 26480 80055 26796
rect 80305 26480 80345 26796
rect 80015 26440 80180 26480
rect 79905 26356 79988 26396
rect 79564 25556 79604 26356
rect 79564 25507 79604 25516
rect 79755 25556 79797 25565
rect 79755 25516 79756 25556
rect 79796 25516 79797 25556
rect 79755 25507 79797 25516
rect 79756 25422 79796 25507
rect 79084 25348 79220 25388
rect 79468 25348 79604 25388
rect 78891 25304 78933 25313
rect 78891 25264 78892 25304
rect 78932 25293 79111 25304
rect 78932 25264 79071 25293
rect 78891 25255 78933 25264
rect 78892 25170 78932 25255
rect 79071 25244 79111 25253
rect 78796 24800 78836 24809
rect 78700 24760 78796 24800
rect 78796 24751 78836 24760
rect 79180 24800 79220 25348
rect 79371 25304 79413 25313
rect 79371 25264 79372 25304
rect 79412 25293 79508 25304
rect 79412 25264 79468 25293
rect 79371 25255 79413 25264
rect 79468 25244 79508 25253
rect 79180 24751 79220 24760
rect 79564 24800 79604 25348
rect 79851 25304 79893 25313
rect 79851 25264 79852 25304
rect 79892 25264 79893 25304
rect 79851 25255 79893 25264
rect 79852 25170 79892 25255
rect 79564 24751 79604 24760
rect 79948 24800 79988 26356
rect 80140 25556 80180 26440
rect 80140 25507 80180 25516
rect 80236 26440 80345 26480
rect 80043 25304 80085 25313
rect 80043 25264 80044 25304
rect 80084 25264 80085 25304
rect 80043 25255 80085 25264
rect 80044 25170 80084 25255
rect 79948 24751 79988 24760
rect 77644 24548 77684 24557
rect 77548 24508 77644 24548
rect 77259 24499 77301 24508
rect 77644 24499 77684 24508
rect 77835 24548 77877 24557
rect 77835 24508 77836 24548
rect 77876 24508 77877 24548
rect 77835 24499 77877 24508
rect 78219 24548 78261 24557
rect 78219 24508 78220 24548
rect 78260 24508 78261 24548
rect 78219 24499 78261 24508
rect 78603 24548 78645 24557
rect 78603 24508 78604 24548
rect 78644 24508 78645 24548
rect 78603 24499 78645 24508
rect 78987 24548 79029 24557
rect 78987 24508 78988 24548
rect 79028 24508 79029 24548
rect 78987 24499 79029 24508
rect 79371 24548 79413 24557
rect 79371 24508 79372 24548
rect 79412 24508 79413 24548
rect 79371 24499 79413 24508
rect 79755 24548 79797 24557
rect 79755 24508 79756 24548
rect 79796 24508 79797 24548
rect 79755 24499 79797 24508
rect 80139 24548 80181 24557
rect 80139 24508 80140 24548
rect 80180 24508 80181 24548
rect 80139 24499 80181 24508
rect 75244 24414 75284 24499
rect 76012 24414 76052 24499
rect 76396 24414 76436 24499
rect 76876 24414 76916 24499
rect 77260 24414 77300 24499
rect 77836 24464 77876 24499
rect 77836 24413 77876 24424
rect 78220 24414 78260 24499
rect 78604 24414 78644 24499
rect 78988 24414 79028 24499
rect 79372 24414 79412 24499
rect 79756 24414 79796 24499
rect 80140 24414 80180 24499
rect 74379 24380 74421 24389
rect 74379 24340 74380 24380
rect 74420 24340 74421 24380
rect 74379 24331 74421 24340
rect 74763 24380 74805 24389
rect 74763 24340 74764 24380
rect 74804 24340 74805 24380
rect 74763 24331 74805 24340
rect 74380 24246 74420 24331
rect 71112 24212 71480 24221
rect 71152 24172 71194 24212
rect 71234 24172 71276 24212
rect 71316 24172 71358 24212
rect 71398 24172 71440 24212
rect 71112 24163 71480 24172
rect 75112 24212 75480 24221
rect 75152 24172 75194 24212
rect 75234 24172 75276 24212
rect 75316 24172 75358 24212
rect 75398 24172 75440 24212
rect 75112 24163 75480 24172
rect 79112 24212 79480 24221
rect 79152 24172 79194 24212
rect 79234 24172 79276 24212
rect 79316 24172 79358 24212
rect 79398 24172 79440 24212
rect 79112 24163 79480 24172
rect 80140 23960 80180 23969
rect 80236 23960 80276 26440
rect 80415 26396 80455 26796
rect 80332 26356 80455 26396
rect 80705 26396 80745 26796
rect 80815 26396 80855 26796
rect 81105 26396 81145 26796
rect 81215 26396 81255 26796
rect 81505 26480 81545 26796
rect 80705 26356 80756 26396
rect 80332 25556 80372 26356
rect 80332 25507 80372 25516
rect 80716 25388 80756 26356
rect 80812 26356 80855 26396
rect 81100 26356 81145 26396
rect 81196 26356 81255 26396
rect 81388 26440 81545 26480
rect 80812 25556 80852 26356
rect 80812 25507 80852 25516
rect 81100 25388 81140 26356
rect 81196 25556 81236 26356
rect 81196 25507 81236 25516
rect 81195 25388 81237 25397
rect 80716 25348 81044 25388
rect 81100 25348 81196 25388
rect 81236 25348 81237 25388
rect 80428 25304 80468 25315
rect 80428 25229 80468 25264
rect 80716 25293 80756 25302
rect 80716 25229 80756 25253
rect 80427 25220 80469 25229
rect 80427 25180 80428 25220
rect 80468 25180 80469 25220
rect 80427 25171 80469 25180
rect 80715 25220 80757 25229
rect 80715 25180 80716 25220
rect 80756 25180 80757 25220
rect 80715 25171 80757 25180
rect 80907 25220 80949 25229
rect 80907 25180 80908 25220
rect 80948 25180 80949 25220
rect 80907 25171 80949 25180
rect 80428 24632 80468 25171
rect 80716 25158 80756 25171
rect 80428 24583 80468 24592
rect 80620 24632 80660 24641
rect 80620 24389 80660 24592
rect 80908 24548 80948 25171
rect 81004 24800 81044 25348
rect 81195 25339 81237 25348
rect 81100 25293 81140 25302
rect 81100 25229 81140 25253
rect 81099 25220 81141 25229
rect 81099 25180 81100 25220
rect 81140 25180 81141 25220
rect 81099 25171 81141 25180
rect 81100 25158 81140 25171
rect 81388 24809 81428 26440
rect 81615 26396 81655 26796
rect 81580 26356 81655 26396
rect 81580 25556 81620 26356
rect 81905 26312 81945 26796
rect 82015 26396 82055 26796
rect 82305 26480 82345 26796
rect 82252 26440 82345 26480
rect 82015 26356 82100 26396
rect 81905 26272 82004 26312
rect 81580 25507 81620 25516
rect 81964 25472 82004 26272
rect 82060 25556 82100 26356
rect 82060 25507 82100 25516
rect 81868 25432 82004 25472
rect 81579 25388 81621 25397
rect 81579 25348 81580 25388
rect 81620 25348 81621 25388
rect 81579 25339 81621 25348
rect 81484 25304 81524 25315
rect 81484 25229 81524 25264
rect 81483 25220 81525 25229
rect 81483 25180 81484 25220
rect 81524 25180 81525 25220
rect 81483 25171 81525 25180
rect 81196 24800 81236 24809
rect 81004 24760 81196 24800
rect 81196 24751 81236 24760
rect 81387 24800 81429 24809
rect 81387 24760 81388 24800
rect 81428 24760 81429 24800
rect 81387 24751 81429 24760
rect 81580 24800 81620 25339
rect 81580 24751 81620 24760
rect 81004 24548 81044 24557
rect 80908 24508 81004 24548
rect 81004 24499 81044 24508
rect 81388 24548 81428 24557
rect 80619 24380 80661 24389
rect 80619 24340 80620 24380
rect 80660 24340 80661 24380
rect 80619 24331 80661 24340
rect 80812 24380 80852 24389
rect 80180 23920 80276 23960
rect 80140 23911 80180 23920
rect 80812 23885 80852 24340
rect 81388 23885 81428 24508
rect 81772 24548 81812 24557
rect 80331 23876 80373 23885
rect 80331 23836 80332 23876
rect 80372 23836 80373 23876
rect 80331 23827 80373 23836
rect 80811 23876 80853 23885
rect 80811 23836 80812 23876
rect 80852 23836 80853 23876
rect 80811 23827 80853 23836
rect 81387 23876 81429 23885
rect 81387 23836 81388 23876
rect 81428 23836 81429 23876
rect 81387 23827 81429 23836
rect 81675 23876 81717 23885
rect 81772 23876 81812 24508
rect 81868 24044 81908 25432
rect 82252 25388 82292 26440
rect 82415 26396 82455 26796
rect 82705 26480 82745 26796
rect 82348 26356 82455 26396
rect 82540 26440 82745 26480
rect 82348 25556 82388 26356
rect 82348 25507 82388 25516
rect 82252 25348 82388 25388
rect 81964 25304 82004 25313
rect 82004 25264 82100 25304
rect 81964 25255 82004 25264
rect 81963 24800 82005 24809
rect 81963 24760 81964 24800
rect 82004 24760 82005 24800
rect 81963 24751 82005 24760
rect 81964 24666 82004 24751
rect 82060 24548 82100 25264
rect 82252 25293 82292 25302
rect 82252 25229 82292 25253
rect 82251 25220 82293 25229
rect 82251 25180 82252 25220
rect 82292 25180 82293 25220
rect 82251 25171 82293 25180
rect 82252 25158 82292 25171
rect 82348 24800 82388 25348
rect 82540 25136 82580 26440
rect 82815 26396 82855 26796
rect 83105 26396 83145 26796
rect 83215 26396 83255 26796
rect 83505 26396 83545 26796
rect 82732 26356 82855 26396
rect 83020 26356 83145 26396
rect 83212 26356 83255 26396
rect 83500 26356 83545 26396
rect 83615 26396 83655 26796
rect 83905 26396 83945 26796
rect 83615 26356 83732 26396
rect 82732 25556 82772 26356
rect 82732 25507 82772 25516
rect 82636 25304 82676 25313
rect 82636 25220 82676 25264
rect 82731 25220 82773 25229
rect 82636 25180 82732 25220
rect 82772 25180 82773 25220
rect 82731 25171 82773 25180
rect 82540 25096 82676 25136
rect 82348 24751 82388 24760
rect 82156 24548 82196 24557
rect 82060 24508 82156 24548
rect 81868 23995 81908 24004
rect 82156 23885 82196 24508
rect 82540 24548 82580 24557
rect 81675 23836 81676 23876
rect 81716 23836 81812 23876
rect 82155 23876 82197 23885
rect 82155 23836 82156 23876
rect 82196 23836 82197 23876
rect 81675 23827 81717 23836
rect 82155 23827 82197 23836
rect 82443 23876 82485 23885
rect 82540 23876 82580 24508
rect 82636 23960 82676 25096
rect 82732 24548 82772 25171
rect 83020 24800 83060 26356
rect 83116 25556 83156 25565
rect 83212 25556 83252 26356
rect 83156 25516 83252 25556
rect 83116 25507 83156 25516
rect 83212 25304 83252 25313
rect 83116 24800 83156 24809
rect 83020 24760 83116 24800
rect 83116 24751 83156 24760
rect 82924 24548 82964 24557
rect 82732 24508 82924 24548
rect 83212 24548 83252 25264
rect 83500 24800 83540 26356
rect 83692 25565 83732 26356
rect 83884 26356 83945 26396
rect 84015 26396 84055 26796
rect 84305 26396 84345 26796
rect 84415 26480 84455 26796
rect 84415 26440 84596 26480
rect 84015 26356 84116 26396
rect 84305 26356 84404 26396
rect 83691 25556 83733 25565
rect 83691 25516 83692 25556
rect 83732 25516 83733 25556
rect 83691 25507 83733 25516
rect 83788 25472 83828 25481
rect 83500 24751 83540 24760
rect 83596 25388 83636 25397
rect 83307 24548 83349 24557
rect 83212 24508 83308 24548
rect 83348 24508 83349 24548
rect 82924 24499 82964 24508
rect 83307 24499 83349 24508
rect 83308 24414 83348 24499
rect 83596 24389 83636 25348
rect 83788 25313 83828 25432
rect 83787 25304 83829 25313
rect 83787 25264 83788 25304
rect 83828 25264 83829 25304
rect 83787 25255 83829 25264
rect 83884 24800 83924 26356
rect 83979 25556 84021 25565
rect 83979 25516 83980 25556
rect 84020 25516 84021 25556
rect 84076 25556 84116 26356
rect 84268 25556 84308 25565
rect 84076 25516 84268 25556
rect 83979 25507 84021 25516
rect 84268 25507 84308 25516
rect 83980 25422 84020 25507
rect 84364 25472 84404 26356
rect 84556 25556 84596 26440
rect 84705 26312 84745 26796
rect 84815 26396 84855 26796
rect 85105 26396 85145 26796
rect 84815 26356 84884 26396
rect 84705 26272 84788 26312
rect 84556 25507 84596 25516
rect 84364 25432 84500 25472
rect 84075 25304 84117 25313
rect 84075 25264 84076 25304
rect 84116 25264 84117 25304
rect 84075 25255 84117 25264
rect 84363 25304 84405 25313
rect 84363 25264 84364 25304
rect 84404 25264 84405 25304
rect 84363 25255 84405 25264
rect 84076 25170 84116 25255
rect 84364 25170 84404 25255
rect 83884 24751 83924 24760
rect 84460 24800 84500 25432
rect 84651 25304 84693 25313
rect 84651 25264 84652 25304
rect 84692 25264 84693 25304
rect 84651 25255 84693 25264
rect 84652 25170 84692 25255
rect 84748 24800 84788 26272
rect 84844 25556 84884 26356
rect 84844 25507 84884 25516
rect 85036 26356 85145 26396
rect 85215 26396 85255 26796
rect 85505 26396 85545 26796
rect 85615 26396 85655 26796
rect 85905 26396 85945 26796
rect 86015 26396 86055 26796
rect 86305 26396 86345 26796
rect 85215 26356 85268 26396
rect 84939 25304 84981 25313
rect 84939 25264 84940 25304
rect 84980 25264 84981 25304
rect 84939 25255 84981 25264
rect 84940 25170 84980 25255
rect 85036 25136 85076 26356
rect 85228 25556 85268 26356
rect 85228 25507 85268 25516
rect 85420 26356 85545 26396
rect 85612 26356 85655 26396
rect 85804 26356 85945 26396
rect 85996 26356 86055 26396
rect 86284 26356 86345 26396
rect 85132 25313 85172 25398
rect 85131 25304 85173 25313
rect 85131 25264 85132 25304
rect 85172 25264 85173 25304
rect 85131 25255 85173 25264
rect 85036 25096 85172 25136
rect 84844 24800 84884 24809
rect 84748 24760 84844 24800
rect 84460 24751 84500 24760
rect 84844 24751 84884 24760
rect 83691 24548 83733 24557
rect 83691 24508 83692 24548
rect 83732 24508 83733 24548
rect 83691 24499 83733 24508
rect 84076 24548 84116 24557
rect 83692 24414 83732 24499
rect 84076 24389 84116 24508
rect 84267 24548 84309 24557
rect 84267 24508 84268 24548
rect 84308 24508 84309 24548
rect 84267 24499 84309 24508
rect 84651 24548 84693 24557
rect 85035 24548 85077 24557
rect 84651 24508 84652 24548
rect 84692 24508 84693 24548
rect 84651 24499 84693 24508
rect 84940 24508 85036 24548
rect 85076 24508 85077 24548
rect 84268 24464 84308 24499
rect 84268 24413 84308 24424
rect 84652 24414 84692 24499
rect 83595 24380 83637 24389
rect 83595 24340 83596 24380
rect 83636 24340 83637 24380
rect 83595 24331 83637 24340
rect 84075 24380 84117 24389
rect 84075 24340 84076 24380
rect 84116 24340 84117 24380
rect 84075 24331 84117 24340
rect 83112 24212 83480 24221
rect 83152 24172 83194 24212
rect 83234 24172 83276 24212
rect 83316 24172 83358 24212
rect 83398 24172 83440 24212
rect 83112 24163 83480 24172
rect 82636 23911 82676 23920
rect 84940 23885 84980 24508
rect 85035 24499 85077 24508
rect 85036 24414 85076 24499
rect 85132 23960 85172 25096
rect 85420 24800 85460 26356
rect 85612 25556 85652 26356
rect 85612 25507 85652 25516
rect 85515 25304 85557 25313
rect 85515 25264 85516 25304
rect 85556 25264 85557 25304
rect 85515 25255 85557 25264
rect 85516 25170 85556 25255
rect 85516 24800 85556 24809
rect 85420 24760 85516 24800
rect 85516 24751 85556 24760
rect 85323 24548 85365 24557
rect 85323 24508 85324 24548
rect 85364 24508 85365 24548
rect 85323 24499 85365 24508
rect 85324 24414 85364 24499
rect 85804 23960 85844 26356
rect 85996 25556 86036 26356
rect 85996 25507 86036 25516
rect 85899 25304 85941 25313
rect 85899 25264 85900 25304
rect 85940 25264 85941 25304
rect 85899 25255 85941 25264
rect 85900 25170 85940 25255
rect 86284 24800 86324 26356
rect 86415 26312 86455 26796
rect 86705 26396 86745 26796
rect 86380 26272 86455 26312
rect 86668 26356 86745 26396
rect 86815 26396 86855 26796
rect 87105 26396 87145 26796
rect 86815 26356 86900 26396
rect 86380 25556 86420 26272
rect 86380 25507 86420 25516
rect 86476 25304 86516 25332
rect 86571 25304 86613 25313
rect 86516 25264 86572 25304
rect 86612 25264 86613 25304
rect 86476 25255 86516 25264
rect 86571 25255 86613 25264
rect 86284 24751 86324 24760
rect 86091 24548 86133 24557
rect 86091 24508 86092 24548
rect 86132 24508 86133 24548
rect 86091 24499 86133 24508
rect 86475 24548 86517 24557
rect 86475 24508 86476 24548
rect 86516 24508 86517 24548
rect 86475 24499 86517 24508
rect 86572 24548 86612 25255
rect 86572 24499 86612 24508
rect 86092 24414 86132 24499
rect 85900 23960 85940 23969
rect 85804 23920 85900 23960
rect 85132 23911 85172 23920
rect 85900 23911 85940 23920
rect 82443 23836 82444 23876
rect 82484 23836 82580 23876
rect 84939 23876 84981 23885
rect 84939 23836 84940 23876
rect 84980 23836 84981 23876
rect 82443 23827 82485 23836
rect 84939 23827 84981 23836
rect 85707 23876 85749 23885
rect 85707 23836 85708 23876
rect 85748 23836 85749 23876
rect 85707 23827 85749 23836
rect 86476 23876 86516 24499
rect 86668 23960 86708 26356
rect 86860 25565 86900 26356
rect 87052 26356 87145 26396
rect 87215 26396 87255 26796
rect 87505 26396 87545 26796
rect 87215 26356 87284 26396
rect 86859 25556 86901 25565
rect 86859 25516 86860 25556
rect 86900 25516 86901 25556
rect 86859 25507 86901 25516
rect 86955 25472 86997 25481
rect 86955 25432 86956 25472
rect 86996 25432 86997 25472
rect 86955 25423 86997 25432
rect 86763 25304 86805 25313
rect 86763 25264 86764 25304
rect 86804 25264 86805 25304
rect 86763 25255 86805 25264
rect 86956 25304 86996 25423
rect 86956 25255 86996 25264
rect 86764 25170 86804 25255
rect 87052 24800 87092 26356
rect 87147 25388 87189 25397
rect 87147 25348 87148 25388
rect 87188 25348 87189 25388
rect 87147 25339 87189 25348
rect 87148 25254 87188 25339
rect 87148 24800 87188 24809
rect 87052 24760 87148 24800
rect 87148 24751 87188 24760
rect 87244 24716 87284 26356
rect 87436 26356 87545 26396
rect 87615 26396 87655 26796
rect 87905 26396 87945 26796
rect 88015 26396 88055 26796
rect 88305 26396 88345 26796
rect 88415 26396 88455 26796
rect 88705 26480 88745 26796
rect 87615 26356 87860 26396
rect 87905 26356 87956 26396
rect 88015 26356 88148 26396
rect 87340 25472 87380 25483
rect 87340 25397 87380 25432
rect 87339 25388 87381 25397
rect 87339 25348 87340 25388
rect 87380 25348 87381 25388
rect 87339 25339 87381 25348
rect 87436 24800 87476 26356
rect 87531 25556 87573 25565
rect 87531 25516 87532 25556
rect 87572 25516 87573 25556
rect 87531 25507 87573 25516
rect 87820 25556 87860 26356
rect 87820 25507 87860 25516
rect 87532 25422 87572 25507
rect 87916 25472 87956 26356
rect 88108 25556 88148 26356
rect 88108 25507 88148 25516
rect 88300 26356 88345 26396
rect 88396 26356 88455 26396
rect 88588 26440 88745 26480
rect 87916 25432 88052 25472
rect 87627 25304 87669 25313
rect 87627 25264 87628 25304
rect 87668 25264 87669 25304
rect 87627 25255 87669 25264
rect 87915 25304 87957 25313
rect 87915 25264 87916 25304
rect 87956 25264 87957 25304
rect 87915 25255 87957 25264
rect 87628 25170 87668 25255
rect 87916 25170 87956 25255
rect 87532 24800 87572 24809
rect 87436 24760 87532 24800
rect 87532 24751 87572 24760
rect 87244 24676 87476 24716
rect 87436 24632 87476 24676
rect 87724 24632 87764 24641
rect 87436 24592 87724 24632
rect 87724 24583 87764 24592
rect 87820 24632 87860 24643
rect 87820 24557 87860 24592
rect 86763 24548 86805 24557
rect 86763 24508 86764 24548
rect 86804 24508 86805 24548
rect 86763 24499 86805 24508
rect 86955 24548 86997 24557
rect 86955 24508 86956 24548
rect 86996 24508 86997 24548
rect 86955 24499 86997 24508
rect 87339 24548 87381 24557
rect 87339 24508 87340 24548
rect 87380 24508 87381 24548
rect 87339 24499 87381 24508
rect 87819 24548 87861 24557
rect 87819 24508 87820 24548
rect 87860 24508 87861 24548
rect 87819 24499 87861 24508
rect 86764 24464 86804 24499
rect 86764 24413 86804 24424
rect 86956 24414 86996 24499
rect 87340 24414 87380 24499
rect 87112 24212 87480 24221
rect 87152 24172 87194 24212
rect 87234 24172 87276 24212
rect 87316 24172 87358 24212
rect 87398 24172 87440 24212
rect 87112 24163 87480 24172
rect 86668 23911 86708 23920
rect 86476 23827 86516 23836
rect 87724 23876 87764 23885
rect 87820 23876 87860 24499
rect 87916 23960 87956 23969
rect 88012 23960 88052 25432
rect 88203 25304 88245 25313
rect 88203 25264 88204 25304
rect 88244 25264 88245 25304
rect 88203 25255 88245 25264
rect 88204 25170 88244 25255
rect 88300 24800 88340 26356
rect 88396 25556 88436 26356
rect 88396 25507 88436 25516
rect 88491 25304 88533 25313
rect 88491 25264 88492 25304
rect 88532 25264 88533 25304
rect 88491 25255 88533 25264
rect 88492 25170 88532 25255
rect 88588 24800 88628 26440
rect 88815 26396 88855 26796
rect 89105 26480 89145 26796
rect 88780 26356 88855 26396
rect 88972 26440 89145 26480
rect 88780 25556 88820 26356
rect 88780 25507 88820 25516
rect 88875 25388 88917 25397
rect 88875 25348 88876 25388
rect 88916 25348 88917 25388
rect 88875 25339 88917 25348
rect 88683 25304 88725 25313
rect 88683 25264 88684 25304
rect 88724 25264 88820 25304
rect 88683 25255 88725 25264
rect 88684 25170 88724 25255
rect 88684 24800 88724 24809
rect 88588 24760 88684 24800
rect 88300 24751 88340 24760
rect 88684 24751 88724 24760
rect 88107 24548 88149 24557
rect 88107 24508 88108 24548
rect 88148 24508 88149 24548
rect 88107 24499 88149 24508
rect 88491 24548 88533 24557
rect 88491 24508 88492 24548
rect 88532 24508 88533 24548
rect 88491 24499 88533 24508
rect 88108 24414 88148 24499
rect 88492 24414 88532 24499
rect 87956 23920 88052 23960
rect 87916 23911 87956 23920
rect 87764 23836 87860 23876
rect 88780 23876 88820 25264
rect 88876 24548 88916 25339
rect 88876 24499 88916 24508
rect 88972 23960 89012 26440
rect 89215 26396 89255 26796
rect 89505 26396 89545 26796
rect 89164 26356 89255 26396
rect 89452 26356 89545 26396
rect 89615 26396 89655 26796
rect 89905 26396 89945 26796
rect 89615 26356 89684 26396
rect 89164 25556 89204 26356
rect 89164 25507 89204 25516
rect 89068 25304 89108 25313
rect 89068 24557 89108 25264
rect 89452 24800 89492 26356
rect 89644 25565 89684 26356
rect 89836 26356 89945 26396
rect 90015 26396 90055 26796
rect 90305 26396 90345 26796
rect 90415 26396 90455 26796
rect 90705 26396 90745 26796
rect 90815 26396 90855 26796
rect 91105 26480 91145 26796
rect 90015 26356 90260 26396
rect 90305 26356 90356 26396
rect 90415 26356 90548 26396
rect 89643 25556 89685 25565
rect 89643 25516 89644 25556
rect 89684 25516 89685 25556
rect 89643 25507 89685 25516
rect 89740 25472 89780 25481
rect 89547 25388 89589 25397
rect 89547 25348 89548 25388
rect 89588 25348 89589 25388
rect 89547 25339 89589 25348
rect 89548 25254 89588 25339
rect 89740 25313 89780 25432
rect 89739 25304 89781 25313
rect 89739 25264 89740 25304
rect 89780 25264 89781 25304
rect 89739 25255 89781 25264
rect 89836 24800 89876 26356
rect 89931 25556 89973 25565
rect 89931 25516 89932 25556
rect 89972 25516 89973 25556
rect 89931 25507 89973 25516
rect 90220 25556 90260 26356
rect 90316 25556 90356 26356
rect 90508 25556 90548 26356
rect 90316 25516 90452 25556
rect 90220 25507 90260 25516
rect 89932 25422 89972 25507
rect 90027 25304 90069 25313
rect 90027 25264 90028 25304
rect 90068 25264 90069 25304
rect 90027 25255 90069 25264
rect 90315 25304 90357 25313
rect 90315 25264 90316 25304
rect 90356 25264 90357 25304
rect 90315 25255 90357 25264
rect 90028 25170 90068 25255
rect 90316 25170 90356 25255
rect 89932 24800 89972 24809
rect 89836 24760 89932 24800
rect 89452 24751 89492 24760
rect 89932 24751 89972 24760
rect 90316 24800 90356 24809
rect 90412 24800 90452 25516
rect 90508 25507 90548 25516
rect 90604 26356 90745 26396
rect 90796 26356 90855 26396
rect 91084 26440 91145 26480
rect 90604 25472 90644 26356
rect 90796 25556 90836 26356
rect 90796 25507 90836 25516
rect 90604 25432 90740 25472
rect 90603 25304 90645 25313
rect 90603 25264 90604 25304
rect 90644 25264 90645 25304
rect 90603 25255 90645 25264
rect 90604 25170 90644 25255
rect 90356 24760 90452 24800
rect 90700 24800 90740 25432
rect 90891 25304 90933 25313
rect 90891 25264 90892 25304
rect 90932 25264 90933 25304
rect 90891 25255 90933 25264
rect 90892 25170 90932 25255
rect 91084 24800 91124 26440
rect 91215 26396 91255 26796
rect 91505 26480 91545 26796
rect 91180 26356 91255 26396
rect 91468 26440 91545 26480
rect 91180 25556 91220 26356
rect 91180 25507 91220 25516
rect 91468 25388 91508 26440
rect 91615 26396 91655 26796
rect 91905 26396 91945 26796
rect 91564 26356 91655 26396
rect 91852 26356 91945 26396
rect 92015 26396 92055 26796
rect 92305 26396 92345 26796
rect 92015 26356 92084 26396
rect 91564 25556 91604 26356
rect 91564 25507 91604 25516
rect 91468 25348 91604 25388
rect 91275 25304 91317 25313
rect 91275 25264 91276 25304
rect 91316 25293 91495 25304
rect 91316 25264 91455 25293
rect 91275 25255 91317 25264
rect 91276 25170 91316 25255
rect 91455 25244 91495 25253
rect 91180 24800 91220 24809
rect 91084 24760 91180 24800
rect 90316 24751 90356 24760
rect 90700 24751 90740 24760
rect 91180 24751 91220 24760
rect 89067 24548 89109 24557
rect 89067 24508 89068 24548
rect 89108 24508 89109 24548
rect 89067 24499 89109 24508
rect 89259 24548 89301 24557
rect 89259 24508 89260 24548
rect 89300 24508 89301 24548
rect 89259 24499 89301 24508
rect 89739 24548 89781 24557
rect 89739 24508 89740 24548
rect 89780 24508 89781 24548
rect 89739 24499 89781 24508
rect 90123 24548 90165 24557
rect 90123 24508 90124 24548
rect 90164 24508 90165 24548
rect 90123 24499 90165 24508
rect 90507 24548 90549 24557
rect 90507 24508 90508 24548
rect 90548 24508 90549 24548
rect 90507 24499 90549 24508
rect 90987 24548 91029 24557
rect 90987 24508 90988 24548
rect 91028 24508 91029 24548
rect 90987 24499 91029 24508
rect 89068 24464 89108 24499
rect 89068 24413 89108 24424
rect 89260 24414 89300 24499
rect 89740 24414 89780 24499
rect 90124 24414 90164 24499
rect 90508 24414 90548 24499
rect 89068 23960 89108 23969
rect 88972 23920 89068 23960
rect 90988 23960 91028 24499
rect 91112 24212 91480 24221
rect 91152 24172 91194 24212
rect 91234 24172 91276 24212
rect 91316 24172 91358 24212
rect 91398 24172 91440 24212
rect 91112 24163 91480 24172
rect 91468 23960 91508 23969
rect 91564 23960 91604 25348
rect 91852 24800 91892 26356
rect 92044 25556 92084 26356
rect 92044 25507 92084 25516
rect 92140 26356 92345 26396
rect 92415 26396 92455 26796
rect 92705 26396 92745 26796
rect 92815 26396 92855 26796
rect 93105 26396 93145 26796
rect 93215 26396 93255 26796
rect 93505 26480 93545 26796
rect 92415 26356 92468 26396
rect 92705 26356 92756 26396
rect 91947 25304 91989 25313
rect 91947 25264 91948 25304
rect 91988 25264 91989 25304
rect 91947 25255 91989 25264
rect 91948 25170 91988 25255
rect 91852 24751 91892 24760
rect 92140 24800 92180 26356
rect 92331 25388 92373 25397
rect 92331 25348 92332 25388
rect 92372 25348 92373 25388
rect 92331 25339 92373 25348
rect 92332 25304 92372 25339
rect 92332 25253 92372 25264
rect 92140 24751 92180 24760
rect 91659 24548 91701 24557
rect 91659 24508 91660 24548
rect 91700 24508 91701 24548
rect 91659 24499 91701 24508
rect 92331 24548 92373 24557
rect 92331 24508 92332 24548
rect 92372 24508 92373 24548
rect 92331 24499 92373 24508
rect 91660 24414 91700 24499
rect 90988 23920 91316 23960
rect 89068 23911 89108 23920
rect 88876 23876 88916 23885
rect 88780 23836 88876 23876
rect 87724 23827 87764 23836
rect 88876 23827 88916 23836
rect 91276 23876 91316 23920
rect 91508 23920 91604 23960
rect 91468 23911 91508 23920
rect 91276 23827 91316 23836
rect 80332 23742 80372 23827
rect 81676 23742 81716 23827
rect 82444 23742 82484 23827
rect 84940 23742 84980 23827
rect 85708 23742 85748 23827
rect 92332 23792 92372 24499
rect 92428 23960 92468 26356
rect 92523 25304 92565 25313
rect 92523 25264 92524 25304
rect 92564 25264 92660 25304
rect 92523 25255 92565 25264
rect 92524 25170 92564 25255
rect 92523 24548 92565 24557
rect 92523 24508 92524 24548
rect 92564 24508 92565 24548
rect 92620 24548 92660 25264
rect 92716 24800 92756 26356
rect 92812 26356 92855 26396
rect 93100 26356 93145 26396
rect 93196 26356 93255 26396
rect 93484 26440 93545 26480
rect 92812 25556 92852 26356
rect 92812 25507 92852 25516
rect 93100 25388 93140 26356
rect 93196 25556 93236 26356
rect 93196 25507 93236 25516
rect 93484 25388 93524 26440
rect 93615 26396 93655 26796
rect 93905 26396 93945 26796
rect 93580 26356 93655 26396
rect 93868 26356 93945 26396
rect 94015 26396 94055 26796
rect 94305 26480 94345 26796
rect 94252 26440 94345 26480
rect 94015 26356 94100 26396
rect 93580 25556 93620 26356
rect 93580 25507 93620 25516
rect 93100 25348 93236 25388
rect 93484 25348 93620 25388
rect 92907 25304 92949 25313
rect 92907 25264 92908 25304
rect 92948 25293 93127 25304
rect 92948 25264 93087 25293
rect 92907 25255 92949 25264
rect 92908 25170 92948 25255
rect 93087 25244 93127 25253
rect 92908 24800 92948 24809
rect 92716 24760 92908 24800
rect 93196 24800 93236 25348
rect 93292 24800 93332 24809
rect 93196 24760 93292 24800
rect 92908 24751 92948 24760
rect 93292 24751 93332 24760
rect 92716 24548 92756 24557
rect 92620 24508 92716 24548
rect 92523 24499 92565 24508
rect 92716 24499 92756 24508
rect 93099 24548 93141 24557
rect 93099 24508 93100 24548
rect 93140 24508 93141 24548
rect 93099 24499 93141 24508
rect 93483 24548 93525 24557
rect 93483 24508 93484 24548
rect 93524 24508 93525 24548
rect 93483 24499 93525 24508
rect 92524 24464 92564 24499
rect 92524 24413 92564 24424
rect 93100 24414 93140 24499
rect 93484 23960 93524 24499
rect 92428 23911 92468 23920
rect 93388 23920 93524 23960
rect 93580 23960 93620 25348
rect 93675 25304 93717 25313
rect 93675 25264 93676 25304
rect 93716 25264 93717 25304
rect 93675 25255 93717 25264
rect 93676 25170 93716 25255
rect 93868 24800 93908 26356
rect 94060 25556 94100 26356
rect 94060 25507 94100 25516
rect 94252 25388 94292 26440
rect 94415 26396 94455 26796
rect 94348 26356 94455 26396
rect 94705 26396 94745 26796
rect 94815 26396 94855 26796
rect 95105 26396 95145 26796
rect 95215 26396 95255 26796
rect 94705 26356 94772 26396
rect 94815 26356 94868 26396
rect 95105 26356 95156 26396
rect 94348 25556 94388 26356
rect 94348 25507 94388 25516
rect 94252 25348 94388 25388
rect 93963 25304 94005 25313
rect 93963 25264 93964 25304
rect 94004 25264 94005 25304
rect 93963 25255 94005 25264
rect 94155 25304 94197 25313
rect 94155 25264 94156 25304
rect 94196 25293 94292 25304
rect 94196 25264 94252 25293
rect 94155 25255 94197 25264
rect 93964 25170 94004 25255
rect 94252 25244 94292 25253
rect 93964 24800 94004 24809
rect 93868 24760 93964 24800
rect 93964 24751 94004 24760
rect 94348 24800 94388 25348
rect 94348 24751 94388 24760
rect 94732 24800 94772 26356
rect 94828 25556 94868 26356
rect 94828 25507 94868 25516
rect 94923 25304 94965 25313
rect 94923 25264 94924 25304
rect 94964 25264 94965 25304
rect 94923 25255 94965 25264
rect 94732 24751 94772 24760
rect 93771 24548 93813 24557
rect 93771 24508 93772 24548
rect 93812 24508 93813 24548
rect 93771 24499 93813 24508
rect 94155 24548 94197 24557
rect 94155 24508 94156 24548
rect 94196 24508 94197 24548
rect 94155 24499 94197 24508
rect 94539 24548 94581 24557
rect 94539 24508 94540 24548
rect 94580 24508 94581 24548
rect 94539 24499 94581 24508
rect 94924 24548 94964 25255
rect 95116 24800 95156 26356
rect 95212 26356 95255 26396
rect 95505 26396 95545 26796
rect 95615 26480 95655 26796
rect 95615 26440 95732 26480
rect 95505 26356 95636 26396
rect 95212 25556 95252 26356
rect 95212 25507 95252 25516
rect 95308 25304 95348 25313
rect 95348 25264 95444 25304
rect 95308 25255 95348 25264
rect 95404 24809 95444 25264
rect 95116 24751 95156 24760
rect 95403 24800 95445 24809
rect 95403 24760 95404 24800
rect 95444 24760 95445 24800
rect 95403 24751 95445 24760
rect 95596 24800 95636 26356
rect 95692 25565 95732 26440
rect 95905 26396 95945 26796
rect 95884 26356 95945 26396
rect 96015 26396 96055 26796
rect 96305 26573 96345 26796
rect 96304 26564 96346 26573
rect 96304 26524 96305 26564
rect 96345 26524 96346 26564
rect 96415 26564 96455 26796
rect 96555 26564 96597 26573
rect 96415 26524 96500 26564
rect 96304 26515 96346 26524
rect 96015 26356 96404 26396
rect 95691 25556 95733 25565
rect 95691 25516 95692 25556
rect 95732 25516 95733 25556
rect 95691 25507 95733 25516
rect 95691 25388 95733 25397
rect 95691 25348 95692 25388
rect 95732 25348 95828 25388
rect 95691 25339 95733 25348
rect 95692 25254 95732 25339
rect 95596 24751 95636 24760
rect 94924 24499 94964 24508
rect 95404 24548 95444 24751
rect 95404 24499 95444 24508
rect 95788 24548 95828 25348
rect 95884 25293 95924 26356
rect 96075 25556 96117 25565
rect 96075 25516 96076 25556
rect 96116 25516 96117 25556
rect 96075 25507 96117 25516
rect 96364 25556 96404 26356
rect 96460 25565 96500 26524
rect 96555 26524 96556 26564
rect 96596 26524 96597 26564
rect 96555 26515 96597 26524
rect 96364 25507 96404 25516
rect 96459 25556 96501 25565
rect 96459 25516 96460 25556
rect 96500 25516 96501 25556
rect 96459 25507 96501 25516
rect 96076 25422 96116 25507
rect 96172 25304 96212 25315
rect 95884 25253 96020 25293
rect 95883 25136 95925 25145
rect 95883 25096 95884 25136
rect 95924 25096 95925 25136
rect 95883 25087 95925 25096
rect 95884 25002 95924 25087
rect 95980 24968 96020 25253
rect 96172 25229 96212 25264
rect 96460 25304 96500 25315
rect 96460 25229 96500 25264
rect 96171 25220 96213 25229
rect 96171 25180 96172 25220
rect 96212 25180 96213 25220
rect 96171 25171 96213 25180
rect 96459 25220 96501 25229
rect 96459 25180 96460 25220
rect 96500 25180 96501 25220
rect 96459 25171 96501 25180
rect 95980 24928 96212 24968
rect 95979 24800 96021 24809
rect 95979 24760 95980 24800
rect 96020 24760 96021 24800
rect 95979 24751 96021 24760
rect 96172 24800 96212 24928
rect 96172 24751 96212 24760
rect 96363 24800 96405 24809
rect 96363 24760 96364 24800
rect 96404 24760 96405 24800
rect 96363 24751 96405 24760
rect 96556 24800 96596 26515
rect 96705 26396 96745 26796
rect 96652 26356 96745 26396
rect 96815 26396 96855 26796
rect 97105 26396 97145 26796
rect 97215 26396 97255 26796
rect 97505 26396 97545 26796
rect 97615 26396 97655 26796
rect 97905 26396 97945 26796
rect 96815 26356 96884 26396
rect 97105 26356 97172 26396
rect 97215 26356 97268 26396
rect 97505 26356 97556 26396
rect 97615 26356 97748 26396
rect 96652 25136 96692 26356
rect 96844 25556 96884 26356
rect 96844 25507 96884 25516
rect 96748 25313 96788 25398
rect 97132 25388 97172 26356
rect 97228 25556 97268 26356
rect 97228 25507 97268 25516
rect 97419 25556 97461 25565
rect 97419 25516 97420 25556
rect 97460 25516 97461 25556
rect 97516 25556 97556 26356
rect 97708 25556 97748 26356
rect 97516 25516 97652 25556
rect 97419 25507 97461 25516
rect 97420 25422 97460 25507
rect 97132 25348 97364 25388
rect 96747 25304 96789 25313
rect 96747 25264 96748 25304
rect 96788 25264 96789 25304
rect 96747 25255 96789 25264
rect 97035 25304 97077 25313
rect 97035 25264 97036 25304
rect 97076 25293 97077 25304
rect 97127 25293 97167 25302
rect 97076 25264 97127 25293
rect 97035 25255 97127 25264
rect 97036 25253 97127 25255
rect 97127 25244 97167 25253
rect 96652 25096 96980 25136
rect 96556 24751 96596 24760
rect 96747 24800 96789 24809
rect 96747 24760 96748 24800
rect 96788 24760 96789 24800
rect 96747 24751 96789 24760
rect 96940 24800 96980 25096
rect 96940 24751 96980 24760
rect 97131 24800 97173 24809
rect 97131 24760 97132 24800
rect 97172 24760 97173 24800
rect 97131 24751 97173 24760
rect 97324 24800 97364 25348
rect 97515 25304 97557 25313
rect 97515 25264 97516 25304
rect 97556 25264 97557 25304
rect 97515 25255 97557 25264
rect 97516 25170 97556 25255
rect 97324 24751 97364 24760
rect 97515 24800 97557 24809
rect 97515 24760 97516 24800
rect 97556 24760 97557 24800
rect 97612 24800 97652 25516
rect 97708 25507 97748 25516
rect 97900 26356 97945 26396
rect 98015 26396 98055 26796
rect 98305 26396 98345 26796
rect 98415 26480 98455 26796
rect 98415 26440 98804 26480
rect 98015 26356 98132 26396
rect 98305 26356 98420 26396
rect 97803 25304 97845 25313
rect 97803 25264 97804 25304
rect 97844 25264 97845 25304
rect 97803 25255 97845 25264
rect 97804 25170 97844 25255
rect 97708 24800 97748 24809
rect 97612 24760 97708 24800
rect 97900 24800 97940 26356
rect 98092 25556 98132 26356
rect 98092 25507 98132 25516
rect 98380 25556 98420 26356
rect 98380 25507 98420 25516
rect 98764 25556 98804 26440
rect 98860 26153 98900 32824
rect 99147 32864 99189 32873
rect 99147 32824 99148 32864
rect 99188 32824 99189 32864
rect 99147 32815 99189 32824
rect 99148 32730 99188 32815
rect 98956 32696 98996 32705
rect 98956 32201 98996 32656
rect 99244 32696 99284 32705
rect 98955 32192 98997 32201
rect 98955 32152 98956 32192
rect 98996 32152 98997 32192
rect 98955 32143 98997 32152
rect 99244 32117 99284 32656
rect 99243 32108 99285 32117
rect 99243 32068 99244 32108
rect 99284 32068 99285 32108
rect 99243 32059 99285 32068
rect 98859 26144 98901 26153
rect 98859 26104 98860 26144
rect 98900 26104 98901 26144
rect 98859 26095 98901 26104
rect 98764 25507 98804 25516
rect 98572 25388 98612 25397
rect 98860 25388 98900 26095
rect 98612 25348 98900 25388
rect 98572 25339 98612 25348
rect 97995 25304 98037 25313
rect 97995 25264 97996 25304
rect 98036 25264 98037 25304
rect 97995 25255 98037 25264
rect 98860 25304 98900 25348
rect 98860 25255 98900 25264
rect 97996 25170 98036 25255
rect 98092 24800 98132 24809
rect 97900 24760 98092 24800
rect 97515 24751 97557 24760
rect 97708 24751 97748 24760
rect 98092 24751 98132 24760
rect 95980 24666 96020 24751
rect 95788 24499 95828 24508
rect 96364 24548 96404 24751
rect 96364 24499 96404 24508
rect 96748 24548 96788 24751
rect 96748 24499 96788 24508
rect 97132 24548 97172 24751
rect 97516 24557 97556 24751
rect 97132 24499 97172 24508
rect 97515 24548 97557 24557
rect 97515 24508 97516 24548
rect 97556 24508 97557 24548
rect 97515 24499 97557 24508
rect 97899 24548 97941 24557
rect 97899 24508 97900 24548
rect 97940 24508 97941 24548
rect 97899 24499 97941 24508
rect 98283 24548 98325 24557
rect 98283 24508 98284 24548
rect 98324 24508 98325 24548
rect 98283 24499 98325 24508
rect 93772 24414 93812 24499
rect 94156 24414 94196 24499
rect 94540 24414 94580 24499
rect 97516 24414 97556 24499
rect 97900 24414 97940 24499
rect 98284 24414 98324 24499
rect 95112 24212 95480 24221
rect 95152 24172 95194 24212
rect 95234 24172 95276 24212
rect 95316 24172 95358 24212
rect 95398 24172 95440 24212
rect 95112 24163 95480 24172
rect 99112 24212 99480 24221
rect 99152 24172 99194 24212
rect 99234 24172 99276 24212
rect 99316 24172 99358 24212
rect 99398 24172 99440 24212
rect 99112 24163 99480 24172
rect 93388 23876 93428 23920
rect 93580 23911 93620 23920
rect 93388 23827 93428 23836
rect 92332 23743 92372 23752
rect 72352 23456 72720 23465
rect 72392 23416 72434 23456
rect 72474 23416 72516 23456
rect 72556 23416 72598 23456
rect 72638 23416 72680 23456
rect 72352 23407 72720 23416
rect 76352 23456 76720 23465
rect 76392 23416 76434 23456
rect 76474 23416 76516 23456
rect 76556 23416 76598 23456
rect 76638 23416 76680 23456
rect 76352 23407 76720 23416
rect 80352 23456 80720 23465
rect 80392 23416 80434 23456
rect 80474 23416 80516 23456
rect 80556 23416 80598 23456
rect 80638 23416 80680 23456
rect 80352 23407 80720 23416
rect 84352 23456 84720 23465
rect 84392 23416 84434 23456
rect 84474 23416 84516 23456
rect 84556 23416 84598 23456
rect 84638 23416 84680 23456
rect 84352 23407 84720 23416
rect 88352 23456 88720 23465
rect 88392 23416 88434 23456
rect 88474 23416 88516 23456
rect 88556 23416 88598 23456
rect 88638 23416 88680 23456
rect 88352 23407 88720 23416
rect 92352 23456 92720 23465
rect 92392 23416 92434 23456
rect 92474 23416 92516 23456
rect 92556 23416 92598 23456
rect 92638 23416 92680 23456
rect 92352 23407 92720 23416
rect 96352 23456 96720 23465
rect 96392 23416 96434 23456
rect 96474 23416 96516 23456
rect 96556 23416 96598 23456
rect 96638 23416 96680 23456
rect 96352 23407 96720 23416
rect 71112 22700 71480 22709
rect 71152 22660 71194 22700
rect 71234 22660 71276 22700
rect 71316 22660 71358 22700
rect 71398 22660 71440 22700
rect 71112 22651 71480 22660
rect 75112 22700 75480 22709
rect 75152 22660 75194 22700
rect 75234 22660 75276 22700
rect 75316 22660 75358 22700
rect 75398 22660 75440 22700
rect 75112 22651 75480 22660
rect 79112 22700 79480 22709
rect 79152 22660 79194 22700
rect 79234 22660 79276 22700
rect 79316 22660 79358 22700
rect 79398 22660 79440 22700
rect 79112 22651 79480 22660
rect 83112 22700 83480 22709
rect 83152 22660 83194 22700
rect 83234 22660 83276 22700
rect 83316 22660 83358 22700
rect 83398 22660 83440 22700
rect 83112 22651 83480 22660
rect 87112 22700 87480 22709
rect 87152 22660 87194 22700
rect 87234 22660 87276 22700
rect 87316 22660 87358 22700
rect 87398 22660 87440 22700
rect 87112 22651 87480 22660
rect 91112 22700 91480 22709
rect 91152 22660 91194 22700
rect 91234 22660 91276 22700
rect 91316 22660 91358 22700
rect 91398 22660 91440 22700
rect 91112 22651 91480 22660
rect 95112 22700 95480 22709
rect 95152 22660 95194 22700
rect 95234 22660 95276 22700
rect 95316 22660 95358 22700
rect 95398 22660 95440 22700
rect 95112 22651 95480 22660
rect 99112 22700 99480 22709
rect 99152 22660 99194 22700
rect 99234 22660 99276 22700
rect 99316 22660 99358 22700
rect 99398 22660 99440 22700
rect 99112 22651 99480 22660
rect 72352 21944 72720 21953
rect 72392 21904 72434 21944
rect 72474 21904 72516 21944
rect 72556 21904 72598 21944
rect 72638 21904 72680 21944
rect 72352 21895 72720 21904
rect 76352 21944 76720 21953
rect 76392 21904 76434 21944
rect 76474 21904 76516 21944
rect 76556 21904 76598 21944
rect 76638 21904 76680 21944
rect 76352 21895 76720 21904
rect 80352 21944 80720 21953
rect 80392 21904 80434 21944
rect 80474 21904 80516 21944
rect 80556 21904 80598 21944
rect 80638 21904 80680 21944
rect 80352 21895 80720 21904
rect 84352 21944 84720 21953
rect 84392 21904 84434 21944
rect 84474 21904 84516 21944
rect 84556 21904 84598 21944
rect 84638 21904 84680 21944
rect 84352 21895 84720 21904
rect 88352 21944 88720 21953
rect 88392 21904 88434 21944
rect 88474 21904 88516 21944
rect 88556 21904 88598 21944
rect 88638 21904 88680 21944
rect 88352 21895 88720 21904
rect 92352 21944 92720 21953
rect 92392 21904 92434 21944
rect 92474 21904 92516 21944
rect 92556 21904 92598 21944
rect 92638 21904 92680 21944
rect 92352 21895 92720 21904
rect 96352 21944 96720 21953
rect 96392 21904 96434 21944
rect 96474 21904 96516 21944
rect 96556 21904 96598 21944
rect 96638 21904 96680 21944
rect 96352 21895 96720 21904
rect 71112 21188 71480 21197
rect 71152 21148 71194 21188
rect 71234 21148 71276 21188
rect 71316 21148 71358 21188
rect 71398 21148 71440 21188
rect 71112 21139 71480 21148
rect 75112 21188 75480 21197
rect 75152 21148 75194 21188
rect 75234 21148 75276 21188
rect 75316 21148 75358 21188
rect 75398 21148 75440 21188
rect 75112 21139 75480 21148
rect 79112 21188 79480 21197
rect 79152 21148 79194 21188
rect 79234 21148 79276 21188
rect 79316 21148 79358 21188
rect 79398 21148 79440 21188
rect 79112 21139 79480 21148
rect 83112 21188 83480 21197
rect 83152 21148 83194 21188
rect 83234 21148 83276 21188
rect 83316 21148 83358 21188
rect 83398 21148 83440 21188
rect 83112 21139 83480 21148
rect 87112 21188 87480 21197
rect 87152 21148 87194 21188
rect 87234 21148 87276 21188
rect 87316 21148 87358 21188
rect 87398 21148 87440 21188
rect 87112 21139 87480 21148
rect 91112 21188 91480 21197
rect 91152 21148 91194 21188
rect 91234 21148 91276 21188
rect 91316 21148 91358 21188
rect 91398 21148 91440 21188
rect 91112 21139 91480 21148
rect 95112 21188 95480 21197
rect 95152 21148 95194 21188
rect 95234 21148 95276 21188
rect 95316 21148 95358 21188
rect 95398 21148 95440 21188
rect 95112 21139 95480 21148
rect 99112 21188 99480 21197
rect 99152 21148 99194 21188
rect 99234 21148 99276 21188
rect 99316 21148 99358 21188
rect 99398 21148 99440 21188
rect 99112 21139 99480 21148
rect 72352 20432 72720 20441
rect 72392 20392 72434 20432
rect 72474 20392 72516 20432
rect 72556 20392 72598 20432
rect 72638 20392 72680 20432
rect 72352 20383 72720 20392
rect 76352 20432 76720 20441
rect 76392 20392 76434 20432
rect 76474 20392 76516 20432
rect 76556 20392 76598 20432
rect 76638 20392 76680 20432
rect 76352 20383 76720 20392
rect 80352 20432 80720 20441
rect 80392 20392 80434 20432
rect 80474 20392 80516 20432
rect 80556 20392 80598 20432
rect 80638 20392 80680 20432
rect 80352 20383 80720 20392
rect 84352 20432 84720 20441
rect 84392 20392 84434 20432
rect 84474 20392 84516 20432
rect 84556 20392 84598 20432
rect 84638 20392 84680 20432
rect 84352 20383 84720 20392
rect 88352 20432 88720 20441
rect 88392 20392 88434 20432
rect 88474 20392 88516 20432
rect 88556 20392 88598 20432
rect 88638 20392 88680 20432
rect 88352 20383 88720 20392
rect 92352 20432 92720 20441
rect 92392 20392 92434 20432
rect 92474 20392 92516 20432
rect 92556 20392 92598 20432
rect 92638 20392 92680 20432
rect 92352 20383 92720 20392
rect 96352 20432 96720 20441
rect 96392 20392 96434 20432
rect 96474 20392 96516 20432
rect 96556 20392 96598 20432
rect 96638 20392 96680 20432
rect 96352 20383 96720 20392
rect 71112 19676 71480 19685
rect 71152 19636 71194 19676
rect 71234 19636 71276 19676
rect 71316 19636 71358 19676
rect 71398 19636 71440 19676
rect 71112 19627 71480 19636
rect 75112 19676 75480 19685
rect 75152 19636 75194 19676
rect 75234 19636 75276 19676
rect 75316 19636 75358 19676
rect 75398 19636 75440 19676
rect 75112 19627 75480 19636
rect 79112 19676 79480 19685
rect 79152 19636 79194 19676
rect 79234 19636 79276 19676
rect 79316 19636 79358 19676
rect 79398 19636 79440 19676
rect 79112 19627 79480 19636
rect 83112 19676 83480 19685
rect 83152 19636 83194 19676
rect 83234 19636 83276 19676
rect 83316 19636 83358 19676
rect 83398 19636 83440 19676
rect 83112 19627 83480 19636
rect 87112 19676 87480 19685
rect 87152 19636 87194 19676
rect 87234 19636 87276 19676
rect 87316 19636 87358 19676
rect 87398 19636 87440 19676
rect 87112 19627 87480 19636
rect 91112 19676 91480 19685
rect 91152 19636 91194 19676
rect 91234 19636 91276 19676
rect 91316 19636 91358 19676
rect 91398 19636 91440 19676
rect 91112 19627 91480 19636
rect 95112 19676 95480 19685
rect 95152 19636 95194 19676
rect 95234 19636 95276 19676
rect 95316 19636 95358 19676
rect 95398 19636 95440 19676
rect 95112 19627 95480 19636
rect 99112 19676 99480 19685
rect 99152 19636 99194 19676
rect 99234 19636 99276 19676
rect 99316 19636 99358 19676
rect 99398 19636 99440 19676
rect 99112 19627 99480 19636
rect 72352 18920 72720 18929
rect 72392 18880 72434 18920
rect 72474 18880 72516 18920
rect 72556 18880 72598 18920
rect 72638 18880 72680 18920
rect 72352 18871 72720 18880
rect 76352 18920 76720 18929
rect 76392 18880 76434 18920
rect 76474 18880 76516 18920
rect 76556 18880 76598 18920
rect 76638 18880 76680 18920
rect 76352 18871 76720 18880
rect 80352 18920 80720 18929
rect 80392 18880 80434 18920
rect 80474 18880 80516 18920
rect 80556 18880 80598 18920
rect 80638 18880 80680 18920
rect 80352 18871 80720 18880
rect 84352 18920 84720 18929
rect 84392 18880 84434 18920
rect 84474 18880 84516 18920
rect 84556 18880 84598 18920
rect 84638 18880 84680 18920
rect 84352 18871 84720 18880
rect 88352 18920 88720 18929
rect 88392 18880 88434 18920
rect 88474 18880 88516 18920
rect 88556 18880 88598 18920
rect 88638 18880 88680 18920
rect 88352 18871 88720 18880
rect 92352 18920 92720 18929
rect 92392 18880 92434 18920
rect 92474 18880 92516 18920
rect 92556 18880 92598 18920
rect 92638 18880 92680 18920
rect 92352 18871 92720 18880
rect 96352 18920 96720 18929
rect 96392 18880 96434 18920
rect 96474 18880 96516 18920
rect 96556 18880 96598 18920
rect 96638 18880 96680 18920
rect 96352 18871 96720 18880
rect 71112 18164 71480 18173
rect 71152 18124 71194 18164
rect 71234 18124 71276 18164
rect 71316 18124 71358 18164
rect 71398 18124 71440 18164
rect 71112 18115 71480 18124
rect 75112 18164 75480 18173
rect 75152 18124 75194 18164
rect 75234 18124 75276 18164
rect 75316 18124 75358 18164
rect 75398 18124 75440 18164
rect 75112 18115 75480 18124
rect 79112 18164 79480 18173
rect 79152 18124 79194 18164
rect 79234 18124 79276 18164
rect 79316 18124 79358 18164
rect 79398 18124 79440 18164
rect 79112 18115 79480 18124
rect 83112 18164 83480 18173
rect 83152 18124 83194 18164
rect 83234 18124 83276 18164
rect 83316 18124 83358 18164
rect 83398 18124 83440 18164
rect 83112 18115 83480 18124
rect 87112 18164 87480 18173
rect 87152 18124 87194 18164
rect 87234 18124 87276 18164
rect 87316 18124 87358 18164
rect 87398 18124 87440 18164
rect 87112 18115 87480 18124
rect 91112 18164 91480 18173
rect 91152 18124 91194 18164
rect 91234 18124 91276 18164
rect 91316 18124 91358 18164
rect 91398 18124 91440 18164
rect 91112 18115 91480 18124
rect 95112 18164 95480 18173
rect 95152 18124 95194 18164
rect 95234 18124 95276 18164
rect 95316 18124 95358 18164
rect 95398 18124 95440 18164
rect 95112 18115 95480 18124
rect 99112 18164 99480 18173
rect 99152 18124 99194 18164
rect 99234 18124 99276 18164
rect 99316 18124 99358 18164
rect 99398 18124 99440 18164
rect 99112 18115 99480 18124
rect 72352 17408 72720 17417
rect 72392 17368 72434 17408
rect 72474 17368 72516 17408
rect 72556 17368 72598 17408
rect 72638 17368 72680 17408
rect 72352 17359 72720 17368
rect 76352 17408 76720 17417
rect 76392 17368 76434 17408
rect 76474 17368 76516 17408
rect 76556 17368 76598 17408
rect 76638 17368 76680 17408
rect 76352 17359 76720 17368
rect 80352 17408 80720 17417
rect 80392 17368 80434 17408
rect 80474 17368 80516 17408
rect 80556 17368 80598 17408
rect 80638 17368 80680 17408
rect 80352 17359 80720 17368
rect 84352 17408 84720 17417
rect 84392 17368 84434 17408
rect 84474 17368 84516 17408
rect 84556 17368 84598 17408
rect 84638 17368 84680 17408
rect 84352 17359 84720 17368
rect 88352 17408 88720 17417
rect 88392 17368 88434 17408
rect 88474 17368 88516 17408
rect 88556 17368 88598 17408
rect 88638 17368 88680 17408
rect 88352 17359 88720 17368
rect 92352 17408 92720 17417
rect 92392 17368 92434 17408
rect 92474 17368 92516 17408
rect 92556 17368 92598 17408
rect 92638 17368 92680 17408
rect 92352 17359 92720 17368
rect 96352 17408 96720 17417
rect 96392 17368 96434 17408
rect 96474 17368 96516 17408
rect 96556 17368 96598 17408
rect 96638 17368 96680 17408
rect 96352 17359 96720 17368
rect 86572 17072 86612 17081
rect 86476 17032 86572 17072
rect 80428 16988 80468 16997
rect 71112 16652 71480 16661
rect 71152 16612 71194 16652
rect 71234 16612 71276 16652
rect 71316 16612 71358 16652
rect 71398 16612 71440 16652
rect 71112 16603 71480 16612
rect 75112 16652 75480 16661
rect 75152 16612 75194 16652
rect 75234 16612 75276 16652
rect 75316 16612 75358 16652
rect 75398 16612 75440 16652
rect 75112 16603 75480 16612
rect 79112 16652 79480 16661
rect 79152 16612 79194 16652
rect 79234 16612 79276 16652
rect 79316 16612 79358 16652
rect 79398 16612 79440 16652
rect 79112 16603 79480 16612
rect 71787 16400 71829 16409
rect 71787 16360 71788 16400
rect 71828 16360 71829 16400
rect 71787 16351 71829 16360
rect 74476 16400 74516 16411
rect 71020 15100 71156 15140
rect 67112 15091 67480 15100
rect 70635 14804 70677 14813
rect 70635 14764 70636 14804
rect 70676 14764 70677 14804
rect 70635 14755 70677 14764
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 8352 14384 8720 14393
rect 8392 14344 8434 14384
rect 8474 14344 8516 14384
rect 8556 14344 8598 14384
rect 8638 14344 8680 14384
rect 8352 14335 8720 14344
rect 12352 14384 12720 14393
rect 12392 14344 12434 14384
rect 12474 14344 12516 14384
rect 12556 14344 12598 14384
rect 12638 14344 12680 14384
rect 12352 14335 12720 14344
rect 16352 14384 16720 14393
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16352 14335 16720 14344
rect 20352 14384 20720 14393
rect 20392 14344 20434 14384
rect 20474 14344 20516 14384
rect 20556 14344 20598 14384
rect 20638 14344 20680 14384
rect 20352 14335 20720 14344
rect 24352 14384 24720 14393
rect 24392 14344 24434 14384
rect 24474 14344 24516 14384
rect 24556 14344 24598 14384
rect 24638 14344 24680 14384
rect 24352 14335 24720 14344
rect 28352 14384 28720 14393
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28352 14335 28720 14344
rect 32352 14384 32720 14393
rect 32392 14344 32434 14384
rect 32474 14344 32516 14384
rect 32556 14344 32598 14384
rect 32638 14344 32680 14384
rect 32352 14335 32720 14344
rect 36352 14384 36720 14393
rect 36392 14344 36434 14384
rect 36474 14344 36516 14384
rect 36556 14344 36598 14384
rect 36638 14344 36680 14384
rect 36352 14335 36720 14344
rect 40352 14384 40720 14393
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40352 14335 40720 14344
rect 44352 14384 44720 14393
rect 44392 14344 44434 14384
rect 44474 14344 44516 14384
rect 44556 14344 44598 14384
rect 44638 14344 44680 14384
rect 44352 14335 44720 14344
rect 48352 14384 48720 14393
rect 48392 14344 48434 14384
rect 48474 14344 48516 14384
rect 48556 14344 48598 14384
rect 48638 14344 48680 14384
rect 48352 14335 48720 14344
rect 52352 14384 52720 14393
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52352 14335 52720 14344
rect 56352 14384 56720 14393
rect 56392 14344 56434 14384
rect 56474 14344 56516 14384
rect 56556 14344 56598 14384
rect 56638 14344 56680 14384
rect 56352 14335 56720 14344
rect 60352 14384 60720 14393
rect 60392 14344 60434 14384
rect 60474 14344 60516 14384
rect 60556 14344 60598 14384
rect 60638 14344 60680 14384
rect 60352 14335 60720 14344
rect 64352 14384 64720 14393
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64352 14335 64720 14344
rect 68352 14384 68720 14393
rect 68392 14344 68434 14384
rect 68474 14344 68516 14384
rect 68556 14344 68598 14384
rect 68638 14344 68680 14384
rect 68352 14335 68720 14344
rect 70539 14048 70581 14057
rect 70539 14008 70540 14048
rect 70580 14008 70581 14048
rect 70539 13999 70581 14008
rect 70636 14048 70676 14755
rect 70636 13999 70676 14008
rect 70827 14048 70869 14057
rect 70827 14008 70828 14048
rect 70868 14008 70869 14048
rect 70827 13999 70869 14008
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 7112 13628 7480 13637
rect 7152 13588 7194 13628
rect 7234 13588 7276 13628
rect 7316 13588 7358 13628
rect 7398 13588 7440 13628
rect 7112 13579 7480 13588
rect 11112 13628 11480 13637
rect 11152 13588 11194 13628
rect 11234 13588 11276 13628
rect 11316 13588 11358 13628
rect 11398 13588 11440 13628
rect 11112 13579 11480 13588
rect 15112 13628 15480 13637
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15112 13579 15480 13588
rect 19112 13628 19480 13637
rect 19152 13588 19194 13628
rect 19234 13588 19276 13628
rect 19316 13588 19358 13628
rect 19398 13588 19440 13628
rect 19112 13579 19480 13588
rect 23112 13628 23480 13637
rect 23152 13588 23194 13628
rect 23234 13588 23276 13628
rect 23316 13588 23358 13628
rect 23398 13588 23440 13628
rect 23112 13579 23480 13588
rect 27112 13628 27480 13637
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27112 13579 27480 13588
rect 31112 13628 31480 13637
rect 31152 13588 31194 13628
rect 31234 13588 31276 13628
rect 31316 13588 31358 13628
rect 31398 13588 31440 13628
rect 31112 13579 31480 13588
rect 35112 13628 35480 13637
rect 35152 13588 35194 13628
rect 35234 13588 35276 13628
rect 35316 13588 35358 13628
rect 35398 13588 35440 13628
rect 35112 13579 35480 13588
rect 39112 13628 39480 13637
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39112 13579 39480 13588
rect 43112 13628 43480 13637
rect 43152 13588 43194 13628
rect 43234 13588 43276 13628
rect 43316 13588 43358 13628
rect 43398 13588 43440 13628
rect 43112 13579 43480 13588
rect 47112 13628 47480 13637
rect 47152 13588 47194 13628
rect 47234 13588 47276 13628
rect 47316 13588 47358 13628
rect 47398 13588 47440 13628
rect 47112 13579 47480 13588
rect 51112 13628 51480 13637
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51112 13579 51480 13588
rect 55112 13628 55480 13637
rect 55152 13588 55194 13628
rect 55234 13588 55276 13628
rect 55316 13588 55358 13628
rect 55398 13588 55440 13628
rect 55112 13579 55480 13588
rect 59112 13628 59480 13637
rect 59152 13588 59194 13628
rect 59234 13588 59276 13628
rect 59316 13588 59358 13628
rect 59398 13588 59440 13628
rect 59112 13579 59480 13588
rect 63112 13628 63480 13637
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63112 13579 63480 13588
rect 67112 13628 67480 13637
rect 67152 13588 67194 13628
rect 67234 13588 67276 13628
rect 67316 13588 67358 13628
rect 67398 13588 67440 13628
rect 67112 13579 67480 13588
rect 70059 13628 70101 13637
rect 70059 13588 70060 13628
rect 70100 13588 70101 13628
rect 70059 13579 70101 13588
rect 70060 13460 70100 13579
rect 70060 13411 70100 13420
rect 69868 13292 69908 13303
rect 69868 13217 69908 13252
rect 69867 13208 69909 13217
rect 69867 13168 69868 13208
rect 69908 13168 69909 13208
rect 69867 13159 69909 13168
rect 70347 13208 70389 13217
rect 70540 13208 70580 13999
rect 70731 13964 70773 13973
rect 70731 13924 70732 13964
rect 70772 13924 70773 13964
rect 70731 13915 70773 13924
rect 70635 13796 70677 13805
rect 70635 13756 70636 13796
rect 70676 13756 70677 13796
rect 70635 13747 70677 13756
rect 70347 13168 70348 13208
rect 70388 13168 70484 13208
rect 70347 13159 70389 13168
rect 70348 13074 70388 13159
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 8352 12872 8720 12881
rect 8392 12832 8434 12872
rect 8474 12832 8516 12872
rect 8556 12832 8598 12872
rect 8638 12832 8680 12872
rect 8352 12823 8720 12832
rect 12352 12872 12720 12881
rect 12392 12832 12434 12872
rect 12474 12832 12516 12872
rect 12556 12832 12598 12872
rect 12638 12832 12680 12872
rect 12352 12823 12720 12832
rect 16352 12872 16720 12881
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16352 12823 16720 12832
rect 20352 12872 20720 12881
rect 20392 12832 20434 12872
rect 20474 12832 20516 12872
rect 20556 12832 20598 12872
rect 20638 12832 20680 12872
rect 20352 12823 20720 12832
rect 24352 12872 24720 12881
rect 24392 12832 24434 12872
rect 24474 12832 24516 12872
rect 24556 12832 24598 12872
rect 24638 12832 24680 12872
rect 24352 12823 24720 12832
rect 28352 12872 28720 12881
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28352 12823 28720 12832
rect 32352 12872 32720 12881
rect 32392 12832 32434 12872
rect 32474 12832 32516 12872
rect 32556 12832 32598 12872
rect 32638 12832 32680 12872
rect 32352 12823 32720 12832
rect 36352 12872 36720 12881
rect 36392 12832 36434 12872
rect 36474 12832 36516 12872
rect 36556 12832 36598 12872
rect 36638 12832 36680 12872
rect 36352 12823 36720 12832
rect 40352 12872 40720 12881
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40352 12823 40720 12832
rect 44352 12872 44720 12881
rect 44392 12832 44434 12872
rect 44474 12832 44516 12872
rect 44556 12832 44598 12872
rect 44638 12832 44680 12872
rect 44352 12823 44720 12832
rect 48352 12872 48720 12881
rect 48392 12832 48434 12872
rect 48474 12832 48516 12872
rect 48556 12832 48598 12872
rect 48638 12832 48680 12872
rect 48352 12823 48720 12832
rect 52352 12872 52720 12881
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52352 12823 52720 12832
rect 56352 12872 56720 12881
rect 56392 12832 56434 12872
rect 56474 12832 56516 12872
rect 56556 12832 56598 12872
rect 56638 12832 56680 12872
rect 56352 12823 56720 12832
rect 60352 12872 60720 12881
rect 60392 12832 60434 12872
rect 60474 12832 60516 12872
rect 60556 12832 60598 12872
rect 60638 12832 60680 12872
rect 60352 12823 60720 12832
rect 64352 12872 64720 12881
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64352 12823 64720 12832
rect 68352 12872 68720 12881
rect 68392 12832 68434 12872
rect 68474 12832 68516 12872
rect 68556 12832 68598 12872
rect 68638 12832 68680 12872
rect 68352 12823 68720 12832
rect 70444 12536 70484 13168
rect 70540 13159 70580 13168
rect 70540 12620 70580 12629
rect 70636 12620 70676 13747
rect 70732 13292 70772 13915
rect 70732 13217 70772 13252
rect 70731 13208 70773 13217
rect 70731 13168 70732 13208
rect 70772 13168 70773 13208
rect 70731 13159 70773 13168
rect 70732 13128 70772 13159
rect 70580 12580 70676 12620
rect 70540 12571 70580 12580
rect 70444 12487 70484 12496
rect 70828 12536 70868 13999
rect 71019 13712 71061 13721
rect 71019 13672 71020 13712
rect 71060 13672 71061 13712
rect 71019 13663 71061 13672
rect 70923 13460 70965 13469
rect 70923 13420 70924 13460
rect 70964 13420 70965 13460
rect 70923 13411 70965 13420
rect 70924 13326 70964 13411
rect 70924 12620 70964 12629
rect 71020 12620 71060 13663
rect 71116 13301 71156 15100
rect 71307 14720 71349 14729
rect 71307 14680 71308 14720
rect 71348 14680 71349 14720
rect 71307 14671 71349 14680
rect 71308 14048 71348 14671
rect 71308 13973 71348 14008
rect 71307 13964 71349 13973
rect 71307 13924 71308 13964
rect 71348 13924 71349 13964
rect 71307 13915 71349 13924
rect 71308 13884 71348 13915
rect 71403 13880 71445 13889
rect 71403 13840 71404 13880
rect 71444 13840 71445 13880
rect 71403 13831 71445 13840
rect 71404 13746 71444 13831
rect 71307 13460 71349 13469
rect 71307 13420 71308 13460
rect 71348 13420 71349 13460
rect 71307 13411 71349 13420
rect 71211 13376 71253 13385
rect 71211 13336 71212 13376
rect 71252 13336 71253 13376
rect 71211 13327 71253 13336
rect 71115 13292 71157 13301
rect 71115 13252 71116 13292
rect 71156 13252 71157 13292
rect 71115 13243 71157 13252
rect 70964 12580 71060 12620
rect 70924 12571 70964 12580
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 7112 12116 7480 12125
rect 7152 12076 7194 12116
rect 7234 12076 7276 12116
rect 7316 12076 7358 12116
rect 7398 12076 7440 12116
rect 7112 12067 7480 12076
rect 11112 12116 11480 12125
rect 11152 12076 11194 12116
rect 11234 12076 11276 12116
rect 11316 12076 11358 12116
rect 11398 12076 11440 12116
rect 11112 12067 11480 12076
rect 15112 12116 15480 12125
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15112 12067 15480 12076
rect 19112 12116 19480 12125
rect 19152 12076 19194 12116
rect 19234 12076 19276 12116
rect 19316 12076 19358 12116
rect 19398 12076 19440 12116
rect 19112 12067 19480 12076
rect 23112 12116 23480 12125
rect 23152 12076 23194 12116
rect 23234 12076 23276 12116
rect 23316 12076 23358 12116
rect 23398 12076 23440 12116
rect 23112 12067 23480 12076
rect 27112 12116 27480 12125
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27112 12067 27480 12076
rect 31112 12116 31480 12125
rect 31152 12076 31194 12116
rect 31234 12076 31276 12116
rect 31316 12076 31358 12116
rect 31398 12076 31440 12116
rect 31112 12067 31480 12076
rect 35112 12116 35480 12125
rect 35152 12076 35194 12116
rect 35234 12076 35276 12116
rect 35316 12076 35358 12116
rect 35398 12076 35440 12116
rect 35112 12067 35480 12076
rect 39112 12116 39480 12125
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39112 12067 39480 12076
rect 43112 12116 43480 12125
rect 43152 12076 43194 12116
rect 43234 12076 43276 12116
rect 43316 12076 43358 12116
rect 43398 12076 43440 12116
rect 43112 12067 43480 12076
rect 47112 12116 47480 12125
rect 47152 12076 47194 12116
rect 47234 12076 47276 12116
rect 47316 12076 47358 12116
rect 47398 12076 47440 12116
rect 47112 12067 47480 12076
rect 51112 12116 51480 12125
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51112 12067 51480 12076
rect 55112 12116 55480 12125
rect 55152 12076 55194 12116
rect 55234 12076 55276 12116
rect 55316 12076 55358 12116
rect 55398 12076 55440 12116
rect 55112 12067 55480 12076
rect 59112 12116 59480 12125
rect 59152 12076 59194 12116
rect 59234 12076 59276 12116
rect 59316 12076 59358 12116
rect 59398 12076 59440 12116
rect 59112 12067 59480 12076
rect 63112 12116 63480 12125
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63112 12067 63480 12076
rect 67112 12116 67480 12125
rect 67152 12076 67194 12116
rect 67234 12076 67276 12116
rect 67316 12076 67358 12116
rect 67398 12076 67440 12116
rect 67112 12067 67480 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 8352 11360 8720 11369
rect 8392 11320 8434 11360
rect 8474 11320 8516 11360
rect 8556 11320 8598 11360
rect 8638 11320 8680 11360
rect 8352 11311 8720 11320
rect 12352 11360 12720 11369
rect 12392 11320 12434 11360
rect 12474 11320 12516 11360
rect 12556 11320 12598 11360
rect 12638 11320 12680 11360
rect 12352 11311 12720 11320
rect 16352 11360 16720 11369
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16352 11311 16720 11320
rect 20352 11360 20720 11369
rect 20392 11320 20434 11360
rect 20474 11320 20516 11360
rect 20556 11320 20598 11360
rect 20638 11320 20680 11360
rect 20352 11311 20720 11320
rect 24352 11360 24720 11369
rect 24392 11320 24434 11360
rect 24474 11320 24516 11360
rect 24556 11320 24598 11360
rect 24638 11320 24680 11360
rect 24352 11311 24720 11320
rect 28352 11360 28720 11369
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28352 11311 28720 11320
rect 32352 11360 32720 11369
rect 32392 11320 32434 11360
rect 32474 11320 32516 11360
rect 32556 11320 32598 11360
rect 32638 11320 32680 11360
rect 32352 11311 32720 11320
rect 36352 11360 36720 11369
rect 36392 11320 36434 11360
rect 36474 11320 36516 11360
rect 36556 11320 36598 11360
rect 36638 11320 36680 11360
rect 36352 11311 36720 11320
rect 40352 11360 40720 11369
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40352 11311 40720 11320
rect 44352 11360 44720 11369
rect 44392 11320 44434 11360
rect 44474 11320 44516 11360
rect 44556 11320 44598 11360
rect 44638 11320 44680 11360
rect 44352 11311 44720 11320
rect 48352 11360 48720 11369
rect 48392 11320 48434 11360
rect 48474 11320 48516 11360
rect 48556 11320 48598 11360
rect 48638 11320 48680 11360
rect 48352 11311 48720 11320
rect 52352 11360 52720 11369
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52352 11311 52720 11320
rect 56352 11360 56720 11369
rect 56392 11320 56434 11360
rect 56474 11320 56516 11360
rect 56556 11320 56598 11360
rect 56638 11320 56680 11360
rect 56352 11311 56720 11320
rect 60352 11360 60720 11369
rect 60392 11320 60434 11360
rect 60474 11320 60516 11360
rect 60556 11320 60598 11360
rect 60638 11320 60680 11360
rect 60352 11311 60720 11320
rect 64352 11360 64720 11369
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64352 11311 64720 11320
rect 68352 11360 68720 11369
rect 68392 11320 68434 11360
rect 68474 11320 68516 11360
rect 68556 11320 68598 11360
rect 68638 11320 68680 11360
rect 68352 11311 68720 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 7112 10604 7480 10613
rect 7152 10564 7194 10604
rect 7234 10564 7276 10604
rect 7316 10564 7358 10604
rect 7398 10564 7440 10604
rect 7112 10555 7480 10564
rect 11112 10604 11480 10613
rect 11152 10564 11194 10604
rect 11234 10564 11276 10604
rect 11316 10564 11358 10604
rect 11398 10564 11440 10604
rect 11112 10555 11480 10564
rect 15112 10604 15480 10613
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15112 10555 15480 10564
rect 19112 10604 19480 10613
rect 19152 10564 19194 10604
rect 19234 10564 19276 10604
rect 19316 10564 19358 10604
rect 19398 10564 19440 10604
rect 19112 10555 19480 10564
rect 23112 10604 23480 10613
rect 23152 10564 23194 10604
rect 23234 10564 23276 10604
rect 23316 10564 23358 10604
rect 23398 10564 23440 10604
rect 23112 10555 23480 10564
rect 27112 10604 27480 10613
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27112 10555 27480 10564
rect 31112 10604 31480 10613
rect 31152 10564 31194 10604
rect 31234 10564 31276 10604
rect 31316 10564 31358 10604
rect 31398 10564 31440 10604
rect 31112 10555 31480 10564
rect 35112 10604 35480 10613
rect 35152 10564 35194 10604
rect 35234 10564 35276 10604
rect 35316 10564 35358 10604
rect 35398 10564 35440 10604
rect 35112 10555 35480 10564
rect 39112 10604 39480 10613
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39112 10555 39480 10564
rect 43112 10604 43480 10613
rect 43152 10564 43194 10604
rect 43234 10564 43276 10604
rect 43316 10564 43358 10604
rect 43398 10564 43440 10604
rect 43112 10555 43480 10564
rect 47112 10604 47480 10613
rect 47152 10564 47194 10604
rect 47234 10564 47276 10604
rect 47316 10564 47358 10604
rect 47398 10564 47440 10604
rect 47112 10555 47480 10564
rect 51112 10604 51480 10613
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51112 10555 51480 10564
rect 55112 10604 55480 10613
rect 55152 10564 55194 10604
rect 55234 10564 55276 10604
rect 55316 10564 55358 10604
rect 55398 10564 55440 10604
rect 55112 10555 55480 10564
rect 59112 10604 59480 10613
rect 59152 10564 59194 10604
rect 59234 10564 59276 10604
rect 59316 10564 59358 10604
rect 59398 10564 59440 10604
rect 59112 10555 59480 10564
rect 63112 10604 63480 10613
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63112 10555 63480 10564
rect 67112 10604 67480 10613
rect 67152 10564 67194 10604
rect 67234 10564 67276 10604
rect 67316 10564 67358 10604
rect 67398 10564 67440 10604
rect 67112 10555 67480 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 8352 9848 8720 9857
rect 8392 9808 8434 9848
rect 8474 9808 8516 9848
rect 8556 9808 8598 9848
rect 8638 9808 8680 9848
rect 8352 9799 8720 9808
rect 12352 9848 12720 9857
rect 12392 9808 12434 9848
rect 12474 9808 12516 9848
rect 12556 9808 12598 9848
rect 12638 9808 12680 9848
rect 12352 9799 12720 9808
rect 16352 9848 16720 9857
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16352 9799 16720 9808
rect 20352 9848 20720 9857
rect 20392 9808 20434 9848
rect 20474 9808 20516 9848
rect 20556 9808 20598 9848
rect 20638 9808 20680 9848
rect 20352 9799 20720 9808
rect 24352 9848 24720 9857
rect 24392 9808 24434 9848
rect 24474 9808 24516 9848
rect 24556 9808 24598 9848
rect 24638 9808 24680 9848
rect 24352 9799 24720 9808
rect 28352 9848 28720 9857
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28352 9799 28720 9808
rect 32352 9848 32720 9857
rect 32392 9808 32434 9848
rect 32474 9808 32516 9848
rect 32556 9808 32598 9848
rect 32638 9808 32680 9848
rect 32352 9799 32720 9808
rect 36352 9848 36720 9857
rect 36392 9808 36434 9848
rect 36474 9808 36516 9848
rect 36556 9808 36598 9848
rect 36638 9808 36680 9848
rect 36352 9799 36720 9808
rect 40352 9848 40720 9857
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40352 9799 40720 9808
rect 44352 9848 44720 9857
rect 44392 9808 44434 9848
rect 44474 9808 44516 9848
rect 44556 9808 44598 9848
rect 44638 9808 44680 9848
rect 44352 9799 44720 9808
rect 48352 9848 48720 9857
rect 48392 9808 48434 9848
rect 48474 9808 48516 9848
rect 48556 9808 48598 9848
rect 48638 9808 48680 9848
rect 48352 9799 48720 9808
rect 52352 9848 52720 9857
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52352 9799 52720 9808
rect 56352 9848 56720 9857
rect 56392 9808 56434 9848
rect 56474 9808 56516 9848
rect 56556 9808 56598 9848
rect 56638 9808 56680 9848
rect 56352 9799 56720 9808
rect 60352 9848 60720 9857
rect 60392 9808 60434 9848
rect 60474 9808 60516 9848
rect 60556 9808 60598 9848
rect 60638 9808 60680 9848
rect 60352 9799 60720 9808
rect 64352 9848 64720 9857
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64352 9799 64720 9808
rect 68352 9848 68720 9857
rect 68392 9808 68434 9848
rect 68474 9808 68516 9848
rect 68556 9808 68598 9848
rect 68638 9808 68680 9848
rect 68352 9799 68720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 7112 9092 7480 9101
rect 7152 9052 7194 9092
rect 7234 9052 7276 9092
rect 7316 9052 7358 9092
rect 7398 9052 7440 9092
rect 7112 9043 7480 9052
rect 11112 9092 11480 9101
rect 11152 9052 11194 9092
rect 11234 9052 11276 9092
rect 11316 9052 11358 9092
rect 11398 9052 11440 9092
rect 11112 9043 11480 9052
rect 15112 9092 15480 9101
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15112 9043 15480 9052
rect 19112 9092 19480 9101
rect 19152 9052 19194 9092
rect 19234 9052 19276 9092
rect 19316 9052 19358 9092
rect 19398 9052 19440 9092
rect 19112 9043 19480 9052
rect 23112 9092 23480 9101
rect 23152 9052 23194 9092
rect 23234 9052 23276 9092
rect 23316 9052 23358 9092
rect 23398 9052 23440 9092
rect 23112 9043 23480 9052
rect 27112 9092 27480 9101
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27112 9043 27480 9052
rect 31112 9092 31480 9101
rect 31152 9052 31194 9092
rect 31234 9052 31276 9092
rect 31316 9052 31358 9092
rect 31398 9052 31440 9092
rect 31112 9043 31480 9052
rect 35112 9092 35480 9101
rect 35152 9052 35194 9092
rect 35234 9052 35276 9092
rect 35316 9052 35358 9092
rect 35398 9052 35440 9092
rect 35112 9043 35480 9052
rect 39112 9092 39480 9101
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39112 9043 39480 9052
rect 43112 9092 43480 9101
rect 43152 9052 43194 9092
rect 43234 9052 43276 9092
rect 43316 9052 43358 9092
rect 43398 9052 43440 9092
rect 43112 9043 43480 9052
rect 47112 9092 47480 9101
rect 47152 9052 47194 9092
rect 47234 9052 47276 9092
rect 47316 9052 47358 9092
rect 47398 9052 47440 9092
rect 47112 9043 47480 9052
rect 51112 9092 51480 9101
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51112 9043 51480 9052
rect 55112 9092 55480 9101
rect 55152 9052 55194 9092
rect 55234 9052 55276 9092
rect 55316 9052 55358 9092
rect 55398 9052 55440 9092
rect 55112 9043 55480 9052
rect 59112 9092 59480 9101
rect 59152 9052 59194 9092
rect 59234 9052 59276 9092
rect 59316 9052 59358 9092
rect 59398 9052 59440 9092
rect 59112 9043 59480 9052
rect 63112 9092 63480 9101
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63112 9043 63480 9052
rect 67112 9092 67480 9101
rect 67152 9052 67194 9092
rect 67234 9052 67276 9092
rect 67316 9052 67358 9092
rect 67398 9052 67440 9092
rect 67112 9043 67480 9052
rect 2092 8707 2132 8716
rect 70828 8672 70868 12496
rect 71116 12536 71156 13243
rect 71212 12620 71252 13327
rect 71308 13326 71348 13411
rect 71212 12571 71252 12580
rect 71116 11612 71156 12496
rect 71116 11572 71252 11612
rect 70924 8672 70964 8681
rect 70828 8632 70924 8672
rect 70924 8623 70964 8632
rect 71116 8672 71156 8681
rect 1900 8504 1940 8513
rect 1324 8464 1900 8504
rect 652 8177 692 8464
rect 651 8168 693 8177
rect 651 8128 652 8168
rect 692 8128 693 8168
rect 651 8119 693 8128
rect 844 7916 884 7925
rect 652 7748 692 7757
rect 652 7337 692 7708
rect 844 7421 884 7876
rect 843 7412 885 7421
rect 843 7372 844 7412
rect 884 7372 885 7412
rect 843 7363 885 7372
rect 1515 7412 1557 7421
rect 1515 7372 1516 7412
rect 1556 7372 1557 7412
rect 1515 7363 1557 7372
rect 651 7328 693 7337
rect 651 7288 652 7328
rect 692 7288 693 7328
rect 651 7279 693 7288
rect 1516 7278 1556 7363
rect 844 7244 884 7253
rect 1708 7244 1748 8464
rect 1900 8455 1940 8464
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 8352 8336 8720 8345
rect 8392 8296 8434 8336
rect 8474 8296 8516 8336
rect 8556 8296 8598 8336
rect 8638 8296 8680 8336
rect 8352 8287 8720 8296
rect 12352 8336 12720 8345
rect 12392 8296 12434 8336
rect 12474 8296 12516 8336
rect 12556 8296 12598 8336
rect 12638 8296 12680 8336
rect 12352 8287 12720 8296
rect 16352 8336 16720 8345
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16352 8287 16720 8296
rect 20352 8336 20720 8345
rect 20392 8296 20434 8336
rect 20474 8296 20516 8336
rect 20556 8296 20598 8336
rect 20638 8296 20680 8336
rect 20352 8287 20720 8296
rect 24352 8336 24720 8345
rect 24392 8296 24434 8336
rect 24474 8296 24516 8336
rect 24556 8296 24598 8336
rect 24638 8296 24680 8336
rect 24352 8287 24720 8296
rect 28352 8336 28720 8345
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28352 8287 28720 8296
rect 32352 8336 32720 8345
rect 32392 8296 32434 8336
rect 32474 8296 32516 8336
rect 32556 8296 32598 8336
rect 32638 8296 32680 8336
rect 32352 8287 32720 8296
rect 36352 8336 36720 8345
rect 36392 8296 36434 8336
rect 36474 8296 36516 8336
rect 36556 8296 36598 8336
rect 36638 8296 36680 8336
rect 36352 8287 36720 8296
rect 40352 8336 40720 8345
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40352 8287 40720 8296
rect 44352 8336 44720 8345
rect 44392 8296 44434 8336
rect 44474 8296 44516 8336
rect 44556 8296 44598 8336
rect 44638 8296 44680 8336
rect 44352 8287 44720 8296
rect 48352 8336 48720 8345
rect 48392 8296 48434 8336
rect 48474 8296 48516 8336
rect 48556 8296 48598 8336
rect 48638 8296 48680 8336
rect 48352 8287 48720 8296
rect 52352 8336 52720 8345
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52352 8287 52720 8296
rect 56352 8336 56720 8345
rect 56392 8296 56434 8336
rect 56474 8296 56516 8336
rect 56556 8296 56598 8336
rect 56638 8296 56680 8336
rect 56352 8287 56720 8296
rect 60352 8336 60720 8345
rect 60392 8296 60434 8336
rect 60474 8296 60516 8336
rect 60556 8296 60598 8336
rect 60638 8296 60680 8336
rect 60352 8287 60720 8296
rect 64352 8336 64720 8345
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64352 8287 64720 8296
rect 68352 8336 68720 8345
rect 68392 8296 68434 8336
rect 68474 8296 68516 8336
rect 68556 8296 68598 8336
rect 68638 8296 68680 8336
rect 68352 8287 68720 8296
rect 71116 8084 71156 8632
rect 70828 8044 71156 8084
rect 70828 7916 70868 8044
rect 70828 7867 70868 7876
rect 71019 7916 71061 7925
rect 71019 7876 71020 7916
rect 71060 7876 71061 7916
rect 71019 7867 71061 7876
rect 71020 7832 71060 7867
rect 71020 7781 71060 7792
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 7112 7580 7480 7589
rect 7152 7540 7194 7580
rect 7234 7540 7276 7580
rect 7316 7540 7358 7580
rect 7398 7540 7440 7580
rect 7112 7531 7480 7540
rect 11112 7580 11480 7589
rect 11152 7540 11194 7580
rect 11234 7540 11276 7580
rect 11316 7540 11358 7580
rect 11398 7540 11440 7580
rect 11112 7531 11480 7540
rect 15112 7580 15480 7589
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15112 7531 15480 7540
rect 19112 7580 19480 7589
rect 19152 7540 19194 7580
rect 19234 7540 19276 7580
rect 19316 7540 19358 7580
rect 19398 7540 19440 7580
rect 19112 7531 19480 7540
rect 23112 7580 23480 7589
rect 23152 7540 23194 7580
rect 23234 7540 23276 7580
rect 23316 7540 23358 7580
rect 23398 7540 23440 7580
rect 23112 7531 23480 7540
rect 27112 7580 27480 7589
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27112 7531 27480 7540
rect 31112 7580 31480 7589
rect 31152 7540 31194 7580
rect 31234 7540 31276 7580
rect 31316 7540 31358 7580
rect 31398 7540 31440 7580
rect 31112 7531 31480 7540
rect 35112 7580 35480 7589
rect 35152 7540 35194 7580
rect 35234 7540 35276 7580
rect 35316 7540 35358 7580
rect 35398 7540 35440 7580
rect 35112 7531 35480 7540
rect 39112 7580 39480 7589
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39112 7531 39480 7540
rect 43112 7580 43480 7589
rect 43152 7540 43194 7580
rect 43234 7540 43276 7580
rect 43316 7540 43358 7580
rect 43398 7540 43440 7580
rect 43112 7531 43480 7540
rect 47112 7580 47480 7589
rect 47152 7540 47194 7580
rect 47234 7540 47276 7580
rect 47316 7540 47358 7580
rect 47398 7540 47440 7580
rect 47112 7531 47480 7540
rect 51112 7580 51480 7589
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51112 7531 51480 7540
rect 55112 7580 55480 7589
rect 55152 7540 55194 7580
rect 55234 7540 55276 7580
rect 55316 7540 55358 7580
rect 55398 7540 55440 7580
rect 55112 7531 55480 7540
rect 59112 7580 59480 7589
rect 59152 7540 59194 7580
rect 59234 7540 59276 7580
rect 59316 7540 59358 7580
rect 59398 7540 59440 7580
rect 59112 7531 59480 7540
rect 63112 7580 63480 7589
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63112 7531 63480 7540
rect 67112 7580 67480 7589
rect 67152 7540 67194 7580
rect 67234 7540 67276 7580
rect 67316 7540 67358 7580
rect 67398 7540 67440 7580
rect 67112 7531 67480 7540
rect 652 6992 692 7001
rect 652 6497 692 6952
rect 844 6665 884 7204
rect 1612 7204 1708 7244
rect 843 6656 885 6665
rect 843 6616 844 6656
rect 884 6616 885 6656
rect 843 6607 885 6616
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 1516 6404 1556 6413
rect 1612 6404 1652 7204
rect 1708 7195 1748 7204
rect 71116 7169 71156 8044
rect 71212 7916 71252 11572
rect 71252 7876 71348 7916
rect 71212 7867 71252 7876
rect 71115 7160 71157 7169
rect 71115 7120 71116 7160
rect 71156 7120 71157 7160
rect 71115 7111 71157 7120
rect 71308 7160 71348 7876
rect 71403 7832 71445 7841
rect 71403 7792 71404 7832
rect 71444 7792 71445 7832
rect 71403 7783 71445 7792
rect 71404 7698 71444 7783
rect 71499 7748 71541 7757
rect 71499 7708 71500 7748
rect 71540 7708 71541 7748
rect 71499 7699 71541 7708
rect 71404 7412 71444 7421
rect 71500 7412 71540 7699
rect 71788 7421 71828 16351
rect 73899 16316 73941 16325
rect 73899 16276 73900 16316
rect 73940 16276 73941 16316
rect 73899 16267 73941 16276
rect 74284 16316 74324 16327
rect 74476 16325 74516 16360
rect 80428 16325 80468 16948
rect 86188 16988 86228 16997
rect 80620 16820 80660 16829
rect 80620 16325 80660 16780
rect 83112 16652 83480 16661
rect 83152 16612 83194 16652
rect 83234 16612 83276 16652
rect 83316 16612 83358 16652
rect 83398 16612 83440 16652
rect 83112 16603 83480 16612
rect 86188 16409 86228 16948
rect 86380 16820 86420 16829
rect 81580 16400 81620 16409
rect 73131 16232 73173 16241
rect 73131 16192 73132 16232
rect 73172 16192 73173 16232
rect 73131 16183 73173 16192
rect 72352 15896 72720 15905
rect 72392 15856 72434 15896
rect 72474 15856 72516 15896
rect 72556 15856 72598 15896
rect 72638 15856 72680 15896
rect 72352 15847 72720 15856
rect 73036 14804 73076 14815
rect 73036 14729 73076 14764
rect 72747 14720 72789 14729
rect 72747 14680 72748 14720
rect 72788 14680 72789 14720
rect 72747 14671 72789 14680
rect 73035 14720 73077 14729
rect 73035 14680 73036 14720
rect 73076 14680 73077 14720
rect 73035 14671 73077 14680
rect 72748 14586 72788 14671
rect 72843 14552 72885 14561
rect 72843 14512 72844 14552
rect 72884 14512 72885 14552
rect 72843 14503 72885 14512
rect 72844 14418 72884 14503
rect 73132 14057 73172 16183
rect 73900 16182 73940 16267
rect 74284 16241 74324 16276
rect 74475 16316 74517 16325
rect 74475 16276 74476 16316
rect 74516 16276 74517 16316
rect 74475 16267 74517 16276
rect 76780 16316 76820 16325
rect 74283 16232 74325 16241
rect 74283 16192 74284 16232
rect 74324 16192 74325 16232
rect 74283 16183 74325 16192
rect 76780 16073 76820 16276
rect 77163 16316 77205 16325
rect 77163 16276 77164 16316
rect 77204 16276 77205 16316
rect 77163 16267 77205 16276
rect 80427 16316 80469 16325
rect 80427 16276 80428 16316
rect 80468 16276 80469 16316
rect 80427 16267 80469 16276
rect 80524 16316 80564 16325
rect 80619 16316 80661 16325
rect 80564 16276 80620 16316
rect 80660 16276 80661 16316
rect 80524 16267 80564 16276
rect 80619 16267 80661 16276
rect 81196 16316 81236 16325
rect 81580 16316 81620 16360
rect 83115 16400 83157 16409
rect 83115 16360 83116 16400
rect 83156 16360 83157 16400
rect 83115 16351 83157 16360
rect 83403 16400 83445 16409
rect 83403 16360 83404 16400
rect 83444 16360 83445 16400
rect 83403 16351 83445 16360
rect 83787 16400 83829 16409
rect 83787 16360 83788 16400
rect 83828 16360 83829 16400
rect 83787 16351 83829 16360
rect 86187 16400 86229 16409
rect 86187 16360 86188 16400
rect 86228 16360 86229 16400
rect 86187 16351 86229 16360
rect 81236 16276 81620 16316
rect 81196 16267 81236 16276
rect 77164 16182 77204 16267
rect 80620 16182 80660 16267
rect 81580 16073 81620 16276
rect 81771 16316 81813 16325
rect 81771 16276 81772 16316
rect 81812 16276 81813 16316
rect 81771 16267 81813 16276
rect 82156 16316 82196 16325
rect 82540 16316 82580 16325
rect 82196 16276 82292 16316
rect 82156 16267 82196 16276
rect 81772 16182 81812 16267
rect 82252 16073 82292 16276
rect 74092 16064 74132 16073
rect 76779 16064 76821 16073
rect 76972 16064 77012 16073
rect 74132 16024 74324 16064
rect 74092 16015 74132 16024
rect 73707 15476 73749 15485
rect 73707 15436 73708 15476
rect 73748 15436 73749 15476
rect 73707 15427 73749 15436
rect 74091 15476 74133 15485
rect 74284 15476 74324 16024
rect 76779 16024 76780 16064
rect 76820 16024 76916 16064
rect 76779 16015 76821 16024
rect 76352 15896 76720 15905
rect 76392 15856 76434 15896
rect 76474 15856 76516 15896
rect 76556 15856 76598 15896
rect 76638 15856 76680 15896
rect 76352 15847 76720 15856
rect 74091 15436 74092 15476
rect 74132 15436 74133 15476
rect 74091 15427 74133 15436
rect 74188 15436 74284 15476
rect 73708 15342 73748 15427
rect 74092 15392 74132 15427
rect 74092 15341 74132 15352
rect 73899 15308 73941 15317
rect 73899 15268 73900 15308
rect 73940 15268 73941 15308
rect 73899 15259 73941 15268
rect 73900 15174 73940 15259
rect 73708 14888 73748 14897
rect 73748 14848 74132 14888
rect 73708 14839 73748 14848
rect 73516 14804 73556 14815
rect 73516 14729 73556 14764
rect 73515 14720 73557 14729
rect 73515 14680 73516 14720
rect 73556 14680 73557 14720
rect 73515 14671 73557 14680
rect 73899 14720 73941 14729
rect 73899 14680 73900 14720
rect 73940 14680 73941 14720
rect 73899 14671 73941 14680
rect 73900 14586 73940 14671
rect 73228 14552 73268 14561
rect 73996 14552 74036 14561
rect 73268 14512 73652 14552
rect 73228 14503 73268 14512
rect 73131 14048 73173 14057
rect 73131 14008 73132 14048
rect 73172 14008 73173 14048
rect 73131 13999 73173 14008
rect 73515 13880 73557 13889
rect 73515 13840 73516 13880
rect 73556 13840 73557 13880
rect 73515 13831 73557 13840
rect 73131 13796 73173 13805
rect 73131 13756 73132 13796
rect 73172 13756 73173 13796
rect 73131 13747 73173 13756
rect 72651 13712 72693 13721
rect 72651 13672 72652 13712
rect 72692 13672 72693 13712
rect 72651 13663 72693 13672
rect 72652 13544 72692 13663
rect 72843 13544 72885 13553
rect 73132 13544 73172 13747
rect 73227 13544 73269 13553
rect 73516 13544 73556 13831
rect 72652 13504 72745 13544
rect 72414 13460 72456 13469
rect 72414 13420 72415 13460
rect 72455 13420 72456 13460
rect 72414 13411 72456 13420
rect 72304 13376 72346 13385
rect 72304 13336 72305 13376
rect 72345 13336 72346 13376
rect 72304 13327 72346 13336
rect 72305 13188 72345 13327
rect 72415 13188 72455 13411
rect 72705 13188 72745 13504
rect 72815 13504 72844 13544
rect 72884 13504 72885 13544
rect 72815 13495 72885 13504
rect 73105 13504 73172 13544
rect 73215 13504 73228 13544
rect 73268 13504 73269 13544
rect 72815 13188 72855 13495
rect 73105 13188 73145 13504
rect 73215 13495 73269 13504
rect 73505 13504 73556 13544
rect 73612 13544 73652 14512
rect 73996 13544 74036 14512
rect 73612 13504 73655 13544
rect 73215 13188 73255 13495
rect 73505 13188 73545 13504
rect 73615 13188 73655 13504
rect 73905 13504 74036 13544
rect 73905 13188 73945 13504
rect 74092 13460 74132 14848
rect 74188 14729 74228 15436
rect 74284 15427 74324 15436
rect 74475 15476 74517 15485
rect 74475 15436 74476 15476
rect 74516 15436 74517 15476
rect 74475 15427 74517 15436
rect 74859 15476 74901 15485
rect 75340 15476 75380 15485
rect 74859 15436 74860 15476
rect 74900 15436 74901 15476
rect 74859 15427 74901 15436
rect 75244 15436 75340 15476
rect 74379 15308 74421 15317
rect 74379 15268 74380 15308
rect 74420 15268 74421 15308
rect 74379 15259 74421 15268
rect 74187 14720 74229 14729
rect 74187 14680 74188 14720
rect 74228 14680 74229 14720
rect 74187 14671 74229 14680
rect 74188 14586 74228 14671
rect 74284 14552 74324 14561
rect 74187 14468 74229 14477
rect 74187 14428 74188 14468
rect 74228 14428 74229 14468
rect 74187 14419 74229 14428
rect 74015 13420 74132 13460
rect 74188 13460 74228 14419
rect 74284 13637 74324 14512
rect 74283 13628 74325 13637
rect 74283 13588 74284 13628
rect 74324 13588 74325 13628
rect 74283 13579 74325 13588
rect 74380 13544 74420 15259
rect 74476 14804 74516 15427
rect 74860 15342 74900 15427
rect 75052 15308 75092 15317
rect 75092 15268 75188 15308
rect 75052 15259 75092 15268
rect 74476 14755 74516 14764
rect 74859 14720 74901 14729
rect 74859 14680 74860 14720
rect 74900 14680 74901 14720
rect 74859 14671 74901 14680
rect 74860 14586 74900 14671
rect 74668 14552 74708 14561
rect 74956 14552 74996 14561
rect 74708 14512 74804 14552
rect 74668 14503 74708 14512
rect 74667 13628 74709 13637
rect 74667 13588 74668 13628
rect 74708 13588 74709 13628
rect 74667 13579 74709 13588
rect 74380 13504 74455 13544
rect 74188 13420 74345 13460
rect 74015 13188 74055 13420
rect 74305 13188 74345 13420
rect 74415 13188 74455 13504
rect 74668 13460 74708 13579
rect 74764 13544 74804 14512
rect 74996 14512 75092 14552
rect 74956 14503 74996 14512
rect 75052 13544 75092 14512
rect 75148 13628 75188 15268
rect 75244 14729 75284 15436
rect 75340 15427 75380 15436
rect 75820 15476 75860 15485
rect 75820 15317 75860 15436
rect 76204 15476 76244 15485
rect 76204 15317 76244 15436
rect 76588 15476 76628 15485
rect 76588 15317 76628 15436
rect 75339 15308 75381 15317
rect 75339 15268 75340 15308
rect 75380 15268 75381 15308
rect 75339 15259 75381 15268
rect 75532 15308 75572 15317
rect 75243 14720 75285 14729
rect 75243 14680 75244 14720
rect 75284 14680 75285 14720
rect 75243 14671 75285 14680
rect 75340 14720 75380 15259
rect 75340 14671 75380 14680
rect 75436 14552 75476 14561
rect 75148 13588 75255 13628
rect 74764 13504 74855 13544
rect 75052 13504 75145 13544
rect 74668 13420 74745 13460
rect 74705 13188 74745 13420
rect 74815 13188 74855 13504
rect 75105 13188 75145 13504
rect 75215 13188 75255 13588
rect 75436 13376 75476 14512
rect 75532 13544 75572 15268
rect 75819 15308 75861 15317
rect 75819 15268 75820 15308
rect 75860 15268 75861 15308
rect 75819 15259 75861 15268
rect 76012 15308 76052 15317
rect 75819 14720 75861 14729
rect 75819 14680 75820 14720
rect 75860 14680 75861 14720
rect 75819 14671 75861 14680
rect 75820 14586 75860 14671
rect 75916 14552 75956 14561
rect 75532 13504 75655 13544
rect 75436 13336 75545 13376
rect 75505 13188 75545 13336
rect 75615 13188 75655 13504
rect 75916 13460 75956 14512
rect 76012 13544 76052 15268
rect 76203 15308 76245 15317
rect 76203 15268 76204 15308
rect 76244 15268 76245 15308
rect 76203 15259 76245 15268
rect 76396 15308 76436 15317
rect 76107 14720 76149 14729
rect 76107 14680 76108 14720
rect 76148 14680 76149 14720
rect 76107 14671 76149 14680
rect 76108 14586 76148 14671
rect 76204 14552 76244 14561
rect 76244 14512 76340 14552
rect 76204 14503 76244 14512
rect 76300 13544 76340 14512
rect 76396 13544 76436 15268
rect 76587 15308 76629 15317
rect 76587 15268 76588 15308
rect 76628 15268 76629 15308
rect 76587 15259 76629 15268
rect 76780 15308 76820 15317
rect 76588 14720 76628 15259
rect 76588 14671 76628 14680
rect 76684 14552 76724 14561
rect 76012 13504 76055 13544
rect 76300 13504 76345 13544
rect 76396 13504 76455 13544
rect 75905 13420 75956 13460
rect 75905 13188 75945 13420
rect 76015 13188 76055 13504
rect 76305 13188 76345 13504
rect 76415 13188 76455 13504
rect 76684 13460 76724 14512
rect 76780 13544 76820 15268
rect 76876 15149 76916 16024
rect 76972 15476 77012 16024
rect 77355 16064 77397 16073
rect 80332 16064 80372 16073
rect 77355 16024 77356 16064
rect 77396 16024 77397 16064
rect 77355 16015 77397 16024
rect 80236 16024 80332 16064
rect 77356 15930 77396 16015
rect 76972 15233 77012 15436
rect 77356 15476 77396 15485
rect 77164 15308 77204 15317
rect 77204 15268 77300 15308
rect 77164 15259 77204 15268
rect 76971 15224 77013 15233
rect 76971 15184 76972 15224
rect 77012 15184 77013 15224
rect 76971 15175 77013 15184
rect 76875 15140 76917 15149
rect 76875 15100 76876 15140
rect 76916 15100 76917 15140
rect 76875 15091 76917 15100
rect 76876 14720 76916 15091
rect 76972 14720 77012 14729
rect 76876 14680 76972 14720
rect 76972 14671 77012 14680
rect 77068 14552 77108 14561
rect 76780 13504 76855 13544
rect 76684 13420 76745 13460
rect 76705 13188 76745 13420
rect 76815 13188 76855 13504
rect 77068 13460 77108 14512
rect 77260 13460 77300 15268
rect 77356 15233 77396 15436
rect 77740 15476 77780 15485
rect 77548 15308 77588 15317
rect 77355 15224 77397 15233
rect 77355 15184 77356 15224
rect 77396 15184 77397 15224
rect 77355 15175 77397 15184
rect 77356 14720 77396 15175
rect 77356 14671 77396 14680
rect 77068 13420 77145 13460
rect 77105 13188 77145 13420
rect 77215 13420 77300 13460
rect 77452 14552 77492 14561
rect 77215 13188 77255 13420
rect 77452 13376 77492 14512
rect 77548 13460 77588 15268
rect 77740 15233 77780 15436
rect 78124 15476 78164 15485
rect 77932 15308 77972 15317
rect 77972 15268 78068 15308
rect 77932 15259 77972 15268
rect 77739 15224 77781 15233
rect 77739 15184 77740 15224
rect 77780 15184 77781 15224
rect 77739 15175 77781 15184
rect 77835 15140 77877 15149
rect 77835 15100 77836 15140
rect 77876 15100 77877 15140
rect 77835 15091 77877 15100
rect 77836 14720 77876 15091
rect 77836 14671 77876 14680
rect 77932 14552 77972 14561
rect 77932 13460 77972 14512
rect 78028 13544 78068 15268
rect 78124 15233 78164 15436
rect 78604 15476 78644 15485
rect 78316 15308 78356 15317
rect 78356 15268 78452 15308
rect 78316 15259 78356 15268
rect 78123 15224 78165 15233
rect 78123 15184 78124 15224
rect 78164 15184 78165 15224
rect 78123 15175 78165 15184
rect 78124 14720 78164 15175
rect 78124 14671 78164 14680
rect 77548 13420 77684 13460
rect 77644 13376 77684 13420
rect 77452 13336 77545 13376
rect 77505 13188 77545 13336
rect 77615 13336 77684 13376
rect 77905 13420 77972 13460
rect 78015 13504 78068 13544
rect 78220 14552 78260 14561
rect 78220 13544 78260 14512
rect 78220 13504 78345 13544
rect 77615 13188 77655 13336
rect 77905 13188 77945 13420
rect 78015 13188 78055 13504
rect 78305 13188 78345 13504
rect 78412 13460 78452 15268
rect 78604 15149 78644 15436
rect 79179 15465 79219 15486
rect 79179 15401 79219 15425
rect 79372 15476 79412 15487
rect 80236 15485 80276 16024
rect 80332 16015 80372 16024
rect 81388 16064 81428 16073
rect 81579 16064 81621 16073
rect 81428 16024 81524 16064
rect 81388 16015 81428 16024
rect 80352 15896 80720 15905
rect 80392 15856 80434 15896
rect 80474 15856 80516 15896
rect 80556 15856 80598 15896
rect 80638 15856 80680 15896
rect 80352 15847 80720 15856
rect 79372 15401 79412 15436
rect 79756 15476 79796 15485
rect 80235 15476 80277 15485
rect 78795 15392 78837 15401
rect 79179 15392 79221 15401
rect 78795 15352 78796 15392
rect 78836 15352 78932 15392
rect 78795 15343 78837 15352
rect 78796 15258 78836 15343
rect 78603 15140 78645 15149
rect 78603 15100 78604 15140
rect 78644 15100 78645 15140
rect 78603 15091 78645 15100
rect 78892 14804 78932 15352
rect 79179 15352 79180 15392
rect 79220 15352 79221 15392
rect 79179 15343 79221 15352
rect 79371 15392 79413 15401
rect 79371 15352 79372 15392
rect 79412 15352 79413 15392
rect 79371 15343 79413 15352
rect 79659 15392 79701 15401
rect 79659 15352 79660 15392
rect 79700 15352 79701 15392
rect 79659 15343 79701 15352
rect 78700 14764 78892 14804
rect 78700 14720 78740 14764
rect 78892 14755 78932 14764
rect 78988 15308 79028 15317
rect 78700 14671 78740 14680
rect 78604 14552 78644 14561
rect 78644 14512 78740 14552
rect 78604 14503 78644 14512
rect 78700 13544 78740 14512
rect 78988 13964 79028 15268
rect 79372 14720 79412 15343
rect 79372 14671 79412 14680
rect 79564 15308 79604 15317
rect 79084 14552 79124 14561
rect 79468 14552 79508 14561
rect 79124 14512 79220 14552
rect 79084 14503 79124 14512
rect 78892 13924 79028 13964
rect 78892 13544 78932 13924
rect 79083 13880 79125 13889
rect 79083 13840 79084 13880
rect 79124 13840 79125 13880
rect 79083 13831 79125 13840
rect 78700 13504 78745 13544
rect 78412 13420 78455 13460
rect 78415 13188 78455 13420
rect 78705 13188 78745 13504
rect 78815 13504 78932 13544
rect 78815 13188 78855 13504
rect 79084 13460 79124 13831
rect 79180 13544 79220 14512
rect 79180 13504 79255 13544
rect 79084 13420 79145 13460
rect 79105 13188 79145 13420
rect 79215 13188 79255 13504
rect 79468 13460 79508 14512
rect 79564 13544 79604 15268
rect 79660 14720 79700 15343
rect 79756 15233 79796 15436
rect 80140 15436 80236 15476
rect 80276 15436 80277 15476
rect 79948 15308 79988 15317
rect 79988 15268 80084 15308
rect 79948 15259 79988 15268
rect 79755 15224 79797 15233
rect 79755 15184 79756 15224
rect 79796 15184 79797 15224
rect 79755 15175 79797 15184
rect 79660 14671 79700 14680
rect 79756 14552 79796 14561
rect 79756 13889 79796 14512
rect 79755 13880 79797 13889
rect 79755 13840 79756 13880
rect 79796 13840 79797 13880
rect 79755 13831 79797 13840
rect 80044 13544 80084 15268
rect 80140 14720 80180 15436
rect 80235 15427 80277 15436
rect 80715 15476 80757 15485
rect 81099 15476 81141 15485
rect 80715 15436 80716 15476
rect 80756 15436 80852 15476
rect 80715 15427 80757 15436
rect 80236 15342 80276 15427
rect 80716 15342 80756 15427
rect 80428 15308 80468 15317
rect 80140 14671 80180 14680
rect 80332 15268 80428 15308
rect 79564 13504 79700 13544
rect 79660 13460 79700 13504
rect 80015 13504 80084 13544
rect 80236 14552 80276 14561
rect 79468 13420 79545 13460
rect 79505 13188 79545 13420
rect 79615 13420 79700 13460
rect 79904 13460 79946 13469
rect 79904 13420 79905 13460
rect 79945 13420 79946 13460
rect 79615 13188 79655 13420
rect 79904 13411 79946 13420
rect 79905 13188 79945 13411
rect 80015 13188 80055 13504
rect 80236 13460 80276 14512
rect 80332 13544 80372 15268
rect 80428 15259 80468 15268
rect 80427 15140 80469 15149
rect 80427 15100 80428 15140
rect 80468 15100 80469 15140
rect 80427 15091 80469 15100
rect 80428 14720 80468 15091
rect 80428 14671 80468 14680
rect 80812 14720 80852 15436
rect 81004 15436 81100 15476
rect 81140 15436 81141 15476
rect 80812 14671 80852 14680
rect 80908 15308 80948 15317
rect 80524 14552 80564 14561
rect 80524 13721 80564 14512
rect 80716 14552 80756 14561
rect 80523 13712 80565 13721
rect 80523 13672 80524 13712
rect 80564 13672 80565 13712
rect 80523 13663 80565 13672
rect 80716 13544 80756 14512
rect 80908 13544 80948 15268
rect 81004 14720 81044 15436
rect 81099 15427 81141 15436
rect 81387 15476 81429 15485
rect 81387 15436 81388 15476
rect 81428 15436 81429 15476
rect 81387 15427 81429 15436
rect 81100 15342 81140 15427
rect 81292 15308 81332 15317
rect 81004 14671 81044 14680
rect 81196 15268 81292 15308
rect 80332 13504 80455 13544
rect 80226 13420 80276 13460
rect 80226 13376 80266 13420
rect 80226 13336 80345 13376
rect 80305 13188 80345 13336
rect 80415 13188 80455 13504
rect 80705 13504 80756 13544
rect 80815 13504 80948 13544
rect 81100 14552 81140 14561
rect 80705 13188 80745 13504
rect 80815 13188 80855 13504
rect 81100 13460 81140 14512
rect 81100 13420 81145 13460
rect 81105 13188 81145 13420
rect 81196 13292 81236 15268
rect 81292 15259 81332 15268
rect 81388 14720 81428 15427
rect 81484 14720 81524 16024
rect 81579 16024 81580 16064
rect 81620 16024 81621 16064
rect 81579 16015 81621 16024
rect 81771 16064 81813 16073
rect 81771 16024 81772 16064
rect 81812 16024 81813 16064
rect 81771 16015 81813 16024
rect 81964 16064 82004 16073
rect 82251 16064 82293 16073
rect 82004 16024 82196 16064
rect 81964 16015 82004 16024
rect 81772 15560 81812 16015
rect 81812 15520 82004 15560
rect 81772 15511 81812 15520
rect 81868 15308 81908 15317
rect 81484 14680 81620 14720
rect 81388 14671 81428 14680
rect 81484 14552 81524 14561
rect 81484 13460 81524 14512
rect 81580 13544 81620 14680
rect 81868 14552 81908 15268
rect 81964 14720 82004 15520
rect 81964 14671 82004 14680
rect 82060 14552 82100 14561
rect 81868 14512 82004 14552
rect 81964 13544 82004 14512
rect 82060 13637 82100 14512
rect 82059 13628 82101 13637
rect 82059 13588 82060 13628
rect 82100 13588 82101 13628
rect 82059 13579 82101 13588
rect 81580 13504 81655 13544
rect 81484 13420 81545 13460
rect 81196 13252 81255 13292
rect 81215 13188 81255 13252
rect 81505 13188 81545 13420
rect 81615 13188 81655 13504
rect 81905 13504 82004 13544
rect 81905 13188 81945 13504
rect 82156 13460 82196 16024
rect 82251 16024 82252 16064
rect 82292 16024 82293 16064
rect 82251 16015 82293 16024
rect 82252 14804 82292 16015
rect 82540 15485 82580 16276
rect 83116 16266 83156 16351
rect 83307 16316 83349 16325
rect 83307 16276 83308 16316
rect 83348 16276 83349 16316
rect 83307 16267 83349 16276
rect 83308 16182 83348 16267
rect 82732 16064 82772 16073
rect 82772 16024 82868 16064
rect 82732 16015 82772 16024
rect 82539 15476 82581 15485
rect 82539 15436 82540 15476
rect 82580 15436 82581 15476
rect 82539 15427 82581 15436
rect 82292 14764 82676 14804
rect 82252 14755 82292 14764
rect 82636 14720 82676 14764
rect 82636 14671 82676 14680
rect 82444 14552 82484 14561
rect 82444 13544 82484 14512
rect 82415 13504 82484 13544
rect 82732 14552 82772 14561
rect 82015 13420 82196 13460
rect 82304 13460 82346 13469
rect 82304 13420 82305 13460
rect 82345 13420 82346 13460
rect 82015 13188 82055 13420
rect 82304 13411 82346 13420
rect 82305 13188 82345 13411
rect 82415 13188 82455 13504
rect 82732 13460 82772 14512
rect 82828 13544 82868 16024
rect 83404 15485 83444 16351
rect 83788 16316 83828 16351
rect 86380 16325 86420 16780
rect 83788 16265 83828 16276
rect 84651 16316 84693 16325
rect 84651 16276 84652 16316
rect 84692 16276 84693 16316
rect 84651 16267 84693 16276
rect 86379 16316 86421 16325
rect 86379 16276 86380 16316
rect 86420 16276 86421 16316
rect 86379 16267 86421 16276
rect 84652 16182 84692 16267
rect 86476 16241 86516 17032
rect 86572 17023 86612 17032
rect 86764 17072 86804 17081
rect 86764 16409 86804 17032
rect 87112 16652 87480 16661
rect 87152 16612 87194 16652
rect 87234 16612 87276 16652
rect 87316 16612 87358 16652
rect 87398 16612 87440 16652
rect 87112 16603 87480 16612
rect 91112 16652 91480 16661
rect 91152 16612 91194 16652
rect 91234 16612 91276 16652
rect 91316 16612 91358 16652
rect 91398 16612 91440 16652
rect 91112 16603 91480 16612
rect 95112 16652 95480 16661
rect 95152 16612 95194 16652
rect 95234 16612 95276 16652
rect 95316 16612 95358 16652
rect 95398 16612 95440 16652
rect 95112 16603 95480 16612
rect 99112 16652 99480 16661
rect 99152 16612 99194 16652
rect 99234 16612 99276 16652
rect 99316 16612 99358 16652
rect 99398 16612 99440 16652
rect 99112 16603 99480 16612
rect 86763 16400 86805 16409
rect 86763 16360 86764 16400
rect 86804 16360 86805 16400
rect 86763 16351 86805 16360
rect 86571 16316 86613 16325
rect 86571 16276 86572 16316
rect 86612 16276 86613 16316
rect 86571 16267 86613 16276
rect 87436 16316 87476 16325
rect 86475 16232 86517 16241
rect 86475 16192 86476 16232
rect 86516 16192 86517 16232
rect 86475 16183 86517 16192
rect 86572 16182 86612 16267
rect 83980 16064 84020 16073
rect 84844 16064 84884 16073
rect 86380 16064 86420 16073
rect 84020 16024 84116 16064
rect 83980 16015 84020 16024
rect 83884 15560 83924 15571
rect 83884 15485 83924 15520
rect 83019 15476 83061 15485
rect 83019 15436 83020 15476
rect 83060 15436 83061 15476
rect 83019 15427 83061 15436
rect 83403 15476 83445 15485
rect 83403 15436 83404 15476
rect 83444 15436 83445 15476
rect 83403 15427 83445 15436
rect 83883 15476 83925 15485
rect 83883 15436 83884 15476
rect 83924 15436 83925 15476
rect 83883 15427 83925 15436
rect 83020 14720 83060 15427
rect 83020 14671 83060 14680
rect 83212 15308 83252 15317
rect 82705 13420 82772 13460
rect 82815 13504 82868 13544
rect 83116 14552 83156 14561
rect 82705 13188 82745 13420
rect 82815 13188 82855 13504
rect 83116 13460 83156 14512
rect 83212 13544 83252 15268
rect 83404 14720 83444 15427
rect 83404 14671 83444 14680
rect 83596 15308 83636 15317
rect 83500 14552 83540 14561
rect 83212 13504 83255 13544
rect 83105 13420 83156 13460
rect 83105 13188 83145 13420
rect 83215 13188 83255 13504
rect 83500 13460 83540 14512
rect 83596 13544 83636 15268
rect 83788 14720 83828 14729
rect 83884 14720 83924 15427
rect 83979 15308 84021 15317
rect 83979 15268 83980 15308
rect 84020 15268 84021 15308
rect 83979 15259 84021 15268
rect 83980 15174 84020 15259
rect 83828 14680 83924 14720
rect 83788 14671 83828 14680
rect 83884 14552 83924 14561
rect 83884 13544 83924 14512
rect 84076 13544 84116 16024
rect 84884 16024 85076 16064
rect 84844 16015 84884 16024
rect 84352 15896 84720 15905
rect 84392 15856 84434 15896
rect 84474 15856 84516 15896
rect 84556 15856 84598 15896
rect 84638 15856 84680 15896
rect 84352 15847 84720 15856
rect 85036 15485 85076 16024
rect 86380 15485 86420 16024
rect 87436 15560 87476 16276
rect 88203 16316 88245 16325
rect 88203 16276 88204 16316
rect 88244 16276 88245 16316
rect 88203 16267 88245 16276
rect 89355 16316 89397 16325
rect 89355 16276 89356 16316
rect 89396 16276 89397 16316
rect 89355 16267 89397 16276
rect 90219 16316 90261 16325
rect 90219 16276 90220 16316
rect 90260 16276 90261 16316
rect 90219 16267 90261 16276
rect 90603 16316 90645 16325
rect 90603 16276 90604 16316
rect 90644 16276 90645 16316
rect 90603 16267 90645 16276
rect 92236 16316 92276 16325
rect 88204 16182 88244 16267
rect 89356 16182 89396 16267
rect 87436 15485 87476 15520
rect 87628 16064 87668 16073
rect 84171 15476 84213 15485
rect 84171 15436 84172 15476
rect 84212 15436 84213 15476
rect 84171 15427 84213 15436
rect 84555 15476 84597 15485
rect 84555 15436 84556 15476
rect 84596 15436 84597 15476
rect 84555 15427 84597 15436
rect 85035 15476 85077 15485
rect 85035 15436 85036 15476
rect 85076 15436 85077 15476
rect 85035 15427 85077 15436
rect 85419 15476 85461 15485
rect 85419 15436 85420 15476
rect 85460 15436 85461 15476
rect 85419 15427 85461 15436
rect 85803 15476 85845 15485
rect 85803 15436 85804 15476
rect 85844 15436 85845 15476
rect 85803 15427 85845 15436
rect 86187 15476 86229 15485
rect 86379 15476 86421 15485
rect 86187 15436 86188 15476
rect 86228 15436 86324 15476
rect 86187 15427 86229 15436
rect 84172 15342 84212 15427
rect 84267 15308 84309 15317
rect 84267 15268 84268 15308
rect 84308 15268 84309 15308
rect 84267 15259 84309 15268
rect 84364 15308 84404 15317
rect 84404 15268 84500 15308
rect 84364 15259 84404 15268
rect 83596 13504 83655 13544
rect 83884 13504 83945 13544
rect 83500 13420 83545 13460
rect 83505 13188 83545 13420
rect 83615 13188 83655 13504
rect 83905 13188 83945 13504
rect 84015 13504 84116 13544
rect 84268 13544 84308 15259
rect 84460 13544 84500 15268
rect 84556 14720 84596 15427
rect 84556 14671 84596 14680
rect 84748 15308 84788 15317
rect 84268 13504 84345 13544
rect 84015 13188 84055 13504
rect 84305 13188 84345 13504
rect 84415 13504 84500 13544
rect 84652 14552 84692 14561
rect 84415 13188 84455 13504
rect 84652 13460 84692 14512
rect 84748 13460 84788 15268
rect 85036 14720 85076 15427
rect 85036 14671 85076 14680
rect 85228 15308 85268 15317
rect 85132 14552 85172 14561
rect 85132 13460 85172 14512
rect 85228 13544 85268 15268
rect 85420 14720 85460 15427
rect 85420 14671 85460 14680
rect 85612 15308 85652 15317
rect 84652 13420 84703 13460
rect 84748 13420 84884 13460
rect 84663 13376 84703 13420
rect 84844 13376 84884 13420
rect 84663 13336 84745 13376
rect 84705 13188 84745 13336
rect 84815 13336 84884 13376
rect 85105 13420 85172 13460
rect 85215 13504 85268 13544
rect 85516 14552 85556 14561
rect 84815 13188 84855 13336
rect 85105 13188 85145 13420
rect 85215 13188 85255 13504
rect 85516 13460 85556 14512
rect 85612 13544 85652 15268
rect 85804 14720 85844 15427
rect 86188 15342 86228 15427
rect 85804 14671 85844 14680
rect 85996 15308 86036 15317
rect 85900 14552 85940 14561
rect 85612 13504 85655 13544
rect 85505 13420 85556 13460
rect 85505 13188 85545 13420
rect 85615 13188 85655 13504
rect 85900 13460 85940 14512
rect 85996 13544 86036 15268
rect 86284 14720 86324 15436
rect 86379 15436 86380 15476
rect 86420 15436 86421 15476
rect 86379 15427 86421 15436
rect 86571 15476 86613 15485
rect 87051 15476 87093 15485
rect 86571 15436 86572 15476
rect 86612 15436 86708 15476
rect 86571 15427 86613 15436
rect 86572 15342 86612 15427
rect 86380 15308 86420 15317
rect 86420 15268 86516 15308
rect 86380 15259 86420 15268
rect 86380 14720 86420 14729
rect 86284 14680 86380 14720
rect 86380 14671 86420 14680
rect 86284 14552 86324 14561
rect 85996 13504 86055 13544
rect 85900 13420 85945 13460
rect 85905 13188 85945 13420
rect 86015 13188 86055 13504
rect 86284 13460 86324 14512
rect 86476 13544 86516 15268
rect 86668 14720 86708 15436
rect 87051 15436 87052 15476
rect 87092 15436 87093 15476
rect 87051 15427 87093 15436
rect 87435 15476 87477 15485
rect 87435 15436 87436 15476
rect 87476 15436 87477 15476
rect 87435 15427 87477 15436
rect 86764 15308 86804 15317
rect 86804 15268 86900 15308
rect 86764 15259 86804 15268
rect 86764 14720 86804 14729
rect 86668 14680 86764 14720
rect 86764 14671 86804 14680
rect 86415 13504 86516 13544
rect 86668 14552 86708 14561
rect 86284 13420 86345 13460
rect 86305 13188 86345 13420
rect 86415 13188 86455 13504
rect 86668 13460 86708 14512
rect 86860 13544 86900 15268
rect 87052 14720 87092 15427
rect 87436 15396 87476 15427
rect 87052 14671 87092 14680
rect 87244 15308 87284 15317
rect 87148 14552 87188 14561
rect 86815 13504 86900 13544
rect 87052 14512 87148 14552
rect 87052 13544 87092 14512
rect 87148 14503 87188 14512
rect 87244 13544 87284 15268
rect 87532 15308 87572 15317
rect 87532 13544 87572 15268
rect 87628 13544 87668 16024
rect 88012 16064 88052 16073
rect 87916 15476 87956 15485
rect 88012 15476 88052 16024
rect 89164 16064 89204 16073
rect 88352 15896 88720 15905
rect 88392 15856 88434 15896
rect 88474 15856 88516 15896
rect 88556 15856 88598 15896
rect 88638 15856 88680 15896
rect 88352 15847 88720 15856
rect 88299 15476 88341 15485
rect 88683 15476 88725 15485
rect 89067 15476 89109 15485
rect 89164 15476 89204 16024
rect 87956 15436 88300 15476
rect 88340 15436 88341 15476
rect 87916 14720 87956 15436
rect 87916 14671 87956 14680
rect 88108 15308 88148 15317
rect 87052 13504 87145 13544
rect 86668 13420 86745 13460
rect 86705 13188 86745 13420
rect 86815 13188 86855 13504
rect 87105 13188 87145 13504
rect 87215 13504 87284 13544
rect 87505 13504 87572 13544
rect 87615 13504 87668 13544
rect 87820 14552 87860 14561
rect 87820 13544 87860 14512
rect 88108 13544 88148 15268
rect 88204 14720 88244 15436
rect 88299 15427 88341 15436
rect 88588 15436 88684 15476
rect 88724 15436 88725 15476
rect 88300 15342 88340 15427
rect 88492 15308 88532 15317
rect 88204 14671 88244 14680
rect 88396 15268 88492 15308
rect 87820 13504 87945 13544
rect 87215 13188 87255 13504
rect 87505 13188 87545 13504
rect 87615 13188 87655 13504
rect 87905 13188 87945 13504
rect 88015 13504 88148 13544
rect 88300 14552 88340 14561
rect 88015 13188 88055 13504
rect 88300 13460 88340 14512
rect 88300 13420 88345 13460
rect 88305 13188 88345 13420
rect 88396 13292 88436 15268
rect 88492 15259 88532 15268
rect 88588 14720 88628 15436
rect 88683 15427 88725 15436
rect 88972 15436 89068 15476
rect 89108 15436 89204 15476
rect 89451 15476 89493 15485
rect 89835 15476 89877 15485
rect 89451 15436 89452 15476
rect 89492 15436 89588 15476
rect 88684 15342 88724 15427
rect 88588 14671 88628 14680
rect 88876 15308 88916 15317
rect 88684 14552 88724 14561
rect 88684 13460 88724 14512
rect 88876 13460 88916 15268
rect 88972 14720 89012 15436
rect 89067 15427 89109 15436
rect 89451 15427 89493 15436
rect 89068 15342 89108 15427
rect 89452 15342 89492 15427
rect 88972 14671 89012 14680
rect 89260 15308 89300 15317
rect 89068 14552 89108 14561
rect 89068 13544 89108 14512
rect 89068 13504 89145 13544
rect 88684 13420 88735 13460
rect 88695 13376 88735 13420
rect 88815 13420 88916 13460
rect 88695 13336 88745 13376
rect 88396 13252 88455 13292
rect 88415 13188 88455 13252
rect 88705 13188 88745 13336
rect 88815 13188 88855 13420
rect 89105 13188 89145 13504
rect 89260 13376 89300 15268
rect 89548 14720 89588 15436
rect 89835 15436 89836 15476
rect 89876 15436 89972 15476
rect 89835 15427 89877 15436
rect 89836 15342 89876 15427
rect 89644 15308 89684 15317
rect 89684 15268 89780 15308
rect 89644 15259 89684 15268
rect 89644 14720 89684 14729
rect 89548 14680 89644 14720
rect 89644 14671 89684 14680
rect 89548 14552 89588 14561
rect 89452 14512 89548 14552
rect 89452 13544 89492 14512
rect 89548 14503 89588 14512
rect 89740 13880 89780 15268
rect 89932 14720 89972 15436
rect 90028 15308 90068 15317
rect 90068 15268 90164 15308
rect 90028 15259 90068 15268
rect 90028 14720 90068 14729
rect 89932 14680 90028 14720
rect 90028 14671 90068 14680
rect 89644 13840 89780 13880
rect 89932 14552 89972 14561
rect 89644 13544 89684 13840
rect 89452 13504 89545 13544
rect 89215 13336 89300 13376
rect 89215 13188 89255 13336
rect 89505 13188 89545 13504
rect 89615 13504 89684 13544
rect 89615 13188 89655 13504
rect 89932 13460 89972 14512
rect 90124 14048 90164 15268
rect 90220 14720 90260 16267
rect 90604 16182 90644 16267
rect 90988 16232 91028 16241
rect 90796 16064 90836 16073
rect 90988 16064 91028 16192
rect 90508 16024 90796 16064
rect 90836 16024 91028 16064
rect 91084 16064 91124 16073
rect 92044 16064 92084 16073
rect 91124 16024 91220 16064
rect 90508 15476 90548 16024
rect 90796 16015 90836 16024
rect 91084 16015 91124 16024
rect 90508 15233 90548 15436
rect 91083 15476 91125 15485
rect 91083 15436 91084 15476
rect 91124 15436 91125 15476
rect 91083 15427 91125 15436
rect 91084 15342 91124 15427
rect 90700 15308 90740 15317
rect 90891 15308 90933 15317
rect 90740 15268 90836 15308
rect 90700 15259 90740 15268
rect 90507 15224 90549 15233
rect 90507 15184 90508 15224
rect 90548 15184 90549 15224
rect 90507 15175 90549 15184
rect 90508 14720 90548 15175
rect 90604 14720 90644 14729
rect 90508 14680 90604 14720
rect 90220 14671 90260 14680
rect 90604 14671 90644 14680
rect 90796 14636 90836 15268
rect 90891 15268 90892 15308
rect 90932 15268 90933 15308
rect 90891 15259 90933 15268
rect 90892 15174 90932 15259
rect 91083 15224 91125 15233
rect 91083 15184 91084 15224
rect 91124 15184 91125 15224
rect 91083 15175 91125 15184
rect 91084 14804 91124 15175
rect 91084 14755 91124 14764
rect 90796 14596 90932 14636
rect 90028 14008 90164 14048
rect 90316 14552 90356 14561
rect 90028 13544 90068 14008
rect 89905 13420 89972 13460
rect 90015 13504 90068 13544
rect 89905 13188 89945 13420
rect 90015 13188 90055 13504
rect 90316 13460 90356 14512
rect 90700 14552 90740 14561
rect 90740 14512 90836 14552
rect 90700 14503 90740 14512
rect 90796 13544 90836 14512
rect 90705 13504 90836 13544
rect 90305 13420 90356 13460
rect 90414 13460 90456 13469
rect 90414 13420 90415 13460
rect 90455 13420 90456 13460
rect 90305 13188 90345 13420
rect 90414 13411 90456 13420
rect 90415 13188 90455 13411
rect 90705 13188 90745 13504
rect 90892 13460 90932 14596
rect 91180 13544 91220 16024
rect 92236 16064 92276 16276
rect 92427 16316 92469 16325
rect 92427 16276 92428 16316
rect 92468 16276 92469 16316
rect 92427 16267 92469 16276
rect 94060 16316 94100 16325
rect 95595 16316 95637 16325
rect 94100 16276 94196 16316
rect 94060 16267 94100 16276
rect 92428 16182 92468 16267
rect 92620 16064 92660 16073
rect 93868 16064 93908 16073
rect 92236 16024 92620 16064
rect 92660 16024 92852 16064
rect 91468 15476 91508 15485
rect 91468 15224 91508 15436
rect 91947 15476 91989 15485
rect 91947 15436 91948 15476
rect 91988 15436 91989 15476
rect 92044 15476 92084 16024
rect 92620 16015 92660 16024
rect 92352 15896 92720 15905
rect 92392 15856 92434 15896
rect 92474 15856 92516 15896
rect 92556 15856 92598 15896
rect 92638 15856 92680 15896
rect 92352 15847 92720 15856
rect 92524 15476 92564 15485
rect 92716 15476 92756 15485
rect 92044 15436 92276 15476
rect 91947 15427 91989 15436
rect 91948 15342 91988 15427
rect 92236 15317 92276 15436
rect 92564 15436 92716 15476
rect 92524 15427 92564 15436
rect 92716 15317 92756 15436
rect 91660 15308 91700 15317
rect 92140 15308 92180 15317
rect 91563 15224 91605 15233
rect 91468 15184 91564 15224
rect 91604 15184 91605 15224
rect 91563 15175 91605 15184
rect 91564 14720 91604 15175
rect 91564 14671 91604 14680
rect 90815 13420 90932 13460
rect 91084 13504 91220 13544
rect 91276 14552 91316 14561
rect 90815 13188 90855 13420
rect 91084 13376 91124 13504
rect 91276 13460 91316 14512
rect 91215 13420 91316 13460
rect 91468 14552 91508 14561
rect 91084 13336 91145 13376
rect 91105 13188 91145 13336
rect 91215 13188 91255 13420
rect 91468 13376 91508 14512
rect 91660 13460 91700 15268
rect 92044 15268 92140 15308
rect 91755 15224 91797 15233
rect 91755 15184 91756 15224
rect 91796 15184 91797 15224
rect 91755 15175 91797 15184
rect 91756 14720 91796 15175
rect 91756 14671 91796 14680
rect 91615 13420 91700 13460
rect 91852 14552 91892 14561
rect 91468 13336 91545 13376
rect 91505 13188 91545 13336
rect 91615 13188 91655 13420
rect 91852 13376 91892 14512
rect 92044 13544 92084 15268
rect 92140 15259 92180 15268
rect 92235 15308 92277 15317
rect 92235 15268 92236 15308
rect 92276 15268 92277 15308
rect 92235 15259 92277 15268
rect 92332 15308 92372 15317
rect 92140 14720 92180 14729
rect 92236 14720 92276 15259
rect 92180 14680 92276 14720
rect 92140 14671 92180 14680
rect 92015 13504 92084 13544
rect 92236 14552 92276 14561
rect 91852 13336 91945 13376
rect 91905 13188 91945 13336
rect 92015 13188 92055 13504
rect 92236 13460 92276 14512
rect 92332 13544 92372 15268
rect 92715 15308 92757 15317
rect 92715 15268 92716 15308
rect 92756 15268 92757 15308
rect 92715 15259 92757 15268
rect 92427 15140 92469 15149
rect 92427 15100 92428 15140
rect 92468 15100 92469 15140
rect 92427 15091 92469 15100
rect 92428 14733 92468 15091
rect 92428 14684 92468 14693
rect 92716 14720 92756 15259
rect 92812 15149 92852 16024
rect 93868 15485 93908 16024
rect 93388 15476 93428 15485
rect 93388 15317 93428 15436
rect 93772 15476 93812 15485
rect 93867 15476 93909 15485
rect 93812 15436 93868 15476
rect 93908 15436 93909 15476
rect 93772 15427 93812 15436
rect 93867 15427 93909 15436
rect 92908 15308 92948 15317
rect 92811 15140 92853 15149
rect 92811 15100 92812 15140
rect 92852 15100 92853 15140
rect 92811 15091 92853 15100
rect 92716 14671 92756 14680
rect 92524 14552 92564 14561
rect 92811 14552 92853 14561
rect 92564 14512 92660 14552
rect 92524 14503 92564 14512
rect 92620 13544 92660 14512
rect 92811 14512 92812 14552
rect 92852 14512 92853 14552
rect 92811 14503 92853 14512
rect 92812 14418 92852 14503
rect 92908 13544 92948 15268
rect 93387 15308 93429 15317
rect 93387 15268 93388 15308
rect 93428 15268 93429 15308
rect 93387 15259 93429 15268
rect 93580 15308 93620 15317
rect 93004 14804 93044 14813
rect 93388 14804 93428 15259
rect 93044 14764 93428 14804
rect 93004 14755 93044 14764
rect 93388 14720 93428 14764
rect 93388 14671 93428 14680
rect 93099 14552 93141 14561
rect 93099 14512 93100 14552
rect 93140 14512 93141 14552
rect 93099 14503 93141 14512
rect 93196 14552 93236 14561
rect 92332 13504 92455 13544
rect 92620 13504 92745 13544
rect 92236 13420 92372 13460
rect 92332 13376 92372 13420
rect 92305 13336 92372 13376
rect 92305 13188 92345 13336
rect 92415 13188 92455 13504
rect 92705 13188 92745 13504
rect 92815 13504 92948 13544
rect 93100 13544 93140 14503
rect 93196 13544 93236 14512
rect 93484 14552 93524 14561
rect 93100 13504 93145 13544
rect 93196 13504 93255 13544
rect 92815 13188 92855 13504
rect 93105 13188 93145 13504
rect 93215 13188 93255 13504
rect 93484 13460 93524 14512
rect 93580 13544 93620 15268
rect 93868 14720 93908 15427
rect 93964 15308 94004 15317
rect 94004 15268 94100 15308
rect 93964 15259 94004 15268
rect 93964 14720 94004 14729
rect 93868 14680 93964 14720
rect 93964 14671 94004 14680
rect 93868 14552 93908 14561
rect 93580 13504 93655 13544
rect 93484 13420 93545 13460
rect 93505 13188 93545 13420
rect 93615 13188 93655 13504
rect 93868 13460 93908 14512
rect 94060 13544 94100 15268
rect 94156 15149 94196 16276
rect 95595 16276 95596 16316
rect 95636 16276 95637 16316
rect 95595 16267 95637 16276
rect 95596 16182 95636 16267
rect 95788 16064 95828 16073
rect 95499 15560 95541 15569
rect 95499 15520 95500 15560
rect 95540 15520 95541 15560
rect 95499 15511 95541 15520
rect 94251 15476 94293 15485
rect 94251 15436 94252 15476
rect 94292 15436 94293 15476
rect 94251 15427 94293 15436
rect 94635 15476 94677 15485
rect 94635 15436 94636 15476
rect 94676 15436 94677 15476
rect 94635 15427 94677 15436
rect 94923 15476 94965 15485
rect 94923 15436 94924 15476
rect 94964 15436 94965 15476
rect 94923 15427 94965 15436
rect 95020 15476 95060 15485
rect 94155 15140 94197 15149
rect 94155 15100 94156 15140
rect 94196 15100 94197 15140
rect 94155 15091 94197 15100
rect 94156 14729 94196 15091
rect 94155 14720 94197 14729
rect 94155 14680 94156 14720
rect 94196 14680 94197 14720
rect 94155 14671 94197 14680
rect 94252 14720 94292 15427
rect 94636 15342 94676 15427
rect 94252 14671 94292 14680
rect 94444 15308 94484 15317
rect 94348 14552 94388 14561
rect 94015 13504 94100 13544
rect 94252 14512 94348 14552
rect 94252 13544 94292 14512
rect 94348 14503 94388 14512
rect 94444 13544 94484 15268
rect 94828 15308 94868 15317
rect 94635 14720 94677 14729
rect 94635 14680 94636 14720
rect 94676 14680 94677 14720
rect 94635 14671 94677 14680
rect 94636 14586 94676 14671
rect 94252 13504 94345 13544
rect 93868 13420 93945 13460
rect 93905 13188 93945 13420
rect 94015 13188 94055 13504
rect 94305 13188 94345 13504
rect 94415 13504 94484 13544
rect 94732 14552 94772 14561
rect 94415 13188 94455 13504
rect 94732 13460 94772 14512
rect 94828 13544 94868 15268
rect 94924 14720 94964 15427
rect 95020 15317 95060 15436
rect 95500 15392 95540 15511
rect 95692 15476 95732 15485
rect 95788 15476 95828 16024
rect 96352 15896 96720 15905
rect 96392 15856 96434 15896
rect 96474 15856 96516 15896
rect 96556 15856 96598 15896
rect 96638 15856 96680 15896
rect 96352 15847 96720 15856
rect 96075 15560 96117 15569
rect 96555 15560 96597 15569
rect 96075 15520 96076 15560
rect 96116 15520 96117 15560
rect 96075 15511 96117 15520
rect 96460 15520 96556 15560
rect 96596 15520 96597 15560
rect 95979 15476 96021 15485
rect 95732 15436 95980 15476
rect 96020 15436 96021 15476
rect 95692 15427 95732 15436
rect 95979 15427 96021 15436
rect 96076 15476 96116 15511
rect 96460 15476 96500 15520
rect 96555 15511 96597 15520
rect 96843 15560 96885 15569
rect 96843 15520 96844 15560
rect 96884 15520 96885 15560
rect 96843 15511 96885 15520
rect 95019 15308 95061 15317
rect 95019 15268 95020 15308
rect 95060 15268 95061 15308
rect 95019 15259 95061 15268
rect 95212 15308 95252 15317
rect 95020 14720 95060 14729
rect 94924 14680 95020 14720
rect 95020 14671 95060 14680
rect 94705 13420 94772 13460
rect 94815 13504 94868 13544
rect 95116 14552 95156 14561
rect 94705 13188 94745 13420
rect 94815 13188 94855 13504
rect 95116 13460 95156 14512
rect 95212 13544 95252 15268
rect 95500 14720 95540 15352
rect 95884 15308 95924 15317
rect 95500 14671 95540 14680
rect 95788 15268 95884 15308
rect 95404 14552 95444 14561
rect 95444 14512 95540 14552
rect 95404 14503 95444 14512
rect 95500 13544 95540 14512
rect 95788 13544 95828 15268
rect 95884 15259 95924 15268
rect 95980 14720 96020 15427
rect 96076 15425 96116 15436
rect 96364 15436 96460 15476
rect 96268 15308 96308 15317
rect 95980 14671 96020 14680
rect 96076 15268 96268 15308
rect 95212 13504 95255 13544
rect 95500 13504 95545 13544
rect 95105 13420 95156 13460
rect 95105 13188 95145 13420
rect 95215 13188 95255 13504
rect 95505 13188 95545 13504
rect 95615 13504 95828 13544
rect 95884 14552 95924 14561
rect 95615 13188 95655 13504
rect 95884 13460 95924 14512
rect 96076 13544 96116 15268
rect 96268 15259 96308 15268
rect 96364 14720 96404 15436
rect 96460 15427 96500 15436
rect 96844 15476 96884 15511
rect 97228 15485 97268 15570
rect 98572 15560 98612 15569
rect 98476 15520 98572 15560
rect 96844 15425 96884 15436
rect 97227 15476 97269 15485
rect 97227 15436 97228 15476
rect 97268 15436 97269 15476
rect 97227 15427 97269 15436
rect 97612 15476 97652 15485
rect 97612 15392 97652 15436
rect 97707 15476 97749 15485
rect 97707 15436 97708 15476
rect 97748 15436 97749 15476
rect 97707 15427 97749 15436
rect 97995 15476 98037 15485
rect 97995 15436 97996 15476
rect 98036 15436 98037 15476
rect 97995 15427 98037 15436
rect 98379 15476 98421 15485
rect 98476 15476 98516 15520
rect 98572 15511 98612 15520
rect 98379 15436 98380 15476
rect 98420 15436 98516 15476
rect 98379 15427 98421 15436
rect 97516 15352 97652 15392
rect 96652 15308 96692 15317
rect 96364 14671 96404 14680
rect 96460 15268 96652 15308
rect 96015 13504 96116 13544
rect 96268 14552 96308 14561
rect 95884 13420 95945 13460
rect 95905 13188 95945 13420
rect 96015 13188 96055 13504
rect 96268 13460 96308 14512
rect 96460 13544 96500 15268
rect 96652 15259 96692 15268
rect 97036 15308 97076 15317
rect 97420 15308 97460 15317
rect 97036 15149 97076 15268
rect 97228 15268 97420 15308
rect 97035 15140 97077 15149
rect 97035 15100 97036 15140
rect 97076 15100 97077 15140
rect 97035 15091 97077 15100
rect 96844 14804 96884 14813
rect 97036 14804 97076 15091
rect 96884 14764 97076 14804
rect 96844 14755 96884 14764
rect 97036 14720 97076 14764
rect 97132 14720 97172 14729
rect 97036 14680 97132 14720
rect 97132 14671 97172 14680
rect 96652 14552 96692 14561
rect 97036 14552 97076 14561
rect 96692 14512 96788 14552
rect 96652 14503 96692 14512
rect 96415 13504 96500 13544
rect 96748 13544 96788 14512
rect 97036 13628 97076 14512
rect 97131 14552 97173 14561
rect 97131 14512 97132 14552
rect 97172 14512 97173 14552
rect 97131 14503 97173 14512
rect 96940 13588 97076 13628
rect 96748 13504 96855 13544
rect 96268 13420 96345 13460
rect 96305 13188 96345 13420
rect 96415 13188 96455 13504
rect 96704 13376 96746 13385
rect 96704 13336 96705 13376
rect 96745 13336 96746 13376
rect 96704 13327 96746 13336
rect 96705 13188 96745 13327
rect 96815 13188 96855 13504
rect 96940 13385 96980 13588
rect 96939 13376 96981 13385
rect 97132 13376 97172 14503
rect 97228 13544 97268 15268
rect 97420 15259 97460 15268
rect 97516 15149 97556 15352
rect 97515 15140 97557 15149
rect 97515 15100 97516 15140
rect 97556 15100 97557 15140
rect 97515 15091 97557 15100
rect 97420 14720 97460 14729
rect 97516 14720 97556 15091
rect 97460 14680 97556 14720
rect 97708 14720 97748 15427
rect 97996 15342 98036 15427
rect 98380 15342 98420 15427
rect 97804 15308 97844 15317
rect 98188 15308 98228 15317
rect 97844 15268 97940 15308
rect 97804 15259 97844 15268
rect 97420 14671 97460 14680
rect 97708 14671 97748 14680
rect 96939 13336 96940 13376
rect 96980 13336 96981 13376
rect 96939 13327 96981 13336
rect 97105 13336 97172 13376
rect 97215 13504 97268 13544
rect 97516 14552 97556 14561
rect 97105 13188 97145 13336
rect 97215 13188 97255 13504
rect 97516 13460 97556 14512
rect 97803 14552 97845 14561
rect 97803 14512 97804 14552
rect 97844 14512 97845 14552
rect 97803 14503 97845 14512
rect 97804 14418 97844 14503
rect 97900 14048 97940 15268
rect 97708 14008 97940 14048
rect 98092 15268 98188 15308
rect 97708 13544 97748 14008
rect 98092 13544 98132 15268
rect 98188 15259 98228 15268
rect 98668 15308 98708 15317
rect 98380 14720 98420 14729
rect 97505 13420 97556 13460
rect 97615 13504 97748 13544
rect 98015 13504 98132 13544
rect 98284 14552 98324 14561
rect 97505 13188 97545 13420
rect 97615 13188 97655 13504
rect 97904 13460 97946 13469
rect 97904 13420 97905 13460
rect 97945 13420 97946 13460
rect 97904 13411 97946 13420
rect 97905 13188 97945 13411
rect 98015 13188 98055 13504
rect 98284 13460 98324 14512
rect 98380 13721 98420 14680
rect 98572 14552 98612 14561
rect 98476 14512 98572 14552
rect 98379 13712 98421 13721
rect 98379 13672 98380 13712
rect 98420 13672 98421 13712
rect 98379 13663 98421 13672
rect 98476 13544 98516 14512
rect 98572 14503 98612 14512
rect 98415 13504 98516 13544
rect 98284 13420 98345 13460
rect 98305 13188 98345 13420
rect 98415 13188 98455 13504
rect 98668 13469 98708 15268
rect 98764 14804 98804 14813
rect 98764 13721 98804 14764
rect 98763 13712 98805 13721
rect 98763 13672 98764 13712
rect 98804 13672 98900 13712
rect 98763 13663 98805 13672
rect 98667 13460 98709 13469
rect 98667 13420 98668 13460
rect 98708 13420 98709 13460
rect 98667 13411 98709 13420
rect 72305 7841 72345 8064
rect 72415 7841 72455 8064
rect 72705 7925 72745 8064
rect 72704 7916 72746 7925
rect 72704 7876 72705 7916
rect 72745 7876 72746 7916
rect 72704 7867 72746 7876
rect 72304 7832 72346 7841
rect 72304 7792 72305 7832
rect 72345 7792 72346 7832
rect 72304 7783 72346 7792
rect 72414 7832 72456 7841
rect 72414 7792 72415 7832
rect 72455 7792 72456 7832
rect 72414 7783 72456 7792
rect 72815 7664 72855 8064
rect 72172 7624 72855 7664
rect 73105 7664 73145 8064
rect 73215 7664 73255 8064
rect 73505 7664 73545 8064
rect 73105 7624 73172 7664
rect 73215 7624 73364 7664
rect 71444 7372 71540 7412
rect 71787 7412 71829 7421
rect 71787 7372 71788 7412
rect 71828 7372 71829 7412
rect 71404 7363 71444 7372
rect 71787 7363 71829 7372
rect 72172 7412 72212 7624
rect 73132 7505 73172 7624
rect 72555 7496 72597 7505
rect 72555 7456 72556 7496
rect 72596 7456 72597 7496
rect 72555 7447 72597 7456
rect 73131 7496 73173 7505
rect 73131 7456 73132 7496
rect 73172 7456 73173 7496
rect 73131 7447 73173 7456
rect 72172 7363 72212 7372
rect 72556 7412 72596 7447
rect 72556 7361 72596 7372
rect 73324 7412 73364 7624
rect 73324 7363 73364 7372
rect 73420 7624 73545 7664
rect 73615 7664 73655 8064
rect 73905 7664 73945 8064
rect 74015 7664 74055 8064
rect 74305 7664 74345 8064
rect 73615 7624 73748 7664
rect 73132 7328 73172 7337
rect 72364 7244 72404 7255
rect 72364 7169 72404 7204
rect 72940 7244 72980 7255
rect 73132 7244 73172 7288
rect 73420 7244 73460 7624
rect 73708 7412 73748 7624
rect 73708 7363 73748 7372
rect 73804 7624 73945 7664
rect 73996 7624 74055 7664
rect 74188 7624 74345 7664
rect 74415 7664 74455 8064
rect 74705 7664 74745 8064
rect 74415 7624 74516 7664
rect 73132 7204 73460 7244
rect 72940 7169 72980 7204
rect 71308 7111 71348 7120
rect 72075 7160 72117 7169
rect 72075 7120 72076 7160
rect 72116 7120 72117 7160
rect 72075 7111 72117 7120
rect 72363 7160 72405 7169
rect 72363 7120 72364 7160
rect 72404 7120 72405 7160
rect 72363 7111 72405 7120
rect 72939 7160 72981 7169
rect 73611 7160 73653 7169
rect 72939 7120 72940 7160
rect 72980 7120 72981 7160
rect 72939 7111 72981 7120
rect 73433 7149 73612 7160
rect 72076 7026 72116 7111
rect 73473 7120 73612 7149
rect 73652 7120 73653 7160
rect 73611 7111 73653 7120
rect 73433 7100 73473 7109
rect 73227 7076 73269 7085
rect 73227 7036 73228 7076
rect 73268 7036 73269 7076
rect 73227 7027 73269 7036
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 8352 6824 8720 6833
rect 8392 6784 8434 6824
rect 8474 6784 8516 6824
rect 8556 6784 8598 6824
rect 8638 6784 8680 6824
rect 8352 6775 8720 6784
rect 12352 6824 12720 6833
rect 12392 6784 12434 6824
rect 12474 6784 12516 6824
rect 12556 6784 12598 6824
rect 12638 6784 12680 6824
rect 12352 6775 12720 6784
rect 16352 6824 16720 6833
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16352 6775 16720 6784
rect 20352 6824 20720 6833
rect 20392 6784 20434 6824
rect 20474 6784 20516 6824
rect 20556 6784 20598 6824
rect 20638 6784 20680 6824
rect 20352 6775 20720 6784
rect 24352 6824 24720 6833
rect 24392 6784 24434 6824
rect 24474 6784 24516 6824
rect 24556 6784 24598 6824
rect 24638 6784 24680 6824
rect 24352 6775 24720 6784
rect 28352 6824 28720 6833
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28352 6775 28720 6784
rect 32352 6824 32720 6833
rect 32392 6784 32434 6824
rect 32474 6784 32516 6824
rect 32556 6784 32598 6824
rect 32638 6784 32680 6824
rect 32352 6775 32720 6784
rect 36352 6824 36720 6833
rect 36392 6784 36434 6824
rect 36474 6784 36516 6824
rect 36556 6784 36598 6824
rect 36638 6784 36680 6824
rect 36352 6775 36720 6784
rect 40352 6824 40720 6833
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40352 6775 40720 6784
rect 44352 6824 44720 6833
rect 44392 6784 44434 6824
rect 44474 6784 44516 6824
rect 44556 6784 44598 6824
rect 44638 6784 44680 6824
rect 44352 6775 44720 6784
rect 48352 6824 48720 6833
rect 48392 6784 48434 6824
rect 48474 6784 48516 6824
rect 48556 6784 48598 6824
rect 48638 6784 48680 6824
rect 48352 6775 48720 6784
rect 52352 6824 52720 6833
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52352 6775 52720 6784
rect 56352 6824 56720 6833
rect 56392 6784 56434 6824
rect 56474 6784 56516 6824
rect 56556 6784 56598 6824
rect 56638 6784 56680 6824
rect 56352 6775 56720 6784
rect 60352 6824 60720 6833
rect 60392 6784 60434 6824
rect 60474 6784 60516 6824
rect 60556 6784 60598 6824
rect 60638 6784 60680 6824
rect 60352 6775 60720 6784
rect 64352 6824 64720 6833
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64352 6775 64720 6784
rect 68352 6824 68720 6833
rect 68392 6784 68434 6824
rect 68474 6784 68516 6824
rect 68556 6784 68598 6824
rect 68638 6784 68680 6824
rect 68352 6775 68720 6784
rect 1707 6656 1749 6665
rect 1707 6616 1708 6656
rect 1748 6616 1749 6656
rect 1707 6607 1749 6616
rect 1708 6522 1748 6607
rect 73228 6488 73268 7027
rect 73612 7026 73652 7111
rect 73708 6656 73748 6665
rect 73804 6656 73844 7624
rect 73996 6740 74036 7624
rect 74091 6992 74133 7001
rect 74091 6952 74092 6992
rect 74132 6952 74133 6992
rect 74091 6943 74133 6952
rect 74092 6858 74132 6943
rect 73748 6616 73844 6656
rect 73900 6700 74036 6740
rect 73708 6607 73748 6616
rect 73324 6572 73364 6581
rect 73364 6532 73652 6572
rect 73324 6523 73364 6532
rect 73612 6488 73652 6532
rect 73900 6488 73940 6700
rect 74188 6656 74228 7624
rect 74283 7328 74325 7337
rect 74283 7288 74284 7328
rect 74324 7288 74325 7328
rect 74283 7279 74325 7288
rect 74284 7244 74324 7279
rect 74476 7253 74516 7624
rect 74572 7624 74745 7664
rect 74815 7664 74855 8064
rect 75105 7664 75145 8064
rect 74815 7624 74900 7664
rect 74284 6992 74324 7204
rect 74475 7244 74517 7253
rect 74475 7204 74476 7244
rect 74516 7204 74517 7244
rect 74475 7195 74517 7204
rect 74476 6992 74516 7001
rect 74284 6952 74476 6992
rect 74476 6943 74516 6952
rect 74188 6607 74228 6616
rect 74572 6656 74612 7624
rect 74860 7421 74900 7624
rect 75052 7624 75145 7664
rect 75215 7664 75255 8064
rect 75505 7664 75545 8064
rect 75615 7673 75655 8064
rect 75215 7624 75284 7664
rect 74667 7412 74709 7421
rect 74667 7372 74668 7412
rect 74708 7372 74709 7412
rect 74667 7363 74709 7372
rect 74859 7412 74901 7421
rect 74859 7372 74860 7412
rect 74900 7372 74901 7412
rect 74859 7363 74901 7372
rect 74668 7244 74708 7363
rect 74668 7195 74708 7204
rect 74859 7244 74901 7253
rect 74859 7204 74860 7244
rect 74900 7204 74901 7244
rect 74859 7195 74901 7204
rect 74860 7110 74900 7195
rect 74956 7160 74996 7169
rect 74956 7001 74996 7120
rect 74955 6992 74997 7001
rect 74572 6607 74612 6616
rect 74860 6952 74956 6992
rect 74996 6952 74997 6992
rect 73612 6448 73940 6488
rect 1900 6404 1940 6413
rect 1556 6364 1900 6404
rect 73228 6404 73268 6448
rect 73996 6413 74036 6498
rect 74380 6413 74420 6498
rect 74860 6413 74900 6952
rect 74955 6943 74997 6952
rect 75052 6656 75092 7624
rect 75244 7505 75284 7624
rect 75436 7624 75545 7664
rect 75614 7664 75656 7673
rect 75905 7664 75945 8064
rect 75614 7624 75615 7664
rect 75655 7624 75656 7664
rect 75243 7496 75285 7505
rect 75243 7456 75244 7496
rect 75284 7456 75285 7496
rect 75243 7447 75285 7456
rect 75147 7412 75189 7421
rect 75147 7372 75148 7412
rect 75188 7372 75189 7412
rect 75147 7363 75189 7372
rect 75148 7278 75188 7363
rect 75244 7160 75284 7169
rect 75244 7001 75284 7120
rect 75243 6992 75285 7001
rect 75243 6952 75244 6992
rect 75284 6952 75285 6992
rect 75243 6943 75285 6952
rect 75052 6607 75092 6616
rect 73516 6404 73556 6413
rect 73228 6364 73516 6404
rect 1324 6320 1364 6329
rect 1516 6320 1556 6364
rect 1900 6355 1940 6364
rect 73516 6355 73556 6364
rect 73995 6404 74037 6413
rect 73995 6364 73996 6404
rect 74036 6364 74037 6404
rect 73995 6355 74037 6364
rect 74379 6404 74421 6413
rect 74379 6364 74380 6404
rect 74420 6364 74421 6404
rect 74379 6355 74421 6364
rect 74859 6404 74901 6413
rect 74859 6364 74860 6404
rect 74900 6364 74901 6404
rect 74859 6355 74901 6364
rect 75244 6404 75284 6943
rect 75436 6656 75476 7624
rect 75614 7615 75656 7624
rect 75820 7624 75945 7664
rect 76015 7664 76055 8064
rect 76203 7664 76245 7673
rect 76015 7624 76148 7664
rect 75531 7328 75573 7337
rect 75531 7288 75532 7328
rect 75572 7288 75573 7328
rect 75531 7279 75573 7288
rect 75532 7244 75572 7279
rect 75532 7193 75572 7204
rect 75723 7160 75765 7169
rect 75723 7120 75724 7160
rect 75764 7120 75765 7160
rect 75723 7111 75765 7120
rect 75436 6607 75476 6616
rect 75724 6992 75764 7111
rect 75244 6355 75284 6364
rect 75628 6404 75668 6413
rect 75724 6404 75764 6952
rect 75820 6656 75860 7624
rect 75915 7496 75957 7505
rect 75915 7456 75916 7496
rect 75956 7456 75957 7496
rect 75915 7447 75957 7456
rect 75916 7412 75956 7447
rect 75916 7361 75956 7372
rect 76108 7253 76148 7624
rect 76203 7624 76204 7664
rect 76244 7624 76245 7664
rect 76305 7664 76345 8064
rect 76415 7748 76455 8064
rect 76415 7708 76532 7748
rect 76305 7624 76436 7664
rect 76203 7615 76245 7624
rect 76204 7412 76244 7615
rect 76204 7363 76244 7372
rect 76107 7244 76149 7253
rect 76107 7204 76108 7244
rect 76148 7204 76149 7244
rect 76107 7195 76149 7204
rect 76012 7160 76052 7169
rect 76012 7001 76052 7120
rect 76299 7160 76341 7169
rect 76299 7120 76300 7160
rect 76340 7120 76341 7160
rect 76299 7111 76341 7120
rect 76300 7026 76340 7111
rect 76011 6992 76053 7001
rect 76011 6952 76012 6992
rect 76052 6952 76053 6992
rect 76011 6943 76053 6952
rect 75820 6607 75860 6616
rect 76204 6656 76244 6665
rect 76396 6656 76436 7624
rect 76492 7421 76532 7708
rect 76705 7664 76745 8064
rect 76684 7624 76745 7664
rect 76491 7412 76533 7421
rect 76491 7372 76492 7412
rect 76532 7372 76533 7412
rect 76491 7363 76533 7372
rect 76491 7244 76533 7253
rect 76491 7204 76492 7244
rect 76532 7204 76533 7244
rect 76491 7195 76533 7204
rect 76492 7110 76532 7195
rect 76587 7160 76629 7169
rect 76587 7120 76588 7160
rect 76628 7120 76629 7160
rect 76587 7111 76629 7120
rect 76588 7026 76628 7111
rect 76491 6992 76533 7001
rect 76491 6952 76492 6992
rect 76532 6952 76533 6992
rect 76491 6943 76533 6952
rect 76244 6616 76436 6656
rect 76204 6607 76244 6616
rect 76012 6404 76052 6413
rect 75668 6364 76012 6404
rect 75628 6355 75668 6364
rect 76012 6355 76052 6364
rect 76492 6404 76532 6943
rect 76684 6656 76724 7624
rect 76815 7580 76855 8064
rect 77105 7664 77145 8064
rect 77068 7624 77145 7664
rect 77215 7664 77255 8064
rect 77505 7664 77545 8064
rect 77215 7624 77300 7664
rect 76815 7540 76916 7580
rect 76779 7412 76821 7421
rect 76779 7372 76780 7412
rect 76820 7372 76821 7412
rect 76779 7363 76821 7372
rect 76780 7278 76820 7363
rect 76876 7337 76916 7540
rect 76875 7328 76917 7337
rect 76875 7288 76876 7328
rect 76916 7288 76917 7328
rect 76875 7279 76917 7288
rect 76875 7160 76917 7169
rect 76875 7120 76876 7160
rect 76916 7120 76917 7160
rect 76875 7111 76917 7120
rect 76876 7026 76916 7111
rect 76684 6607 76724 6616
rect 77068 6656 77108 7624
rect 77260 7421 77300 7624
rect 77452 7624 77545 7664
rect 77615 7664 77655 8064
rect 77905 7664 77945 8064
rect 77615 7624 77684 7664
rect 77259 7412 77301 7421
rect 77259 7372 77260 7412
rect 77300 7372 77301 7412
rect 77259 7363 77301 7372
rect 77355 7244 77397 7253
rect 77355 7204 77356 7244
rect 77396 7204 77397 7244
rect 77355 7195 77397 7204
rect 77356 7110 77396 7195
rect 77164 6992 77204 7001
rect 77204 6952 77300 6992
rect 77164 6943 77204 6952
rect 77068 6607 77108 6616
rect 76876 6413 76916 6498
rect 77260 6413 77300 6952
rect 77452 6656 77492 7624
rect 77644 7505 77684 7624
rect 77740 7624 77945 7664
rect 78015 7664 78055 8064
rect 78305 7664 78345 8064
rect 78415 7673 78455 8064
rect 78414 7664 78456 7673
rect 78705 7664 78745 8064
rect 78815 7664 78855 8064
rect 79105 7664 79145 8064
rect 79215 7832 79255 8064
rect 78015 7624 78068 7664
rect 78305 7624 78356 7664
rect 77643 7496 77685 7505
rect 77643 7456 77644 7496
rect 77684 7456 77685 7496
rect 77643 7447 77685 7456
rect 77643 7328 77685 7337
rect 77643 7288 77644 7328
rect 77684 7288 77685 7328
rect 77643 7279 77685 7288
rect 77644 7194 77684 7279
rect 77547 7160 77589 7169
rect 77547 7120 77548 7160
rect 77588 7120 77589 7160
rect 77547 7111 77589 7120
rect 77548 7026 77588 7111
rect 77740 6656 77780 7624
rect 78028 7421 78068 7624
rect 78123 7496 78165 7505
rect 78123 7456 78124 7496
rect 78164 7456 78165 7496
rect 78123 7447 78165 7456
rect 77835 7412 77877 7421
rect 77835 7372 77836 7412
rect 77876 7372 77877 7412
rect 77835 7363 77877 7372
rect 78027 7412 78069 7421
rect 78027 7372 78028 7412
rect 78068 7372 78069 7412
rect 78027 7363 78069 7372
rect 78124 7412 78164 7447
rect 77836 7278 77876 7363
rect 78124 7361 78164 7372
rect 77931 7160 77973 7169
rect 77931 7120 77932 7160
rect 77972 7120 77973 7160
rect 77931 7111 77973 7120
rect 78219 7160 78261 7169
rect 78219 7120 78220 7160
rect 78260 7120 78261 7160
rect 78219 7111 78261 7120
rect 77932 7026 77972 7111
rect 77836 6656 77876 6665
rect 77740 6616 77836 6656
rect 77452 6607 77492 6616
rect 77836 6607 77876 6616
rect 77644 6413 77684 6498
rect 78124 6413 78164 6498
rect 76492 6355 76532 6364
rect 76875 6404 76917 6413
rect 76875 6364 76876 6404
rect 76916 6364 76917 6404
rect 76875 6355 76917 6364
rect 77259 6404 77301 6413
rect 77259 6364 77260 6404
rect 77300 6364 77301 6404
rect 77259 6355 77301 6364
rect 77643 6404 77685 6413
rect 77643 6364 77644 6404
rect 77684 6364 77685 6404
rect 77643 6355 77685 6364
rect 78123 6404 78165 6413
rect 78220 6404 78260 7111
rect 78316 6656 78356 7624
rect 78414 7624 78415 7664
rect 78455 7624 78456 7664
rect 78414 7615 78456 7624
rect 78700 7624 78745 7664
rect 78796 7624 78855 7664
rect 79084 7624 79145 7664
rect 79188 7792 79255 7832
rect 78411 7412 78453 7421
rect 78411 7372 78412 7412
rect 78452 7372 78453 7412
rect 78411 7363 78453 7372
rect 78412 7278 78452 7363
rect 78507 7160 78549 7169
rect 78507 7120 78508 7160
rect 78548 7120 78549 7160
rect 78507 7111 78549 7120
rect 78508 7026 78548 7111
rect 78316 6607 78356 6616
rect 78700 6656 78740 7624
rect 78796 7421 78836 7624
rect 78795 7412 78837 7421
rect 78795 7372 78796 7412
rect 78836 7372 78837 7412
rect 78795 7363 78837 7372
rect 78795 7244 78837 7253
rect 78795 7204 78796 7244
rect 78836 7204 78837 7244
rect 78795 7195 78837 7204
rect 78796 7110 78836 7195
rect 78987 6992 79029 7001
rect 78987 6952 78988 6992
rect 79028 6952 79029 6992
rect 78987 6943 79029 6952
rect 78988 6858 79028 6943
rect 78700 6607 78740 6616
rect 79084 6656 79124 7624
rect 79188 7580 79228 7792
rect 79275 7664 79317 7673
rect 79505 7664 79545 8064
rect 79275 7624 79276 7664
rect 79316 7624 79317 7664
rect 79275 7615 79317 7624
rect 79372 7624 79545 7664
rect 79615 7664 79655 8064
rect 79905 7664 79945 8064
rect 79615 7624 79700 7664
rect 79180 7540 79228 7580
rect 79180 7337 79220 7540
rect 79276 7412 79316 7615
rect 79276 7363 79316 7372
rect 79179 7328 79221 7337
rect 79179 7288 79180 7328
rect 79220 7288 79221 7328
rect 79179 7279 79221 7288
rect 79179 7160 79221 7169
rect 79179 7120 79180 7160
rect 79220 7120 79221 7160
rect 79179 7111 79221 7120
rect 79180 7026 79220 7111
rect 79372 6656 79412 7624
rect 79467 7412 79509 7421
rect 79467 7372 79468 7412
rect 79508 7372 79509 7412
rect 79467 7363 79509 7372
rect 79468 7278 79508 7363
rect 79564 7160 79604 7169
rect 79564 7001 79604 7120
rect 79563 6992 79605 7001
rect 79563 6952 79564 6992
rect 79604 6952 79605 6992
rect 79563 6943 79605 6952
rect 79660 6917 79700 7624
rect 79852 7624 79945 7664
rect 80015 7664 80055 8064
rect 80305 7664 80345 8064
rect 80015 7624 80084 7664
rect 79756 7253 79796 7338
rect 79755 7244 79797 7253
rect 79755 7204 79756 7244
rect 79796 7204 79797 7244
rect 79755 7195 79797 7204
rect 79755 6992 79797 7001
rect 79755 6952 79756 6992
rect 79796 6952 79797 6992
rect 79755 6943 79797 6952
rect 79659 6908 79701 6917
rect 79659 6868 79660 6908
rect 79700 6868 79701 6908
rect 79659 6859 79701 6868
rect 79468 6656 79508 6665
rect 79372 6616 79468 6656
rect 79084 6607 79124 6616
rect 79468 6607 79508 6616
rect 78508 6413 78548 6498
rect 78892 6413 78932 6498
rect 79276 6413 79316 6498
rect 79756 6413 79796 6943
rect 79852 6656 79892 7624
rect 80044 7421 80084 7624
rect 80236 7624 80345 7664
rect 80415 7664 80455 8064
rect 80705 7664 80745 8064
rect 80815 7664 80855 8064
rect 81105 7664 81145 8064
rect 81215 7664 81255 8064
rect 81505 7664 81545 8064
rect 80415 7624 80468 7664
rect 80705 7624 80756 7664
rect 80815 7624 80948 7664
rect 80043 7412 80085 7421
rect 80043 7372 80044 7412
rect 80084 7372 80085 7412
rect 80043 7363 80085 7372
rect 80140 7328 80180 7339
rect 80140 7253 80180 7288
rect 80139 7244 80181 7253
rect 80139 7204 80140 7244
rect 80180 7204 80181 7244
rect 80139 7195 80181 7204
rect 79948 6992 79988 7001
rect 79988 6952 80084 6992
rect 79948 6943 79988 6952
rect 79948 6656 79988 6665
rect 79852 6616 79948 6656
rect 79948 6607 79988 6616
rect 78123 6364 78124 6404
rect 78164 6364 78260 6404
rect 78507 6404 78549 6413
rect 78507 6364 78508 6404
rect 78548 6364 78549 6404
rect 78123 6355 78165 6364
rect 78507 6355 78549 6364
rect 78891 6404 78933 6413
rect 78891 6364 78892 6404
rect 78932 6364 78933 6404
rect 78891 6355 78933 6364
rect 79275 6404 79317 6413
rect 79275 6364 79276 6404
rect 79316 6364 79317 6404
rect 79275 6355 79317 6364
rect 79755 6404 79797 6413
rect 79755 6364 79756 6404
rect 79796 6364 79797 6404
rect 80044 6404 80084 6952
rect 80236 6656 80276 7624
rect 80331 7496 80373 7505
rect 80331 7456 80332 7496
rect 80372 7456 80373 7496
rect 80331 7447 80373 7456
rect 80332 7244 80372 7447
rect 80332 7195 80372 7204
rect 80428 6665 80468 7624
rect 80523 7328 80565 7337
rect 80523 7288 80524 7328
rect 80564 7288 80565 7328
rect 80523 7279 80565 7288
rect 80524 7194 80564 7279
rect 80620 7160 80660 7169
rect 80620 7001 80660 7120
rect 80619 6992 80661 7001
rect 80619 6952 80620 6992
rect 80660 6952 80661 6992
rect 80619 6943 80661 6952
rect 80332 6656 80372 6665
rect 80236 6616 80332 6656
rect 80332 6607 80372 6616
rect 80427 6656 80469 6665
rect 80427 6616 80428 6656
rect 80468 6616 80469 6656
rect 80427 6607 80469 6616
rect 80716 6656 80756 7624
rect 80908 7169 80948 7624
rect 81004 7624 81145 7664
rect 81196 7624 81255 7664
rect 81484 7624 81545 7664
rect 81615 7664 81655 8064
rect 81905 7664 81945 8064
rect 82015 7748 82055 8064
rect 82015 7708 82100 7748
rect 81615 7624 81716 7664
rect 81905 7624 82004 7664
rect 80812 7160 80852 7169
rect 80812 7001 80852 7120
rect 80907 7160 80949 7169
rect 80907 7120 80908 7160
rect 80948 7120 80949 7160
rect 80907 7111 80949 7120
rect 80811 6992 80853 7001
rect 80811 6952 80812 6992
rect 80852 6952 80853 6992
rect 80811 6943 80853 6952
rect 80908 6992 80948 7003
rect 80908 6917 80948 6952
rect 80907 6908 80949 6917
rect 80907 6868 80908 6908
rect 80948 6868 80949 6908
rect 80907 6859 80949 6868
rect 81004 6824 81044 7624
rect 81196 7505 81236 7624
rect 81195 7496 81237 7505
rect 81195 7456 81196 7496
rect 81236 7456 81237 7496
rect 81195 7447 81237 7456
rect 81099 7412 81141 7421
rect 81099 7372 81100 7412
rect 81140 7372 81141 7412
rect 81099 7363 81141 7372
rect 81100 7278 81140 7363
rect 81195 7160 81237 7169
rect 81195 7120 81196 7160
rect 81236 7120 81237 7160
rect 81195 7111 81237 7120
rect 81004 6784 81140 6824
rect 80716 6607 80756 6616
rect 80907 6656 80949 6665
rect 80907 6616 80908 6656
rect 80948 6616 80949 6656
rect 80907 6607 80949 6616
rect 80908 6522 80948 6607
rect 80140 6413 80180 6498
rect 80524 6413 80564 6498
rect 81004 6488 81044 6499
rect 81004 6413 81044 6448
rect 80139 6404 80181 6413
rect 80044 6364 80140 6404
rect 80180 6364 80181 6404
rect 79755 6355 79797 6364
rect 80139 6355 80181 6364
rect 80523 6404 80565 6413
rect 80523 6364 80524 6404
rect 80564 6364 80565 6404
rect 80523 6355 80565 6364
rect 81003 6404 81045 6413
rect 81003 6364 81004 6404
rect 81044 6364 81045 6404
rect 81003 6355 81045 6364
rect 844 6280 1324 6320
rect 844 5732 884 6280
rect 1324 6271 1364 6280
rect 1420 6280 1556 6320
rect 844 5683 884 5692
rect 651 5648 693 5657
rect 651 5608 652 5648
rect 692 5608 693 5648
rect 651 5599 693 5608
rect 652 5480 692 5599
rect 652 5431 692 5440
rect 1420 4901 1460 6280
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 7112 6068 7480 6077
rect 7152 6028 7194 6068
rect 7234 6028 7276 6068
rect 7316 6028 7358 6068
rect 7398 6028 7440 6068
rect 7112 6019 7480 6028
rect 11112 6068 11480 6077
rect 11152 6028 11194 6068
rect 11234 6028 11276 6068
rect 11316 6028 11358 6068
rect 11398 6028 11440 6068
rect 11112 6019 11480 6028
rect 15112 6068 15480 6077
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15112 6019 15480 6028
rect 19112 6068 19480 6077
rect 19152 6028 19194 6068
rect 19234 6028 19276 6068
rect 19316 6028 19358 6068
rect 19398 6028 19440 6068
rect 19112 6019 19480 6028
rect 23112 6068 23480 6077
rect 23152 6028 23194 6068
rect 23234 6028 23276 6068
rect 23316 6028 23358 6068
rect 23398 6028 23440 6068
rect 23112 6019 23480 6028
rect 27112 6068 27480 6077
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27112 6019 27480 6028
rect 31112 6068 31480 6077
rect 31152 6028 31194 6068
rect 31234 6028 31276 6068
rect 31316 6028 31358 6068
rect 31398 6028 31440 6068
rect 31112 6019 31480 6028
rect 35112 6068 35480 6077
rect 35152 6028 35194 6068
rect 35234 6028 35276 6068
rect 35316 6028 35358 6068
rect 35398 6028 35440 6068
rect 35112 6019 35480 6028
rect 39112 6068 39480 6077
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39112 6019 39480 6028
rect 43112 6068 43480 6077
rect 43152 6028 43194 6068
rect 43234 6028 43276 6068
rect 43316 6028 43358 6068
rect 43398 6028 43440 6068
rect 43112 6019 43480 6028
rect 47112 6068 47480 6077
rect 47152 6028 47194 6068
rect 47234 6028 47276 6068
rect 47316 6028 47358 6068
rect 47398 6028 47440 6068
rect 47112 6019 47480 6028
rect 51112 6068 51480 6077
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51112 6019 51480 6028
rect 55112 6068 55480 6077
rect 55152 6028 55194 6068
rect 55234 6028 55276 6068
rect 55316 6028 55358 6068
rect 55398 6028 55440 6068
rect 55112 6019 55480 6028
rect 59112 6068 59480 6077
rect 59152 6028 59194 6068
rect 59234 6028 59276 6068
rect 59316 6028 59358 6068
rect 59398 6028 59440 6068
rect 59112 6019 59480 6028
rect 63112 6068 63480 6077
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63112 6019 63480 6028
rect 67112 6068 67480 6077
rect 67152 6028 67194 6068
rect 67234 6028 67276 6068
rect 67316 6028 67358 6068
rect 67398 6028 67440 6068
rect 67112 6019 67480 6028
rect 80908 5732 80948 5741
rect 81004 5732 81044 6355
rect 81100 5900 81140 6784
rect 81196 6413 81236 7111
rect 81484 6656 81524 7624
rect 81676 7421 81716 7624
rect 81675 7412 81717 7421
rect 81675 7372 81676 7412
rect 81716 7372 81717 7412
rect 81675 7363 81717 7372
rect 81579 7244 81621 7253
rect 81579 7204 81580 7244
rect 81620 7204 81621 7244
rect 81579 7195 81621 7204
rect 81580 7110 81620 7195
rect 81964 7160 82004 7624
rect 82060 7589 82100 7708
rect 82305 7664 82345 8064
rect 82156 7624 82345 7664
rect 82415 7664 82455 8064
rect 82705 7664 82745 8064
rect 82815 7916 82855 8064
rect 82815 7876 82964 7916
rect 82415 7624 82484 7664
rect 82705 7624 82772 7664
rect 82059 7580 82101 7589
rect 82059 7540 82060 7580
rect 82100 7540 82101 7580
rect 82059 7531 82101 7540
rect 81868 7120 82004 7160
rect 82059 7160 82101 7169
rect 82059 7120 82060 7160
rect 82100 7120 82101 7160
rect 81484 6607 81524 6616
rect 81772 6992 81812 7001
rect 81195 6404 81237 6413
rect 81292 6404 81332 6432
rect 81195 6364 81196 6404
rect 81236 6364 81292 6404
rect 81195 6355 81237 6364
rect 81292 6355 81332 6364
rect 81676 6404 81716 6432
rect 81772 6413 81812 6952
rect 81868 6656 81908 7120
rect 82059 7111 82101 7120
rect 82060 7026 82100 7111
rect 81963 6992 82005 7001
rect 81963 6952 81964 6992
rect 82004 6952 82005 6992
rect 81963 6943 82005 6952
rect 81964 6858 82004 6943
rect 82156 6656 82196 7624
rect 82347 7496 82389 7505
rect 82347 7456 82348 7496
rect 82388 7456 82389 7496
rect 82347 7447 82389 7456
rect 82348 7412 82388 7447
rect 82348 7361 82388 7372
rect 82444 7337 82484 7624
rect 82539 7412 82581 7421
rect 82539 7372 82540 7412
rect 82580 7372 82581 7412
rect 82539 7363 82581 7372
rect 82443 7328 82485 7337
rect 82443 7288 82444 7328
rect 82484 7288 82485 7328
rect 82443 7279 82485 7288
rect 82540 7278 82580 7363
rect 82251 7160 82293 7169
rect 82251 7120 82252 7160
rect 82292 7120 82293 7160
rect 82251 7111 82293 7120
rect 82635 7160 82677 7169
rect 82635 7120 82636 7160
rect 82676 7120 82677 7160
rect 82635 7111 82677 7120
rect 82252 7026 82292 7111
rect 82252 6656 82292 6665
rect 82156 6616 82252 6656
rect 81868 6607 81908 6616
rect 82252 6607 82292 6616
rect 82060 6413 82100 6498
rect 82540 6413 82580 6498
rect 81771 6404 81813 6413
rect 81716 6364 81772 6404
rect 81812 6364 81813 6404
rect 81676 6355 81716 6364
rect 81771 6355 81813 6364
rect 82059 6404 82101 6413
rect 82059 6364 82060 6404
rect 82100 6364 82101 6404
rect 82059 6355 82101 6364
rect 82539 6404 82581 6413
rect 82636 6404 82676 7111
rect 82732 6656 82772 7624
rect 82827 7580 82869 7589
rect 82827 7540 82828 7580
rect 82868 7540 82869 7580
rect 82827 7531 82869 7540
rect 82828 7412 82868 7531
rect 82924 7505 82964 7876
rect 83105 7664 83145 8064
rect 83215 7664 83255 8064
rect 83505 7664 83545 8064
rect 83615 7673 83655 8064
rect 83105 7624 83156 7664
rect 83215 7624 83348 7664
rect 82923 7496 82965 7505
rect 82923 7456 82924 7496
rect 82964 7456 82965 7496
rect 82923 7447 82965 7456
rect 82828 7363 82868 7372
rect 82923 7160 82965 7169
rect 82923 7120 82924 7160
rect 82964 7120 82965 7160
rect 82923 7111 82965 7120
rect 82732 6607 82772 6616
rect 82539 6364 82540 6404
rect 82580 6364 82676 6404
rect 82924 6404 82964 7111
rect 83116 6656 83156 7624
rect 83211 7244 83253 7253
rect 83211 7204 83212 7244
rect 83252 7204 83253 7244
rect 83211 7195 83253 7204
rect 83212 7110 83252 7195
rect 83116 6607 83156 6616
rect 83308 6656 83348 7624
rect 83500 7624 83545 7664
rect 83614 7664 83656 7673
rect 83905 7664 83945 8064
rect 83614 7624 83615 7664
rect 83655 7624 83656 7664
rect 83308 6607 83348 6616
rect 83404 6992 83444 7001
rect 83404 6488 83444 6952
rect 83404 6413 83444 6448
rect 83403 6404 83445 6413
rect 82539 6355 82581 6364
rect 82924 6355 82964 6364
rect 83308 6364 83404 6404
rect 83444 6364 83445 6404
rect 81100 5851 81140 5860
rect 80948 5692 81044 5732
rect 83308 5732 83348 6364
rect 83403 6355 83445 6364
rect 83500 5900 83540 7624
rect 83614 7615 83656 7624
rect 83788 7624 83945 7664
rect 84015 7664 84055 8064
rect 84171 7664 84213 7673
rect 84015 7624 84116 7664
rect 83595 7328 83637 7337
rect 83595 7288 83596 7328
rect 83636 7288 83637 7328
rect 83595 7279 83637 7288
rect 83596 7194 83636 7279
rect 83691 7160 83733 7169
rect 83691 7120 83692 7160
rect 83732 7120 83733 7160
rect 83691 7111 83733 7120
rect 83692 7026 83732 7111
rect 83788 6656 83828 7624
rect 83979 7496 84021 7505
rect 83979 7456 83980 7496
rect 84020 7456 84021 7496
rect 83979 7447 84021 7456
rect 83980 7412 84020 7447
rect 84076 7421 84116 7624
rect 84171 7624 84172 7664
rect 84212 7624 84213 7664
rect 84305 7664 84345 8064
rect 84415 7841 84455 8064
rect 84414 7832 84456 7841
rect 84414 7792 84415 7832
rect 84455 7792 84456 7832
rect 84414 7783 84456 7792
rect 84705 7664 84745 8064
rect 84305 7624 84404 7664
rect 84171 7615 84213 7624
rect 83980 7361 84020 7372
rect 84075 7412 84117 7421
rect 84075 7372 84076 7412
rect 84116 7372 84117 7412
rect 84075 7363 84117 7372
rect 84172 7412 84212 7615
rect 84172 7363 84212 7372
rect 83883 7160 83925 7169
rect 83883 7120 83884 7160
rect 83924 7120 83925 7160
rect 83883 7111 83925 7120
rect 84268 7160 84308 7169
rect 83884 7026 83924 7111
rect 84268 7001 84308 7120
rect 84267 6992 84309 7001
rect 84267 6952 84268 6992
rect 84308 6952 84309 6992
rect 84267 6943 84309 6952
rect 83884 6656 83924 6665
rect 83788 6616 83884 6656
rect 83884 6607 83924 6616
rect 84268 6656 84308 6665
rect 84364 6656 84404 7624
rect 84652 7624 84745 7664
rect 84815 7664 84855 8064
rect 85105 7664 85145 8064
rect 85215 7748 85255 8064
rect 85323 7832 85365 7841
rect 85323 7792 85324 7832
rect 85364 7792 85365 7832
rect 85323 7783 85365 7792
rect 85215 7708 85268 7748
rect 84815 7624 84884 7664
rect 85105 7624 85172 7664
rect 84459 7412 84501 7421
rect 84459 7372 84460 7412
rect 84500 7372 84501 7412
rect 84459 7363 84501 7372
rect 84460 7278 84500 7363
rect 84556 7160 84596 7169
rect 84556 7001 84596 7120
rect 84555 6992 84597 7001
rect 84555 6952 84556 6992
rect 84596 6952 84597 6992
rect 84555 6943 84597 6952
rect 84308 6616 84404 6656
rect 84268 6607 84308 6616
rect 83692 6413 83732 6498
rect 84076 6413 84116 6498
rect 84460 6413 84500 6498
rect 83691 6404 83733 6413
rect 83691 6364 83692 6404
rect 83732 6364 83733 6404
rect 83691 6355 83733 6364
rect 84075 6404 84117 6413
rect 84075 6364 84076 6404
rect 84116 6364 84117 6404
rect 84075 6355 84117 6364
rect 84459 6404 84501 6413
rect 84556 6404 84596 6943
rect 84652 6656 84692 7624
rect 84844 7505 84884 7624
rect 84843 7496 84885 7505
rect 84843 7456 84844 7496
rect 84884 7456 84885 7496
rect 84843 7447 84885 7456
rect 84843 7244 84885 7253
rect 84843 7204 84844 7244
rect 84884 7204 84885 7244
rect 84843 7195 84885 7204
rect 84844 7110 84884 7195
rect 85035 7160 85077 7169
rect 85035 7120 85036 7160
rect 85076 7120 85077 7160
rect 85035 7111 85077 7120
rect 85036 6992 85076 7111
rect 85036 6943 85076 6952
rect 84652 6607 84692 6616
rect 85036 6656 85076 6665
rect 85132 6656 85172 7624
rect 85228 7421 85268 7708
rect 85227 7412 85269 7421
rect 85227 7372 85228 7412
rect 85268 7372 85269 7412
rect 85227 7363 85269 7372
rect 85324 7412 85364 7783
rect 85505 7664 85545 8064
rect 85615 7664 85655 8064
rect 85324 7363 85364 7372
rect 85420 7624 85545 7664
rect 85612 7624 85655 7664
rect 85905 7664 85945 8064
rect 86015 7748 86055 8064
rect 86015 7708 86228 7748
rect 85905 7624 86036 7664
rect 85228 7160 85268 7169
rect 85228 7001 85268 7120
rect 85227 6992 85269 7001
rect 85227 6952 85228 6992
rect 85268 6952 85269 6992
rect 85227 6943 85269 6952
rect 85076 6616 85172 6656
rect 85420 6656 85460 7624
rect 85515 7496 85557 7505
rect 85515 7456 85516 7496
rect 85556 7456 85557 7496
rect 85515 7447 85557 7456
rect 85516 7412 85556 7447
rect 85516 7361 85556 7372
rect 85612 7328 85652 7624
rect 85803 7412 85845 7421
rect 85803 7372 85804 7412
rect 85844 7372 85845 7412
rect 85803 7363 85845 7372
rect 85707 7328 85749 7337
rect 85612 7288 85708 7328
rect 85748 7288 85749 7328
rect 85707 7279 85749 7288
rect 85804 7278 85844 7363
rect 85611 7160 85653 7169
rect 85611 7120 85612 7160
rect 85652 7120 85653 7160
rect 85611 7111 85653 7120
rect 85899 7160 85941 7169
rect 85899 7120 85900 7160
rect 85940 7120 85941 7160
rect 85899 7111 85941 7120
rect 85516 6656 85556 6665
rect 85420 6616 85516 6656
rect 85036 6607 85076 6616
rect 85516 6607 85556 6616
rect 84844 6413 84884 6498
rect 85324 6413 85364 6498
rect 84459 6364 84460 6404
rect 84500 6364 84596 6404
rect 84843 6404 84885 6413
rect 84843 6364 84844 6404
rect 84884 6364 84885 6404
rect 84459 6355 84501 6364
rect 84843 6355 84885 6364
rect 85323 6404 85365 6413
rect 85612 6404 85652 7111
rect 85900 7026 85940 7111
rect 85900 6656 85940 6665
rect 85996 6656 86036 7624
rect 86188 7085 86228 7708
rect 86305 7664 86345 8064
rect 86415 7748 86455 8064
rect 86415 7708 86516 7748
rect 86305 7624 86420 7664
rect 86283 7244 86325 7253
rect 86283 7204 86284 7244
rect 86324 7204 86325 7244
rect 86283 7195 86325 7204
rect 86284 7110 86324 7195
rect 86187 7076 86229 7085
rect 86187 7036 86188 7076
rect 86228 7036 86229 7076
rect 86187 7027 86229 7036
rect 85940 6616 86036 6656
rect 86092 6992 86132 7001
rect 85900 6607 85940 6616
rect 86092 6413 86132 6952
rect 86284 6656 86324 6665
rect 86380 6656 86420 7624
rect 86476 7421 86516 7708
rect 86705 7664 86745 8064
rect 86815 7748 86855 8064
rect 86815 7708 86900 7748
rect 86705 7624 86804 7664
rect 86667 7496 86709 7505
rect 86667 7456 86668 7496
rect 86708 7456 86709 7496
rect 86667 7447 86709 7456
rect 86475 7412 86517 7421
rect 86475 7372 86476 7412
rect 86516 7372 86517 7412
rect 86475 7363 86517 7372
rect 86475 7244 86517 7253
rect 86475 7204 86476 7244
rect 86516 7204 86517 7244
rect 86475 7195 86517 7204
rect 86668 7244 86708 7447
rect 86476 6992 86516 7195
rect 86476 6943 86516 6952
rect 86668 6917 86708 7204
rect 86667 6908 86709 6917
rect 86667 6868 86668 6908
rect 86708 6868 86709 6908
rect 86667 6859 86709 6868
rect 86324 6616 86420 6656
rect 86668 6656 86708 6665
rect 86764 6656 86804 7624
rect 86860 7505 86900 7708
rect 87105 7664 87145 8064
rect 87052 7624 87145 7664
rect 87215 7664 87255 8064
rect 87505 7664 87545 8064
rect 87615 7748 87655 8064
rect 87615 7708 87860 7748
rect 87215 7624 87284 7664
rect 87505 7624 87668 7664
rect 86859 7496 86901 7505
rect 86859 7456 86860 7496
rect 86900 7456 86901 7496
rect 86859 7447 86901 7456
rect 86859 7328 86901 7337
rect 86859 7288 86860 7328
rect 86900 7288 86901 7328
rect 86859 7279 86901 7288
rect 86860 7194 86900 7279
rect 86955 7160 86997 7169
rect 86955 7120 86956 7160
rect 86996 7120 86997 7160
rect 86955 7111 86997 7120
rect 86956 7026 86996 7111
rect 86708 6616 86804 6656
rect 87052 6656 87092 7624
rect 87244 7337 87284 7624
rect 87435 7412 87477 7421
rect 87435 7372 87436 7412
rect 87476 7372 87477 7412
rect 87435 7363 87477 7372
rect 87243 7328 87285 7337
rect 87243 7288 87244 7328
rect 87284 7288 87285 7328
rect 87243 7279 87285 7288
rect 87436 7278 87476 7363
rect 87147 7160 87189 7169
rect 87147 7120 87148 7160
rect 87188 7120 87189 7160
rect 87147 7111 87189 7120
rect 87339 7160 87381 7169
rect 87339 7120 87340 7160
rect 87380 7120 87381 7160
rect 87339 7111 87381 7120
rect 87531 7160 87573 7169
rect 87531 7120 87532 7160
rect 87572 7120 87573 7160
rect 87531 7111 87573 7120
rect 87148 7026 87188 7111
rect 87243 7076 87285 7085
rect 87243 7036 87244 7076
rect 87284 7036 87285 7076
rect 87243 7027 87285 7036
rect 87244 6942 87284 7027
rect 86284 6607 86324 6616
rect 86668 6607 86708 6616
rect 87052 6607 87092 6616
rect 86476 6413 86516 6498
rect 86860 6413 86900 6498
rect 87340 6413 87380 7111
rect 87532 7026 87572 7111
rect 87532 6656 87572 6665
rect 87628 6656 87668 7624
rect 87820 7589 87860 7708
rect 87905 7664 87945 8064
rect 88015 7664 88055 8064
rect 88305 7664 88345 8064
rect 88415 7664 88455 8064
rect 88705 7664 88745 8064
rect 88815 7748 88855 8064
rect 88815 7708 88916 7748
rect 87905 7624 87956 7664
rect 87819 7580 87861 7589
rect 87819 7540 87820 7580
rect 87860 7540 87861 7580
rect 87819 7531 87861 7540
rect 87723 7496 87765 7505
rect 87723 7456 87724 7496
rect 87764 7456 87765 7496
rect 87723 7447 87765 7456
rect 87724 7412 87764 7447
rect 87724 7361 87764 7372
rect 87819 7160 87861 7169
rect 87819 7120 87820 7160
rect 87860 7120 87861 7160
rect 87819 7111 87861 7120
rect 87820 7026 87860 7111
rect 87572 6616 87668 6656
rect 87724 6656 87764 6665
rect 87916 6656 87956 7624
rect 88012 7624 88055 7664
rect 88300 7624 88345 7664
rect 88396 7624 88455 7664
rect 88588 7624 88745 7664
rect 88012 7421 88052 7624
rect 88011 7412 88053 7421
rect 88011 7372 88012 7412
rect 88052 7372 88053 7412
rect 88011 7363 88053 7372
rect 88203 7244 88245 7253
rect 88203 7204 88204 7244
rect 88244 7204 88245 7244
rect 88203 7195 88245 7204
rect 88204 7110 88244 7195
rect 88012 6992 88052 7001
rect 88052 6952 88148 6992
rect 88012 6943 88052 6952
rect 87764 6616 87956 6656
rect 87532 6607 87572 6616
rect 87724 6607 87764 6616
rect 87916 6413 87956 6498
rect 88108 6413 88148 6952
rect 88300 6656 88340 7624
rect 88396 7505 88436 7624
rect 88395 7496 88437 7505
rect 88395 7456 88396 7496
rect 88436 7456 88437 7496
rect 88395 7447 88437 7456
rect 88395 7328 88437 7337
rect 88395 7288 88396 7328
rect 88436 7288 88437 7328
rect 88395 7279 88437 7288
rect 88396 7194 88436 7279
rect 88491 7160 88533 7169
rect 88491 7120 88492 7160
rect 88532 7120 88533 7160
rect 88491 7111 88533 7120
rect 88492 7026 88532 7111
rect 88588 6656 88628 7624
rect 88779 7580 88821 7589
rect 88779 7540 88780 7580
rect 88820 7540 88821 7580
rect 88779 7531 88821 7540
rect 88780 7412 88820 7531
rect 88780 7363 88820 7372
rect 88876 7337 88916 7708
rect 89105 7664 89145 8064
rect 89215 7748 89255 8064
rect 89215 7708 89300 7748
rect 89105 7624 89204 7664
rect 88971 7412 89013 7421
rect 88971 7372 88972 7412
rect 89012 7372 89013 7412
rect 88971 7363 89013 7372
rect 88875 7328 88917 7337
rect 88875 7288 88876 7328
rect 88916 7288 88917 7328
rect 88875 7279 88917 7288
rect 88972 7278 89012 7363
rect 88683 7160 88725 7169
rect 88683 7120 88684 7160
rect 88724 7120 88725 7160
rect 88683 7111 88725 7120
rect 88875 7160 88917 7169
rect 88875 7120 88876 7160
rect 88916 7120 88917 7160
rect 88875 7111 88917 7120
rect 89067 7160 89109 7169
rect 89067 7120 89068 7160
rect 89108 7120 89109 7160
rect 89067 7111 89109 7120
rect 88684 7026 88724 7111
rect 88684 6656 88724 6665
rect 88588 6616 88684 6656
rect 88300 6607 88340 6616
rect 88684 6607 88724 6616
rect 88492 6413 88532 6498
rect 88876 6413 88916 7111
rect 89068 7026 89108 7111
rect 89068 6656 89108 6665
rect 89164 6656 89204 7624
rect 89260 7421 89300 7708
rect 89505 7664 89545 8064
rect 89615 7757 89655 8064
rect 89614 7748 89656 7757
rect 89614 7708 89615 7748
rect 89655 7708 89656 7748
rect 89614 7699 89656 7708
rect 89905 7664 89945 8064
rect 89505 7624 89588 7664
rect 89259 7412 89301 7421
rect 89259 7372 89260 7412
rect 89300 7372 89301 7412
rect 89259 7363 89301 7372
rect 89259 7244 89301 7253
rect 89259 7204 89260 7244
rect 89300 7204 89301 7244
rect 89259 7195 89301 7204
rect 89260 7110 89300 7195
rect 89451 7076 89493 7085
rect 89451 7036 89452 7076
rect 89492 7036 89493 7076
rect 89451 7027 89493 7036
rect 89452 6992 89492 7027
rect 89452 6941 89492 6952
rect 89108 6616 89204 6656
rect 89452 6656 89492 6665
rect 89548 6656 89588 7624
rect 89836 7624 89945 7664
rect 90015 7664 90055 8064
rect 90305 7664 90345 8064
rect 90415 7916 90455 8064
rect 90415 7876 90644 7916
rect 90507 7748 90549 7757
rect 90507 7708 90508 7748
rect 90548 7708 90549 7748
rect 90507 7699 90549 7708
rect 90015 7624 90068 7664
rect 90305 7624 90452 7664
rect 89643 7496 89685 7505
rect 89643 7456 89644 7496
rect 89684 7456 89685 7496
rect 89643 7447 89685 7456
rect 89644 7412 89684 7447
rect 89644 7361 89684 7372
rect 89739 7160 89781 7169
rect 89739 7120 89740 7160
rect 89780 7120 89781 7160
rect 89739 7111 89781 7120
rect 89740 7026 89780 7111
rect 89492 6616 89588 6656
rect 89836 6656 89876 7624
rect 90028 7505 90068 7624
rect 90027 7496 90069 7505
rect 90027 7456 90028 7496
rect 90068 7456 90069 7496
rect 90027 7447 90069 7456
rect 90219 7412 90261 7421
rect 90219 7372 90220 7412
rect 90260 7372 90261 7412
rect 90219 7363 90261 7372
rect 90027 7328 90069 7337
rect 90027 7288 90028 7328
rect 90068 7288 90069 7328
rect 90027 7279 90069 7288
rect 90028 7194 90068 7279
rect 90220 7278 90260 7363
rect 89931 7160 89973 7169
rect 89931 7120 89932 7160
rect 89972 7120 89973 7160
rect 89931 7111 89973 7120
rect 90315 7160 90357 7169
rect 90315 7120 90316 7160
rect 90356 7120 90357 7160
rect 90315 7111 90357 7120
rect 89932 7026 89972 7111
rect 90316 7026 90356 7111
rect 89932 6656 89972 6665
rect 89836 6616 89932 6656
rect 89068 6607 89108 6616
rect 89452 6607 89492 6616
rect 89932 6607 89972 6616
rect 90316 6656 90356 6665
rect 90412 6656 90452 7624
rect 90508 7412 90548 7699
rect 90604 7421 90644 7876
rect 90508 7363 90548 7372
rect 90603 7412 90645 7421
rect 90705 7412 90745 8064
rect 90815 7673 90855 8064
rect 90987 7748 91029 7757
rect 90987 7708 90988 7748
rect 91028 7708 91029 7748
rect 90987 7699 91029 7708
rect 90814 7664 90856 7673
rect 90814 7624 90815 7664
rect 90855 7624 90856 7664
rect 90814 7615 90856 7624
rect 90603 7372 90604 7412
rect 90644 7372 90645 7412
rect 90603 7363 90645 7372
rect 90700 7372 90745 7412
rect 90603 7160 90645 7169
rect 90603 7120 90604 7160
rect 90644 7120 90645 7160
rect 90603 7111 90645 7120
rect 90356 6616 90452 6656
rect 90316 6607 90356 6616
rect 89260 6413 89300 6498
rect 89740 6413 89780 6498
rect 90124 6413 90164 6498
rect 90508 6413 90548 6498
rect 85708 6404 85748 6413
rect 85323 6364 85324 6404
rect 85364 6364 85708 6404
rect 85323 6355 85365 6364
rect 85708 6336 85748 6364
rect 86091 6404 86133 6413
rect 86091 6364 86092 6404
rect 86132 6364 86133 6404
rect 86091 6355 86133 6364
rect 86475 6404 86517 6413
rect 86475 6364 86476 6404
rect 86516 6364 86517 6404
rect 86475 6355 86517 6364
rect 86859 6404 86901 6413
rect 86859 6364 86860 6404
rect 86900 6364 86901 6404
rect 86859 6355 86901 6364
rect 87339 6404 87381 6413
rect 87339 6364 87340 6404
rect 87380 6364 87381 6404
rect 87339 6355 87381 6364
rect 87915 6404 87957 6413
rect 87915 6364 87916 6404
rect 87956 6364 87957 6404
rect 87915 6355 87957 6364
rect 88107 6404 88149 6413
rect 88107 6364 88108 6404
rect 88148 6364 88149 6404
rect 88107 6355 88149 6364
rect 88491 6404 88533 6413
rect 88491 6364 88492 6404
rect 88532 6364 88533 6404
rect 88491 6355 88533 6364
rect 88875 6404 88917 6413
rect 88875 6364 88876 6404
rect 88916 6364 88917 6404
rect 88875 6355 88917 6364
rect 89259 6404 89301 6413
rect 89259 6364 89260 6404
rect 89300 6364 89301 6404
rect 89259 6355 89301 6364
rect 89739 6404 89781 6413
rect 89739 6364 89740 6404
rect 89780 6364 89781 6404
rect 89739 6355 89781 6364
rect 90123 6404 90165 6413
rect 90123 6364 90124 6404
rect 90164 6364 90165 6404
rect 90123 6355 90165 6364
rect 90507 6404 90549 6413
rect 90604 6404 90644 7111
rect 90700 6656 90740 7372
rect 90988 7253 91028 7699
rect 91105 7664 91145 8064
rect 91215 7757 91255 8064
rect 91214 7748 91256 7757
rect 91214 7708 91215 7748
rect 91255 7708 91256 7748
rect 91214 7699 91256 7708
rect 91505 7664 91545 8064
rect 91084 7624 91145 7664
rect 91372 7624 91545 7664
rect 91615 7664 91655 8064
rect 91755 7664 91797 7673
rect 91615 7624 91700 7664
rect 90795 7244 90837 7253
rect 90795 7204 90796 7244
rect 90836 7204 90837 7244
rect 90795 7195 90837 7204
rect 90987 7244 91029 7253
rect 90987 7204 90988 7244
rect 91028 7204 91029 7244
rect 90987 7195 91029 7204
rect 90796 7110 90836 7195
rect 90700 6607 90740 6616
rect 90988 6992 91028 7001
rect 90507 6364 90508 6404
rect 90548 6364 90644 6404
rect 90892 6404 90932 6432
rect 90988 6413 91028 6952
rect 91084 6656 91124 7624
rect 91180 7412 91220 7421
rect 91275 7412 91317 7421
rect 91220 7372 91276 7412
rect 91316 7372 91317 7412
rect 91180 7363 91220 7372
rect 91275 7363 91317 7372
rect 91179 7244 91221 7253
rect 91179 7204 91180 7244
rect 91220 7204 91221 7244
rect 91179 7195 91221 7204
rect 91084 6607 91124 6616
rect 90987 6404 91029 6413
rect 90932 6364 90988 6404
rect 91028 6364 91029 6404
rect 90507 6355 90549 6364
rect 90892 6355 90932 6364
rect 90987 6355 91029 6364
rect 83500 5851 83540 5860
rect 80908 5683 80948 5692
rect 83308 5683 83348 5692
rect 90988 5648 91028 6355
rect 91180 5900 91220 7195
rect 91275 7160 91317 7169
rect 91275 7120 91276 7160
rect 91316 7120 91317 7160
rect 91275 7111 91317 7120
rect 91276 7026 91316 7111
rect 91372 6656 91412 7624
rect 91563 7328 91605 7337
rect 91563 7288 91564 7328
rect 91604 7288 91605 7328
rect 91563 7279 91605 7288
rect 91564 7194 91604 7279
rect 91660 7253 91700 7624
rect 91755 7624 91756 7664
rect 91796 7624 91797 7664
rect 91905 7664 91945 8064
rect 92015 7748 92055 8064
rect 92015 7708 92084 7748
rect 91905 7624 91988 7664
rect 91755 7615 91797 7624
rect 91756 7412 91796 7615
rect 91756 7363 91796 7372
rect 91851 7328 91893 7337
rect 91851 7288 91852 7328
rect 91892 7288 91893 7328
rect 91851 7279 91893 7288
rect 91659 7244 91701 7253
rect 91659 7204 91660 7244
rect 91700 7204 91701 7244
rect 91659 7195 91701 7204
rect 91467 7160 91509 7169
rect 91467 7120 91468 7160
rect 91508 7120 91509 7160
rect 91467 7111 91509 7120
rect 91852 7160 91892 7279
rect 91468 7026 91508 7111
rect 91468 6656 91508 6665
rect 91372 6616 91468 6656
rect 91468 6607 91508 6616
rect 91275 6404 91317 6413
rect 91275 6364 91276 6404
rect 91316 6364 91317 6404
rect 91275 6355 91317 6364
rect 91755 6404 91797 6413
rect 91852 6404 91892 7120
rect 91755 6364 91756 6404
rect 91796 6364 91892 6404
rect 91755 6355 91797 6364
rect 91276 6270 91316 6355
rect 91756 6270 91796 6355
rect 91948 6320 91988 7624
rect 92044 7001 92084 7708
rect 92305 7664 92345 8064
rect 92236 7624 92345 7664
rect 92415 7664 92455 8064
rect 92705 7664 92745 8064
rect 92815 7664 92855 8064
rect 93105 7664 93145 8064
rect 92415 7624 92468 7664
rect 92043 6992 92085 7001
rect 92043 6952 92044 6992
rect 92084 6952 92085 6992
rect 92043 6943 92085 6952
rect 92140 6992 92180 7001
rect 92140 6413 92180 6952
rect 92236 6656 92276 7624
rect 92428 7505 92468 7624
rect 92620 7624 92745 7664
rect 92812 7624 92855 7664
rect 93100 7624 93145 7664
rect 92427 7496 92469 7505
rect 92427 7456 92428 7496
rect 92468 7456 92469 7496
rect 92427 7447 92469 7456
rect 92332 7244 92372 7253
rect 92332 7085 92372 7204
rect 92331 7076 92373 7085
rect 92331 7036 92332 7076
rect 92372 7036 92373 7076
rect 92331 7027 92373 7036
rect 92523 7076 92565 7085
rect 92523 7036 92524 7076
rect 92564 7036 92565 7076
rect 92523 7027 92565 7036
rect 92524 6992 92564 7027
rect 92524 6941 92564 6952
rect 92332 6656 92372 6665
rect 92236 6616 92332 6656
rect 92620 6656 92660 7624
rect 92812 7421 92852 7624
rect 92811 7412 92853 7421
rect 92811 7372 92812 7412
rect 92852 7372 92853 7412
rect 92811 7363 92853 7372
rect 93003 7328 93045 7337
rect 93003 7288 93004 7328
rect 93044 7288 93045 7328
rect 93003 7279 93045 7288
rect 92716 7244 92756 7253
rect 92716 6917 92756 7204
rect 92907 7244 92949 7253
rect 92907 7204 92908 7244
rect 92948 7204 92949 7244
rect 92907 7195 92949 7204
rect 92908 7110 92948 7195
rect 93004 7160 93044 7279
rect 93004 7111 93044 7120
rect 92715 6908 92757 6917
rect 92715 6868 92716 6908
rect 92756 6868 92757 6908
rect 92715 6859 92757 6868
rect 92716 6656 92756 6665
rect 92620 6616 92716 6656
rect 92332 6607 92372 6616
rect 92716 6607 92756 6616
rect 93100 6656 93140 7624
rect 93215 7580 93255 8064
rect 93505 7664 93545 8064
rect 93615 7748 93655 8064
rect 93905 7841 93945 8064
rect 93904 7832 93946 7841
rect 93904 7792 93905 7832
rect 93945 7792 93946 7832
rect 93904 7783 93946 7792
rect 93615 7708 93812 7748
rect 93505 7624 93716 7664
rect 93215 7540 93332 7580
rect 93195 7328 93237 7337
rect 93195 7288 93196 7328
rect 93236 7288 93237 7328
rect 93195 7279 93237 7288
rect 93196 7160 93236 7279
rect 93292 7169 93332 7540
rect 93483 7496 93525 7505
rect 93483 7456 93484 7496
rect 93524 7456 93525 7496
rect 93483 7447 93525 7456
rect 93484 7412 93524 7447
rect 93484 7361 93524 7372
rect 93579 7328 93621 7337
rect 93579 7288 93580 7328
rect 93620 7288 93621 7328
rect 93579 7279 93621 7288
rect 93196 7111 93236 7120
rect 93291 7160 93333 7169
rect 93580 7160 93620 7279
rect 93291 7120 93292 7160
rect 93332 7120 93333 7160
rect 93291 7111 93333 7120
rect 93388 7120 93580 7160
rect 93291 6992 93333 7001
rect 93291 6952 93292 6992
rect 93332 6952 93333 6992
rect 93291 6943 93333 6952
rect 93292 6858 93332 6943
rect 93100 6607 93140 6616
rect 93388 6413 93428 7120
rect 93580 7111 93620 7120
rect 93580 6656 93620 6665
rect 93676 6656 93716 7624
rect 93772 7589 93812 7708
rect 94015 7664 94055 8064
rect 93964 7624 94055 7664
rect 94305 7664 94345 8064
rect 94415 7748 94455 8064
rect 94415 7708 94484 7748
rect 94305 7624 94388 7664
rect 93771 7580 93813 7589
rect 93771 7540 93772 7580
rect 93812 7540 93813 7580
rect 93771 7531 93813 7540
rect 93771 7412 93813 7421
rect 93771 7372 93772 7412
rect 93812 7372 93813 7412
rect 93771 7363 93813 7372
rect 93772 7278 93812 7363
rect 93867 7328 93909 7337
rect 93867 7288 93868 7328
rect 93908 7288 93909 7328
rect 93867 7279 93909 7288
rect 93868 7160 93908 7279
rect 93868 7111 93908 7120
rect 93964 6740 94004 7624
rect 94252 7244 94292 7253
rect 94252 7085 94292 7204
rect 94251 7076 94293 7085
rect 94251 7036 94252 7076
rect 94292 7036 94293 7076
rect 94251 7027 94293 7036
rect 94060 6992 94100 7001
rect 94100 6952 94196 6992
rect 94060 6943 94100 6952
rect 93964 6700 94100 6740
rect 93620 6616 93716 6656
rect 93771 6656 93813 6665
rect 93771 6616 93772 6656
rect 93812 6616 93813 6656
rect 93580 6607 93620 6616
rect 93771 6607 93813 6616
rect 93772 6522 93812 6607
rect 93963 6488 94005 6497
rect 93963 6448 93964 6488
rect 94004 6448 94005 6488
rect 93963 6439 94005 6448
rect 92139 6404 92181 6413
rect 92139 6364 92140 6404
rect 92180 6364 92181 6404
rect 92139 6355 92181 6364
rect 92523 6404 92565 6413
rect 92523 6364 92524 6404
rect 92564 6364 92565 6404
rect 92523 6355 92565 6364
rect 92907 6404 92949 6413
rect 92907 6364 92908 6404
rect 92948 6364 92949 6404
rect 92907 6355 92949 6364
rect 93387 6404 93429 6413
rect 93387 6364 93388 6404
rect 93428 6364 93429 6404
rect 93387 6355 93429 6364
rect 93964 6404 94004 6439
rect 91948 6271 91988 6280
rect 92140 6270 92180 6355
rect 92524 6270 92564 6355
rect 92908 6270 92948 6355
rect 93388 6270 93428 6355
rect 91180 5851 91220 5860
rect 91084 5648 91124 5657
rect 90988 5608 91084 5648
rect 91084 5599 91124 5608
rect 93964 5648 94004 6364
rect 94060 5900 94100 6700
rect 94156 6497 94196 6952
rect 94252 6917 94292 7027
rect 94251 6908 94293 6917
rect 94251 6868 94252 6908
rect 94292 6868 94293 6908
rect 94251 6859 94293 6868
rect 94348 6656 94388 7624
rect 94444 7253 94484 7708
rect 94705 7664 94745 8064
rect 94636 7624 94745 7664
rect 94815 7664 94855 8064
rect 95105 7664 95145 8064
rect 95215 7664 95255 8064
rect 95505 7664 95545 8064
rect 95615 7664 95655 8064
rect 94815 7624 94868 7664
rect 95105 7624 95156 7664
rect 95215 7624 95348 7664
rect 94539 7328 94581 7337
rect 94539 7288 94540 7328
rect 94580 7288 94581 7328
rect 94539 7279 94581 7288
rect 94443 7244 94485 7253
rect 94443 7204 94444 7244
rect 94484 7204 94485 7244
rect 94443 7195 94485 7204
rect 94540 7169 94580 7279
rect 94539 7160 94581 7169
rect 94539 7120 94540 7160
rect 94580 7120 94581 7160
rect 94539 7111 94581 7120
rect 94443 7076 94485 7085
rect 94443 7036 94444 7076
rect 94484 7036 94485 7076
rect 94443 7027 94485 7036
rect 94444 6942 94484 7027
rect 94540 7026 94580 7111
rect 94636 6656 94676 7624
rect 94828 7337 94868 7624
rect 94923 7580 94965 7589
rect 94923 7540 94924 7580
rect 94964 7540 94965 7580
rect 94923 7531 94965 7540
rect 94827 7328 94869 7337
rect 94827 7288 94828 7328
rect 94868 7288 94869 7328
rect 94827 7279 94869 7288
rect 94731 7160 94773 7169
rect 94731 7120 94732 7160
rect 94772 7120 94773 7160
rect 94731 7111 94773 7120
rect 94828 7160 94868 7169
rect 94924 7160 94964 7531
rect 94868 7120 94964 7160
rect 94828 7111 94868 7120
rect 94732 7026 94772 7111
rect 94732 6656 94772 6665
rect 94636 6616 94732 6656
rect 94348 6607 94388 6616
rect 94732 6607 94772 6616
rect 95116 6656 95156 7624
rect 95212 7244 95252 7253
rect 95212 6917 95252 7204
rect 95308 7169 95348 7624
rect 95500 7624 95545 7664
rect 95596 7624 95655 7664
rect 95905 7664 95945 8064
rect 96015 7748 96055 8064
rect 96015 7708 96212 7748
rect 95905 7624 96116 7664
rect 95307 7160 95349 7169
rect 95307 7120 95308 7160
rect 95348 7120 95349 7160
rect 95307 7111 95349 7120
rect 95404 6992 95444 7001
rect 95211 6908 95253 6917
rect 95211 6868 95212 6908
rect 95252 6868 95253 6908
rect 95211 6859 95253 6868
rect 95116 6607 95156 6616
rect 94155 6488 94197 6497
rect 94155 6448 94156 6488
rect 94196 6448 94197 6488
rect 94155 6439 94197 6448
rect 94539 6488 94581 6497
rect 94539 6448 94540 6488
rect 94580 6448 94581 6488
rect 94539 6439 94581 6448
rect 94923 6488 94965 6497
rect 94923 6448 94924 6488
rect 94964 6448 94965 6488
rect 94923 6439 94965 6448
rect 94156 6404 94196 6439
rect 94156 6353 94196 6364
rect 94540 6404 94580 6439
rect 94540 6353 94580 6364
rect 94924 6404 94964 6439
rect 95404 6413 95444 6952
rect 95500 6656 95540 7624
rect 95596 7421 95636 7624
rect 95595 7412 95637 7421
rect 95595 7372 95596 7412
rect 95636 7372 95637 7412
rect 95595 7363 95637 7372
rect 95979 7328 96021 7337
rect 95979 7288 95980 7328
rect 96020 7288 96021 7328
rect 95979 7279 96021 7288
rect 95595 7244 95637 7253
rect 95595 7204 95596 7244
rect 95636 7204 95637 7244
rect 95595 7195 95637 7204
rect 95596 7110 95636 7195
rect 95980 7194 96020 7279
rect 95692 7160 95732 7169
rect 95884 7160 95924 7169
rect 95732 7120 95884 7160
rect 95596 6656 95636 6665
rect 95500 6616 95596 6656
rect 95596 6607 95636 6616
rect 95692 6497 95732 7120
rect 95884 7111 95924 7120
rect 95980 6656 96020 6665
rect 96076 6656 96116 7624
rect 96172 7580 96212 7708
rect 96305 7664 96345 8064
rect 96415 7748 96455 8064
rect 96415 7708 96596 7748
rect 96305 7624 96404 7664
rect 96172 7540 96308 7580
rect 96172 7253 96212 7338
rect 96268 7337 96308 7540
rect 96267 7328 96309 7337
rect 96267 7288 96268 7328
rect 96308 7288 96309 7328
rect 96267 7279 96309 7288
rect 96171 7244 96213 7253
rect 96171 7204 96172 7244
rect 96212 7204 96213 7244
rect 96171 7195 96213 7204
rect 96268 7160 96308 7171
rect 96268 7085 96308 7120
rect 96267 7076 96309 7085
rect 96020 6616 96116 6656
rect 96172 7036 96268 7076
rect 96308 7036 96309 7076
rect 95980 6607 96020 6616
rect 95691 6488 95733 6497
rect 95691 6448 95692 6488
rect 95732 6448 95733 6488
rect 95691 6439 95733 6448
rect 96172 6413 96212 7036
rect 96267 7027 96309 7036
rect 96364 6656 96404 7624
rect 96556 7496 96596 7708
rect 96705 7664 96745 8064
rect 96815 7748 96855 8064
rect 96815 7708 96884 7748
rect 96705 7624 96788 7664
rect 96556 7456 96692 7496
rect 96459 7412 96501 7421
rect 96459 7372 96460 7412
rect 96500 7372 96501 7412
rect 96459 7363 96501 7372
rect 96460 7278 96500 7363
rect 96555 7244 96597 7253
rect 96555 7204 96556 7244
rect 96596 7204 96597 7244
rect 96555 7195 96597 7204
rect 96556 7160 96596 7195
rect 96556 7085 96596 7120
rect 96555 7076 96597 7085
rect 96555 7036 96556 7076
rect 96596 7036 96597 7076
rect 96555 7027 96597 7036
rect 96364 6607 96404 6616
rect 94924 6353 94964 6364
rect 95403 6404 95445 6413
rect 95403 6364 95404 6404
rect 95444 6364 95445 6404
rect 95403 6355 95445 6364
rect 95787 6404 95829 6413
rect 95787 6364 95788 6404
rect 95828 6364 95829 6404
rect 95787 6355 95829 6364
rect 96171 6404 96213 6413
rect 96171 6364 96172 6404
rect 96212 6364 96213 6404
rect 96171 6355 96213 6364
rect 96556 6404 96596 7027
rect 96652 7001 96692 7456
rect 96651 6992 96693 7001
rect 96651 6952 96652 6992
rect 96692 6952 96693 6992
rect 96651 6943 96693 6952
rect 96748 6656 96788 7624
rect 96844 7421 96884 7708
rect 97105 7664 97145 8064
rect 97215 7664 97255 8064
rect 97505 7673 97545 8064
rect 97504 7664 97546 7673
rect 97615 7664 97655 8064
rect 97105 7624 97172 7664
rect 97215 7624 97268 7664
rect 96843 7412 96885 7421
rect 96843 7372 96844 7412
rect 96884 7372 96885 7412
rect 96843 7363 96885 7372
rect 96844 7244 96884 7253
rect 96844 6917 96884 7204
rect 97036 6992 97076 7001
rect 96843 6908 96885 6917
rect 96843 6868 96844 6908
rect 96884 6868 96885 6908
rect 96843 6859 96885 6868
rect 97036 6833 97076 6952
rect 97035 6824 97077 6833
rect 97035 6784 97036 6824
rect 97076 6784 97077 6824
rect 97035 6775 97077 6784
rect 96748 6607 96788 6616
rect 97036 6656 97076 6665
rect 97132 6656 97172 7624
rect 97228 7337 97268 7624
rect 97504 7624 97505 7664
rect 97545 7624 97546 7664
rect 97504 7615 97546 7624
rect 97612 7624 97655 7664
rect 97707 7664 97749 7673
rect 97707 7624 97708 7664
rect 97748 7624 97749 7664
rect 97905 7664 97945 8064
rect 98015 7748 98055 8064
rect 98305 7748 98345 8064
rect 98015 7708 98132 7748
rect 97905 7624 98036 7664
rect 97227 7328 97269 7337
rect 97227 7288 97228 7328
rect 97268 7288 97269 7328
rect 97227 7279 97269 7288
rect 97324 7253 97364 7338
rect 97323 7244 97365 7253
rect 97323 7204 97324 7244
rect 97364 7204 97556 7244
rect 97323 7195 97365 7204
rect 97324 7173 97364 7195
rect 97227 7160 97269 7169
rect 97227 7120 97228 7160
rect 97268 7120 97269 7160
rect 97324 7124 97364 7133
rect 97516 7160 97556 7204
rect 97612 7169 97652 7624
rect 97707 7615 97749 7624
rect 97227 7111 97269 7120
rect 97516 7111 97556 7120
rect 97611 7160 97653 7169
rect 97611 7120 97612 7160
rect 97652 7120 97653 7160
rect 97611 7111 97653 7120
rect 97228 7026 97268 7111
rect 97611 6992 97653 7001
rect 97611 6952 97612 6992
rect 97652 6952 97653 6992
rect 97611 6943 97653 6952
rect 97612 6858 97652 6943
rect 97227 6824 97269 6833
rect 97227 6784 97228 6824
rect 97268 6784 97269 6824
rect 97227 6775 97269 6784
rect 97076 6616 97172 6656
rect 97036 6607 97076 6616
rect 97228 6413 97268 6775
rect 97516 6656 97556 6665
rect 97708 6656 97748 7615
rect 97803 7412 97845 7421
rect 97803 7372 97804 7412
rect 97844 7372 97845 7412
rect 97803 7363 97845 7372
rect 97804 7278 97844 7363
rect 97900 7160 97940 7169
rect 97556 6616 97748 6656
rect 97804 7120 97900 7160
rect 97516 6607 97556 6616
rect 96556 6355 96596 6364
rect 97227 6404 97269 6413
rect 97227 6364 97228 6404
rect 97268 6364 97269 6404
rect 97227 6355 97269 6364
rect 97707 6404 97749 6413
rect 97804 6404 97844 7120
rect 97900 7111 97940 7120
rect 97900 6656 97940 6665
rect 97996 6656 98036 7624
rect 98092 7505 98132 7708
rect 98284 7708 98345 7748
rect 98091 7496 98133 7505
rect 98091 7456 98092 7496
rect 98132 7456 98133 7496
rect 98091 7447 98133 7456
rect 98284 7421 98324 7708
rect 98415 7664 98455 8064
rect 98380 7624 98455 7664
rect 98283 7412 98325 7421
rect 98283 7372 98284 7412
rect 98324 7372 98325 7412
rect 98283 7363 98325 7372
rect 98091 7328 98133 7337
rect 98091 7288 98092 7328
rect 98132 7288 98133 7328
rect 98091 7279 98133 7288
rect 98092 7194 98132 7279
rect 98188 7160 98228 7169
rect 98188 7001 98228 7120
rect 98187 6992 98229 7001
rect 98187 6952 98188 6992
rect 98228 6952 98229 6992
rect 98187 6943 98229 6952
rect 97940 6616 98036 6656
rect 97900 6607 97940 6616
rect 97707 6364 97708 6404
rect 97748 6364 97844 6404
rect 98091 6404 98133 6413
rect 98188 6404 98228 6943
rect 98380 6656 98420 7624
rect 98475 7412 98517 7421
rect 98475 7372 98476 7412
rect 98516 7372 98517 7412
rect 98475 7363 98517 7372
rect 98476 7278 98516 7363
rect 98668 7244 98708 7253
rect 98860 7244 98900 13672
rect 99243 7496 99285 7505
rect 99243 7456 99244 7496
rect 99284 7456 99285 7496
rect 99243 7447 99285 7456
rect 99244 7412 99284 7447
rect 99244 7361 99284 7372
rect 98380 6607 98420 6616
rect 98572 7204 98668 7244
rect 98708 7204 98900 7244
rect 98476 6488 98516 6497
rect 98572 6488 98612 7204
rect 98668 7195 98708 7204
rect 98956 7160 98996 7169
rect 99148 7160 99188 7169
rect 98996 7120 99148 7160
rect 98859 7076 98901 7085
rect 98859 7036 98860 7076
rect 98900 7036 98901 7076
rect 98859 7027 98901 7036
rect 98860 6942 98900 7027
rect 98956 7001 98996 7120
rect 99148 7111 99188 7120
rect 98955 6992 98997 7001
rect 98955 6952 98956 6992
rect 98996 6952 98997 6992
rect 98955 6943 98997 6952
rect 98516 6448 98612 6488
rect 98476 6439 98516 6448
rect 98091 6364 98092 6404
rect 98132 6364 98228 6404
rect 97707 6355 97749 6364
rect 98091 6355 98133 6364
rect 95404 6270 95444 6355
rect 95788 6270 95828 6355
rect 96172 6270 96212 6355
rect 97228 6270 97268 6355
rect 97708 6270 97748 6355
rect 98092 6270 98132 6355
rect 94060 5851 94100 5860
rect 93964 5599 94004 5608
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 8352 5312 8720 5321
rect 8392 5272 8434 5312
rect 8474 5272 8516 5312
rect 8556 5272 8598 5312
rect 8638 5272 8680 5312
rect 8352 5263 8720 5272
rect 12352 5312 12720 5321
rect 12392 5272 12434 5312
rect 12474 5272 12516 5312
rect 12556 5272 12598 5312
rect 12638 5272 12680 5312
rect 12352 5263 12720 5272
rect 16352 5312 16720 5321
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16352 5263 16720 5272
rect 20352 5312 20720 5321
rect 20392 5272 20434 5312
rect 20474 5272 20516 5312
rect 20556 5272 20598 5312
rect 20638 5272 20680 5312
rect 20352 5263 20720 5272
rect 24352 5312 24720 5321
rect 24392 5272 24434 5312
rect 24474 5272 24516 5312
rect 24556 5272 24598 5312
rect 24638 5272 24680 5312
rect 24352 5263 24720 5272
rect 28352 5312 28720 5321
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28352 5263 28720 5272
rect 32352 5312 32720 5321
rect 32392 5272 32434 5312
rect 32474 5272 32516 5312
rect 32556 5272 32598 5312
rect 32638 5272 32680 5312
rect 32352 5263 32720 5272
rect 36352 5312 36720 5321
rect 36392 5272 36434 5312
rect 36474 5272 36516 5312
rect 36556 5272 36598 5312
rect 36638 5272 36680 5312
rect 36352 5263 36720 5272
rect 40352 5312 40720 5321
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40352 5263 40720 5272
rect 44352 5312 44720 5321
rect 44392 5272 44434 5312
rect 44474 5272 44516 5312
rect 44556 5272 44598 5312
rect 44638 5272 44680 5312
rect 44352 5263 44720 5272
rect 48352 5312 48720 5321
rect 48392 5272 48434 5312
rect 48474 5272 48516 5312
rect 48556 5272 48598 5312
rect 48638 5272 48680 5312
rect 48352 5263 48720 5272
rect 52352 5312 52720 5321
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52352 5263 52720 5272
rect 56352 5312 56720 5321
rect 56392 5272 56434 5312
rect 56474 5272 56516 5312
rect 56556 5272 56598 5312
rect 56638 5272 56680 5312
rect 56352 5263 56720 5272
rect 60352 5312 60720 5321
rect 60392 5272 60434 5312
rect 60474 5272 60516 5312
rect 60556 5272 60598 5312
rect 60638 5272 60680 5312
rect 60352 5263 60720 5272
rect 64352 5312 64720 5321
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64352 5263 64720 5272
rect 68352 5312 68720 5321
rect 68392 5272 68434 5312
rect 68474 5272 68516 5312
rect 68556 5272 68598 5312
rect 68638 5272 68680 5312
rect 68352 5263 68720 5272
rect 72352 5312 72720 5321
rect 72392 5272 72434 5312
rect 72474 5272 72516 5312
rect 72556 5272 72598 5312
rect 72638 5272 72680 5312
rect 72352 5263 72720 5272
rect 76352 5312 76720 5321
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76352 5263 76720 5272
rect 80352 5312 80720 5321
rect 80392 5272 80434 5312
rect 80474 5272 80516 5312
rect 80556 5272 80598 5312
rect 80638 5272 80680 5312
rect 80352 5263 80720 5272
rect 84352 5312 84720 5321
rect 84392 5272 84434 5312
rect 84474 5272 84516 5312
rect 84556 5272 84598 5312
rect 84638 5272 84680 5312
rect 84352 5263 84720 5272
rect 88352 5312 88720 5321
rect 88392 5272 88434 5312
rect 88474 5272 88516 5312
rect 88556 5272 88598 5312
rect 88638 5272 88680 5312
rect 88352 5263 88720 5272
rect 92352 5312 92720 5321
rect 92392 5272 92434 5312
rect 92474 5272 92516 5312
rect 92556 5272 92598 5312
rect 92638 5272 92680 5312
rect 92352 5263 92720 5272
rect 96352 5312 96720 5321
rect 96392 5272 96434 5312
rect 96474 5272 96516 5312
rect 96556 5272 96598 5312
rect 96638 5272 96680 5312
rect 96352 5263 96720 5272
rect 1035 4892 1077 4901
rect 1035 4852 1036 4892
rect 1076 4852 1077 4892
rect 1035 4843 1077 4852
rect 1419 4892 1461 4901
rect 1419 4852 1420 4892
rect 1460 4852 1461 4892
rect 1419 4843 1461 4852
rect 1803 4892 1845 4901
rect 1803 4852 1804 4892
rect 1844 4852 1845 4892
rect 1803 4843 1845 4852
rect 2187 4892 2229 4901
rect 2187 4852 2188 4892
rect 2228 4852 2229 4892
rect 2187 4843 2229 4852
rect 651 4808 693 4817
rect 651 4768 652 4808
rect 692 4768 693 4808
rect 651 4759 693 4768
rect 652 4388 692 4759
rect 1036 4758 1076 4843
rect 1420 4758 1460 4843
rect 1804 4758 1844 4843
rect 2188 4758 2228 4843
rect 747 4724 789 4733
rect 747 4684 748 4724
rect 788 4684 789 4724
rect 747 4675 789 4684
rect 844 4724 884 4733
rect 1228 4724 1268 4733
rect 884 4684 980 4724
rect 844 4675 884 4684
rect 652 4339 692 4348
rect 651 3212 693 3221
rect 651 3172 652 3212
rect 692 3172 693 3212
rect 651 3163 693 3172
rect 652 3078 692 3163
rect 748 2708 788 4675
rect 843 4220 885 4229
rect 843 4180 844 4220
rect 884 4180 885 4220
rect 843 4171 885 4180
rect 844 4086 884 4171
rect 844 3380 884 3389
rect 940 3380 980 4684
rect 1228 4220 1268 4684
rect 1612 4724 1652 4733
rect 1612 4229 1652 4684
rect 1995 4724 2037 4733
rect 1995 4684 1996 4724
rect 2036 4684 2037 4724
rect 1995 4675 2037 4684
rect 1996 4590 2036 4675
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 7112 4556 7480 4565
rect 7152 4516 7194 4556
rect 7234 4516 7276 4556
rect 7316 4516 7358 4556
rect 7398 4516 7440 4556
rect 7112 4507 7480 4516
rect 11112 4556 11480 4565
rect 11152 4516 11194 4556
rect 11234 4516 11276 4556
rect 11316 4516 11358 4556
rect 11398 4516 11440 4556
rect 11112 4507 11480 4516
rect 15112 4556 15480 4565
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15112 4507 15480 4516
rect 19112 4556 19480 4565
rect 19152 4516 19194 4556
rect 19234 4516 19276 4556
rect 19316 4516 19358 4556
rect 19398 4516 19440 4556
rect 19112 4507 19480 4516
rect 23112 4556 23480 4565
rect 23152 4516 23194 4556
rect 23234 4516 23276 4556
rect 23316 4516 23358 4556
rect 23398 4516 23440 4556
rect 23112 4507 23480 4516
rect 27112 4556 27480 4565
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27112 4507 27480 4516
rect 31112 4556 31480 4565
rect 31152 4516 31194 4556
rect 31234 4516 31276 4556
rect 31316 4516 31358 4556
rect 31398 4516 31440 4556
rect 31112 4507 31480 4516
rect 35112 4556 35480 4565
rect 35152 4516 35194 4556
rect 35234 4516 35276 4556
rect 35316 4516 35358 4556
rect 35398 4516 35440 4556
rect 35112 4507 35480 4516
rect 39112 4556 39480 4565
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39112 4507 39480 4516
rect 43112 4556 43480 4565
rect 43152 4516 43194 4556
rect 43234 4516 43276 4556
rect 43316 4516 43358 4556
rect 43398 4516 43440 4556
rect 43112 4507 43480 4516
rect 47112 4556 47480 4565
rect 47152 4516 47194 4556
rect 47234 4516 47276 4556
rect 47316 4516 47358 4556
rect 47398 4516 47440 4556
rect 47112 4507 47480 4516
rect 51112 4556 51480 4565
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51112 4507 51480 4516
rect 55112 4556 55480 4565
rect 55152 4516 55194 4556
rect 55234 4516 55276 4556
rect 55316 4516 55358 4556
rect 55398 4516 55440 4556
rect 55112 4507 55480 4516
rect 59112 4556 59480 4565
rect 59152 4516 59194 4556
rect 59234 4516 59276 4556
rect 59316 4516 59358 4556
rect 59398 4516 59440 4556
rect 59112 4507 59480 4516
rect 63112 4556 63480 4565
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63112 4507 63480 4516
rect 67112 4556 67480 4565
rect 67152 4516 67194 4556
rect 67234 4516 67276 4556
rect 67316 4516 67358 4556
rect 67398 4516 67440 4556
rect 67112 4507 67480 4516
rect 71112 4556 71480 4565
rect 71152 4516 71194 4556
rect 71234 4516 71276 4556
rect 71316 4516 71358 4556
rect 71398 4516 71440 4556
rect 71112 4507 71480 4516
rect 75112 4556 75480 4565
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75112 4507 75480 4516
rect 79112 4556 79480 4565
rect 79152 4516 79194 4556
rect 79234 4516 79276 4556
rect 79316 4516 79358 4556
rect 79398 4516 79440 4556
rect 79112 4507 79480 4516
rect 83112 4556 83480 4565
rect 83152 4516 83194 4556
rect 83234 4516 83276 4556
rect 83316 4516 83358 4556
rect 83398 4516 83440 4556
rect 83112 4507 83480 4516
rect 87112 4556 87480 4565
rect 87152 4516 87194 4556
rect 87234 4516 87276 4556
rect 87316 4516 87358 4556
rect 87398 4516 87440 4556
rect 87112 4507 87480 4516
rect 91112 4556 91480 4565
rect 91152 4516 91194 4556
rect 91234 4516 91276 4556
rect 91316 4516 91358 4556
rect 91398 4516 91440 4556
rect 91112 4507 91480 4516
rect 95112 4556 95480 4565
rect 95152 4516 95194 4556
rect 95234 4516 95276 4556
rect 95316 4516 95358 4556
rect 95398 4516 95440 4556
rect 95112 4507 95480 4516
rect 99112 4556 99480 4565
rect 99152 4516 99194 4556
rect 99234 4516 99276 4556
rect 99316 4516 99358 4556
rect 99398 4516 99440 4556
rect 99112 4507 99480 4516
rect 1228 4171 1268 4180
rect 1611 4220 1653 4229
rect 1611 4180 1612 4220
rect 1652 4180 1653 4220
rect 1611 4171 1653 4180
rect 1035 3968 1077 3977
rect 1035 3928 1036 3968
rect 1076 3928 1077 3968
rect 1035 3919 1077 3928
rect 1036 3834 1076 3919
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 8352 3800 8720 3809
rect 8392 3760 8434 3800
rect 8474 3760 8516 3800
rect 8556 3760 8598 3800
rect 8638 3760 8680 3800
rect 8352 3751 8720 3760
rect 12352 3800 12720 3809
rect 12392 3760 12434 3800
rect 12474 3760 12516 3800
rect 12556 3760 12598 3800
rect 12638 3760 12680 3800
rect 12352 3751 12720 3760
rect 16352 3800 16720 3809
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16352 3751 16720 3760
rect 20352 3800 20720 3809
rect 20392 3760 20434 3800
rect 20474 3760 20516 3800
rect 20556 3760 20598 3800
rect 20638 3760 20680 3800
rect 20352 3751 20720 3760
rect 24352 3800 24720 3809
rect 24392 3760 24434 3800
rect 24474 3760 24516 3800
rect 24556 3760 24598 3800
rect 24638 3760 24680 3800
rect 24352 3751 24720 3760
rect 28352 3800 28720 3809
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28352 3751 28720 3760
rect 32352 3800 32720 3809
rect 32392 3760 32434 3800
rect 32474 3760 32516 3800
rect 32556 3760 32598 3800
rect 32638 3760 32680 3800
rect 32352 3751 32720 3760
rect 36352 3800 36720 3809
rect 36392 3760 36434 3800
rect 36474 3760 36516 3800
rect 36556 3760 36598 3800
rect 36638 3760 36680 3800
rect 36352 3751 36720 3760
rect 40352 3800 40720 3809
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40352 3751 40720 3760
rect 44352 3800 44720 3809
rect 44392 3760 44434 3800
rect 44474 3760 44516 3800
rect 44556 3760 44598 3800
rect 44638 3760 44680 3800
rect 44352 3751 44720 3760
rect 48352 3800 48720 3809
rect 48392 3760 48434 3800
rect 48474 3760 48516 3800
rect 48556 3760 48598 3800
rect 48638 3760 48680 3800
rect 48352 3751 48720 3760
rect 52352 3800 52720 3809
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52352 3751 52720 3760
rect 56352 3800 56720 3809
rect 56392 3760 56434 3800
rect 56474 3760 56516 3800
rect 56556 3760 56598 3800
rect 56638 3760 56680 3800
rect 56352 3751 56720 3760
rect 60352 3800 60720 3809
rect 60392 3760 60434 3800
rect 60474 3760 60516 3800
rect 60556 3760 60598 3800
rect 60638 3760 60680 3800
rect 60352 3751 60720 3760
rect 64352 3800 64720 3809
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64352 3751 64720 3760
rect 68352 3800 68720 3809
rect 68392 3760 68434 3800
rect 68474 3760 68516 3800
rect 68556 3760 68598 3800
rect 68638 3760 68680 3800
rect 68352 3751 68720 3760
rect 72352 3800 72720 3809
rect 72392 3760 72434 3800
rect 72474 3760 72516 3800
rect 72556 3760 72598 3800
rect 72638 3760 72680 3800
rect 72352 3751 72720 3760
rect 76352 3800 76720 3809
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76352 3751 76720 3760
rect 80352 3800 80720 3809
rect 80392 3760 80434 3800
rect 80474 3760 80516 3800
rect 80556 3760 80598 3800
rect 80638 3760 80680 3800
rect 80352 3751 80720 3760
rect 84352 3800 84720 3809
rect 84392 3760 84434 3800
rect 84474 3760 84516 3800
rect 84556 3760 84598 3800
rect 84638 3760 84680 3800
rect 84352 3751 84720 3760
rect 88352 3800 88720 3809
rect 88392 3760 88434 3800
rect 88474 3760 88516 3800
rect 88556 3760 88598 3800
rect 88638 3760 88680 3800
rect 88352 3751 88720 3760
rect 92352 3800 92720 3809
rect 92392 3760 92434 3800
rect 92474 3760 92516 3800
rect 92556 3760 92598 3800
rect 92638 3760 92680 3800
rect 92352 3751 92720 3760
rect 96352 3800 96720 3809
rect 96392 3760 96434 3800
rect 96474 3760 96516 3800
rect 96556 3760 96598 3800
rect 96638 3760 96680 3800
rect 96352 3751 96720 3760
rect 884 3340 980 3380
rect 844 3331 884 3340
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 7112 3044 7480 3053
rect 7152 3004 7194 3044
rect 7234 3004 7276 3044
rect 7316 3004 7358 3044
rect 7398 3004 7440 3044
rect 7112 2995 7480 3004
rect 11112 3044 11480 3053
rect 11152 3004 11194 3044
rect 11234 3004 11276 3044
rect 11316 3004 11358 3044
rect 11398 3004 11440 3044
rect 11112 2995 11480 3004
rect 15112 3044 15480 3053
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15112 2995 15480 3004
rect 19112 3044 19480 3053
rect 19152 3004 19194 3044
rect 19234 3004 19276 3044
rect 19316 3004 19358 3044
rect 19398 3004 19440 3044
rect 19112 2995 19480 3004
rect 23112 3044 23480 3053
rect 23152 3004 23194 3044
rect 23234 3004 23276 3044
rect 23316 3004 23358 3044
rect 23398 3004 23440 3044
rect 23112 2995 23480 3004
rect 27112 3044 27480 3053
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27112 2995 27480 3004
rect 31112 3044 31480 3053
rect 31152 3004 31194 3044
rect 31234 3004 31276 3044
rect 31316 3004 31358 3044
rect 31398 3004 31440 3044
rect 31112 2995 31480 3004
rect 35112 3044 35480 3053
rect 35152 3004 35194 3044
rect 35234 3004 35276 3044
rect 35316 3004 35358 3044
rect 35398 3004 35440 3044
rect 35112 2995 35480 3004
rect 39112 3044 39480 3053
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39112 2995 39480 3004
rect 43112 3044 43480 3053
rect 43152 3004 43194 3044
rect 43234 3004 43276 3044
rect 43316 3004 43358 3044
rect 43398 3004 43440 3044
rect 43112 2995 43480 3004
rect 47112 3044 47480 3053
rect 47152 3004 47194 3044
rect 47234 3004 47276 3044
rect 47316 3004 47358 3044
rect 47398 3004 47440 3044
rect 47112 2995 47480 3004
rect 51112 3044 51480 3053
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51112 2995 51480 3004
rect 55112 3044 55480 3053
rect 55152 3004 55194 3044
rect 55234 3004 55276 3044
rect 55316 3004 55358 3044
rect 55398 3004 55440 3044
rect 55112 2995 55480 3004
rect 59112 3044 59480 3053
rect 59152 3004 59194 3044
rect 59234 3004 59276 3044
rect 59316 3004 59358 3044
rect 59398 3004 59440 3044
rect 59112 2995 59480 3004
rect 63112 3044 63480 3053
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63112 2995 63480 3004
rect 67112 3044 67480 3053
rect 67152 3004 67194 3044
rect 67234 3004 67276 3044
rect 67316 3004 67358 3044
rect 67398 3004 67440 3044
rect 67112 2995 67480 3004
rect 71112 3044 71480 3053
rect 71152 3004 71194 3044
rect 71234 3004 71276 3044
rect 71316 3004 71358 3044
rect 71398 3004 71440 3044
rect 71112 2995 71480 3004
rect 75112 3044 75480 3053
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75112 2995 75480 3004
rect 79112 3044 79480 3053
rect 79152 3004 79194 3044
rect 79234 3004 79276 3044
rect 79316 3004 79358 3044
rect 79398 3004 79440 3044
rect 79112 2995 79480 3004
rect 83112 3044 83480 3053
rect 83152 3004 83194 3044
rect 83234 3004 83276 3044
rect 83316 3004 83358 3044
rect 83398 3004 83440 3044
rect 83112 2995 83480 3004
rect 87112 3044 87480 3053
rect 87152 3004 87194 3044
rect 87234 3004 87276 3044
rect 87316 3004 87358 3044
rect 87398 3004 87440 3044
rect 87112 2995 87480 3004
rect 91112 3044 91480 3053
rect 91152 3004 91194 3044
rect 91234 3004 91276 3044
rect 91316 3004 91358 3044
rect 91398 3004 91440 3044
rect 91112 2995 91480 3004
rect 95112 3044 95480 3053
rect 95152 3004 95194 3044
rect 95234 3004 95276 3044
rect 95316 3004 95358 3044
rect 95398 3004 95440 3044
rect 95112 2995 95480 3004
rect 99112 3044 99480 3053
rect 99152 3004 99194 3044
rect 99234 3004 99276 3044
rect 99316 3004 99358 3044
rect 99398 3004 99440 3044
rect 99112 2995 99480 3004
rect 844 2708 884 2717
rect 748 2668 844 2708
rect 844 2659 884 2668
rect 652 2456 692 2465
rect 652 2297 692 2416
rect 651 2288 693 2297
rect 651 2248 652 2288
rect 692 2248 693 2288
rect 651 2239 693 2248
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 8352 2288 8720 2297
rect 8392 2248 8434 2288
rect 8474 2248 8516 2288
rect 8556 2248 8598 2288
rect 8638 2248 8680 2288
rect 8352 2239 8720 2248
rect 12352 2288 12720 2297
rect 12392 2248 12434 2288
rect 12474 2248 12516 2288
rect 12556 2248 12598 2288
rect 12638 2248 12680 2288
rect 12352 2239 12720 2248
rect 16352 2288 16720 2297
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16352 2239 16720 2248
rect 20352 2288 20720 2297
rect 20392 2248 20434 2288
rect 20474 2248 20516 2288
rect 20556 2248 20598 2288
rect 20638 2248 20680 2288
rect 20352 2239 20720 2248
rect 24352 2288 24720 2297
rect 24392 2248 24434 2288
rect 24474 2248 24516 2288
rect 24556 2248 24598 2288
rect 24638 2248 24680 2288
rect 24352 2239 24720 2248
rect 28352 2288 28720 2297
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28352 2239 28720 2248
rect 32352 2288 32720 2297
rect 32392 2248 32434 2288
rect 32474 2248 32516 2288
rect 32556 2248 32598 2288
rect 32638 2248 32680 2288
rect 32352 2239 32720 2248
rect 36352 2288 36720 2297
rect 36392 2248 36434 2288
rect 36474 2248 36516 2288
rect 36556 2248 36598 2288
rect 36638 2248 36680 2288
rect 36352 2239 36720 2248
rect 40352 2288 40720 2297
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40352 2239 40720 2248
rect 44352 2288 44720 2297
rect 44392 2248 44434 2288
rect 44474 2248 44516 2288
rect 44556 2248 44598 2288
rect 44638 2248 44680 2288
rect 44352 2239 44720 2248
rect 48352 2288 48720 2297
rect 48392 2248 48434 2288
rect 48474 2248 48516 2288
rect 48556 2248 48598 2288
rect 48638 2248 48680 2288
rect 48352 2239 48720 2248
rect 52352 2288 52720 2297
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52352 2239 52720 2248
rect 56352 2288 56720 2297
rect 56392 2248 56434 2288
rect 56474 2248 56516 2288
rect 56556 2248 56598 2288
rect 56638 2248 56680 2288
rect 56352 2239 56720 2248
rect 60352 2288 60720 2297
rect 60392 2248 60434 2288
rect 60474 2248 60516 2288
rect 60556 2248 60598 2288
rect 60638 2248 60680 2288
rect 60352 2239 60720 2248
rect 64352 2288 64720 2297
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64352 2239 64720 2248
rect 68352 2288 68720 2297
rect 68392 2248 68434 2288
rect 68474 2248 68516 2288
rect 68556 2248 68598 2288
rect 68638 2248 68680 2288
rect 68352 2239 68720 2248
rect 72352 2288 72720 2297
rect 72392 2248 72434 2288
rect 72474 2248 72516 2288
rect 72556 2248 72598 2288
rect 72638 2248 72680 2288
rect 72352 2239 72720 2248
rect 76352 2288 76720 2297
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76352 2239 76720 2248
rect 80352 2288 80720 2297
rect 80392 2248 80434 2288
rect 80474 2248 80516 2288
rect 80556 2248 80598 2288
rect 80638 2248 80680 2288
rect 80352 2239 80720 2248
rect 84352 2288 84720 2297
rect 84392 2248 84434 2288
rect 84474 2248 84516 2288
rect 84556 2248 84598 2288
rect 84638 2248 84680 2288
rect 84352 2239 84720 2248
rect 88352 2288 88720 2297
rect 88392 2248 88434 2288
rect 88474 2248 88516 2288
rect 88556 2248 88598 2288
rect 88638 2248 88680 2288
rect 88352 2239 88720 2248
rect 92352 2288 92720 2297
rect 92392 2248 92434 2288
rect 92474 2248 92516 2288
rect 92556 2248 92598 2288
rect 92638 2248 92680 2288
rect 92352 2239 92720 2248
rect 96352 2288 96720 2297
rect 96392 2248 96434 2288
rect 96474 2248 96516 2288
rect 96556 2248 96598 2288
rect 96638 2248 96680 2288
rect 96352 2239 96720 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 7112 1532 7480 1541
rect 7152 1492 7194 1532
rect 7234 1492 7276 1532
rect 7316 1492 7358 1532
rect 7398 1492 7440 1532
rect 7112 1483 7480 1492
rect 11112 1532 11480 1541
rect 11152 1492 11194 1532
rect 11234 1492 11276 1532
rect 11316 1492 11358 1532
rect 11398 1492 11440 1532
rect 11112 1483 11480 1492
rect 15112 1532 15480 1541
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15112 1483 15480 1492
rect 19112 1532 19480 1541
rect 19152 1492 19194 1532
rect 19234 1492 19276 1532
rect 19316 1492 19358 1532
rect 19398 1492 19440 1532
rect 19112 1483 19480 1492
rect 23112 1532 23480 1541
rect 23152 1492 23194 1532
rect 23234 1492 23276 1532
rect 23316 1492 23358 1532
rect 23398 1492 23440 1532
rect 23112 1483 23480 1492
rect 27112 1532 27480 1541
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27112 1483 27480 1492
rect 31112 1532 31480 1541
rect 31152 1492 31194 1532
rect 31234 1492 31276 1532
rect 31316 1492 31358 1532
rect 31398 1492 31440 1532
rect 31112 1483 31480 1492
rect 35112 1532 35480 1541
rect 35152 1492 35194 1532
rect 35234 1492 35276 1532
rect 35316 1492 35358 1532
rect 35398 1492 35440 1532
rect 35112 1483 35480 1492
rect 39112 1532 39480 1541
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39112 1483 39480 1492
rect 43112 1532 43480 1541
rect 43152 1492 43194 1532
rect 43234 1492 43276 1532
rect 43316 1492 43358 1532
rect 43398 1492 43440 1532
rect 43112 1483 43480 1492
rect 47112 1532 47480 1541
rect 47152 1492 47194 1532
rect 47234 1492 47276 1532
rect 47316 1492 47358 1532
rect 47398 1492 47440 1532
rect 47112 1483 47480 1492
rect 51112 1532 51480 1541
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51112 1483 51480 1492
rect 55112 1532 55480 1541
rect 55152 1492 55194 1532
rect 55234 1492 55276 1532
rect 55316 1492 55358 1532
rect 55398 1492 55440 1532
rect 55112 1483 55480 1492
rect 59112 1532 59480 1541
rect 59152 1492 59194 1532
rect 59234 1492 59276 1532
rect 59316 1492 59358 1532
rect 59398 1492 59440 1532
rect 59112 1483 59480 1492
rect 63112 1532 63480 1541
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63112 1483 63480 1492
rect 67112 1532 67480 1541
rect 67152 1492 67194 1532
rect 67234 1492 67276 1532
rect 67316 1492 67358 1532
rect 67398 1492 67440 1532
rect 67112 1483 67480 1492
rect 71112 1532 71480 1541
rect 71152 1492 71194 1532
rect 71234 1492 71276 1532
rect 71316 1492 71358 1532
rect 71398 1492 71440 1532
rect 71112 1483 71480 1492
rect 75112 1532 75480 1541
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75112 1483 75480 1492
rect 79112 1532 79480 1541
rect 79152 1492 79194 1532
rect 79234 1492 79276 1532
rect 79316 1492 79358 1532
rect 79398 1492 79440 1532
rect 79112 1483 79480 1492
rect 83112 1532 83480 1541
rect 83152 1492 83194 1532
rect 83234 1492 83276 1532
rect 83316 1492 83358 1532
rect 83398 1492 83440 1532
rect 83112 1483 83480 1492
rect 87112 1532 87480 1541
rect 87152 1492 87194 1532
rect 87234 1492 87276 1532
rect 87316 1492 87358 1532
rect 87398 1492 87440 1532
rect 87112 1483 87480 1492
rect 91112 1532 91480 1541
rect 91152 1492 91194 1532
rect 91234 1492 91276 1532
rect 91316 1492 91358 1532
rect 91398 1492 91440 1532
rect 91112 1483 91480 1492
rect 95112 1532 95480 1541
rect 95152 1492 95194 1532
rect 95234 1492 95276 1532
rect 95316 1492 95358 1532
rect 95398 1492 95440 1532
rect 95112 1483 95480 1492
rect 99112 1532 99480 1541
rect 99152 1492 99194 1532
rect 99234 1492 99276 1532
rect 99316 1492 99358 1532
rect 99398 1492 99440 1532
rect 99112 1483 99480 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 8352 776 8720 785
rect 8392 736 8434 776
rect 8474 736 8516 776
rect 8556 736 8598 776
rect 8638 736 8680 776
rect 8352 727 8720 736
rect 12352 776 12720 785
rect 12392 736 12434 776
rect 12474 736 12516 776
rect 12556 736 12598 776
rect 12638 736 12680 776
rect 12352 727 12720 736
rect 16352 776 16720 785
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16352 727 16720 736
rect 20352 776 20720 785
rect 20392 736 20434 776
rect 20474 736 20516 776
rect 20556 736 20598 776
rect 20638 736 20680 776
rect 20352 727 20720 736
rect 24352 776 24720 785
rect 24392 736 24434 776
rect 24474 736 24516 776
rect 24556 736 24598 776
rect 24638 736 24680 776
rect 24352 727 24720 736
rect 28352 776 28720 785
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28352 727 28720 736
rect 32352 776 32720 785
rect 32392 736 32434 776
rect 32474 736 32516 776
rect 32556 736 32598 776
rect 32638 736 32680 776
rect 32352 727 32720 736
rect 36352 776 36720 785
rect 36392 736 36434 776
rect 36474 736 36516 776
rect 36556 736 36598 776
rect 36638 736 36680 776
rect 36352 727 36720 736
rect 40352 776 40720 785
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40352 727 40720 736
rect 44352 776 44720 785
rect 44392 736 44434 776
rect 44474 736 44516 776
rect 44556 736 44598 776
rect 44638 736 44680 776
rect 44352 727 44720 736
rect 48352 776 48720 785
rect 48392 736 48434 776
rect 48474 736 48516 776
rect 48556 736 48598 776
rect 48638 736 48680 776
rect 48352 727 48720 736
rect 52352 776 52720 785
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52352 727 52720 736
rect 56352 776 56720 785
rect 56392 736 56434 776
rect 56474 736 56516 776
rect 56556 736 56598 776
rect 56638 736 56680 776
rect 56352 727 56720 736
rect 60352 776 60720 785
rect 60392 736 60434 776
rect 60474 736 60516 776
rect 60556 736 60598 776
rect 60638 736 60680 776
rect 60352 727 60720 736
rect 64352 776 64720 785
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64352 727 64720 736
rect 68352 776 68720 785
rect 68392 736 68434 776
rect 68474 736 68516 776
rect 68556 736 68598 776
rect 68638 736 68680 776
rect 68352 727 68720 736
rect 72352 776 72720 785
rect 72392 736 72434 776
rect 72474 736 72516 776
rect 72556 736 72598 776
rect 72638 736 72680 776
rect 72352 727 72720 736
rect 76352 776 76720 785
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76352 727 76720 736
rect 80352 776 80720 785
rect 80392 736 80434 776
rect 80474 736 80516 776
rect 80556 736 80598 776
rect 80638 736 80680 776
rect 80352 727 80720 736
rect 84352 776 84720 785
rect 84392 736 84434 776
rect 84474 736 84516 776
rect 84556 736 84598 776
rect 84638 736 84680 776
rect 84352 727 84720 736
rect 88352 776 88720 785
rect 88392 736 88434 776
rect 88474 736 88516 776
rect 88556 736 88598 776
rect 88638 736 88680 776
rect 88352 727 88720 736
rect 92352 776 92720 785
rect 92392 736 92434 776
rect 92474 736 92516 776
rect 92556 736 92598 776
rect 92638 736 92680 776
rect 92352 727 92720 736
rect 96352 776 96720 785
rect 96392 736 96434 776
rect 96474 736 96516 776
rect 96556 736 96598 776
rect 96638 736 96680 776
rect 96352 727 96720 736
<< via2 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 8352 38536 8392 38576
rect 8434 38536 8474 38576
rect 8516 38536 8556 38576
rect 8598 38536 8638 38576
rect 8680 38536 8720 38576
rect 12352 38536 12392 38576
rect 12434 38536 12474 38576
rect 12516 38536 12556 38576
rect 12598 38536 12638 38576
rect 12680 38536 12720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 20352 38536 20392 38576
rect 20434 38536 20474 38576
rect 20516 38536 20556 38576
rect 20598 38536 20638 38576
rect 20680 38536 20720 38576
rect 24352 38536 24392 38576
rect 24434 38536 24474 38576
rect 24516 38536 24556 38576
rect 24598 38536 24638 38576
rect 24680 38536 24720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 32352 38536 32392 38576
rect 32434 38536 32474 38576
rect 32516 38536 32556 38576
rect 32598 38536 32638 38576
rect 32680 38536 32720 38576
rect 36352 38536 36392 38576
rect 36434 38536 36474 38576
rect 36516 38536 36556 38576
rect 36598 38536 36638 38576
rect 36680 38536 36720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 44352 38536 44392 38576
rect 44434 38536 44474 38576
rect 44516 38536 44556 38576
rect 44598 38536 44638 38576
rect 44680 38536 44720 38576
rect 48352 38536 48392 38576
rect 48434 38536 48474 38576
rect 48516 38536 48556 38576
rect 48598 38536 48638 38576
rect 48680 38536 48720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 56352 38536 56392 38576
rect 56434 38536 56474 38576
rect 56516 38536 56556 38576
rect 56598 38536 56638 38576
rect 56680 38536 56720 38576
rect 60352 38536 60392 38576
rect 60434 38536 60474 38576
rect 60516 38536 60556 38576
rect 60598 38536 60638 38576
rect 60680 38536 60720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 68352 38536 68392 38576
rect 68434 38536 68474 38576
rect 68516 38536 68556 38576
rect 68598 38536 68638 38576
rect 68680 38536 68720 38576
rect 72352 38536 72392 38576
rect 72434 38536 72474 38576
rect 72516 38536 72556 38576
rect 72598 38536 72638 38576
rect 72680 38536 72720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 80352 38536 80392 38576
rect 80434 38536 80474 38576
rect 80516 38536 80556 38576
rect 80598 38536 80638 38576
rect 80680 38536 80720 38576
rect 84352 38536 84392 38576
rect 84434 38536 84474 38576
rect 84516 38536 84556 38576
rect 84598 38536 84638 38576
rect 84680 38536 84720 38576
rect 88352 38536 88392 38576
rect 88434 38536 88474 38576
rect 88516 38536 88556 38576
rect 88598 38536 88638 38576
rect 88680 38536 88720 38576
rect 92352 38536 92392 38576
rect 92434 38536 92474 38576
rect 92516 38536 92556 38576
rect 92598 38536 92638 38576
rect 92680 38536 92720 38576
rect 96352 38536 96392 38576
rect 96434 38536 96474 38576
rect 96516 38536 96556 38576
rect 96598 38536 96638 38576
rect 96680 38536 96720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 7112 37780 7152 37820
rect 7194 37780 7234 37820
rect 7276 37780 7316 37820
rect 7358 37780 7398 37820
rect 7440 37780 7480 37820
rect 11112 37780 11152 37820
rect 11194 37780 11234 37820
rect 11276 37780 11316 37820
rect 11358 37780 11398 37820
rect 11440 37780 11480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 19112 37780 19152 37820
rect 19194 37780 19234 37820
rect 19276 37780 19316 37820
rect 19358 37780 19398 37820
rect 19440 37780 19480 37820
rect 23112 37780 23152 37820
rect 23194 37780 23234 37820
rect 23276 37780 23316 37820
rect 23358 37780 23398 37820
rect 23440 37780 23480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 31112 37780 31152 37820
rect 31194 37780 31234 37820
rect 31276 37780 31316 37820
rect 31358 37780 31398 37820
rect 31440 37780 31480 37820
rect 35112 37780 35152 37820
rect 35194 37780 35234 37820
rect 35276 37780 35316 37820
rect 35358 37780 35398 37820
rect 35440 37780 35480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 43112 37780 43152 37820
rect 43194 37780 43234 37820
rect 43276 37780 43316 37820
rect 43358 37780 43398 37820
rect 43440 37780 43480 37820
rect 47112 37780 47152 37820
rect 47194 37780 47234 37820
rect 47276 37780 47316 37820
rect 47358 37780 47398 37820
rect 47440 37780 47480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 55112 37780 55152 37820
rect 55194 37780 55234 37820
rect 55276 37780 55316 37820
rect 55358 37780 55398 37820
rect 55440 37780 55480 37820
rect 59112 37780 59152 37820
rect 59194 37780 59234 37820
rect 59276 37780 59316 37820
rect 59358 37780 59398 37820
rect 59440 37780 59480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 67112 37780 67152 37820
rect 67194 37780 67234 37820
rect 67276 37780 67316 37820
rect 67358 37780 67398 37820
rect 67440 37780 67480 37820
rect 71112 37780 71152 37820
rect 71194 37780 71234 37820
rect 71276 37780 71316 37820
rect 71358 37780 71398 37820
rect 71440 37780 71480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 79112 37780 79152 37820
rect 79194 37780 79234 37820
rect 79276 37780 79316 37820
rect 79358 37780 79398 37820
rect 79440 37780 79480 37820
rect 83112 37780 83152 37820
rect 83194 37780 83234 37820
rect 83276 37780 83316 37820
rect 83358 37780 83398 37820
rect 83440 37780 83480 37820
rect 87112 37780 87152 37820
rect 87194 37780 87234 37820
rect 87276 37780 87316 37820
rect 87358 37780 87398 37820
rect 87440 37780 87480 37820
rect 91112 37780 91152 37820
rect 91194 37780 91234 37820
rect 91276 37780 91316 37820
rect 91358 37780 91398 37820
rect 91440 37780 91480 37820
rect 95112 37780 95152 37820
rect 95194 37780 95234 37820
rect 95276 37780 95316 37820
rect 95358 37780 95398 37820
rect 95440 37780 95480 37820
rect 99112 37780 99152 37820
rect 99194 37780 99234 37820
rect 99276 37780 99316 37820
rect 99358 37780 99398 37820
rect 99440 37780 99480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 8352 37024 8392 37064
rect 8434 37024 8474 37064
rect 8516 37024 8556 37064
rect 8598 37024 8638 37064
rect 8680 37024 8720 37064
rect 12352 37024 12392 37064
rect 12434 37024 12474 37064
rect 12516 37024 12556 37064
rect 12598 37024 12638 37064
rect 12680 37024 12720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 20352 37024 20392 37064
rect 20434 37024 20474 37064
rect 20516 37024 20556 37064
rect 20598 37024 20638 37064
rect 20680 37024 20720 37064
rect 24352 37024 24392 37064
rect 24434 37024 24474 37064
rect 24516 37024 24556 37064
rect 24598 37024 24638 37064
rect 24680 37024 24720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 32352 37024 32392 37064
rect 32434 37024 32474 37064
rect 32516 37024 32556 37064
rect 32598 37024 32638 37064
rect 32680 37024 32720 37064
rect 36352 37024 36392 37064
rect 36434 37024 36474 37064
rect 36516 37024 36556 37064
rect 36598 37024 36638 37064
rect 36680 37024 36720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 44352 37024 44392 37064
rect 44434 37024 44474 37064
rect 44516 37024 44556 37064
rect 44598 37024 44638 37064
rect 44680 37024 44720 37064
rect 48352 37024 48392 37064
rect 48434 37024 48474 37064
rect 48516 37024 48556 37064
rect 48598 37024 48638 37064
rect 48680 37024 48720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 56352 37024 56392 37064
rect 56434 37024 56474 37064
rect 56516 37024 56556 37064
rect 56598 37024 56638 37064
rect 56680 37024 56720 37064
rect 60352 37024 60392 37064
rect 60434 37024 60474 37064
rect 60516 37024 60556 37064
rect 60598 37024 60638 37064
rect 60680 37024 60720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 68352 37024 68392 37064
rect 68434 37024 68474 37064
rect 68516 37024 68556 37064
rect 68598 37024 68638 37064
rect 68680 37024 68720 37064
rect 72352 37024 72392 37064
rect 72434 37024 72474 37064
rect 72516 37024 72556 37064
rect 72598 37024 72638 37064
rect 72680 37024 72720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 80352 37024 80392 37064
rect 80434 37024 80474 37064
rect 80516 37024 80556 37064
rect 80598 37024 80638 37064
rect 80680 37024 80720 37064
rect 84352 37024 84392 37064
rect 84434 37024 84474 37064
rect 84516 37024 84556 37064
rect 84598 37024 84638 37064
rect 84680 37024 84720 37064
rect 88352 37024 88392 37064
rect 88434 37024 88474 37064
rect 88516 37024 88556 37064
rect 88598 37024 88638 37064
rect 88680 37024 88720 37064
rect 92352 37024 92392 37064
rect 92434 37024 92474 37064
rect 92516 37024 92556 37064
rect 92598 37024 92638 37064
rect 92680 37024 92720 37064
rect 96352 37024 96392 37064
rect 96434 37024 96474 37064
rect 96516 37024 96556 37064
rect 96598 37024 96638 37064
rect 96680 37024 96720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 7112 36268 7152 36308
rect 7194 36268 7234 36308
rect 7276 36268 7316 36308
rect 7358 36268 7398 36308
rect 7440 36268 7480 36308
rect 11112 36268 11152 36308
rect 11194 36268 11234 36308
rect 11276 36268 11316 36308
rect 11358 36268 11398 36308
rect 11440 36268 11480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 19112 36268 19152 36308
rect 19194 36268 19234 36308
rect 19276 36268 19316 36308
rect 19358 36268 19398 36308
rect 19440 36268 19480 36308
rect 23112 36268 23152 36308
rect 23194 36268 23234 36308
rect 23276 36268 23316 36308
rect 23358 36268 23398 36308
rect 23440 36268 23480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 31112 36268 31152 36308
rect 31194 36268 31234 36308
rect 31276 36268 31316 36308
rect 31358 36268 31398 36308
rect 31440 36268 31480 36308
rect 35112 36268 35152 36308
rect 35194 36268 35234 36308
rect 35276 36268 35316 36308
rect 35358 36268 35398 36308
rect 35440 36268 35480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 43112 36268 43152 36308
rect 43194 36268 43234 36308
rect 43276 36268 43316 36308
rect 43358 36268 43398 36308
rect 43440 36268 43480 36308
rect 47112 36268 47152 36308
rect 47194 36268 47234 36308
rect 47276 36268 47316 36308
rect 47358 36268 47398 36308
rect 47440 36268 47480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 55112 36268 55152 36308
rect 55194 36268 55234 36308
rect 55276 36268 55316 36308
rect 55358 36268 55398 36308
rect 55440 36268 55480 36308
rect 59112 36268 59152 36308
rect 59194 36268 59234 36308
rect 59276 36268 59316 36308
rect 59358 36268 59398 36308
rect 59440 36268 59480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 67112 36268 67152 36308
rect 67194 36268 67234 36308
rect 67276 36268 67316 36308
rect 67358 36268 67398 36308
rect 67440 36268 67480 36308
rect 71112 36268 71152 36308
rect 71194 36268 71234 36308
rect 71276 36268 71316 36308
rect 71358 36268 71398 36308
rect 71440 36268 71480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 79112 36268 79152 36308
rect 79194 36268 79234 36308
rect 79276 36268 79316 36308
rect 79358 36268 79398 36308
rect 79440 36268 79480 36308
rect 83112 36268 83152 36308
rect 83194 36268 83234 36308
rect 83276 36268 83316 36308
rect 83358 36268 83398 36308
rect 83440 36268 83480 36308
rect 87112 36268 87152 36308
rect 87194 36268 87234 36308
rect 87276 36268 87316 36308
rect 87358 36268 87398 36308
rect 87440 36268 87480 36308
rect 91112 36268 91152 36308
rect 91194 36268 91234 36308
rect 91276 36268 91316 36308
rect 91358 36268 91398 36308
rect 91440 36268 91480 36308
rect 95112 36268 95152 36308
rect 95194 36268 95234 36308
rect 95276 36268 95316 36308
rect 95358 36268 95398 36308
rect 95440 36268 95480 36308
rect 99112 36268 99152 36308
rect 99194 36268 99234 36308
rect 99276 36268 99316 36308
rect 99358 36268 99398 36308
rect 99440 36268 99480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 8352 35512 8392 35552
rect 8434 35512 8474 35552
rect 8516 35512 8556 35552
rect 8598 35512 8638 35552
rect 8680 35512 8720 35552
rect 12352 35512 12392 35552
rect 12434 35512 12474 35552
rect 12516 35512 12556 35552
rect 12598 35512 12638 35552
rect 12680 35512 12720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 20352 35512 20392 35552
rect 20434 35512 20474 35552
rect 20516 35512 20556 35552
rect 20598 35512 20638 35552
rect 20680 35512 20720 35552
rect 24352 35512 24392 35552
rect 24434 35512 24474 35552
rect 24516 35512 24556 35552
rect 24598 35512 24638 35552
rect 24680 35512 24720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 32352 35512 32392 35552
rect 32434 35512 32474 35552
rect 32516 35512 32556 35552
rect 32598 35512 32638 35552
rect 32680 35512 32720 35552
rect 36352 35512 36392 35552
rect 36434 35512 36474 35552
rect 36516 35512 36556 35552
rect 36598 35512 36638 35552
rect 36680 35512 36720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 44352 35512 44392 35552
rect 44434 35512 44474 35552
rect 44516 35512 44556 35552
rect 44598 35512 44638 35552
rect 44680 35512 44720 35552
rect 48352 35512 48392 35552
rect 48434 35512 48474 35552
rect 48516 35512 48556 35552
rect 48598 35512 48638 35552
rect 48680 35512 48720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 56352 35512 56392 35552
rect 56434 35512 56474 35552
rect 56516 35512 56556 35552
rect 56598 35512 56638 35552
rect 56680 35512 56720 35552
rect 60352 35512 60392 35552
rect 60434 35512 60474 35552
rect 60516 35512 60556 35552
rect 60598 35512 60638 35552
rect 60680 35512 60720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 68352 35512 68392 35552
rect 68434 35512 68474 35552
rect 68516 35512 68556 35552
rect 68598 35512 68638 35552
rect 68680 35512 68720 35552
rect 72352 35512 72392 35552
rect 72434 35512 72474 35552
rect 72516 35512 72556 35552
rect 72598 35512 72638 35552
rect 72680 35512 72720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 80352 35512 80392 35552
rect 80434 35512 80474 35552
rect 80516 35512 80556 35552
rect 80598 35512 80638 35552
rect 80680 35512 80720 35552
rect 84352 35512 84392 35552
rect 84434 35512 84474 35552
rect 84516 35512 84556 35552
rect 84598 35512 84638 35552
rect 84680 35512 84720 35552
rect 88352 35512 88392 35552
rect 88434 35512 88474 35552
rect 88516 35512 88556 35552
rect 88598 35512 88638 35552
rect 88680 35512 88720 35552
rect 92352 35512 92392 35552
rect 92434 35512 92474 35552
rect 92516 35512 92556 35552
rect 92598 35512 92638 35552
rect 92680 35512 92720 35552
rect 96352 35512 96392 35552
rect 96434 35512 96474 35552
rect 96516 35512 96556 35552
rect 96598 35512 96638 35552
rect 96680 35512 96720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 7112 34756 7152 34796
rect 7194 34756 7234 34796
rect 7276 34756 7316 34796
rect 7358 34756 7398 34796
rect 7440 34756 7480 34796
rect 11112 34756 11152 34796
rect 11194 34756 11234 34796
rect 11276 34756 11316 34796
rect 11358 34756 11398 34796
rect 11440 34756 11480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 19112 34756 19152 34796
rect 19194 34756 19234 34796
rect 19276 34756 19316 34796
rect 19358 34756 19398 34796
rect 19440 34756 19480 34796
rect 23112 34756 23152 34796
rect 23194 34756 23234 34796
rect 23276 34756 23316 34796
rect 23358 34756 23398 34796
rect 23440 34756 23480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 31112 34756 31152 34796
rect 31194 34756 31234 34796
rect 31276 34756 31316 34796
rect 31358 34756 31398 34796
rect 31440 34756 31480 34796
rect 35112 34756 35152 34796
rect 35194 34756 35234 34796
rect 35276 34756 35316 34796
rect 35358 34756 35398 34796
rect 35440 34756 35480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 43112 34756 43152 34796
rect 43194 34756 43234 34796
rect 43276 34756 43316 34796
rect 43358 34756 43398 34796
rect 43440 34756 43480 34796
rect 47112 34756 47152 34796
rect 47194 34756 47234 34796
rect 47276 34756 47316 34796
rect 47358 34756 47398 34796
rect 47440 34756 47480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 55112 34756 55152 34796
rect 55194 34756 55234 34796
rect 55276 34756 55316 34796
rect 55358 34756 55398 34796
rect 55440 34756 55480 34796
rect 59112 34756 59152 34796
rect 59194 34756 59234 34796
rect 59276 34756 59316 34796
rect 59358 34756 59398 34796
rect 59440 34756 59480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 67112 34756 67152 34796
rect 67194 34756 67234 34796
rect 67276 34756 67316 34796
rect 67358 34756 67398 34796
rect 67440 34756 67480 34796
rect 71112 34756 71152 34796
rect 71194 34756 71234 34796
rect 71276 34756 71316 34796
rect 71358 34756 71398 34796
rect 71440 34756 71480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 79112 34756 79152 34796
rect 79194 34756 79234 34796
rect 79276 34756 79316 34796
rect 79358 34756 79398 34796
rect 79440 34756 79480 34796
rect 83112 34756 83152 34796
rect 83194 34756 83234 34796
rect 83276 34756 83316 34796
rect 83358 34756 83398 34796
rect 83440 34756 83480 34796
rect 87112 34756 87152 34796
rect 87194 34756 87234 34796
rect 87276 34756 87316 34796
rect 87358 34756 87398 34796
rect 87440 34756 87480 34796
rect 91112 34756 91152 34796
rect 91194 34756 91234 34796
rect 91276 34756 91316 34796
rect 91358 34756 91398 34796
rect 91440 34756 91480 34796
rect 95112 34756 95152 34796
rect 95194 34756 95234 34796
rect 95276 34756 95316 34796
rect 95358 34756 95398 34796
rect 95440 34756 95480 34796
rect 99112 34756 99152 34796
rect 99194 34756 99234 34796
rect 99276 34756 99316 34796
rect 99358 34756 99398 34796
rect 99440 34756 99480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 8352 34000 8392 34040
rect 8434 34000 8474 34040
rect 8516 34000 8556 34040
rect 8598 34000 8638 34040
rect 8680 34000 8720 34040
rect 12352 34000 12392 34040
rect 12434 34000 12474 34040
rect 12516 34000 12556 34040
rect 12598 34000 12638 34040
rect 12680 34000 12720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 20352 34000 20392 34040
rect 20434 34000 20474 34040
rect 20516 34000 20556 34040
rect 20598 34000 20638 34040
rect 20680 34000 20720 34040
rect 24352 34000 24392 34040
rect 24434 34000 24474 34040
rect 24516 34000 24556 34040
rect 24598 34000 24638 34040
rect 24680 34000 24720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 32352 34000 32392 34040
rect 32434 34000 32474 34040
rect 32516 34000 32556 34040
rect 32598 34000 32638 34040
rect 32680 34000 32720 34040
rect 36352 34000 36392 34040
rect 36434 34000 36474 34040
rect 36516 34000 36556 34040
rect 36598 34000 36638 34040
rect 36680 34000 36720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 44352 34000 44392 34040
rect 44434 34000 44474 34040
rect 44516 34000 44556 34040
rect 44598 34000 44638 34040
rect 44680 34000 44720 34040
rect 48352 34000 48392 34040
rect 48434 34000 48474 34040
rect 48516 34000 48556 34040
rect 48598 34000 48638 34040
rect 48680 34000 48720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 56352 34000 56392 34040
rect 56434 34000 56474 34040
rect 56516 34000 56556 34040
rect 56598 34000 56638 34040
rect 56680 34000 56720 34040
rect 60352 34000 60392 34040
rect 60434 34000 60474 34040
rect 60516 34000 60556 34040
rect 60598 34000 60638 34040
rect 60680 34000 60720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 68352 34000 68392 34040
rect 68434 34000 68474 34040
rect 68516 34000 68556 34040
rect 68598 34000 68638 34040
rect 68680 34000 68720 34040
rect 91276 33748 91316 33788
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 7112 33244 7152 33284
rect 7194 33244 7234 33284
rect 7276 33244 7316 33284
rect 7358 33244 7398 33284
rect 7440 33244 7480 33284
rect 11112 33244 11152 33284
rect 11194 33244 11234 33284
rect 11276 33244 11316 33284
rect 11358 33244 11398 33284
rect 11440 33244 11480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 19112 33244 19152 33284
rect 19194 33244 19234 33284
rect 19276 33244 19316 33284
rect 19358 33244 19398 33284
rect 19440 33244 19480 33284
rect 23112 33244 23152 33284
rect 23194 33244 23234 33284
rect 23276 33244 23316 33284
rect 23358 33244 23398 33284
rect 23440 33244 23480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 31112 33244 31152 33284
rect 31194 33244 31234 33284
rect 31276 33244 31316 33284
rect 31358 33244 31398 33284
rect 31440 33244 31480 33284
rect 35112 33244 35152 33284
rect 35194 33244 35234 33284
rect 35276 33244 35316 33284
rect 35358 33244 35398 33284
rect 35440 33244 35480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 43112 33244 43152 33284
rect 43194 33244 43234 33284
rect 43276 33244 43316 33284
rect 43358 33244 43398 33284
rect 43440 33244 43480 33284
rect 47112 33244 47152 33284
rect 47194 33244 47234 33284
rect 47276 33244 47316 33284
rect 47358 33244 47398 33284
rect 47440 33244 47480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 55112 33244 55152 33284
rect 55194 33244 55234 33284
rect 55276 33244 55316 33284
rect 55358 33244 55398 33284
rect 55440 33244 55480 33284
rect 59112 33244 59152 33284
rect 59194 33244 59234 33284
rect 59276 33244 59316 33284
rect 59358 33244 59398 33284
rect 59440 33244 59480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 67112 33244 67152 33284
rect 67194 33244 67234 33284
rect 67276 33244 67316 33284
rect 67358 33244 67398 33284
rect 67440 33244 67480 33284
rect 71788 33244 71828 33284
rect 70732 32908 70772 32948
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 8352 32488 8392 32528
rect 8434 32488 8474 32528
rect 8516 32488 8556 32528
rect 8598 32488 8638 32528
rect 8680 32488 8720 32528
rect 12352 32488 12392 32528
rect 12434 32488 12474 32528
rect 12516 32488 12556 32528
rect 12598 32488 12638 32528
rect 12680 32488 12720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 20352 32488 20392 32528
rect 20434 32488 20474 32528
rect 20516 32488 20556 32528
rect 20598 32488 20638 32528
rect 20680 32488 20720 32528
rect 24352 32488 24392 32528
rect 24434 32488 24474 32528
rect 24516 32488 24556 32528
rect 24598 32488 24638 32528
rect 24680 32488 24720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 32352 32488 32392 32528
rect 32434 32488 32474 32528
rect 32516 32488 32556 32528
rect 32598 32488 32638 32528
rect 32680 32488 32720 32528
rect 36352 32488 36392 32528
rect 36434 32488 36474 32528
rect 36516 32488 36556 32528
rect 36598 32488 36638 32528
rect 36680 32488 36720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 44352 32488 44392 32528
rect 44434 32488 44474 32528
rect 44516 32488 44556 32528
rect 44598 32488 44638 32528
rect 44680 32488 44720 32528
rect 48352 32488 48392 32528
rect 48434 32488 48474 32528
rect 48516 32488 48556 32528
rect 48598 32488 48638 32528
rect 48680 32488 48720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 56352 32488 56392 32528
rect 56434 32488 56474 32528
rect 56516 32488 56556 32528
rect 56598 32488 56638 32528
rect 56680 32488 56720 32528
rect 60352 32488 60392 32528
rect 60434 32488 60474 32528
rect 60516 32488 60556 32528
rect 60598 32488 60638 32528
rect 60680 32488 60720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 68352 32488 68392 32528
rect 68434 32488 68474 32528
rect 68516 32488 68556 32528
rect 68598 32488 68638 32528
rect 68680 32488 68720 32528
rect 71596 32824 71636 32864
rect 70828 32152 70868 32192
rect 70540 32068 70580 32108
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 7112 31732 7152 31772
rect 7194 31732 7234 31772
rect 7276 31732 7316 31772
rect 7358 31732 7398 31772
rect 7440 31732 7480 31772
rect 11112 31732 11152 31772
rect 11194 31732 11234 31772
rect 11276 31732 11316 31772
rect 11358 31732 11398 31772
rect 11440 31732 11480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 19112 31732 19152 31772
rect 19194 31732 19234 31772
rect 19276 31732 19316 31772
rect 19358 31732 19398 31772
rect 19440 31732 19480 31772
rect 23112 31732 23152 31772
rect 23194 31732 23234 31772
rect 23276 31732 23316 31772
rect 23358 31732 23398 31772
rect 23440 31732 23480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 31112 31732 31152 31772
rect 31194 31732 31234 31772
rect 31276 31732 31316 31772
rect 31358 31732 31398 31772
rect 31440 31732 31480 31772
rect 35112 31732 35152 31772
rect 35194 31732 35234 31772
rect 35276 31732 35316 31772
rect 35358 31732 35398 31772
rect 35440 31732 35480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 43112 31732 43152 31772
rect 43194 31732 43234 31772
rect 43276 31732 43316 31772
rect 43358 31732 43398 31772
rect 43440 31732 43480 31772
rect 47112 31732 47152 31772
rect 47194 31732 47234 31772
rect 47276 31732 47316 31772
rect 47358 31732 47398 31772
rect 47440 31732 47480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 55112 31732 55152 31772
rect 55194 31732 55234 31772
rect 55276 31732 55316 31772
rect 55358 31732 55398 31772
rect 55440 31732 55480 31772
rect 59112 31732 59152 31772
rect 59194 31732 59234 31772
rect 59276 31732 59316 31772
rect 59358 31732 59398 31772
rect 59440 31732 59480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 67112 31732 67152 31772
rect 67194 31732 67234 31772
rect 67276 31732 67316 31772
rect 67358 31732 67398 31772
rect 67440 31732 67480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 8352 30976 8392 31016
rect 8434 30976 8474 31016
rect 8516 30976 8556 31016
rect 8598 30976 8638 31016
rect 8680 30976 8720 31016
rect 12352 30976 12392 31016
rect 12434 30976 12474 31016
rect 12516 30976 12556 31016
rect 12598 30976 12638 31016
rect 12680 30976 12720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 20352 30976 20392 31016
rect 20434 30976 20474 31016
rect 20516 30976 20556 31016
rect 20598 30976 20638 31016
rect 20680 30976 20720 31016
rect 24352 30976 24392 31016
rect 24434 30976 24474 31016
rect 24516 30976 24556 31016
rect 24598 30976 24638 31016
rect 24680 30976 24720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 32352 30976 32392 31016
rect 32434 30976 32474 31016
rect 32516 30976 32556 31016
rect 32598 30976 32638 31016
rect 32680 30976 32720 31016
rect 36352 30976 36392 31016
rect 36434 30976 36474 31016
rect 36516 30976 36556 31016
rect 36598 30976 36638 31016
rect 36680 30976 36720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 44352 30976 44392 31016
rect 44434 30976 44474 31016
rect 44516 30976 44556 31016
rect 44598 30976 44638 31016
rect 44680 30976 44720 31016
rect 48352 30976 48392 31016
rect 48434 30976 48474 31016
rect 48516 30976 48556 31016
rect 48598 30976 48638 31016
rect 48680 30976 48720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 56352 30976 56392 31016
rect 56434 30976 56474 31016
rect 56516 30976 56556 31016
rect 56598 30976 56638 31016
rect 56680 30976 56720 31016
rect 60352 30976 60392 31016
rect 60434 30976 60474 31016
rect 60516 30976 60556 31016
rect 60598 30976 60638 31016
rect 60680 30976 60720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 68352 30976 68392 31016
rect 68434 30976 68474 31016
rect 68516 30976 68556 31016
rect 68598 30976 68638 31016
rect 68680 30976 68720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 7112 30220 7152 30260
rect 7194 30220 7234 30260
rect 7276 30220 7316 30260
rect 7358 30220 7398 30260
rect 7440 30220 7480 30260
rect 11112 30220 11152 30260
rect 11194 30220 11234 30260
rect 11276 30220 11316 30260
rect 11358 30220 11398 30260
rect 11440 30220 11480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 19112 30220 19152 30260
rect 19194 30220 19234 30260
rect 19276 30220 19316 30260
rect 19358 30220 19398 30260
rect 19440 30220 19480 30260
rect 23112 30220 23152 30260
rect 23194 30220 23234 30260
rect 23276 30220 23316 30260
rect 23358 30220 23398 30260
rect 23440 30220 23480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 31112 30220 31152 30260
rect 31194 30220 31234 30260
rect 31276 30220 31316 30260
rect 31358 30220 31398 30260
rect 31440 30220 31480 30260
rect 35112 30220 35152 30260
rect 35194 30220 35234 30260
rect 35276 30220 35316 30260
rect 35358 30220 35398 30260
rect 35440 30220 35480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 43112 30220 43152 30260
rect 43194 30220 43234 30260
rect 43276 30220 43316 30260
rect 43358 30220 43398 30260
rect 43440 30220 43480 30260
rect 47112 30220 47152 30260
rect 47194 30220 47234 30260
rect 47276 30220 47316 30260
rect 47358 30220 47398 30260
rect 47440 30220 47480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 55112 30220 55152 30260
rect 55194 30220 55234 30260
rect 55276 30220 55316 30260
rect 55358 30220 55398 30260
rect 55440 30220 55480 30260
rect 59112 30220 59152 30260
rect 59194 30220 59234 30260
rect 59276 30220 59316 30260
rect 59358 30220 59398 30260
rect 59440 30220 59480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 67112 30220 67152 30260
rect 67194 30220 67234 30260
rect 67276 30220 67316 30260
rect 67358 30220 67398 30260
rect 67440 30220 67480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 8352 29464 8392 29504
rect 8434 29464 8474 29504
rect 8516 29464 8556 29504
rect 8598 29464 8638 29504
rect 8680 29464 8720 29504
rect 12352 29464 12392 29504
rect 12434 29464 12474 29504
rect 12516 29464 12556 29504
rect 12598 29464 12638 29504
rect 12680 29464 12720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 20352 29464 20392 29504
rect 20434 29464 20474 29504
rect 20516 29464 20556 29504
rect 20598 29464 20638 29504
rect 20680 29464 20720 29504
rect 24352 29464 24392 29504
rect 24434 29464 24474 29504
rect 24516 29464 24556 29504
rect 24598 29464 24638 29504
rect 24680 29464 24720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 32352 29464 32392 29504
rect 32434 29464 32474 29504
rect 32516 29464 32556 29504
rect 32598 29464 32638 29504
rect 32680 29464 32720 29504
rect 36352 29464 36392 29504
rect 36434 29464 36474 29504
rect 36516 29464 36556 29504
rect 36598 29464 36638 29504
rect 36680 29464 36720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 44352 29464 44392 29504
rect 44434 29464 44474 29504
rect 44516 29464 44556 29504
rect 44598 29464 44638 29504
rect 44680 29464 44720 29504
rect 48352 29464 48392 29504
rect 48434 29464 48474 29504
rect 48516 29464 48556 29504
rect 48598 29464 48638 29504
rect 48680 29464 48720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 56352 29464 56392 29504
rect 56434 29464 56474 29504
rect 56516 29464 56556 29504
rect 56598 29464 56638 29504
rect 56680 29464 56720 29504
rect 60352 29464 60392 29504
rect 60434 29464 60474 29504
rect 60516 29464 60556 29504
rect 60598 29464 60638 29504
rect 60680 29464 60720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 68352 29464 68392 29504
rect 68434 29464 68474 29504
rect 68516 29464 68556 29504
rect 68598 29464 68638 29504
rect 68680 29464 68720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 7112 28708 7152 28748
rect 7194 28708 7234 28748
rect 7276 28708 7316 28748
rect 7358 28708 7398 28748
rect 7440 28708 7480 28748
rect 11112 28708 11152 28748
rect 11194 28708 11234 28748
rect 11276 28708 11316 28748
rect 11358 28708 11398 28748
rect 11440 28708 11480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 19112 28708 19152 28748
rect 19194 28708 19234 28748
rect 19276 28708 19316 28748
rect 19358 28708 19398 28748
rect 19440 28708 19480 28748
rect 23112 28708 23152 28748
rect 23194 28708 23234 28748
rect 23276 28708 23316 28748
rect 23358 28708 23398 28748
rect 23440 28708 23480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 31112 28708 31152 28748
rect 31194 28708 31234 28748
rect 31276 28708 31316 28748
rect 31358 28708 31398 28748
rect 31440 28708 31480 28748
rect 35112 28708 35152 28748
rect 35194 28708 35234 28748
rect 35276 28708 35316 28748
rect 35358 28708 35398 28748
rect 35440 28708 35480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 43112 28708 43152 28748
rect 43194 28708 43234 28748
rect 43276 28708 43316 28748
rect 43358 28708 43398 28748
rect 43440 28708 43480 28748
rect 47112 28708 47152 28748
rect 47194 28708 47234 28748
rect 47276 28708 47316 28748
rect 47358 28708 47398 28748
rect 47440 28708 47480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 55112 28708 55152 28748
rect 55194 28708 55234 28748
rect 55276 28708 55316 28748
rect 55358 28708 55398 28748
rect 55440 28708 55480 28748
rect 59112 28708 59152 28748
rect 59194 28708 59234 28748
rect 59276 28708 59316 28748
rect 59358 28708 59398 28748
rect 59440 28708 59480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 67112 28708 67152 28748
rect 67194 28708 67234 28748
rect 67276 28708 67316 28748
rect 67358 28708 67398 28748
rect 67440 28708 67480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 8352 27952 8392 27992
rect 8434 27952 8474 27992
rect 8516 27952 8556 27992
rect 8598 27952 8638 27992
rect 8680 27952 8720 27992
rect 12352 27952 12392 27992
rect 12434 27952 12474 27992
rect 12516 27952 12556 27992
rect 12598 27952 12638 27992
rect 12680 27952 12720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 20352 27952 20392 27992
rect 20434 27952 20474 27992
rect 20516 27952 20556 27992
rect 20598 27952 20638 27992
rect 20680 27952 20720 27992
rect 24352 27952 24392 27992
rect 24434 27952 24474 27992
rect 24516 27952 24556 27992
rect 24598 27952 24638 27992
rect 24680 27952 24720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 32352 27952 32392 27992
rect 32434 27952 32474 27992
rect 32516 27952 32556 27992
rect 32598 27952 32638 27992
rect 32680 27952 32720 27992
rect 36352 27952 36392 27992
rect 36434 27952 36474 27992
rect 36516 27952 36556 27992
rect 36598 27952 36638 27992
rect 36680 27952 36720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 44352 27952 44392 27992
rect 44434 27952 44474 27992
rect 44516 27952 44556 27992
rect 44598 27952 44638 27992
rect 44680 27952 44720 27992
rect 48352 27952 48392 27992
rect 48434 27952 48474 27992
rect 48516 27952 48556 27992
rect 48598 27952 48638 27992
rect 48680 27952 48720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 56352 27952 56392 27992
rect 56434 27952 56474 27992
rect 56516 27952 56556 27992
rect 56598 27952 56638 27992
rect 56680 27952 56720 27992
rect 60352 27952 60392 27992
rect 60434 27952 60474 27992
rect 60516 27952 60556 27992
rect 60598 27952 60638 27992
rect 60680 27952 60720 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 68352 27952 68392 27992
rect 68434 27952 68474 27992
rect 68516 27952 68556 27992
rect 68598 27952 68638 27992
rect 68680 27952 68720 27992
rect 70924 32068 70964 32108
rect 71116 32068 71156 32108
rect 71404 32320 71444 32360
rect 69964 27616 70004 27656
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 7112 27196 7152 27236
rect 7194 27196 7234 27236
rect 7276 27196 7316 27236
rect 7358 27196 7398 27236
rect 7440 27196 7480 27236
rect 11112 27196 11152 27236
rect 11194 27196 11234 27236
rect 11276 27196 11316 27236
rect 11358 27196 11398 27236
rect 11440 27196 11480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 19112 27196 19152 27236
rect 19194 27196 19234 27236
rect 19276 27196 19316 27236
rect 19358 27196 19398 27236
rect 19440 27196 19480 27236
rect 23112 27196 23152 27236
rect 23194 27196 23234 27236
rect 23276 27196 23316 27236
rect 23358 27196 23398 27236
rect 23440 27196 23480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 31112 27196 31152 27236
rect 31194 27196 31234 27236
rect 31276 27196 31316 27236
rect 31358 27196 31398 27236
rect 31440 27196 31480 27236
rect 35112 27196 35152 27236
rect 35194 27196 35234 27236
rect 35276 27196 35316 27236
rect 35358 27196 35398 27236
rect 35440 27196 35480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 43112 27196 43152 27236
rect 43194 27196 43234 27236
rect 43276 27196 43316 27236
rect 43358 27196 43398 27236
rect 43440 27196 43480 27236
rect 47112 27196 47152 27236
rect 47194 27196 47234 27236
rect 47276 27196 47316 27236
rect 47358 27196 47398 27236
rect 47440 27196 47480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 55112 27196 55152 27236
rect 55194 27196 55234 27236
rect 55276 27196 55316 27236
rect 55358 27196 55398 27236
rect 55440 27196 55480 27236
rect 59112 27196 59152 27236
rect 59194 27196 59234 27236
rect 59276 27196 59316 27236
rect 59358 27196 59398 27236
rect 59440 27196 59480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 67112 27196 67152 27236
rect 67194 27196 67234 27236
rect 67276 27196 67316 27236
rect 67358 27196 67398 27236
rect 67440 27196 67480 27236
rect 69772 26776 69812 26816
rect 70348 26776 70388 26816
rect 69964 26692 70004 26732
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 8352 26440 8392 26480
rect 8434 26440 8474 26480
rect 8516 26440 8556 26480
rect 8598 26440 8638 26480
rect 8680 26440 8720 26480
rect 12352 26440 12392 26480
rect 12434 26440 12474 26480
rect 12516 26440 12556 26480
rect 12598 26440 12638 26480
rect 12680 26440 12720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 20352 26440 20392 26480
rect 20434 26440 20474 26480
rect 20516 26440 20556 26480
rect 20598 26440 20638 26480
rect 20680 26440 20720 26480
rect 24352 26440 24392 26480
rect 24434 26440 24474 26480
rect 24516 26440 24556 26480
rect 24598 26440 24638 26480
rect 24680 26440 24720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 32352 26440 32392 26480
rect 32434 26440 32474 26480
rect 32516 26440 32556 26480
rect 32598 26440 32638 26480
rect 32680 26440 32720 26480
rect 36352 26440 36392 26480
rect 36434 26440 36474 26480
rect 36516 26440 36556 26480
rect 36598 26440 36638 26480
rect 36680 26440 36720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 44352 26440 44392 26480
rect 44434 26440 44474 26480
rect 44516 26440 44556 26480
rect 44598 26440 44638 26480
rect 44680 26440 44720 26480
rect 48352 26440 48392 26480
rect 48434 26440 48474 26480
rect 48516 26440 48556 26480
rect 48598 26440 48638 26480
rect 48680 26440 48720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 56352 26440 56392 26480
rect 56434 26440 56474 26480
rect 56516 26440 56556 26480
rect 56598 26440 56638 26480
rect 56680 26440 56720 26480
rect 60352 26440 60392 26480
rect 60434 26440 60474 26480
rect 60516 26440 60556 26480
rect 60598 26440 60638 26480
rect 60680 26440 60720 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 68352 26440 68392 26480
rect 68434 26440 68474 26480
rect 68516 26440 68556 26480
rect 68598 26440 68638 26480
rect 68680 26440 68720 26480
rect 70540 26356 70580 26396
rect 69292 26272 69332 26312
rect 70444 26272 70484 26312
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 7112 25684 7152 25724
rect 7194 25684 7234 25724
rect 7276 25684 7316 25724
rect 7358 25684 7398 25724
rect 7440 25684 7480 25724
rect 11112 25684 11152 25724
rect 11194 25684 11234 25724
rect 11276 25684 11316 25724
rect 11358 25684 11398 25724
rect 11440 25684 11480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 19112 25684 19152 25724
rect 19194 25684 19234 25724
rect 19276 25684 19316 25724
rect 19358 25684 19398 25724
rect 19440 25684 19480 25724
rect 23112 25684 23152 25724
rect 23194 25684 23234 25724
rect 23276 25684 23316 25724
rect 23358 25684 23398 25724
rect 23440 25684 23480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 31112 25684 31152 25724
rect 31194 25684 31234 25724
rect 31276 25684 31316 25724
rect 31358 25684 31398 25724
rect 31440 25684 31480 25724
rect 35112 25684 35152 25724
rect 35194 25684 35234 25724
rect 35276 25684 35316 25724
rect 35358 25684 35398 25724
rect 35440 25684 35480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 43112 25684 43152 25724
rect 43194 25684 43234 25724
rect 43276 25684 43316 25724
rect 43358 25684 43398 25724
rect 43440 25684 43480 25724
rect 47112 25684 47152 25724
rect 47194 25684 47234 25724
rect 47276 25684 47316 25724
rect 47358 25684 47398 25724
rect 47440 25684 47480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 55112 25684 55152 25724
rect 55194 25684 55234 25724
rect 55276 25684 55316 25724
rect 55358 25684 55398 25724
rect 55440 25684 55480 25724
rect 59112 25684 59152 25724
rect 59194 25684 59234 25724
rect 59276 25684 59316 25724
rect 59358 25684 59398 25724
rect 59440 25684 59480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 67112 25684 67152 25724
rect 67194 25684 67234 25724
rect 67276 25684 67316 25724
rect 67358 25684 67398 25724
rect 67440 25684 67480 25724
rect 844 25264 884 25304
rect 652 24928 692 24968
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 8352 24928 8392 24968
rect 8434 24928 8474 24968
rect 8516 24928 8556 24968
rect 8598 24928 8638 24968
rect 8680 24928 8720 24968
rect 12352 24928 12392 24968
rect 12434 24928 12474 24968
rect 12516 24928 12556 24968
rect 12598 24928 12638 24968
rect 12680 24928 12720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 20352 24928 20392 24968
rect 20434 24928 20474 24968
rect 20516 24928 20556 24968
rect 20598 24928 20638 24968
rect 20680 24928 20720 24968
rect 24352 24928 24392 24968
rect 24434 24928 24474 24968
rect 24516 24928 24556 24968
rect 24598 24928 24638 24968
rect 24680 24928 24720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 32352 24928 32392 24968
rect 32434 24928 32474 24968
rect 32516 24928 32556 24968
rect 32598 24928 32638 24968
rect 32680 24928 32720 24968
rect 36352 24928 36392 24968
rect 36434 24928 36474 24968
rect 36516 24928 36556 24968
rect 36598 24928 36638 24968
rect 36680 24928 36720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 44352 24928 44392 24968
rect 44434 24928 44474 24968
rect 44516 24928 44556 24968
rect 44598 24928 44638 24968
rect 44680 24928 44720 24968
rect 48352 24928 48392 24968
rect 48434 24928 48474 24968
rect 48516 24928 48556 24968
rect 48598 24928 48638 24968
rect 48680 24928 48720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 56352 24928 56392 24968
rect 56434 24928 56474 24968
rect 56516 24928 56556 24968
rect 56598 24928 56638 24968
rect 56680 24928 56720 24968
rect 60352 24928 60392 24968
rect 60434 24928 60474 24968
rect 60516 24928 60556 24968
rect 60598 24928 60638 24968
rect 60680 24928 60720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 68352 24928 68392 24968
rect 68434 24928 68474 24968
rect 68516 24928 68556 24968
rect 68598 24928 68638 24968
rect 68680 24928 68720 24968
rect 844 24592 884 24632
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 7112 24172 7152 24212
rect 7194 24172 7234 24212
rect 7276 24172 7316 24212
rect 7358 24172 7398 24212
rect 7440 24172 7480 24212
rect 11112 24172 11152 24212
rect 11194 24172 11234 24212
rect 11276 24172 11316 24212
rect 11358 24172 11398 24212
rect 11440 24172 11480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 19112 24172 19152 24212
rect 19194 24172 19234 24212
rect 19276 24172 19316 24212
rect 19358 24172 19398 24212
rect 19440 24172 19480 24212
rect 23112 24172 23152 24212
rect 23194 24172 23234 24212
rect 23276 24172 23316 24212
rect 23358 24172 23398 24212
rect 23440 24172 23480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 31112 24172 31152 24212
rect 31194 24172 31234 24212
rect 31276 24172 31316 24212
rect 31358 24172 31398 24212
rect 31440 24172 31480 24212
rect 35112 24172 35152 24212
rect 35194 24172 35234 24212
rect 35276 24172 35316 24212
rect 35358 24172 35398 24212
rect 35440 24172 35480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 43112 24172 43152 24212
rect 43194 24172 43234 24212
rect 43276 24172 43316 24212
rect 43358 24172 43398 24212
rect 43440 24172 43480 24212
rect 47112 24172 47152 24212
rect 47194 24172 47234 24212
rect 47276 24172 47316 24212
rect 47358 24172 47398 24212
rect 47440 24172 47480 24212
rect 51112 24172 51152 24212
rect 51194 24172 51234 24212
rect 51276 24172 51316 24212
rect 51358 24172 51398 24212
rect 51440 24172 51480 24212
rect 55112 24172 55152 24212
rect 55194 24172 55234 24212
rect 55276 24172 55316 24212
rect 55358 24172 55398 24212
rect 55440 24172 55480 24212
rect 59112 24172 59152 24212
rect 59194 24172 59234 24212
rect 59276 24172 59316 24212
rect 59358 24172 59398 24212
rect 59440 24172 59480 24212
rect 63112 24172 63152 24212
rect 63194 24172 63234 24212
rect 63276 24172 63316 24212
rect 63358 24172 63398 24212
rect 63440 24172 63480 24212
rect 67112 24172 67152 24212
rect 67194 24172 67234 24212
rect 67276 24172 67316 24212
rect 67358 24172 67398 24212
rect 67440 24172 67480 24212
rect 652 24088 692 24128
rect 844 23752 884 23792
rect 2092 23752 2132 23792
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 8352 23416 8392 23456
rect 8434 23416 8474 23456
rect 8516 23416 8556 23456
rect 8598 23416 8638 23456
rect 8680 23416 8720 23456
rect 12352 23416 12392 23456
rect 12434 23416 12474 23456
rect 12516 23416 12556 23456
rect 12598 23416 12638 23456
rect 12680 23416 12720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 20352 23416 20392 23456
rect 20434 23416 20474 23456
rect 20516 23416 20556 23456
rect 20598 23416 20638 23456
rect 20680 23416 20720 23456
rect 24352 23416 24392 23456
rect 24434 23416 24474 23456
rect 24516 23416 24556 23456
rect 24598 23416 24638 23456
rect 24680 23416 24720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 32352 23416 32392 23456
rect 32434 23416 32474 23456
rect 32516 23416 32556 23456
rect 32598 23416 32638 23456
rect 32680 23416 32720 23456
rect 36352 23416 36392 23456
rect 36434 23416 36474 23456
rect 36516 23416 36556 23456
rect 36598 23416 36638 23456
rect 36680 23416 36720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 44352 23416 44392 23456
rect 44434 23416 44474 23456
rect 44516 23416 44556 23456
rect 44598 23416 44638 23456
rect 44680 23416 44720 23456
rect 48352 23416 48392 23456
rect 48434 23416 48474 23456
rect 48516 23416 48556 23456
rect 48598 23416 48638 23456
rect 48680 23416 48720 23456
rect 52352 23416 52392 23456
rect 52434 23416 52474 23456
rect 52516 23416 52556 23456
rect 52598 23416 52638 23456
rect 52680 23416 52720 23456
rect 56352 23416 56392 23456
rect 56434 23416 56474 23456
rect 56516 23416 56556 23456
rect 56598 23416 56638 23456
rect 56680 23416 56720 23456
rect 60352 23416 60392 23456
rect 60434 23416 60474 23456
rect 60516 23416 60556 23456
rect 60598 23416 60638 23456
rect 60680 23416 60720 23456
rect 64352 23416 64392 23456
rect 64434 23416 64474 23456
rect 64516 23416 64556 23456
rect 64598 23416 64638 23456
rect 64680 23416 64720 23456
rect 68352 23416 68392 23456
rect 68434 23416 68474 23456
rect 68516 23416 68556 23456
rect 68598 23416 68638 23456
rect 68680 23416 68720 23456
rect 70924 27616 70964 27656
rect 70732 26776 70772 26816
rect 71116 26776 71156 26816
rect 71020 26272 71060 26312
rect 70828 26188 70868 26228
rect 70636 26104 70676 26144
rect 70924 26104 70964 26144
rect 71116 26104 71156 26144
rect 71404 26608 71444 26648
rect 71308 26524 71348 26564
rect 71404 26440 71444 26480
rect 70444 25348 70484 25388
rect 71308 25936 71348 25976
rect 70924 25264 70964 25304
rect 71308 25180 71348 25220
rect 72364 32908 72404 32948
rect 72652 32908 72692 32948
rect 73036 32908 73076 32948
rect 73228 32908 73268 32948
rect 72268 32824 72308 32864
rect 72460 32488 72500 32528
rect 73132 32488 73172 32528
rect 72415 32320 72455 32360
rect 72844 32320 72884 32360
rect 72815 32152 72855 32192
rect 72705 32068 72745 32108
rect 73215 32320 73255 32360
rect 74188 33580 74228 33620
rect 74476 33580 74516 33620
rect 74860 33580 74900 33620
rect 75340 33580 75380 33620
rect 73612 32824 73652 32864
rect 73996 32824 74036 32864
rect 73900 32656 73940 32696
rect 74188 32824 74228 32864
rect 74188 32656 74228 32696
rect 74668 33244 74708 33284
rect 74380 32908 74420 32948
rect 74668 32656 74708 32696
rect 74860 32908 74900 32948
rect 75148 32908 75188 32948
rect 75052 32656 75092 32696
rect 75820 33580 75860 33620
rect 76204 33580 76244 33620
rect 75436 33160 75476 33200
rect 75436 32656 75476 32696
rect 76012 32992 76052 33032
rect 75820 32908 75860 32948
rect 75105 32068 75145 32108
rect 75340 32068 75380 32108
rect 75905 32236 75945 32276
rect 77068 33580 77108 33620
rect 77452 33580 77492 33620
rect 77836 33580 77876 33620
rect 76300 33160 76340 33200
rect 76204 33076 76244 33116
rect 76204 32824 76244 32864
rect 76300 32656 76340 32696
rect 76588 32992 76628 33032
rect 76588 32824 76628 32864
rect 76876 32992 76916 33032
rect 76876 32824 76916 32864
rect 76972 32740 77012 32780
rect 76780 32656 76820 32696
rect 76492 32236 76532 32276
rect 76705 32068 76745 32108
rect 77452 32992 77492 33032
rect 77260 32908 77300 32948
rect 77548 32824 77588 32864
rect 77505 32320 77545 32360
rect 77068 32152 77108 32192
rect 76972 32068 77012 32108
rect 77836 32992 77876 33032
rect 77836 32656 77876 32696
rect 77740 32152 77780 32192
rect 78604 33580 78644 33620
rect 78988 33580 79028 33620
rect 79372 33580 79412 33620
rect 78124 32992 78164 33032
rect 78412 32992 78452 33032
rect 78316 32824 78356 32864
rect 78028 32404 78068 32444
rect 78305 32236 78345 32276
rect 78700 32908 78740 32948
rect 78700 32740 78740 32780
rect 79084 32992 79124 33032
rect 78988 32824 79028 32864
rect 79180 32236 79220 32276
rect 79372 32908 79412 32948
rect 79756 33580 79796 33620
rect 80332 33580 80372 33620
rect 79468 32656 79508 32696
rect 80524 33496 80564 33536
rect 80908 33496 80948 33536
rect 79756 32908 79796 32948
rect 79660 32824 79700 32864
rect 79756 32320 79796 32360
rect 80044 32908 80084 32948
rect 80236 32908 80276 32948
rect 80620 32908 80660 32948
rect 81292 33580 81332 33620
rect 82444 33580 82484 33620
rect 83116 33580 83156 33620
rect 81676 33496 81716 33536
rect 82060 33496 82100 33536
rect 82252 33496 82292 33536
rect 81100 33244 81140 33284
rect 81100 32908 81140 32948
rect 81004 32824 81044 32864
rect 79948 32656 79988 32696
rect 80236 32656 80276 32696
rect 80332 32320 80372 32360
rect 80705 32320 80745 32360
rect 81105 32236 81145 32276
rect 81388 32908 81428 32948
rect 81484 32740 81524 32780
rect 81292 32320 81332 32360
rect 81580 32236 81620 32276
rect 82828 33496 82868 33536
rect 82252 32908 82292 32948
rect 82348 32824 82388 32864
rect 82305 32320 82345 32360
rect 81905 32068 81945 32108
rect 82636 32656 82676 32696
rect 82828 32320 82868 32360
rect 83212 33496 83252 33536
rect 83500 33496 83540 33536
rect 83116 33160 83156 33200
rect 83308 32992 83348 33032
rect 83116 32740 83156 32780
rect 82540 32068 82580 32108
rect 83596 33076 83636 33116
rect 83596 32908 83636 32948
rect 83505 32320 83545 32360
rect 83884 32992 83924 33032
rect 83788 32824 83828 32864
rect 83884 32656 83924 32696
rect 84172 32992 84212 33032
rect 84460 32992 84500 33032
rect 84268 32740 84308 32780
rect 84076 32320 84116 32360
rect 84364 32656 84404 32696
rect 84652 33160 84692 33200
rect 84748 32992 84788 33032
rect 84844 32908 84884 32948
rect 85132 33076 85172 33116
rect 85036 32992 85076 33032
rect 85132 32824 85172 32864
rect 85105 32320 85145 32360
rect 84705 32068 84745 32108
rect 85900 33580 85940 33620
rect 86284 33580 86324 33620
rect 86668 33580 86708 33620
rect 85420 32824 85460 32864
rect 85420 32656 85460 32696
rect 85324 32068 85364 32108
rect 87436 33580 87476 33620
rect 85900 32992 85940 33032
rect 85708 32824 85748 32864
rect 85996 32824 86036 32864
rect 85900 32740 85940 32780
rect 85612 32320 85652 32360
rect 85905 32320 85945 32360
rect 86284 33244 86324 33284
rect 86284 32740 86324 32780
rect 87052 33412 87092 33452
rect 86860 33244 86900 33284
rect 86476 33160 86516 33200
rect 87052 33160 87092 33200
rect 86860 33076 86900 33116
rect 86668 32992 86708 33032
rect 86668 32656 86708 32696
rect 86764 32320 86804 32360
rect 86956 32908 86996 32948
rect 87820 33580 87860 33620
rect 87340 33160 87380 33200
rect 87244 33076 87284 33116
rect 87244 32824 87284 32864
rect 87105 32320 87145 32360
rect 87628 33160 87668 33200
rect 87628 32656 87668 32696
rect 87532 32320 87572 32360
rect 87916 33244 87956 33284
rect 88588 33580 88628 33620
rect 88972 33580 89012 33620
rect 89356 33580 89396 33620
rect 88300 33160 88340 33200
rect 88012 33076 88052 33116
rect 87916 32740 87956 32780
rect 88108 32992 88148 33032
rect 88396 33076 88436 33116
rect 88396 32908 88436 32948
rect 88684 32992 88724 33032
rect 88588 32824 88628 32864
rect 88780 32824 88820 32864
rect 88305 32068 88345 32108
rect 88972 33244 89012 33284
rect 89548 33580 89588 33620
rect 89548 33244 89588 33284
rect 90124 33580 90164 33620
rect 90508 33580 90548 33620
rect 90892 33580 90932 33620
rect 91180 33580 91220 33620
rect 89740 33160 89780 33200
rect 89452 32992 89492 33032
rect 89740 32992 89780 33032
rect 89068 32908 89108 32948
rect 89644 32824 89684 32864
rect 89932 32992 89972 33032
rect 90028 32908 90068 32948
rect 89932 32656 89972 32696
rect 89356 32068 89396 32108
rect 89505 32068 89545 32108
rect 90316 33244 90356 33284
rect 90412 32824 90452 32864
rect 90220 32068 90260 32108
rect 90700 33160 90740 33200
rect 90892 33076 90932 33116
rect 90796 32656 90836 32696
rect 91180 32992 91220 33032
rect 91084 32908 91124 32948
rect 91468 32992 91508 33032
rect 91372 32824 91412 32864
rect 91468 32572 91508 32612
rect 91105 32236 91145 32276
rect 91660 33748 91700 33788
rect 91852 33580 91892 33620
rect 91756 33076 91796 33116
rect 91852 32908 91892 32948
rect 91660 32656 91700 32696
rect 92524 33496 92564 33536
rect 92332 33160 92372 33200
rect 92332 32824 92372 32864
rect 91852 32236 91892 32276
rect 93196 33580 93236 33620
rect 93388 33580 93428 33620
rect 92812 33496 92852 33536
rect 92620 33412 92660 33452
rect 92812 33076 92852 33116
rect 92716 32992 92756 33032
rect 92620 32740 92660 32780
rect 93004 33076 93044 33116
rect 93100 32908 93140 32948
rect 93004 32656 93044 32696
rect 93388 33160 93428 33200
rect 93292 32824 93332 32864
rect 95500 33748 95540 33788
rect 95308 33664 95348 33704
rect 93580 33580 93620 33620
rect 94252 33580 94292 33620
rect 93772 33496 93812 33536
rect 93676 33160 93716 33200
rect 93772 32992 93812 33032
rect 93580 32740 93620 32780
rect 93505 32068 93545 32108
rect 93868 32740 93908 32780
rect 93772 32068 93812 32108
rect 94636 33580 94676 33620
rect 96076 33664 96116 33704
rect 96460 33664 96500 33704
rect 94348 33160 94388 33200
rect 94156 32908 94196 32948
rect 94252 32824 94292 32864
rect 95692 33580 95732 33620
rect 94636 33076 94676 33116
rect 94540 32740 94580 32780
rect 94828 33160 94868 33200
rect 95212 33076 95252 33116
rect 94924 32992 94964 33032
rect 95116 32908 95156 32948
rect 95020 32824 95060 32864
rect 94705 32068 94745 32108
rect 95500 33076 95540 33116
rect 95500 32656 95540 32696
rect 95404 32068 95444 32108
rect 95692 33076 95732 33116
rect 96748 33580 96788 33620
rect 96940 33580 96980 33620
rect 95788 32824 95828 32864
rect 96076 32824 96116 32864
rect 95980 32740 96020 32780
rect 95905 32236 95945 32276
rect 96364 32824 96404 32864
rect 96940 32824 96980 32864
rect 97228 33412 97268 33452
rect 97132 32824 97172 32864
rect 96268 32236 96308 32276
rect 96305 32068 96345 32108
rect 96705 32152 96745 32192
rect 97516 32824 97556 32864
rect 97132 32236 97172 32276
rect 97105 32068 97145 32108
rect 97516 32656 97556 32696
rect 97420 32152 97460 32192
rect 97804 32824 97844 32864
rect 98380 33580 98420 33620
rect 98092 32824 98132 32864
rect 97996 32656 98036 32696
rect 97708 32068 97748 32108
rect 97905 32068 97945 32108
rect 98305 32152 98345 32192
rect 71884 26692 71924 26732
rect 72305 26608 72345 26648
rect 72705 26524 72745 26564
rect 72415 26440 72455 26480
rect 73105 26440 73145 26480
rect 72844 26272 72884 26312
rect 71884 26020 71924 26060
rect 73132 25684 73172 25724
rect 72748 25516 72788 25556
rect 73420 26188 73460 26228
rect 73612 26104 73652 26144
rect 73228 25516 73268 25556
rect 73804 25684 73844 25724
rect 72940 25348 72980 25388
rect 72652 25264 72692 25304
rect 73324 25264 73364 25304
rect 73324 24928 73364 24968
rect 73516 24760 73556 24800
rect 71788 24676 71828 24716
rect 71020 24592 71060 24632
rect 73228 24592 73268 24632
rect 652 23248 692 23288
rect 2092 23248 2132 23288
rect 69292 23248 69332 23288
rect 844 23080 884 23120
rect 1996 23080 2036 23120
rect 556 22408 596 22448
rect 652 21568 692 21608
rect 652 20728 692 20768
rect 652 19888 692 19928
rect 652 19048 692 19088
rect 652 18208 692 18248
rect 652 17368 692 17408
rect 652 16528 692 16568
rect 652 15688 692 15728
rect 844 14932 884 14972
rect 1420 14932 1460 14972
rect 652 14848 692 14888
rect 1996 14764 2036 14804
rect 652 14008 692 14048
rect 1228 13924 1268 13964
rect 1804 13924 1844 13964
rect 844 13336 884 13376
rect 1612 13336 1652 13376
rect 652 13168 692 13208
rect 652 12328 692 12368
rect 652 11488 692 11528
rect 652 10732 692 10772
rect 844 10480 884 10520
rect 1420 10480 1460 10520
rect 1228 10228 1268 10268
rect 1612 10228 1652 10268
rect 652 9808 692 9848
rect 652 8968 692 9008
rect 748 8800 788 8840
rect 1516 8800 1556 8840
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 7112 22660 7152 22700
rect 7194 22660 7234 22700
rect 7276 22660 7316 22700
rect 7358 22660 7398 22700
rect 7440 22660 7480 22700
rect 11112 22660 11152 22700
rect 11194 22660 11234 22700
rect 11276 22660 11316 22700
rect 11358 22660 11398 22700
rect 11440 22660 11480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 19112 22660 19152 22700
rect 19194 22660 19234 22700
rect 19276 22660 19316 22700
rect 19358 22660 19398 22700
rect 19440 22660 19480 22700
rect 23112 22660 23152 22700
rect 23194 22660 23234 22700
rect 23276 22660 23316 22700
rect 23358 22660 23398 22700
rect 23440 22660 23480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 31112 22660 31152 22700
rect 31194 22660 31234 22700
rect 31276 22660 31316 22700
rect 31358 22660 31398 22700
rect 31440 22660 31480 22700
rect 35112 22660 35152 22700
rect 35194 22660 35234 22700
rect 35276 22660 35316 22700
rect 35358 22660 35398 22700
rect 35440 22660 35480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 43112 22660 43152 22700
rect 43194 22660 43234 22700
rect 43276 22660 43316 22700
rect 43358 22660 43398 22700
rect 43440 22660 43480 22700
rect 47112 22660 47152 22700
rect 47194 22660 47234 22700
rect 47276 22660 47316 22700
rect 47358 22660 47398 22700
rect 47440 22660 47480 22700
rect 51112 22660 51152 22700
rect 51194 22660 51234 22700
rect 51276 22660 51316 22700
rect 51358 22660 51398 22700
rect 51440 22660 51480 22700
rect 55112 22660 55152 22700
rect 55194 22660 55234 22700
rect 55276 22660 55316 22700
rect 55358 22660 55398 22700
rect 55440 22660 55480 22700
rect 59112 22660 59152 22700
rect 59194 22660 59234 22700
rect 59276 22660 59316 22700
rect 59358 22660 59398 22700
rect 59440 22660 59480 22700
rect 63112 22660 63152 22700
rect 63194 22660 63234 22700
rect 63276 22660 63316 22700
rect 63358 22660 63398 22700
rect 63440 22660 63480 22700
rect 67112 22660 67152 22700
rect 67194 22660 67234 22700
rect 67276 22660 67316 22700
rect 67358 22660 67398 22700
rect 67440 22660 67480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 8352 21904 8392 21944
rect 8434 21904 8474 21944
rect 8516 21904 8556 21944
rect 8598 21904 8638 21944
rect 8680 21904 8720 21944
rect 12352 21904 12392 21944
rect 12434 21904 12474 21944
rect 12516 21904 12556 21944
rect 12598 21904 12638 21944
rect 12680 21904 12720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 20352 21904 20392 21944
rect 20434 21904 20474 21944
rect 20516 21904 20556 21944
rect 20598 21904 20638 21944
rect 20680 21904 20720 21944
rect 24352 21904 24392 21944
rect 24434 21904 24474 21944
rect 24516 21904 24556 21944
rect 24598 21904 24638 21944
rect 24680 21904 24720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 32352 21904 32392 21944
rect 32434 21904 32474 21944
rect 32516 21904 32556 21944
rect 32598 21904 32638 21944
rect 32680 21904 32720 21944
rect 36352 21904 36392 21944
rect 36434 21904 36474 21944
rect 36516 21904 36556 21944
rect 36598 21904 36638 21944
rect 36680 21904 36720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 44352 21904 44392 21944
rect 44434 21904 44474 21944
rect 44516 21904 44556 21944
rect 44598 21904 44638 21944
rect 44680 21904 44720 21944
rect 48352 21904 48392 21944
rect 48434 21904 48474 21944
rect 48516 21904 48556 21944
rect 48598 21904 48638 21944
rect 48680 21904 48720 21944
rect 52352 21904 52392 21944
rect 52434 21904 52474 21944
rect 52516 21904 52556 21944
rect 52598 21904 52638 21944
rect 52680 21904 52720 21944
rect 56352 21904 56392 21944
rect 56434 21904 56474 21944
rect 56516 21904 56556 21944
rect 56598 21904 56638 21944
rect 56680 21904 56720 21944
rect 60352 21904 60392 21944
rect 60434 21904 60474 21944
rect 60516 21904 60556 21944
rect 60598 21904 60638 21944
rect 60680 21904 60720 21944
rect 64352 21904 64392 21944
rect 64434 21904 64474 21944
rect 64516 21904 64556 21944
rect 64598 21904 64638 21944
rect 64680 21904 64720 21944
rect 68352 21904 68392 21944
rect 68434 21904 68474 21944
rect 68516 21904 68556 21944
rect 68598 21904 68638 21944
rect 68680 21904 68720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 7112 21148 7152 21188
rect 7194 21148 7234 21188
rect 7276 21148 7316 21188
rect 7358 21148 7398 21188
rect 7440 21148 7480 21188
rect 11112 21148 11152 21188
rect 11194 21148 11234 21188
rect 11276 21148 11316 21188
rect 11358 21148 11398 21188
rect 11440 21148 11480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 19112 21148 19152 21188
rect 19194 21148 19234 21188
rect 19276 21148 19316 21188
rect 19358 21148 19398 21188
rect 19440 21148 19480 21188
rect 23112 21148 23152 21188
rect 23194 21148 23234 21188
rect 23276 21148 23316 21188
rect 23358 21148 23398 21188
rect 23440 21148 23480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 31112 21148 31152 21188
rect 31194 21148 31234 21188
rect 31276 21148 31316 21188
rect 31358 21148 31398 21188
rect 31440 21148 31480 21188
rect 35112 21148 35152 21188
rect 35194 21148 35234 21188
rect 35276 21148 35316 21188
rect 35358 21148 35398 21188
rect 35440 21148 35480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 43112 21148 43152 21188
rect 43194 21148 43234 21188
rect 43276 21148 43316 21188
rect 43358 21148 43398 21188
rect 43440 21148 43480 21188
rect 47112 21148 47152 21188
rect 47194 21148 47234 21188
rect 47276 21148 47316 21188
rect 47358 21148 47398 21188
rect 47440 21148 47480 21188
rect 51112 21148 51152 21188
rect 51194 21148 51234 21188
rect 51276 21148 51316 21188
rect 51358 21148 51398 21188
rect 51440 21148 51480 21188
rect 55112 21148 55152 21188
rect 55194 21148 55234 21188
rect 55276 21148 55316 21188
rect 55358 21148 55398 21188
rect 55440 21148 55480 21188
rect 59112 21148 59152 21188
rect 59194 21148 59234 21188
rect 59276 21148 59316 21188
rect 59358 21148 59398 21188
rect 59440 21148 59480 21188
rect 63112 21148 63152 21188
rect 63194 21148 63234 21188
rect 63276 21148 63316 21188
rect 63358 21148 63398 21188
rect 63440 21148 63480 21188
rect 67112 21148 67152 21188
rect 67194 21148 67234 21188
rect 67276 21148 67316 21188
rect 67358 21148 67398 21188
rect 67440 21148 67480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 8352 20392 8392 20432
rect 8434 20392 8474 20432
rect 8516 20392 8556 20432
rect 8598 20392 8638 20432
rect 8680 20392 8720 20432
rect 12352 20392 12392 20432
rect 12434 20392 12474 20432
rect 12516 20392 12556 20432
rect 12598 20392 12638 20432
rect 12680 20392 12720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 20352 20392 20392 20432
rect 20434 20392 20474 20432
rect 20516 20392 20556 20432
rect 20598 20392 20638 20432
rect 20680 20392 20720 20432
rect 24352 20392 24392 20432
rect 24434 20392 24474 20432
rect 24516 20392 24556 20432
rect 24598 20392 24638 20432
rect 24680 20392 24720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 32352 20392 32392 20432
rect 32434 20392 32474 20432
rect 32516 20392 32556 20432
rect 32598 20392 32638 20432
rect 32680 20392 32720 20432
rect 36352 20392 36392 20432
rect 36434 20392 36474 20432
rect 36516 20392 36556 20432
rect 36598 20392 36638 20432
rect 36680 20392 36720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 44352 20392 44392 20432
rect 44434 20392 44474 20432
rect 44516 20392 44556 20432
rect 44598 20392 44638 20432
rect 44680 20392 44720 20432
rect 48352 20392 48392 20432
rect 48434 20392 48474 20432
rect 48516 20392 48556 20432
rect 48598 20392 48638 20432
rect 48680 20392 48720 20432
rect 52352 20392 52392 20432
rect 52434 20392 52474 20432
rect 52516 20392 52556 20432
rect 52598 20392 52638 20432
rect 52680 20392 52720 20432
rect 56352 20392 56392 20432
rect 56434 20392 56474 20432
rect 56516 20392 56556 20432
rect 56598 20392 56638 20432
rect 56680 20392 56720 20432
rect 60352 20392 60392 20432
rect 60434 20392 60474 20432
rect 60516 20392 60556 20432
rect 60598 20392 60638 20432
rect 60680 20392 60720 20432
rect 64352 20392 64392 20432
rect 64434 20392 64474 20432
rect 64516 20392 64556 20432
rect 64598 20392 64638 20432
rect 64680 20392 64720 20432
rect 68352 20392 68392 20432
rect 68434 20392 68474 20432
rect 68516 20392 68556 20432
rect 68598 20392 68638 20432
rect 68680 20392 68720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 7112 19636 7152 19676
rect 7194 19636 7234 19676
rect 7276 19636 7316 19676
rect 7358 19636 7398 19676
rect 7440 19636 7480 19676
rect 11112 19636 11152 19676
rect 11194 19636 11234 19676
rect 11276 19636 11316 19676
rect 11358 19636 11398 19676
rect 11440 19636 11480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 19112 19636 19152 19676
rect 19194 19636 19234 19676
rect 19276 19636 19316 19676
rect 19358 19636 19398 19676
rect 19440 19636 19480 19676
rect 23112 19636 23152 19676
rect 23194 19636 23234 19676
rect 23276 19636 23316 19676
rect 23358 19636 23398 19676
rect 23440 19636 23480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 31112 19636 31152 19676
rect 31194 19636 31234 19676
rect 31276 19636 31316 19676
rect 31358 19636 31398 19676
rect 31440 19636 31480 19676
rect 35112 19636 35152 19676
rect 35194 19636 35234 19676
rect 35276 19636 35316 19676
rect 35358 19636 35398 19676
rect 35440 19636 35480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 43112 19636 43152 19676
rect 43194 19636 43234 19676
rect 43276 19636 43316 19676
rect 43358 19636 43398 19676
rect 43440 19636 43480 19676
rect 47112 19636 47152 19676
rect 47194 19636 47234 19676
rect 47276 19636 47316 19676
rect 47358 19636 47398 19676
rect 47440 19636 47480 19676
rect 51112 19636 51152 19676
rect 51194 19636 51234 19676
rect 51276 19636 51316 19676
rect 51358 19636 51398 19676
rect 51440 19636 51480 19676
rect 55112 19636 55152 19676
rect 55194 19636 55234 19676
rect 55276 19636 55316 19676
rect 55358 19636 55398 19676
rect 55440 19636 55480 19676
rect 59112 19636 59152 19676
rect 59194 19636 59234 19676
rect 59276 19636 59316 19676
rect 59358 19636 59398 19676
rect 59440 19636 59480 19676
rect 63112 19636 63152 19676
rect 63194 19636 63234 19676
rect 63276 19636 63316 19676
rect 63358 19636 63398 19676
rect 63440 19636 63480 19676
rect 67112 19636 67152 19676
rect 67194 19636 67234 19676
rect 67276 19636 67316 19676
rect 67358 19636 67398 19676
rect 67440 19636 67480 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 8352 18880 8392 18920
rect 8434 18880 8474 18920
rect 8516 18880 8556 18920
rect 8598 18880 8638 18920
rect 8680 18880 8720 18920
rect 12352 18880 12392 18920
rect 12434 18880 12474 18920
rect 12516 18880 12556 18920
rect 12598 18880 12638 18920
rect 12680 18880 12720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 20352 18880 20392 18920
rect 20434 18880 20474 18920
rect 20516 18880 20556 18920
rect 20598 18880 20638 18920
rect 20680 18880 20720 18920
rect 24352 18880 24392 18920
rect 24434 18880 24474 18920
rect 24516 18880 24556 18920
rect 24598 18880 24638 18920
rect 24680 18880 24720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 32352 18880 32392 18920
rect 32434 18880 32474 18920
rect 32516 18880 32556 18920
rect 32598 18880 32638 18920
rect 32680 18880 32720 18920
rect 36352 18880 36392 18920
rect 36434 18880 36474 18920
rect 36516 18880 36556 18920
rect 36598 18880 36638 18920
rect 36680 18880 36720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 44352 18880 44392 18920
rect 44434 18880 44474 18920
rect 44516 18880 44556 18920
rect 44598 18880 44638 18920
rect 44680 18880 44720 18920
rect 48352 18880 48392 18920
rect 48434 18880 48474 18920
rect 48516 18880 48556 18920
rect 48598 18880 48638 18920
rect 48680 18880 48720 18920
rect 52352 18880 52392 18920
rect 52434 18880 52474 18920
rect 52516 18880 52556 18920
rect 52598 18880 52638 18920
rect 52680 18880 52720 18920
rect 56352 18880 56392 18920
rect 56434 18880 56474 18920
rect 56516 18880 56556 18920
rect 56598 18880 56638 18920
rect 56680 18880 56720 18920
rect 60352 18880 60392 18920
rect 60434 18880 60474 18920
rect 60516 18880 60556 18920
rect 60598 18880 60638 18920
rect 60680 18880 60720 18920
rect 64352 18880 64392 18920
rect 64434 18880 64474 18920
rect 64516 18880 64556 18920
rect 64598 18880 64638 18920
rect 64680 18880 64720 18920
rect 68352 18880 68392 18920
rect 68434 18880 68474 18920
rect 68516 18880 68556 18920
rect 68598 18880 68638 18920
rect 68680 18880 68720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 7112 18124 7152 18164
rect 7194 18124 7234 18164
rect 7276 18124 7316 18164
rect 7358 18124 7398 18164
rect 7440 18124 7480 18164
rect 11112 18124 11152 18164
rect 11194 18124 11234 18164
rect 11276 18124 11316 18164
rect 11358 18124 11398 18164
rect 11440 18124 11480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 19112 18124 19152 18164
rect 19194 18124 19234 18164
rect 19276 18124 19316 18164
rect 19358 18124 19398 18164
rect 19440 18124 19480 18164
rect 23112 18124 23152 18164
rect 23194 18124 23234 18164
rect 23276 18124 23316 18164
rect 23358 18124 23398 18164
rect 23440 18124 23480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 31112 18124 31152 18164
rect 31194 18124 31234 18164
rect 31276 18124 31316 18164
rect 31358 18124 31398 18164
rect 31440 18124 31480 18164
rect 35112 18124 35152 18164
rect 35194 18124 35234 18164
rect 35276 18124 35316 18164
rect 35358 18124 35398 18164
rect 35440 18124 35480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 43112 18124 43152 18164
rect 43194 18124 43234 18164
rect 43276 18124 43316 18164
rect 43358 18124 43398 18164
rect 43440 18124 43480 18164
rect 47112 18124 47152 18164
rect 47194 18124 47234 18164
rect 47276 18124 47316 18164
rect 47358 18124 47398 18164
rect 47440 18124 47480 18164
rect 51112 18124 51152 18164
rect 51194 18124 51234 18164
rect 51276 18124 51316 18164
rect 51358 18124 51398 18164
rect 51440 18124 51480 18164
rect 55112 18124 55152 18164
rect 55194 18124 55234 18164
rect 55276 18124 55316 18164
rect 55358 18124 55398 18164
rect 55440 18124 55480 18164
rect 59112 18124 59152 18164
rect 59194 18124 59234 18164
rect 59276 18124 59316 18164
rect 59358 18124 59398 18164
rect 59440 18124 59480 18164
rect 63112 18124 63152 18164
rect 63194 18124 63234 18164
rect 63276 18124 63316 18164
rect 63358 18124 63398 18164
rect 63440 18124 63480 18164
rect 67112 18124 67152 18164
rect 67194 18124 67234 18164
rect 67276 18124 67316 18164
rect 67358 18124 67398 18164
rect 67440 18124 67480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 8352 17368 8392 17408
rect 8434 17368 8474 17408
rect 8516 17368 8556 17408
rect 8598 17368 8638 17408
rect 8680 17368 8720 17408
rect 12352 17368 12392 17408
rect 12434 17368 12474 17408
rect 12516 17368 12556 17408
rect 12598 17368 12638 17408
rect 12680 17368 12720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 20352 17368 20392 17408
rect 20434 17368 20474 17408
rect 20516 17368 20556 17408
rect 20598 17368 20638 17408
rect 20680 17368 20720 17408
rect 24352 17368 24392 17408
rect 24434 17368 24474 17408
rect 24516 17368 24556 17408
rect 24598 17368 24638 17408
rect 24680 17368 24720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 32352 17368 32392 17408
rect 32434 17368 32474 17408
rect 32516 17368 32556 17408
rect 32598 17368 32638 17408
rect 32680 17368 32720 17408
rect 36352 17368 36392 17408
rect 36434 17368 36474 17408
rect 36516 17368 36556 17408
rect 36598 17368 36638 17408
rect 36680 17368 36720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 44352 17368 44392 17408
rect 44434 17368 44474 17408
rect 44516 17368 44556 17408
rect 44598 17368 44638 17408
rect 44680 17368 44720 17408
rect 48352 17368 48392 17408
rect 48434 17368 48474 17408
rect 48516 17368 48556 17408
rect 48598 17368 48638 17408
rect 48680 17368 48720 17408
rect 52352 17368 52392 17408
rect 52434 17368 52474 17408
rect 52516 17368 52556 17408
rect 52598 17368 52638 17408
rect 52680 17368 52720 17408
rect 56352 17368 56392 17408
rect 56434 17368 56474 17408
rect 56516 17368 56556 17408
rect 56598 17368 56638 17408
rect 56680 17368 56720 17408
rect 60352 17368 60392 17408
rect 60434 17368 60474 17408
rect 60516 17368 60556 17408
rect 60598 17368 60638 17408
rect 60680 17368 60720 17408
rect 64352 17368 64392 17408
rect 64434 17368 64474 17408
rect 64516 17368 64556 17408
rect 64598 17368 64638 17408
rect 64680 17368 64720 17408
rect 68352 17368 68392 17408
rect 68434 17368 68474 17408
rect 68516 17368 68556 17408
rect 68598 17368 68638 17408
rect 68680 17368 68720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 7112 16612 7152 16652
rect 7194 16612 7234 16652
rect 7276 16612 7316 16652
rect 7358 16612 7398 16652
rect 7440 16612 7480 16652
rect 11112 16612 11152 16652
rect 11194 16612 11234 16652
rect 11276 16612 11316 16652
rect 11358 16612 11398 16652
rect 11440 16612 11480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 19112 16612 19152 16652
rect 19194 16612 19234 16652
rect 19276 16612 19316 16652
rect 19358 16612 19398 16652
rect 19440 16612 19480 16652
rect 23112 16612 23152 16652
rect 23194 16612 23234 16652
rect 23276 16612 23316 16652
rect 23358 16612 23398 16652
rect 23440 16612 23480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 31112 16612 31152 16652
rect 31194 16612 31234 16652
rect 31276 16612 31316 16652
rect 31358 16612 31398 16652
rect 31440 16612 31480 16652
rect 35112 16612 35152 16652
rect 35194 16612 35234 16652
rect 35276 16612 35316 16652
rect 35358 16612 35398 16652
rect 35440 16612 35480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 43112 16612 43152 16652
rect 43194 16612 43234 16652
rect 43276 16612 43316 16652
rect 43358 16612 43398 16652
rect 43440 16612 43480 16652
rect 47112 16612 47152 16652
rect 47194 16612 47234 16652
rect 47276 16612 47316 16652
rect 47358 16612 47398 16652
rect 47440 16612 47480 16652
rect 51112 16612 51152 16652
rect 51194 16612 51234 16652
rect 51276 16612 51316 16652
rect 51358 16612 51398 16652
rect 51440 16612 51480 16652
rect 55112 16612 55152 16652
rect 55194 16612 55234 16652
rect 55276 16612 55316 16652
rect 55358 16612 55398 16652
rect 55440 16612 55480 16652
rect 59112 16612 59152 16652
rect 59194 16612 59234 16652
rect 59276 16612 59316 16652
rect 59358 16612 59398 16652
rect 59440 16612 59480 16652
rect 63112 16612 63152 16652
rect 63194 16612 63234 16652
rect 63276 16612 63316 16652
rect 63358 16612 63398 16652
rect 63440 16612 63480 16652
rect 67112 16612 67152 16652
rect 67194 16612 67234 16652
rect 67276 16612 67316 16652
rect 67358 16612 67398 16652
rect 67440 16612 67480 16652
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 8352 15856 8392 15896
rect 8434 15856 8474 15896
rect 8516 15856 8556 15896
rect 8598 15856 8638 15896
rect 8680 15856 8720 15896
rect 12352 15856 12392 15896
rect 12434 15856 12474 15896
rect 12516 15856 12556 15896
rect 12598 15856 12638 15896
rect 12680 15856 12720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 20352 15856 20392 15896
rect 20434 15856 20474 15896
rect 20516 15856 20556 15896
rect 20598 15856 20638 15896
rect 20680 15856 20720 15896
rect 24352 15856 24392 15896
rect 24434 15856 24474 15896
rect 24516 15856 24556 15896
rect 24598 15856 24638 15896
rect 24680 15856 24720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 32352 15856 32392 15896
rect 32434 15856 32474 15896
rect 32516 15856 32556 15896
rect 32598 15856 32638 15896
rect 32680 15856 32720 15896
rect 36352 15856 36392 15896
rect 36434 15856 36474 15896
rect 36516 15856 36556 15896
rect 36598 15856 36638 15896
rect 36680 15856 36720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 44352 15856 44392 15896
rect 44434 15856 44474 15896
rect 44516 15856 44556 15896
rect 44598 15856 44638 15896
rect 44680 15856 44720 15896
rect 48352 15856 48392 15896
rect 48434 15856 48474 15896
rect 48516 15856 48556 15896
rect 48598 15856 48638 15896
rect 48680 15856 48720 15896
rect 52352 15856 52392 15896
rect 52434 15856 52474 15896
rect 52516 15856 52556 15896
rect 52598 15856 52638 15896
rect 52680 15856 52720 15896
rect 56352 15856 56392 15896
rect 56434 15856 56474 15896
rect 56516 15856 56556 15896
rect 56598 15856 56638 15896
rect 56680 15856 56720 15896
rect 60352 15856 60392 15896
rect 60434 15856 60474 15896
rect 60516 15856 60556 15896
rect 60598 15856 60638 15896
rect 60680 15856 60720 15896
rect 64352 15856 64392 15896
rect 64434 15856 64474 15896
rect 64516 15856 64556 15896
rect 64598 15856 64638 15896
rect 64680 15856 64720 15896
rect 68352 15856 68392 15896
rect 68434 15856 68474 15896
rect 68516 15856 68556 15896
rect 68598 15856 68638 15896
rect 68680 15856 68720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 7112 15100 7152 15140
rect 7194 15100 7234 15140
rect 7276 15100 7316 15140
rect 7358 15100 7398 15140
rect 7440 15100 7480 15140
rect 11112 15100 11152 15140
rect 11194 15100 11234 15140
rect 11276 15100 11316 15140
rect 11358 15100 11398 15140
rect 11440 15100 11480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 19112 15100 19152 15140
rect 19194 15100 19234 15140
rect 19276 15100 19316 15140
rect 19358 15100 19398 15140
rect 19440 15100 19480 15140
rect 23112 15100 23152 15140
rect 23194 15100 23234 15140
rect 23276 15100 23316 15140
rect 23358 15100 23398 15140
rect 23440 15100 23480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 31112 15100 31152 15140
rect 31194 15100 31234 15140
rect 31276 15100 31316 15140
rect 31358 15100 31398 15140
rect 31440 15100 31480 15140
rect 35112 15100 35152 15140
rect 35194 15100 35234 15140
rect 35276 15100 35316 15140
rect 35358 15100 35398 15140
rect 35440 15100 35480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 43112 15100 43152 15140
rect 43194 15100 43234 15140
rect 43276 15100 43316 15140
rect 43358 15100 43398 15140
rect 43440 15100 43480 15140
rect 47112 15100 47152 15140
rect 47194 15100 47234 15140
rect 47276 15100 47316 15140
rect 47358 15100 47398 15140
rect 47440 15100 47480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 55112 15100 55152 15140
rect 55194 15100 55234 15140
rect 55276 15100 55316 15140
rect 55358 15100 55398 15140
rect 55440 15100 55480 15140
rect 59112 15100 59152 15140
rect 59194 15100 59234 15140
rect 59276 15100 59316 15140
rect 59358 15100 59398 15140
rect 59440 15100 59480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 67112 15100 67152 15140
rect 67194 15100 67234 15140
rect 67276 15100 67316 15140
rect 67358 15100 67398 15140
rect 67440 15100 67480 15140
rect 73612 24508 73652 24548
rect 73900 25096 73940 25136
rect 75215 26440 75255 26480
rect 74284 25096 74324 25136
rect 73996 24928 74036 24968
rect 73996 24676 74036 24716
rect 74188 24676 74228 24716
rect 74668 26020 74708 26060
rect 76204 26440 76244 26480
rect 74860 25516 74900 25556
rect 74476 25348 74516 25388
rect 74668 25348 74708 25388
rect 74380 24760 74420 24800
rect 74284 24508 74324 24548
rect 74668 24508 74708 24548
rect 75244 25432 75284 25472
rect 75052 25348 75092 25388
rect 75532 25432 75572 25472
rect 75532 25264 75572 25304
rect 75916 25516 75956 25556
rect 76012 25432 76052 25472
rect 76012 25264 76052 25304
rect 76300 25264 76340 25304
rect 76492 25600 76532 25640
rect 76492 25432 76532 25472
rect 76588 25264 76628 25304
rect 77215 26440 77255 26480
rect 76876 25600 76916 25640
rect 76780 25516 76820 25556
rect 76780 25264 76820 25304
rect 76876 24928 76916 24968
rect 75724 24676 75764 24716
rect 77164 25516 77204 25556
rect 77068 24928 77108 24968
rect 77644 25516 77684 25556
rect 77548 25348 77588 25388
rect 75244 24508 75284 24548
rect 76012 24508 76052 24548
rect 76396 24508 76436 24548
rect 76876 24508 76916 24548
rect 77260 24508 77300 24548
rect 77740 25264 77780 25304
rect 78508 26440 78548 26480
rect 77932 25516 77972 25556
rect 78028 25264 78068 25304
rect 78316 25264 78356 25304
rect 78604 25516 78644 25556
rect 79756 25516 79796 25556
rect 78892 25264 78932 25304
rect 79372 25264 79412 25304
rect 79852 25264 79892 25304
rect 80044 25264 80084 25304
rect 77836 24508 77876 24548
rect 78220 24508 78260 24548
rect 78604 24508 78644 24548
rect 78988 24508 79028 24548
rect 79372 24508 79412 24548
rect 79756 24508 79796 24548
rect 80140 24508 80180 24548
rect 74380 24340 74420 24380
rect 74764 24340 74804 24380
rect 71112 24172 71152 24212
rect 71194 24172 71234 24212
rect 71276 24172 71316 24212
rect 71358 24172 71398 24212
rect 71440 24172 71480 24212
rect 75112 24172 75152 24212
rect 75194 24172 75234 24212
rect 75276 24172 75316 24212
rect 75358 24172 75398 24212
rect 75440 24172 75480 24212
rect 79112 24172 79152 24212
rect 79194 24172 79234 24212
rect 79276 24172 79316 24212
rect 79358 24172 79398 24212
rect 79440 24172 79480 24212
rect 81196 25348 81236 25388
rect 80428 25180 80468 25220
rect 80716 25180 80756 25220
rect 80908 25180 80948 25220
rect 81100 25180 81140 25220
rect 81580 25348 81620 25388
rect 81484 25180 81524 25220
rect 81388 24760 81428 24800
rect 80620 24340 80660 24380
rect 80332 23836 80372 23876
rect 80812 23836 80852 23876
rect 81388 23836 81428 23876
rect 81964 24760 82004 24800
rect 82252 25180 82292 25220
rect 82732 25180 82772 25220
rect 81676 23836 81716 23876
rect 82156 23836 82196 23876
rect 83692 25516 83732 25556
rect 83308 24508 83348 24548
rect 83788 25264 83828 25304
rect 83980 25516 84020 25556
rect 84076 25264 84116 25304
rect 84364 25264 84404 25304
rect 84652 25264 84692 25304
rect 84940 25264 84980 25304
rect 85132 25264 85172 25304
rect 83692 24508 83732 24548
rect 84268 24508 84308 24548
rect 84652 24508 84692 24548
rect 85036 24508 85076 24548
rect 83596 24340 83636 24380
rect 84076 24340 84116 24380
rect 83112 24172 83152 24212
rect 83194 24172 83234 24212
rect 83276 24172 83316 24212
rect 83358 24172 83398 24212
rect 83440 24172 83480 24212
rect 85516 25264 85556 25304
rect 85324 24508 85364 24548
rect 85900 25264 85940 25304
rect 86572 25264 86612 25304
rect 86092 24508 86132 24548
rect 86476 24508 86516 24548
rect 82444 23836 82484 23876
rect 84940 23836 84980 23876
rect 85708 23836 85748 23876
rect 86860 25516 86900 25556
rect 86956 25432 86996 25472
rect 86764 25264 86804 25304
rect 87148 25348 87188 25388
rect 87340 25348 87380 25388
rect 87532 25516 87572 25556
rect 87628 25264 87668 25304
rect 87916 25264 87956 25304
rect 86764 24508 86804 24548
rect 86956 24508 86996 24548
rect 87340 24508 87380 24548
rect 87820 24508 87860 24548
rect 87112 24172 87152 24212
rect 87194 24172 87234 24212
rect 87276 24172 87316 24212
rect 87358 24172 87398 24212
rect 87440 24172 87480 24212
rect 88204 25264 88244 25304
rect 88492 25264 88532 25304
rect 88876 25348 88916 25388
rect 88684 25264 88724 25304
rect 88108 24508 88148 24548
rect 88492 24508 88532 24548
rect 89644 25516 89684 25556
rect 89548 25348 89588 25388
rect 89740 25264 89780 25304
rect 89932 25516 89972 25556
rect 90028 25264 90068 25304
rect 90316 25264 90356 25304
rect 90604 25264 90644 25304
rect 90892 25264 90932 25304
rect 91276 25264 91316 25304
rect 89068 24508 89108 24548
rect 89260 24508 89300 24548
rect 89740 24508 89780 24548
rect 90124 24508 90164 24548
rect 90508 24508 90548 24548
rect 90988 24508 91028 24548
rect 91112 24172 91152 24212
rect 91194 24172 91234 24212
rect 91276 24172 91316 24212
rect 91358 24172 91398 24212
rect 91440 24172 91480 24212
rect 91948 25264 91988 25304
rect 92332 25348 92372 25388
rect 91660 24508 91700 24548
rect 92332 24508 92372 24548
rect 92524 25264 92564 25304
rect 92524 24508 92564 24548
rect 92908 25264 92948 25304
rect 93100 24508 93140 24548
rect 93484 24508 93524 24548
rect 93676 25264 93716 25304
rect 93964 25264 94004 25304
rect 94156 25264 94196 25304
rect 94924 25264 94964 25304
rect 93772 24508 93812 24548
rect 94156 24508 94196 24548
rect 94540 24508 94580 24548
rect 95404 24760 95444 24800
rect 96305 26524 96345 26564
rect 95692 25516 95732 25556
rect 95692 25348 95732 25388
rect 96076 25516 96116 25556
rect 96556 26524 96596 26564
rect 96460 25516 96500 25556
rect 95884 25096 95924 25136
rect 96172 25180 96212 25220
rect 96460 25180 96500 25220
rect 95980 24760 96020 24800
rect 96364 24760 96404 24800
rect 97420 25516 97460 25556
rect 96748 25264 96788 25304
rect 97036 25264 97076 25304
rect 96748 24760 96788 24800
rect 97132 24760 97172 24800
rect 97516 25264 97556 25304
rect 97516 24760 97556 24800
rect 97804 25264 97844 25304
rect 99148 32824 99188 32864
rect 98956 32152 98996 32192
rect 99244 32068 99284 32108
rect 98860 26104 98900 26144
rect 97996 25264 98036 25304
rect 97516 24508 97556 24548
rect 97900 24508 97940 24548
rect 98284 24508 98324 24548
rect 95112 24172 95152 24212
rect 95194 24172 95234 24212
rect 95276 24172 95316 24212
rect 95358 24172 95398 24212
rect 95440 24172 95480 24212
rect 99112 24172 99152 24212
rect 99194 24172 99234 24212
rect 99276 24172 99316 24212
rect 99358 24172 99398 24212
rect 99440 24172 99480 24212
rect 72352 23416 72392 23456
rect 72434 23416 72474 23456
rect 72516 23416 72556 23456
rect 72598 23416 72638 23456
rect 72680 23416 72720 23456
rect 76352 23416 76392 23456
rect 76434 23416 76474 23456
rect 76516 23416 76556 23456
rect 76598 23416 76638 23456
rect 76680 23416 76720 23456
rect 80352 23416 80392 23456
rect 80434 23416 80474 23456
rect 80516 23416 80556 23456
rect 80598 23416 80638 23456
rect 80680 23416 80720 23456
rect 84352 23416 84392 23456
rect 84434 23416 84474 23456
rect 84516 23416 84556 23456
rect 84598 23416 84638 23456
rect 84680 23416 84720 23456
rect 88352 23416 88392 23456
rect 88434 23416 88474 23456
rect 88516 23416 88556 23456
rect 88598 23416 88638 23456
rect 88680 23416 88720 23456
rect 92352 23416 92392 23456
rect 92434 23416 92474 23456
rect 92516 23416 92556 23456
rect 92598 23416 92638 23456
rect 92680 23416 92720 23456
rect 96352 23416 96392 23456
rect 96434 23416 96474 23456
rect 96516 23416 96556 23456
rect 96598 23416 96638 23456
rect 96680 23416 96720 23456
rect 71112 22660 71152 22700
rect 71194 22660 71234 22700
rect 71276 22660 71316 22700
rect 71358 22660 71398 22700
rect 71440 22660 71480 22700
rect 75112 22660 75152 22700
rect 75194 22660 75234 22700
rect 75276 22660 75316 22700
rect 75358 22660 75398 22700
rect 75440 22660 75480 22700
rect 79112 22660 79152 22700
rect 79194 22660 79234 22700
rect 79276 22660 79316 22700
rect 79358 22660 79398 22700
rect 79440 22660 79480 22700
rect 83112 22660 83152 22700
rect 83194 22660 83234 22700
rect 83276 22660 83316 22700
rect 83358 22660 83398 22700
rect 83440 22660 83480 22700
rect 87112 22660 87152 22700
rect 87194 22660 87234 22700
rect 87276 22660 87316 22700
rect 87358 22660 87398 22700
rect 87440 22660 87480 22700
rect 91112 22660 91152 22700
rect 91194 22660 91234 22700
rect 91276 22660 91316 22700
rect 91358 22660 91398 22700
rect 91440 22660 91480 22700
rect 95112 22660 95152 22700
rect 95194 22660 95234 22700
rect 95276 22660 95316 22700
rect 95358 22660 95398 22700
rect 95440 22660 95480 22700
rect 99112 22660 99152 22700
rect 99194 22660 99234 22700
rect 99276 22660 99316 22700
rect 99358 22660 99398 22700
rect 99440 22660 99480 22700
rect 72352 21904 72392 21944
rect 72434 21904 72474 21944
rect 72516 21904 72556 21944
rect 72598 21904 72638 21944
rect 72680 21904 72720 21944
rect 76352 21904 76392 21944
rect 76434 21904 76474 21944
rect 76516 21904 76556 21944
rect 76598 21904 76638 21944
rect 76680 21904 76720 21944
rect 80352 21904 80392 21944
rect 80434 21904 80474 21944
rect 80516 21904 80556 21944
rect 80598 21904 80638 21944
rect 80680 21904 80720 21944
rect 84352 21904 84392 21944
rect 84434 21904 84474 21944
rect 84516 21904 84556 21944
rect 84598 21904 84638 21944
rect 84680 21904 84720 21944
rect 88352 21904 88392 21944
rect 88434 21904 88474 21944
rect 88516 21904 88556 21944
rect 88598 21904 88638 21944
rect 88680 21904 88720 21944
rect 92352 21904 92392 21944
rect 92434 21904 92474 21944
rect 92516 21904 92556 21944
rect 92598 21904 92638 21944
rect 92680 21904 92720 21944
rect 96352 21904 96392 21944
rect 96434 21904 96474 21944
rect 96516 21904 96556 21944
rect 96598 21904 96638 21944
rect 96680 21904 96720 21944
rect 71112 21148 71152 21188
rect 71194 21148 71234 21188
rect 71276 21148 71316 21188
rect 71358 21148 71398 21188
rect 71440 21148 71480 21188
rect 75112 21148 75152 21188
rect 75194 21148 75234 21188
rect 75276 21148 75316 21188
rect 75358 21148 75398 21188
rect 75440 21148 75480 21188
rect 79112 21148 79152 21188
rect 79194 21148 79234 21188
rect 79276 21148 79316 21188
rect 79358 21148 79398 21188
rect 79440 21148 79480 21188
rect 83112 21148 83152 21188
rect 83194 21148 83234 21188
rect 83276 21148 83316 21188
rect 83358 21148 83398 21188
rect 83440 21148 83480 21188
rect 87112 21148 87152 21188
rect 87194 21148 87234 21188
rect 87276 21148 87316 21188
rect 87358 21148 87398 21188
rect 87440 21148 87480 21188
rect 91112 21148 91152 21188
rect 91194 21148 91234 21188
rect 91276 21148 91316 21188
rect 91358 21148 91398 21188
rect 91440 21148 91480 21188
rect 95112 21148 95152 21188
rect 95194 21148 95234 21188
rect 95276 21148 95316 21188
rect 95358 21148 95398 21188
rect 95440 21148 95480 21188
rect 99112 21148 99152 21188
rect 99194 21148 99234 21188
rect 99276 21148 99316 21188
rect 99358 21148 99398 21188
rect 99440 21148 99480 21188
rect 72352 20392 72392 20432
rect 72434 20392 72474 20432
rect 72516 20392 72556 20432
rect 72598 20392 72638 20432
rect 72680 20392 72720 20432
rect 76352 20392 76392 20432
rect 76434 20392 76474 20432
rect 76516 20392 76556 20432
rect 76598 20392 76638 20432
rect 76680 20392 76720 20432
rect 80352 20392 80392 20432
rect 80434 20392 80474 20432
rect 80516 20392 80556 20432
rect 80598 20392 80638 20432
rect 80680 20392 80720 20432
rect 84352 20392 84392 20432
rect 84434 20392 84474 20432
rect 84516 20392 84556 20432
rect 84598 20392 84638 20432
rect 84680 20392 84720 20432
rect 88352 20392 88392 20432
rect 88434 20392 88474 20432
rect 88516 20392 88556 20432
rect 88598 20392 88638 20432
rect 88680 20392 88720 20432
rect 92352 20392 92392 20432
rect 92434 20392 92474 20432
rect 92516 20392 92556 20432
rect 92598 20392 92638 20432
rect 92680 20392 92720 20432
rect 96352 20392 96392 20432
rect 96434 20392 96474 20432
rect 96516 20392 96556 20432
rect 96598 20392 96638 20432
rect 96680 20392 96720 20432
rect 71112 19636 71152 19676
rect 71194 19636 71234 19676
rect 71276 19636 71316 19676
rect 71358 19636 71398 19676
rect 71440 19636 71480 19676
rect 75112 19636 75152 19676
rect 75194 19636 75234 19676
rect 75276 19636 75316 19676
rect 75358 19636 75398 19676
rect 75440 19636 75480 19676
rect 79112 19636 79152 19676
rect 79194 19636 79234 19676
rect 79276 19636 79316 19676
rect 79358 19636 79398 19676
rect 79440 19636 79480 19676
rect 83112 19636 83152 19676
rect 83194 19636 83234 19676
rect 83276 19636 83316 19676
rect 83358 19636 83398 19676
rect 83440 19636 83480 19676
rect 87112 19636 87152 19676
rect 87194 19636 87234 19676
rect 87276 19636 87316 19676
rect 87358 19636 87398 19676
rect 87440 19636 87480 19676
rect 91112 19636 91152 19676
rect 91194 19636 91234 19676
rect 91276 19636 91316 19676
rect 91358 19636 91398 19676
rect 91440 19636 91480 19676
rect 95112 19636 95152 19676
rect 95194 19636 95234 19676
rect 95276 19636 95316 19676
rect 95358 19636 95398 19676
rect 95440 19636 95480 19676
rect 99112 19636 99152 19676
rect 99194 19636 99234 19676
rect 99276 19636 99316 19676
rect 99358 19636 99398 19676
rect 99440 19636 99480 19676
rect 72352 18880 72392 18920
rect 72434 18880 72474 18920
rect 72516 18880 72556 18920
rect 72598 18880 72638 18920
rect 72680 18880 72720 18920
rect 76352 18880 76392 18920
rect 76434 18880 76474 18920
rect 76516 18880 76556 18920
rect 76598 18880 76638 18920
rect 76680 18880 76720 18920
rect 80352 18880 80392 18920
rect 80434 18880 80474 18920
rect 80516 18880 80556 18920
rect 80598 18880 80638 18920
rect 80680 18880 80720 18920
rect 84352 18880 84392 18920
rect 84434 18880 84474 18920
rect 84516 18880 84556 18920
rect 84598 18880 84638 18920
rect 84680 18880 84720 18920
rect 88352 18880 88392 18920
rect 88434 18880 88474 18920
rect 88516 18880 88556 18920
rect 88598 18880 88638 18920
rect 88680 18880 88720 18920
rect 92352 18880 92392 18920
rect 92434 18880 92474 18920
rect 92516 18880 92556 18920
rect 92598 18880 92638 18920
rect 92680 18880 92720 18920
rect 96352 18880 96392 18920
rect 96434 18880 96474 18920
rect 96516 18880 96556 18920
rect 96598 18880 96638 18920
rect 96680 18880 96720 18920
rect 71112 18124 71152 18164
rect 71194 18124 71234 18164
rect 71276 18124 71316 18164
rect 71358 18124 71398 18164
rect 71440 18124 71480 18164
rect 75112 18124 75152 18164
rect 75194 18124 75234 18164
rect 75276 18124 75316 18164
rect 75358 18124 75398 18164
rect 75440 18124 75480 18164
rect 79112 18124 79152 18164
rect 79194 18124 79234 18164
rect 79276 18124 79316 18164
rect 79358 18124 79398 18164
rect 79440 18124 79480 18164
rect 83112 18124 83152 18164
rect 83194 18124 83234 18164
rect 83276 18124 83316 18164
rect 83358 18124 83398 18164
rect 83440 18124 83480 18164
rect 87112 18124 87152 18164
rect 87194 18124 87234 18164
rect 87276 18124 87316 18164
rect 87358 18124 87398 18164
rect 87440 18124 87480 18164
rect 91112 18124 91152 18164
rect 91194 18124 91234 18164
rect 91276 18124 91316 18164
rect 91358 18124 91398 18164
rect 91440 18124 91480 18164
rect 95112 18124 95152 18164
rect 95194 18124 95234 18164
rect 95276 18124 95316 18164
rect 95358 18124 95398 18164
rect 95440 18124 95480 18164
rect 99112 18124 99152 18164
rect 99194 18124 99234 18164
rect 99276 18124 99316 18164
rect 99358 18124 99398 18164
rect 99440 18124 99480 18164
rect 72352 17368 72392 17408
rect 72434 17368 72474 17408
rect 72516 17368 72556 17408
rect 72598 17368 72638 17408
rect 72680 17368 72720 17408
rect 76352 17368 76392 17408
rect 76434 17368 76474 17408
rect 76516 17368 76556 17408
rect 76598 17368 76638 17408
rect 76680 17368 76720 17408
rect 80352 17368 80392 17408
rect 80434 17368 80474 17408
rect 80516 17368 80556 17408
rect 80598 17368 80638 17408
rect 80680 17368 80720 17408
rect 84352 17368 84392 17408
rect 84434 17368 84474 17408
rect 84516 17368 84556 17408
rect 84598 17368 84638 17408
rect 84680 17368 84720 17408
rect 88352 17368 88392 17408
rect 88434 17368 88474 17408
rect 88516 17368 88556 17408
rect 88598 17368 88638 17408
rect 88680 17368 88720 17408
rect 92352 17368 92392 17408
rect 92434 17368 92474 17408
rect 92516 17368 92556 17408
rect 92598 17368 92638 17408
rect 92680 17368 92720 17408
rect 96352 17368 96392 17408
rect 96434 17368 96474 17408
rect 96516 17368 96556 17408
rect 96598 17368 96638 17408
rect 96680 17368 96720 17408
rect 71112 16612 71152 16652
rect 71194 16612 71234 16652
rect 71276 16612 71316 16652
rect 71358 16612 71398 16652
rect 71440 16612 71480 16652
rect 75112 16612 75152 16652
rect 75194 16612 75234 16652
rect 75276 16612 75316 16652
rect 75358 16612 75398 16652
rect 75440 16612 75480 16652
rect 79112 16612 79152 16652
rect 79194 16612 79234 16652
rect 79276 16612 79316 16652
rect 79358 16612 79398 16652
rect 79440 16612 79480 16652
rect 71788 16360 71828 16400
rect 70636 14764 70676 14804
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 8352 14344 8392 14384
rect 8434 14344 8474 14384
rect 8516 14344 8556 14384
rect 8598 14344 8638 14384
rect 8680 14344 8720 14384
rect 12352 14344 12392 14384
rect 12434 14344 12474 14384
rect 12516 14344 12556 14384
rect 12598 14344 12638 14384
rect 12680 14344 12720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 20352 14344 20392 14384
rect 20434 14344 20474 14384
rect 20516 14344 20556 14384
rect 20598 14344 20638 14384
rect 20680 14344 20720 14384
rect 24352 14344 24392 14384
rect 24434 14344 24474 14384
rect 24516 14344 24556 14384
rect 24598 14344 24638 14384
rect 24680 14344 24720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 32352 14344 32392 14384
rect 32434 14344 32474 14384
rect 32516 14344 32556 14384
rect 32598 14344 32638 14384
rect 32680 14344 32720 14384
rect 36352 14344 36392 14384
rect 36434 14344 36474 14384
rect 36516 14344 36556 14384
rect 36598 14344 36638 14384
rect 36680 14344 36720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 44352 14344 44392 14384
rect 44434 14344 44474 14384
rect 44516 14344 44556 14384
rect 44598 14344 44638 14384
rect 44680 14344 44720 14384
rect 48352 14344 48392 14384
rect 48434 14344 48474 14384
rect 48516 14344 48556 14384
rect 48598 14344 48638 14384
rect 48680 14344 48720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 56352 14344 56392 14384
rect 56434 14344 56474 14384
rect 56516 14344 56556 14384
rect 56598 14344 56638 14384
rect 56680 14344 56720 14384
rect 60352 14344 60392 14384
rect 60434 14344 60474 14384
rect 60516 14344 60556 14384
rect 60598 14344 60638 14384
rect 60680 14344 60720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 68352 14344 68392 14384
rect 68434 14344 68474 14384
rect 68516 14344 68556 14384
rect 68598 14344 68638 14384
rect 68680 14344 68720 14384
rect 70540 14008 70580 14048
rect 70828 14008 70868 14048
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 7112 13588 7152 13628
rect 7194 13588 7234 13628
rect 7276 13588 7316 13628
rect 7358 13588 7398 13628
rect 7440 13588 7480 13628
rect 11112 13588 11152 13628
rect 11194 13588 11234 13628
rect 11276 13588 11316 13628
rect 11358 13588 11398 13628
rect 11440 13588 11480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 19112 13588 19152 13628
rect 19194 13588 19234 13628
rect 19276 13588 19316 13628
rect 19358 13588 19398 13628
rect 19440 13588 19480 13628
rect 23112 13588 23152 13628
rect 23194 13588 23234 13628
rect 23276 13588 23316 13628
rect 23358 13588 23398 13628
rect 23440 13588 23480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 31112 13588 31152 13628
rect 31194 13588 31234 13628
rect 31276 13588 31316 13628
rect 31358 13588 31398 13628
rect 31440 13588 31480 13628
rect 35112 13588 35152 13628
rect 35194 13588 35234 13628
rect 35276 13588 35316 13628
rect 35358 13588 35398 13628
rect 35440 13588 35480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 43112 13588 43152 13628
rect 43194 13588 43234 13628
rect 43276 13588 43316 13628
rect 43358 13588 43398 13628
rect 43440 13588 43480 13628
rect 47112 13588 47152 13628
rect 47194 13588 47234 13628
rect 47276 13588 47316 13628
rect 47358 13588 47398 13628
rect 47440 13588 47480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 55112 13588 55152 13628
rect 55194 13588 55234 13628
rect 55276 13588 55316 13628
rect 55358 13588 55398 13628
rect 55440 13588 55480 13628
rect 59112 13588 59152 13628
rect 59194 13588 59234 13628
rect 59276 13588 59316 13628
rect 59358 13588 59398 13628
rect 59440 13588 59480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 67112 13588 67152 13628
rect 67194 13588 67234 13628
rect 67276 13588 67316 13628
rect 67358 13588 67398 13628
rect 67440 13588 67480 13628
rect 70060 13588 70100 13628
rect 69868 13168 69908 13208
rect 70732 13924 70772 13964
rect 70636 13756 70676 13796
rect 70348 13168 70388 13208
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 8352 12832 8392 12872
rect 8434 12832 8474 12872
rect 8516 12832 8556 12872
rect 8598 12832 8638 12872
rect 8680 12832 8720 12872
rect 12352 12832 12392 12872
rect 12434 12832 12474 12872
rect 12516 12832 12556 12872
rect 12598 12832 12638 12872
rect 12680 12832 12720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 20352 12832 20392 12872
rect 20434 12832 20474 12872
rect 20516 12832 20556 12872
rect 20598 12832 20638 12872
rect 20680 12832 20720 12872
rect 24352 12832 24392 12872
rect 24434 12832 24474 12872
rect 24516 12832 24556 12872
rect 24598 12832 24638 12872
rect 24680 12832 24720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 32352 12832 32392 12872
rect 32434 12832 32474 12872
rect 32516 12832 32556 12872
rect 32598 12832 32638 12872
rect 32680 12832 32720 12872
rect 36352 12832 36392 12872
rect 36434 12832 36474 12872
rect 36516 12832 36556 12872
rect 36598 12832 36638 12872
rect 36680 12832 36720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 44352 12832 44392 12872
rect 44434 12832 44474 12872
rect 44516 12832 44556 12872
rect 44598 12832 44638 12872
rect 44680 12832 44720 12872
rect 48352 12832 48392 12872
rect 48434 12832 48474 12872
rect 48516 12832 48556 12872
rect 48598 12832 48638 12872
rect 48680 12832 48720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 56352 12832 56392 12872
rect 56434 12832 56474 12872
rect 56516 12832 56556 12872
rect 56598 12832 56638 12872
rect 56680 12832 56720 12872
rect 60352 12832 60392 12872
rect 60434 12832 60474 12872
rect 60516 12832 60556 12872
rect 60598 12832 60638 12872
rect 60680 12832 60720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 68352 12832 68392 12872
rect 68434 12832 68474 12872
rect 68516 12832 68556 12872
rect 68598 12832 68638 12872
rect 68680 12832 68720 12872
rect 70732 13168 70772 13208
rect 71020 13672 71060 13712
rect 70924 13420 70964 13460
rect 71308 14680 71348 14720
rect 71308 13924 71348 13964
rect 71404 13840 71444 13880
rect 71308 13420 71348 13460
rect 71212 13336 71252 13376
rect 71116 13252 71156 13292
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 7112 12076 7152 12116
rect 7194 12076 7234 12116
rect 7276 12076 7316 12116
rect 7358 12076 7398 12116
rect 7440 12076 7480 12116
rect 11112 12076 11152 12116
rect 11194 12076 11234 12116
rect 11276 12076 11316 12116
rect 11358 12076 11398 12116
rect 11440 12076 11480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 19112 12076 19152 12116
rect 19194 12076 19234 12116
rect 19276 12076 19316 12116
rect 19358 12076 19398 12116
rect 19440 12076 19480 12116
rect 23112 12076 23152 12116
rect 23194 12076 23234 12116
rect 23276 12076 23316 12116
rect 23358 12076 23398 12116
rect 23440 12076 23480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 31112 12076 31152 12116
rect 31194 12076 31234 12116
rect 31276 12076 31316 12116
rect 31358 12076 31398 12116
rect 31440 12076 31480 12116
rect 35112 12076 35152 12116
rect 35194 12076 35234 12116
rect 35276 12076 35316 12116
rect 35358 12076 35398 12116
rect 35440 12076 35480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 43112 12076 43152 12116
rect 43194 12076 43234 12116
rect 43276 12076 43316 12116
rect 43358 12076 43398 12116
rect 43440 12076 43480 12116
rect 47112 12076 47152 12116
rect 47194 12076 47234 12116
rect 47276 12076 47316 12116
rect 47358 12076 47398 12116
rect 47440 12076 47480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 55112 12076 55152 12116
rect 55194 12076 55234 12116
rect 55276 12076 55316 12116
rect 55358 12076 55398 12116
rect 55440 12076 55480 12116
rect 59112 12076 59152 12116
rect 59194 12076 59234 12116
rect 59276 12076 59316 12116
rect 59358 12076 59398 12116
rect 59440 12076 59480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 67112 12076 67152 12116
rect 67194 12076 67234 12116
rect 67276 12076 67316 12116
rect 67358 12076 67398 12116
rect 67440 12076 67480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 8352 11320 8392 11360
rect 8434 11320 8474 11360
rect 8516 11320 8556 11360
rect 8598 11320 8638 11360
rect 8680 11320 8720 11360
rect 12352 11320 12392 11360
rect 12434 11320 12474 11360
rect 12516 11320 12556 11360
rect 12598 11320 12638 11360
rect 12680 11320 12720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 20352 11320 20392 11360
rect 20434 11320 20474 11360
rect 20516 11320 20556 11360
rect 20598 11320 20638 11360
rect 20680 11320 20720 11360
rect 24352 11320 24392 11360
rect 24434 11320 24474 11360
rect 24516 11320 24556 11360
rect 24598 11320 24638 11360
rect 24680 11320 24720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 32352 11320 32392 11360
rect 32434 11320 32474 11360
rect 32516 11320 32556 11360
rect 32598 11320 32638 11360
rect 32680 11320 32720 11360
rect 36352 11320 36392 11360
rect 36434 11320 36474 11360
rect 36516 11320 36556 11360
rect 36598 11320 36638 11360
rect 36680 11320 36720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 44352 11320 44392 11360
rect 44434 11320 44474 11360
rect 44516 11320 44556 11360
rect 44598 11320 44638 11360
rect 44680 11320 44720 11360
rect 48352 11320 48392 11360
rect 48434 11320 48474 11360
rect 48516 11320 48556 11360
rect 48598 11320 48638 11360
rect 48680 11320 48720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 56352 11320 56392 11360
rect 56434 11320 56474 11360
rect 56516 11320 56556 11360
rect 56598 11320 56638 11360
rect 56680 11320 56720 11360
rect 60352 11320 60392 11360
rect 60434 11320 60474 11360
rect 60516 11320 60556 11360
rect 60598 11320 60638 11360
rect 60680 11320 60720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 68352 11320 68392 11360
rect 68434 11320 68474 11360
rect 68516 11320 68556 11360
rect 68598 11320 68638 11360
rect 68680 11320 68720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 7112 10564 7152 10604
rect 7194 10564 7234 10604
rect 7276 10564 7316 10604
rect 7358 10564 7398 10604
rect 7440 10564 7480 10604
rect 11112 10564 11152 10604
rect 11194 10564 11234 10604
rect 11276 10564 11316 10604
rect 11358 10564 11398 10604
rect 11440 10564 11480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 19112 10564 19152 10604
rect 19194 10564 19234 10604
rect 19276 10564 19316 10604
rect 19358 10564 19398 10604
rect 19440 10564 19480 10604
rect 23112 10564 23152 10604
rect 23194 10564 23234 10604
rect 23276 10564 23316 10604
rect 23358 10564 23398 10604
rect 23440 10564 23480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 31112 10564 31152 10604
rect 31194 10564 31234 10604
rect 31276 10564 31316 10604
rect 31358 10564 31398 10604
rect 31440 10564 31480 10604
rect 35112 10564 35152 10604
rect 35194 10564 35234 10604
rect 35276 10564 35316 10604
rect 35358 10564 35398 10604
rect 35440 10564 35480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 43112 10564 43152 10604
rect 43194 10564 43234 10604
rect 43276 10564 43316 10604
rect 43358 10564 43398 10604
rect 43440 10564 43480 10604
rect 47112 10564 47152 10604
rect 47194 10564 47234 10604
rect 47276 10564 47316 10604
rect 47358 10564 47398 10604
rect 47440 10564 47480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 55112 10564 55152 10604
rect 55194 10564 55234 10604
rect 55276 10564 55316 10604
rect 55358 10564 55398 10604
rect 55440 10564 55480 10604
rect 59112 10564 59152 10604
rect 59194 10564 59234 10604
rect 59276 10564 59316 10604
rect 59358 10564 59398 10604
rect 59440 10564 59480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 67112 10564 67152 10604
rect 67194 10564 67234 10604
rect 67276 10564 67316 10604
rect 67358 10564 67398 10604
rect 67440 10564 67480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 8352 9808 8392 9848
rect 8434 9808 8474 9848
rect 8516 9808 8556 9848
rect 8598 9808 8638 9848
rect 8680 9808 8720 9848
rect 12352 9808 12392 9848
rect 12434 9808 12474 9848
rect 12516 9808 12556 9848
rect 12598 9808 12638 9848
rect 12680 9808 12720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 20352 9808 20392 9848
rect 20434 9808 20474 9848
rect 20516 9808 20556 9848
rect 20598 9808 20638 9848
rect 20680 9808 20720 9848
rect 24352 9808 24392 9848
rect 24434 9808 24474 9848
rect 24516 9808 24556 9848
rect 24598 9808 24638 9848
rect 24680 9808 24720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 32352 9808 32392 9848
rect 32434 9808 32474 9848
rect 32516 9808 32556 9848
rect 32598 9808 32638 9848
rect 32680 9808 32720 9848
rect 36352 9808 36392 9848
rect 36434 9808 36474 9848
rect 36516 9808 36556 9848
rect 36598 9808 36638 9848
rect 36680 9808 36720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 44352 9808 44392 9848
rect 44434 9808 44474 9848
rect 44516 9808 44556 9848
rect 44598 9808 44638 9848
rect 44680 9808 44720 9848
rect 48352 9808 48392 9848
rect 48434 9808 48474 9848
rect 48516 9808 48556 9848
rect 48598 9808 48638 9848
rect 48680 9808 48720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 56352 9808 56392 9848
rect 56434 9808 56474 9848
rect 56516 9808 56556 9848
rect 56598 9808 56638 9848
rect 56680 9808 56720 9848
rect 60352 9808 60392 9848
rect 60434 9808 60474 9848
rect 60516 9808 60556 9848
rect 60598 9808 60638 9848
rect 60680 9808 60720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 68352 9808 68392 9848
rect 68434 9808 68474 9848
rect 68516 9808 68556 9848
rect 68598 9808 68638 9848
rect 68680 9808 68720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 7112 9052 7152 9092
rect 7194 9052 7234 9092
rect 7276 9052 7316 9092
rect 7358 9052 7398 9092
rect 7440 9052 7480 9092
rect 11112 9052 11152 9092
rect 11194 9052 11234 9092
rect 11276 9052 11316 9092
rect 11358 9052 11398 9092
rect 11440 9052 11480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 19112 9052 19152 9092
rect 19194 9052 19234 9092
rect 19276 9052 19316 9092
rect 19358 9052 19398 9092
rect 19440 9052 19480 9092
rect 23112 9052 23152 9092
rect 23194 9052 23234 9092
rect 23276 9052 23316 9092
rect 23358 9052 23398 9092
rect 23440 9052 23480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 31112 9052 31152 9092
rect 31194 9052 31234 9092
rect 31276 9052 31316 9092
rect 31358 9052 31398 9092
rect 31440 9052 31480 9092
rect 35112 9052 35152 9092
rect 35194 9052 35234 9092
rect 35276 9052 35316 9092
rect 35358 9052 35398 9092
rect 35440 9052 35480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 43112 9052 43152 9092
rect 43194 9052 43234 9092
rect 43276 9052 43316 9092
rect 43358 9052 43398 9092
rect 43440 9052 43480 9092
rect 47112 9052 47152 9092
rect 47194 9052 47234 9092
rect 47276 9052 47316 9092
rect 47358 9052 47398 9092
rect 47440 9052 47480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 55112 9052 55152 9092
rect 55194 9052 55234 9092
rect 55276 9052 55316 9092
rect 55358 9052 55398 9092
rect 55440 9052 55480 9092
rect 59112 9052 59152 9092
rect 59194 9052 59234 9092
rect 59276 9052 59316 9092
rect 59358 9052 59398 9092
rect 59440 9052 59480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 67112 9052 67152 9092
rect 67194 9052 67234 9092
rect 67276 9052 67316 9092
rect 67358 9052 67398 9092
rect 67440 9052 67480 9092
rect 652 8128 692 8168
rect 844 7372 884 7412
rect 1516 7372 1556 7412
rect 652 7288 692 7328
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 8352 8296 8392 8336
rect 8434 8296 8474 8336
rect 8516 8296 8556 8336
rect 8598 8296 8638 8336
rect 8680 8296 8720 8336
rect 12352 8296 12392 8336
rect 12434 8296 12474 8336
rect 12516 8296 12556 8336
rect 12598 8296 12638 8336
rect 12680 8296 12720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 20352 8296 20392 8336
rect 20434 8296 20474 8336
rect 20516 8296 20556 8336
rect 20598 8296 20638 8336
rect 20680 8296 20720 8336
rect 24352 8296 24392 8336
rect 24434 8296 24474 8336
rect 24516 8296 24556 8336
rect 24598 8296 24638 8336
rect 24680 8296 24720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 32352 8296 32392 8336
rect 32434 8296 32474 8336
rect 32516 8296 32556 8336
rect 32598 8296 32638 8336
rect 32680 8296 32720 8336
rect 36352 8296 36392 8336
rect 36434 8296 36474 8336
rect 36516 8296 36556 8336
rect 36598 8296 36638 8336
rect 36680 8296 36720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 44352 8296 44392 8336
rect 44434 8296 44474 8336
rect 44516 8296 44556 8336
rect 44598 8296 44638 8336
rect 44680 8296 44720 8336
rect 48352 8296 48392 8336
rect 48434 8296 48474 8336
rect 48516 8296 48556 8336
rect 48598 8296 48638 8336
rect 48680 8296 48720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 56352 8296 56392 8336
rect 56434 8296 56474 8336
rect 56516 8296 56556 8336
rect 56598 8296 56638 8336
rect 56680 8296 56720 8336
rect 60352 8296 60392 8336
rect 60434 8296 60474 8336
rect 60516 8296 60556 8336
rect 60598 8296 60638 8336
rect 60680 8296 60720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 68352 8296 68392 8336
rect 68434 8296 68474 8336
rect 68516 8296 68556 8336
rect 68598 8296 68638 8336
rect 68680 8296 68720 8336
rect 71020 7876 71060 7916
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 7112 7540 7152 7580
rect 7194 7540 7234 7580
rect 7276 7540 7316 7580
rect 7358 7540 7398 7580
rect 7440 7540 7480 7580
rect 11112 7540 11152 7580
rect 11194 7540 11234 7580
rect 11276 7540 11316 7580
rect 11358 7540 11398 7580
rect 11440 7540 11480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 19112 7540 19152 7580
rect 19194 7540 19234 7580
rect 19276 7540 19316 7580
rect 19358 7540 19398 7580
rect 19440 7540 19480 7580
rect 23112 7540 23152 7580
rect 23194 7540 23234 7580
rect 23276 7540 23316 7580
rect 23358 7540 23398 7580
rect 23440 7540 23480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 31112 7540 31152 7580
rect 31194 7540 31234 7580
rect 31276 7540 31316 7580
rect 31358 7540 31398 7580
rect 31440 7540 31480 7580
rect 35112 7540 35152 7580
rect 35194 7540 35234 7580
rect 35276 7540 35316 7580
rect 35358 7540 35398 7580
rect 35440 7540 35480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 43112 7540 43152 7580
rect 43194 7540 43234 7580
rect 43276 7540 43316 7580
rect 43358 7540 43398 7580
rect 43440 7540 43480 7580
rect 47112 7540 47152 7580
rect 47194 7540 47234 7580
rect 47276 7540 47316 7580
rect 47358 7540 47398 7580
rect 47440 7540 47480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 55112 7540 55152 7580
rect 55194 7540 55234 7580
rect 55276 7540 55316 7580
rect 55358 7540 55398 7580
rect 55440 7540 55480 7580
rect 59112 7540 59152 7580
rect 59194 7540 59234 7580
rect 59276 7540 59316 7580
rect 59358 7540 59398 7580
rect 59440 7540 59480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 67112 7540 67152 7580
rect 67194 7540 67234 7580
rect 67276 7540 67316 7580
rect 67358 7540 67398 7580
rect 67440 7540 67480 7580
rect 844 6616 884 6656
rect 652 6448 692 6488
rect 71116 7120 71156 7160
rect 71404 7792 71444 7832
rect 71500 7708 71540 7748
rect 73900 16276 73940 16316
rect 83112 16612 83152 16652
rect 83194 16612 83234 16652
rect 83276 16612 83316 16652
rect 83358 16612 83398 16652
rect 83440 16612 83480 16652
rect 73132 16192 73172 16232
rect 72352 15856 72392 15896
rect 72434 15856 72474 15896
rect 72516 15856 72556 15896
rect 72598 15856 72638 15896
rect 72680 15856 72720 15896
rect 72748 14680 72788 14720
rect 73036 14680 73076 14720
rect 72844 14512 72884 14552
rect 74476 16276 74516 16316
rect 74284 16192 74324 16232
rect 77164 16276 77204 16316
rect 80428 16276 80468 16316
rect 80620 16276 80660 16316
rect 83116 16360 83156 16400
rect 83404 16360 83444 16400
rect 83788 16360 83828 16400
rect 86188 16360 86228 16400
rect 81772 16276 81812 16316
rect 73708 15436 73748 15476
rect 76780 16024 76820 16064
rect 76352 15856 76392 15896
rect 76434 15856 76474 15896
rect 76516 15856 76556 15896
rect 76598 15856 76638 15896
rect 76680 15856 76720 15896
rect 74092 15436 74132 15476
rect 73900 15268 73940 15308
rect 73516 14680 73556 14720
rect 73900 14680 73940 14720
rect 73132 14008 73172 14048
rect 73516 13840 73556 13880
rect 73132 13756 73172 13796
rect 72652 13672 72692 13712
rect 72415 13420 72455 13460
rect 72305 13336 72345 13376
rect 72844 13504 72884 13544
rect 73228 13504 73268 13544
rect 74476 15436 74516 15476
rect 74860 15436 74900 15476
rect 74380 15268 74420 15308
rect 74188 14680 74228 14720
rect 74188 14428 74228 14468
rect 74284 13588 74324 13628
rect 74860 14680 74900 14720
rect 74668 13588 74708 13628
rect 75340 15268 75380 15308
rect 75244 14680 75284 14720
rect 75820 15268 75860 15308
rect 75820 14680 75860 14720
rect 76204 15268 76244 15308
rect 76108 14680 76148 14720
rect 76588 15268 76628 15308
rect 77356 16024 77396 16064
rect 76972 15184 77012 15224
rect 76876 15100 76916 15140
rect 77356 15184 77396 15224
rect 77740 15184 77780 15224
rect 77836 15100 77876 15140
rect 78124 15184 78164 15224
rect 80352 15856 80392 15896
rect 80434 15856 80474 15896
rect 80516 15856 80556 15896
rect 80598 15856 80638 15896
rect 80680 15856 80720 15896
rect 78796 15352 78836 15392
rect 78604 15100 78644 15140
rect 79180 15352 79220 15392
rect 79372 15352 79412 15392
rect 79660 15352 79700 15392
rect 79084 13840 79124 13880
rect 80236 15436 80276 15476
rect 79756 15184 79796 15224
rect 79756 13840 79796 13880
rect 80716 15436 80756 15476
rect 79905 13420 79945 13460
rect 80428 15100 80468 15140
rect 81100 15436 81140 15476
rect 80524 13672 80564 13712
rect 81388 15436 81428 15476
rect 81580 16024 81620 16064
rect 81772 16024 81812 16064
rect 82060 13588 82100 13628
rect 82252 16024 82292 16064
rect 83308 16276 83348 16316
rect 82540 15436 82580 15476
rect 82305 13420 82345 13460
rect 84652 16276 84692 16316
rect 86380 16276 86420 16316
rect 87112 16612 87152 16652
rect 87194 16612 87234 16652
rect 87276 16612 87316 16652
rect 87358 16612 87398 16652
rect 87440 16612 87480 16652
rect 91112 16612 91152 16652
rect 91194 16612 91234 16652
rect 91276 16612 91316 16652
rect 91358 16612 91398 16652
rect 91440 16612 91480 16652
rect 95112 16612 95152 16652
rect 95194 16612 95234 16652
rect 95276 16612 95316 16652
rect 95358 16612 95398 16652
rect 95440 16612 95480 16652
rect 99112 16612 99152 16652
rect 99194 16612 99234 16652
rect 99276 16612 99316 16652
rect 99358 16612 99398 16652
rect 99440 16612 99480 16652
rect 86764 16360 86804 16400
rect 86572 16276 86612 16316
rect 86476 16192 86516 16232
rect 83020 15436 83060 15476
rect 83404 15436 83444 15476
rect 83884 15436 83924 15476
rect 83980 15268 84020 15308
rect 84352 15856 84392 15896
rect 84434 15856 84474 15896
rect 84516 15856 84556 15896
rect 84598 15856 84638 15896
rect 84680 15856 84720 15896
rect 88204 16276 88244 16316
rect 89356 16276 89396 16316
rect 90220 16276 90260 16316
rect 90604 16276 90644 16316
rect 84172 15436 84212 15476
rect 84556 15436 84596 15476
rect 85036 15436 85076 15476
rect 85420 15436 85460 15476
rect 85804 15436 85844 15476
rect 86188 15436 86228 15476
rect 84268 15268 84308 15308
rect 86380 15436 86420 15476
rect 86572 15436 86612 15476
rect 87052 15436 87092 15476
rect 87436 15436 87476 15476
rect 88352 15856 88392 15896
rect 88434 15856 88474 15896
rect 88516 15856 88556 15896
rect 88598 15856 88638 15896
rect 88680 15856 88720 15896
rect 88300 15436 88340 15476
rect 88684 15436 88724 15476
rect 89068 15436 89108 15476
rect 89452 15436 89492 15476
rect 89836 15436 89876 15476
rect 91084 15436 91124 15476
rect 90508 15184 90548 15224
rect 90892 15268 90932 15308
rect 91084 15184 91124 15224
rect 90415 13420 90455 13460
rect 92428 16276 92468 16316
rect 91948 15436 91988 15476
rect 92352 15856 92392 15896
rect 92434 15856 92474 15896
rect 92516 15856 92556 15896
rect 92598 15856 92638 15896
rect 92680 15856 92720 15896
rect 91564 15184 91604 15224
rect 91756 15184 91796 15224
rect 92236 15268 92276 15308
rect 92716 15268 92756 15308
rect 92428 15100 92468 15140
rect 93868 15436 93908 15476
rect 92812 15100 92852 15140
rect 92812 14512 92852 14552
rect 93388 15268 93428 15308
rect 93100 14512 93140 14552
rect 95596 16276 95636 16316
rect 95500 15520 95540 15560
rect 94252 15436 94292 15476
rect 94636 15436 94676 15476
rect 94924 15436 94964 15476
rect 94156 15100 94196 15140
rect 94156 14680 94196 14720
rect 94636 14680 94676 14720
rect 96352 15856 96392 15896
rect 96434 15856 96474 15896
rect 96516 15856 96556 15896
rect 96598 15856 96638 15896
rect 96680 15856 96720 15896
rect 96076 15520 96116 15560
rect 96556 15520 96596 15560
rect 95980 15436 96020 15476
rect 96844 15520 96884 15560
rect 95020 15268 95060 15308
rect 97228 15436 97268 15476
rect 97708 15436 97748 15476
rect 97996 15436 98036 15476
rect 98380 15436 98420 15476
rect 97036 15100 97076 15140
rect 97132 14512 97172 14552
rect 96705 13336 96745 13376
rect 97516 15100 97556 15140
rect 96940 13336 96980 13376
rect 97804 14512 97844 14552
rect 97905 13420 97945 13460
rect 98380 13672 98420 13712
rect 98764 13672 98804 13712
rect 98668 13420 98708 13460
rect 72705 7876 72745 7916
rect 72305 7792 72345 7832
rect 72415 7792 72455 7832
rect 71788 7372 71828 7412
rect 72556 7456 72596 7496
rect 73132 7456 73172 7496
rect 72076 7120 72116 7160
rect 72364 7120 72404 7160
rect 72940 7120 72980 7160
rect 73612 7120 73652 7160
rect 73228 7036 73268 7076
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 8352 6784 8392 6824
rect 8434 6784 8474 6824
rect 8516 6784 8556 6824
rect 8598 6784 8638 6824
rect 8680 6784 8720 6824
rect 12352 6784 12392 6824
rect 12434 6784 12474 6824
rect 12516 6784 12556 6824
rect 12598 6784 12638 6824
rect 12680 6784 12720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 20352 6784 20392 6824
rect 20434 6784 20474 6824
rect 20516 6784 20556 6824
rect 20598 6784 20638 6824
rect 20680 6784 20720 6824
rect 24352 6784 24392 6824
rect 24434 6784 24474 6824
rect 24516 6784 24556 6824
rect 24598 6784 24638 6824
rect 24680 6784 24720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 32352 6784 32392 6824
rect 32434 6784 32474 6824
rect 32516 6784 32556 6824
rect 32598 6784 32638 6824
rect 32680 6784 32720 6824
rect 36352 6784 36392 6824
rect 36434 6784 36474 6824
rect 36516 6784 36556 6824
rect 36598 6784 36638 6824
rect 36680 6784 36720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 44352 6784 44392 6824
rect 44434 6784 44474 6824
rect 44516 6784 44556 6824
rect 44598 6784 44638 6824
rect 44680 6784 44720 6824
rect 48352 6784 48392 6824
rect 48434 6784 48474 6824
rect 48516 6784 48556 6824
rect 48598 6784 48638 6824
rect 48680 6784 48720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 56352 6784 56392 6824
rect 56434 6784 56474 6824
rect 56516 6784 56556 6824
rect 56598 6784 56638 6824
rect 56680 6784 56720 6824
rect 60352 6784 60392 6824
rect 60434 6784 60474 6824
rect 60516 6784 60556 6824
rect 60598 6784 60638 6824
rect 60680 6784 60720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 68352 6784 68392 6824
rect 68434 6784 68474 6824
rect 68516 6784 68556 6824
rect 68598 6784 68638 6824
rect 68680 6784 68720 6824
rect 1708 6616 1748 6656
rect 74092 6952 74132 6992
rect 74284 7288 74324 7328
rect 74476 7204 74516 7244
rect 74668 7372 74708 7412
rect 74860 7372 74900 7412
rect 74860 7204 74900 7244
rect 74956 6952 74996 6992
rect 75615 7624 75655 7664
rect 75244 7456 75284 7496
rect 75148 7372 75188 7412
rect 75244 6952 75284 6992
rect 73996 6364 74036 6404
rect 74380 6364 74420 6404
rect 74860 6364 74900 6404
rect 75532 7288 75572 7328
rect 75724 7120 75764 7160
rect 75916 7456 75956 7496
rect 76204 7624 76244 7664
rect 76108 7204 76148 7244
rect 76300 7120 76340 7160
rect 76012 6952 76052 6992
rect 76492 7372 76532 7412
rect 76492 7204 76532 7244
rect 76588 7120 76628 7160
rect 76492 6952 76532 6992
rect 76780 7372 76820 7412
rect 76876 7288 76916 7328
rect 76876 7120 76916 7160
rect 77260 7372 77300 7412
rect 77356 7204 77396 7244
rect 77644 7456 77684 7496
rect 77644 7288 77684 7328
rect 77548 7120 77588 7160
rect 78124 7456 78164 7496
rect 77836 7372 77876 7412
rect 78028 7372 78068 7412
rect 77932 7120 77972 7160
rect 78220 7120 78260 7160
rect 76876 6364 76916 6404
rect 77260 6364 77300 6404
rect 77644 6364 77684 6404
rect 78415 7624 78455 7664
rect 78412 7372 78452 7412
rect 78508 7120 78548 7160
rect 78796 7372 78836 7412
rect 78796 7204 78836 7244
rect 78988 6952 79028 6992
rect 79276 7624 79316 7664
rect 79180 7288 79220 7328
rect 79180 7120 79220 7160
rect 79468 7372 79508 7412
rect 79564 6952 79604 6992
rect 79756 7204 79796 7244
rect 79756 6952 79796 6992
rect 79660 6868 79700 6908
rect 80044 7372 80084 7412
rect 80140 7204 80180 7244
rect 78124 6364 78164 6404
rect 78508 6364 78548 6404
rect 78892 6364 78932 6404
rect 79276 6364 79316 6404
rect 79756 6364 79796 6404
rect 80332 7456 80372 7496
rect 80524 7288 80564 7328
rect 80620 6952 80660 6992
rect 80428 6616 80468 6656
rect 80908 7120 80948 7160
rect 80812 6952 80852 6992
rect 80908 6868 80948 6908
rect 81196 7456 81236 7496
rect 81100 7372 81140 7412
rect 81196 7120 81236 7160
rect 80908 6616 80948 6656
rect 80140 6364 80180 6404
rect 80524 6364 80564 6404
rect 81004 6364 81044 6404
rect 652 5608 692 5648
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 7112 6028 7152 6068
rect 7194 6028 7234 6068
rect 7276 6028 7316 6068
rect 7358 6028 7398 6068
rect 7440 6028 7480 6068
rect 11112 6028 11152 6068
rect 11194 6028 11234 6068
rect 11276 6028 11316 6068
rect 11358 6028 11398 6068
rect 11440 6028 11480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 19112 6028 19152 6068
rect 19194 6028 19234 6068
rect 19276 6028 19316 6068
rect 19358 6028 19398 6068
rect 19440 6028 19480 6068
rect 23112 6028 23152 6068
rect 23194 6028 23234 6068
rect 23276 6028 23316 6068
rect 23358 6028 23398 6068
rect 23440 6028 23480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 31112 6028 31152 6068
rect 31194 6028 31234 6068
rect 31276 6028 31316 6068
rect 31358 6028 31398 6068
rect 31440 6028 31480 6068
rect 35112 6028 35152 6068
rect 35194 6028 35234 6068
rect 35276 6028 35316 6068
rect 35358 6028 35398 6068
rect 35440 6028 35480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 43112 6028 43152 6068
rect 43194 6028 43234 6068
rect 43276 6028 43316 6068
rect 43358 6028 43398 6068
rect 43440 6028 43480 6068
rect 47112 6028 47152 6068
rect 47194 6028 47234 6068
rect 47276 6028 47316 6068
rect 47358 6028 47398 6068
rect 47440 6028 47480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 55112 6028 55152 6068
rect 55194 6028 55234 6068
rect 55276 6028 55316 6068
rect 55358 6028 55398 6068
rect 55440 6028 55480 6068
rect 59112 6028 59152 6068
rect 59194 6028 59234 6068
rect 59276 6028 59316 6068
rect 59358 6028 59398 6068
rect 59440 6028 59480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 67112 6028 67152 6068
rect 67194 6028 67234 6068
rect 67276 6028 67316 6068
rect 67358 6028 67398 6068
rect 67440 6028 67480 6068
rect 81676 7372 81716 7412
rect 81580 7204 81620 7244
rect 82060 7540 82100 7580
rect 82060 7120 82100 7160
rect 81196 6364 81236 6404
rect 81964 6952 82004 6992
rect 82348 7456 82388 7496
rect 82540 7372 82580 7412
rect 82444 7288 82484 7328
rect 82252 7120 82292 7160
rect 82636 7120 82676 7160
rect 81772 6364 81812 6404
rect 82060 6364 82100 6404
rect 82828 7540 82868 7580
rect 82924 7456 82964 7496
rect 82924 7120 82964 7160
rect 82540 6364 82580 6404
rect 83212 7204 83252 7244
rect 83615 7624 83655 7664
rect 83404 6364 83444 6404
rect 83596 7288 83636 7328
rect 83692 7120 83732 7160
rect 83980 7456 84020 7496
rect 84172 7624 84212 7664
rect 84415 7792 84455 7832
rect 84076 7372 84116 7412
rect 83884 7120 83924 7160
rect 84268 6952 84308 6992
rect 85324 7792 85364 7832
rect 84460 7372 84500 7412
rect 84556 6952 84596 6992
rect 83692 6364 83732 6404
rect 84076 6364 84116 6404
rect 84844 7456 84884 7496
rect 84844 7204 84884 7244
rect 85036 7120 85076 7160
rect 85228 7372 85268 7412
rect 85228 6952 85268 6992
rect 85516 7456 85556 7496
rect 85804 7372 85844 7412
rect 85708 7288 85748 7328
rect 85612 7120 85652 7160
rect 85900 7120 85940 7160
rect 84460 6364 84500 6404
rect 84844 6364 84884 6404
rect 86284 7204 86324 7244
rect 86188 7036 86228 7076
rect 86668 7456 86708 7496
rect 86476 7372 86516 7412
rect 86476 7204 86516 7244
rect 86668 6868 86708 6908
rect 86860 7456 86900 7496
rect 86860 7288 86900 7328
rect 86956 7120 86996 7160
rect 87436 7372 87476 7412
rect 87244 7288 87284 7328
rect 87148 7120 87188 7160
rect 87340 7120 87380 7160
rect 87532 7120 87572 7160
rect 87244 7036 87284 7076
rect 87820 7540 87860 7580
rect 87724 7456 87764 7496
rect 87820 7120 87860 7160
rect 88012 7372 88052 7412
rect 88204 7204 88244 7244
rect 88396 7456 88436 7496
rect 88396 7288 88436 7328
rect 88492 7120 88532 7160
rect 88780 7540 88820 7580
rect 88972 7372 89012 7412
rect 88876 7288 88916 7328
rect 88684 7120 88724 7160
rect 88876 7120 88916 7160
rect 89068 7120 89108 7160
rect 89615 7708 89655 7748
rect 89260 7372 89300 7412
rect 89260 7204 89300 7244
rect 89452 7036 89492 7076
rect 90508 7708 90548 7748
rect 89644 7456 89684 7496
rect 89740 7120 89780 7160
rect 90028 7456 90068 7496
rect 90220 7372 90260 7412
rect 90028 7288 90068 7328
rect 89932 7120 89972 7160
rect 90316 7120 90356 7160
rect 90988 7708 91028 7748
rect 90815 7624 90855 7664
rect 90604 7372 90644 7412
rect 90604 7120 90644 7160
rect 85324 6364 85364 6404
rect 86092 6364 86132 6404
rect 86476 6364 86516 6404
rect 86860 6364 86900 6404
rect 87340 6364 87380 6404
rect 87916 6364 87956 6404
rect 88108 6364 88148 6404
rect 88492 6364 88532 6404
rect 88876 6364 88916 6404
rect 89260 6364 89300 6404
rect 89740 6364 89780 6404
rect 90124 6364 90164 6404
rect 91215 7708 91255 7748
rect 90796 7204 90836 7244
rect 90988 7204 91028 7244
rect 90508 6364 90548 6404
rect 91276 7372 91316 7412
rect 91180 7204 91220 7244
rect 90988 6364 91028 6404
rect 91276 7120 91316 7160
rect 91564 7288 91604 7328
rect 91756 7624 91796 7664
rect 91852 7288 91892 7328
rect 91660 7204 91700 7244
rect 91468 7120 91508 7160
rect 91276 6364 91316 6404
rect 91756 6364 91796 6404
rect 92044 6952 92084 6992
rect 92428 7456 92468 7496
rect 92332 7036 92372 7076
rect 92524 7036 92564 7076
rect 92812 7372 92852 7412
rect 93004 7288 93044 7328
rect 92908 7204 92948 7244
rect 92716 6868 92756 6908
rect 93905 7792 93945 7832
rect 93196 7288 93236 7328
rect 93484 7456 93524 7496
rect 93580 7288 93620 7328
rect 93292 7120 93332 7160
rect 93292 6952 93332 6992
rect 93772 7540 93812 7580
rect 93772 7372 93812 7412
rect 93868 7288 93908 7328
rect 94252 7036 94292 7076
rect 93772 6616 93812 6656
rect 93964 6448 94004 6488
rect 92140 6364 92180 6404
rect 92524 6364 92564 6404
rect 92908 6364 92948 6404
rect 93388 6364 93428 6404
rect 94252 6868 94292 6908
rect 94540 7288 94580 7328
rect 94444 7204 94484 7244
rect 94540 7120 94580 7160
rect 94444 7036 94484 7076
rect 94924 7540 94964 7580
rect 94828 7288 94868 7328
rect 94732 7120 94772 7160
rect 95308 7120 95348 7160
rect 95212 6868 95252 6908
rect 94156 6448 94196 6488
rect 94540 6448 94580 6488
rect 94924 6448 94964 6488
rect 95596 7372 95636 7412
rect 95980 7288 96020 7328
rect 95596 7204 95636 7244
rect 96268 7288 96308 7328
rect 96172 7204 96212 7244
rect 96268 7036 96308 7076
rect 95692 6448 95732 6488
rect 96460 7372 96500 7412
rect 96556 7204 96596 7244
rect 96556 7036 96596 7076
rect 95404 6364 95444 6404
rect 95788 6364 95828 6404
rect 96172 6364 96212 6404
rect 96652 6952 96692 6992
rect 96844 7372 96884 7412
rect 96844 6868 96884 6908
rect 97036 6784 97076 6824
rect 97505 7624 97545 7664
rect 97708 7624 97748 7664
rect 97228 7288 97268 7328
rect 97324 7204 97364 7244
rect 97228 7120 97268 7160
rect 97612 7120 97652 7160
rect 97612 6952 97652 6992
rect 97228 6784 97268 6824
rect 97804 7372 97844 7412
rect 97228 6364 97268 6404
rect 98092 7456 98132 7496
rect 98284 7372 98324 7412
rect 98092 7288 98132 7328
rect 98188 6952 98228 6992
rect 97708 6364 97748 6404
rect 98476 7372 98516 7412
rect 99244 7456 99284 7496
rect 98860 7036 98900 7076
rect 98956 6952 98996 6992
rect 98092 6364 98132 6404
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 8352 5272 8392 5312
rect 8434 5272 8474 5312
rect 8516 5272 8556 5312
rect 8598 5272 8638 5312
rect 8680 5272 8720 5312
rect 12352 5272 12392 5312
rect 12434 5272 12474 5312
rect 12516 5272 12556 5312
rect 12598 5272 12638 5312
rect 12680 5272 12720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 20352 5272 20392 5312
rect 20434 5272 20474 5312
rect 20516 5272 20556 5312
rect 20598 5272 20638 5312
rect 20680 5272 20720 5312
rect 24352 5272 24392 5312
rect 24434 5272 24474 5312
rect 24516 5272 24556 5312
rect 24598 5272 24638 5312
rect 24680 5272 24720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 32352 5272 32392 5312
rect 32434 5272 32474 5312
rect 32516 5272 32556 5312
rect 32598 5272 32638 5312
rect 32680 5272 32720 5312
rect 36352 5272 36392 5312
rect 36434 5272 36474 5312
rect 36516 5272 36556 5312
rect 36598 5272 36638 5312
rect 36680 5272 36720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 44352 5272 44392 5312
rect 44434 5272 44474 5312
rect 44516 5272 44556 5312
rect 44598 5272 44638 5312
rect 44680 5272 44720 5312
rect 48352 5272 48392 5312
rect 48434 5272 48474 5312
rect 48516 5272 48556 5312
rect 48598 5272 48638 5312
rect 48680 5272 48720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 56352 5272 56392 5312
rect 56434 5272 56474 5312
rect 56516 5272 56556 5312
rect 56598 5272 56638 5312
rect 56680 5272 56720 5312
rect 60352 5272 60392 5312
rect 60434 5272 60474 5312
rect 60516 5272 60556 5312
rect 60598 5272 60638 5312
rect 60680 5272 60720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 68352 5272 68392 5312
rect 68434 5272 68474 5312
rect 68516 5272 68556 5312
rect 68598 5272 68638 5312
rect 68680 5272 68720 5312
rect 72352 5272 72392 5312
rect 72434 5272 72474 5312
rect 72516 5272 72556 5312
rect 72598 5272 72638 5312
rect 72680 5272 72720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 80352 5272 80392 5312
rect 80434 5272 80474 5312
rect 80516 5272 80556 5312
rect 80598 5272 80638 5312
rect 80680 5272 80720 5312
rect 84352 5272 84392 5312
rect 84434 5272 84474 5312
rect 84516 5272 84556 5312
rect 84598 5272 84638 5312
rect 84680 5272 84720 5312
rect 88352 5272 88392 5312
rect 88434 5272 88474 5312
rect 88516 5272 88556 5312
rect 88598 5272 88638 5312
rect 88680 5272 88720 5312
rect 92352 5272 92392 5312
rect 92434 5272 92474 5312
rect 92516 5272 92556 5312
rect 92598 5272 92638 5312
rect 92680 5272 92720 5312
rect 96352 5272 96392 5312
rect 96434 5272 96474 5312
rect 96516 5272 96556 5312
rect 96598 5272 96638 5312
rect 96680 5272 96720 5312
rect 1036 4852 1076 4892
rect 1420 4852 1460 4892
rect 1804 4852 1844 4892
rect 2188 4852 2228 4892
rect 652 4768 692 4808
rect 748 4684 788 4724
rect 652 3172 692 3212
rect 844 4180 884 4220
rect 1996 4684 2036 4724
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 7112 4516 7152 4556
rect 7194 4516 7234 4556
rect 7276 4516 7316 4556
rect 7358 4516 7398 4556
rect 7440 4516 7480 4556
rect 11112 4516 11152 4556
rect 11194 4516 11234 4556
rect 11276 4516 11316 4556
rect 11358 4516 11398 4556
rect 11440 4516 11480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 19112 4516 19152 4556
rect 19194 4516 19234 4556
rect 19276 4516 19316 4556
rect 19358 4516 19398 4556
rect 19440 4516 19480 4556
rect 23112 4516 23152 4556
rect 23194 4516 23234 4556
rect 23276 4516 23316 4556
rect 23358 4516 23398 4556
rect 23440 4516 23480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 31112 4516 31152 4556
rect 31194 4516 31234 4556
rect 31276 4516 31316 4556
rect 31358 4516 31398 4556
rect 31440 4516 31480 4556
rect 35112 4516 35152 4556
rect 35194 4516 35234 4556
rect 35276 4516 35316 4556
rect 35358 4516 35398 4556
rect 35440 4516 35480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 43112 4516 43152 4556
rect 43194 4516 43234 4556
rect 43276 4516 43316 4556
rect 43358 4516 43398 4556
rect 43440 4516 43480 4556
rect 47112 4516 47152 4556
rect 47194 4516 47234 4556
rect 47276 4516 47316 4556
rect 47358 4516 47398 4556
rect 47440 4516 47480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 55112 4516 55152 4556
rect 55194 4516 55234 4556
rect 55276 4516 55316 4556
rect 55358 4516 55398 4556
rect 55440 4516 55480 4556
rect 59112 4516 59152 4556
rect 59194 4516 59234 4556
rect 59276 4516 59316 4556
rect 59358 4516 59398 4556
rect 59440 4516 59480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 67112 4516 67152 4556
rect 67194 4516 67234 4556
rect 67276 4516 67316 4556
rect 67358 4516 67398 4556
rect 67440 4516 67480 4556
rect 71112 4516 71152 4556
rect 71194 4516 71234 4556
rect 71276 4516 71316 4556
rect 71358 4516 71398 4556
rect 71440 4516 71480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 79112 4516 79152 4556
rect 79194 4516 79234 4556
rect 79276 4516 79316 4556
rect 79358 4516 79398 4556
rect 79440 4516 79480 4556
rect 83112 4516 83152 4556
rect 83194 4516 83234 4556
rect 83276 4516 83316 4556
rect 83358 4516 83398 4556
rect 83440 4516 83480 4556
rect 87112 4516 87152 4556
rect 87194 4516 87234 4556
rect 87276 4516 87316 4556
rect 87358 4516 87398 4556
rect 87440 4516 87480 4556
rect 91112 4516 91152 4556
rect 91194 4516 91234 4556
rect 91276 4516 91316 4556
rect 91358 4516 91398 4556
rect 91440 4516 91480 4556
rect 95112 4516 95152 4556
rect 95194 4516 95234 4556
rect 95276 4516 95316 4556
rect 95358 4516 95398 4556
rect 95440 4516 95480 4556
rect 99112 4516 99152 4556
rect 99194 4516 99234 4556
rect 99276 4516 99316 4556
rect 99358 4516 99398 4556
rect 99440 4516 99480 4556
rect 1612 4180 1652 4220
rect 1036 3928 1076 3968
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 8352 3760 8392 3800
rect 8434 3760 8474 3800
rect 8516 3760 8556 3800
rect 8598 3760 8638 3800
rect 8680 3760 8720 3800
rect 12352 3760 12392 3800
rect 12434 3760 12474 3800
rect 12516 3760 12556 3800
rect 12598 3760 12638 3800
rect 12680 3760 12720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 20352 3760 20392 3800
rect 20434 3760 20474 3800
rect 20516 3760 20556 3800
rect 20598 3760 20638 3800
rect 20680 3760 20720 3800
rect 24352 3760 24392 3800
rect 24434 3760 24474 3800
rect 24516 3760 24556 3800
rect 24598 3760 24638 3800
rect 24680 3760 24720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 32352 3760 32392 3800
rect 32434 3760 32474 3800
rect 32516 3760 32556 3800
rect 32598 3760 32638 3800
rect 32680 3760 32720 3800
rect 36352 3760 36392 3800
rect 36434 3760 36474 3800
rect 36516 3760 36556 3800
rect 36598 3760 36638 3800
rect 36680 3760 36720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 44352 3760 44392 3800
rect 44434 3760 44474 3800
rect 44516 3760 44556 3800
rect 44598 3760 44638 3800
rect 44680 3760 44720 3800
rect 48352 3760 48392 3800
rect 48434 3760 48474 3800
rect 48516 3760 48556 3800
rect 48598 3760 48638 3800
rect 48680 3760 48720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 56352 3760 56392 3800
rect 56434 3760 56474 3800
rect 56516 3760 56556 3800
rect 56598 3760 56638 3800
rect 56680 3760 56720 3800
rect 60352 3760 60392 3800
rect 60434 3760 60474 3800
rect 60516 3760 60556 3800
rect 60598 3760 60638 3800
rect 60680 3760 60720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 68352 3760 68392 3800
rect 68434 3760 68474 3800
rect 68516 3760 68556 3800
rect 68598 3760 68638 3800
rect 68680 3760 68720 3800
rect 72352 3760 72392 3800
rect 72434 3760 72474 3800
rect 72516 3760 72556 3800
rect 72598 3760 72638 3800
rect 72680 3760 72720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 80352 3760 80392 3800
rect 80434 3760 80474 3800
rect 80516 3760 80556 3800
rect 80598 3760 80638 3800
rect 80680 3760 80720 3800
rect 84352 3760 84392 3800
rect 84434 3760 84474 3800
rect 84516 3760 84556 3800
rect 84598 3760 84638 3800
rect 84680 3760 84720 3800
rect 88352 3760 88392 3800
rect 88434 3760 88474 3800
rect 88516 3760 88556 3800
rect 88598 3760 88638 3800
rect 88680 3760 88720 3800
rect 92352 3760 92392 3800
rect 92434 3760 92474 3800
rect 92516 3760 92556 3800
rect 92598 3760 92638 3800
rect 92680 3760 92720 3800
rect 96352 3760 96392 3800
rect 96434 3760 96474 3800
rect 96516 3760 96556 3800
rect 96598 3760 96638 3800
rect 96680 3760 96720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 7112 3004 7152 3044
rect 7194 3004 7234 3044
rect 7276 3004 7316 3044
rect 7358 3004 7398 3044
rect 7440 3004 7480 3044
rect 11112 3004 11152 3044
rect 11194 3004 11234 3044
rect 11276 3004 11316 3044
rect 11358 3004 11398 3044
rect 11440 3004 11480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 19112 3004 19152 3044
rect 19194 3004 19234 3044
rect 19276 3004 19316 3044
rect 19358 3004 19398 3044
rect 19440 3004 19480 3044
rect 23112 3004 23152 3044
rect 23194 3004 23234 3044
rect 23276 3004 23316 3044
rect 23358 3004 23398 3044
rect 23440 3004 23480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 31112 3004 31152 3044
rect 31194 3004 31234 3044
rect 31276 3004 31316 3044
rect 31358 3004 31398 3044
rect 31440 3004 31480 3044
rect 35112 3004 35152 3044
rect 35194 3004 35234 3044
rect 35276 3004 35316 3044
rect 35358 3004 35398 3044
rect 35440 3004 35480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 43112 3004 43152 3044
rect 43194 3004 43234 3044
rect 43276 3004 43316 3044
rect 43358 3004 43398 3044
rect 43440 3004 43480 3044
rect 47112 3004 47152 3044
rect 47194 3004 47234 3044
rect 47276 3004 47316 3044
rect 47358 3004 47398 3044
rect 47440 3004 47480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 55112 3004 55152 3044
rect 55194 3004 55234 3044
rect 55276 3004 55316 3044
rect 55358 3004 55398 3044
rect 55440 3004 55480 3044
rect 59112 3004 59152 3044
rect 59194 3004 59234 3044
rect 59276 3004 59316 3044
rect 59358 3004 59398 3044
rect 59440 3004 59480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 67112 3004 67152 3044
rect 67194 3004 67234 3044
rect 67276 3004 67316 3044
rect 67358 3004 67398 3044
rect 67440 3004 67480 3044
rect 71112 3004 71152 3044
rect 71194 3004 71234 3044
rect 71276 3004 71316 3044
rect 71358 3004 71398 3044
rect 71440 3004 71480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 79112 3004 79152 3044
rect 79194 3004 79234 3044
rect 79276 3004 79316 3044
rect 79358 3004 79398 3044
rect 79440 3004 79480 3044
rect 83112 3004 83152 3044
rect 83194 3004 83234 3044
rect 83276 3004 83316 3044
rect 83358 3004 83398 3044
rect 83440 3004 83480 3044
rect 87112 3004 87152 3044
rect 87194 3004 87234 3044
rect 87276 3004 87316 3044
rect 87358 3004 87398 3044
rect 87440 3004 87480 3044
rect 91112 3004 91152 3044
rect 91194 3004 91234 3044
rect 91276 3004 91316 3044
rect 91358 3004 91398 3044
rect 91440 3004 91480 3044
rect 95112 3004 95152 3044
rect 95194 3004 95234 3044
rect 95276 3004 95316 3044
rect 95358 3004 95398 3044
rect 95440 3004 95480 3044
rect 99112 3004 99152 3044
rect 99194 3004 99234 3044
rect 99276 3004 99316 3044
rect 99358 3004 99398 3044
rect 99440 3004 99480 3044
rect 652 2248 692 2288
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 8352 2248 8392 2288
rect 8434 2248 8474 2288
rect 8516 2248 8556 2288
rect 8598 2248 8638 2288
rect 8680 2248 8720 2288
rect 12352 2248 12392 2288
rect 12434 2248 12474 2288
rect 12516 2248 12556 2288
rect 12598 2248 12638 2288
rect 12680 2248 12720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 20352 2248 20392 2288
rect 20434 2248 20474 2288
rect 20516 2248 20556 2288
rect 20598 2248 20638 2288
rect 20680 2248 20720 2288
rect 24352 2248 24392 2288
rect 24434 2248 24474 2288
rect 24516 2248 24556 2288
rect 24598 2248 24638 2288
rect 24680 2248 24720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 32352 2248 32392 2288
rect 32434 2248 32474 2288
rect 32516 2248 32556 2288
rect 32598 2248 32638 2288
rect 32680 2248 32720 2288
rect 36352 2248 36392 2288
rect 36434 2248 36474 2288
rect 36516 2248 36556 2288
rect 36598 2248 36638 2288
rect 36680 2248 36720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 44352 2248 44392 2288
rect 44434 2248 44474 2288
rect 44516 2248 44556 2288
rect 44598 2248 44638 2288
rect 44680 2248 44720 2288
rect 48352 2248 48392 2288
rect 48434 2248 48474 2288
rect 48516 2248 48556 2288
rect 48598 2248 48638 2288
rect 48680 2248 48720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 56352 2248 56392 2288
rect 56434 2248 56474 2288
rect 56516 2248 56556 2288
rect 56598 2248 56638 2288
rect 56680 2248 56720 2288
rect 60352 2248 60392 2288
rect 60434 2248 60474 2288
rect 60516 2248 60556 2288
rect 60598 2248 60638 2288
rect 60680 2248 60720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 68352 2248 68392 2288
rect 68434 2248 68474 2288
rect 68516 2248 68556 2288
rect 68598 2248 68638 2288
rect 68680 2248 68720 2288
rect 72352 2248 72392 2288
rect 72434 2248 72474 2288
rect 72516 2248 72556 2288
rect 72598 2248 72638 2288
rect 72680 2248 72720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 80352 2248 80392 2288
rect 80434 2248 80474 2288
rect 80516 2248 80556 2288
rect 80598 2248 80638 2288
rect 80680 2248 80720 2288
rect 84352 2248 84392 2288
rect 84434 2248 84474 2288
rect 84516 2248 84556 2288
rect 84598 2248 84638 2288
rect 84680 2248 84720 2288
rect 88352 2248 88392 2288
rect 88434 2248 88474 2288
rect 88516 2248 88556 2288
rect 88598 2248 88638 2288
rect 88680 2248 88720 2288
rect 92352 2248 92392 2288
rect 92434 2248 92474 2288
rect 92516 2248 92556 2288
rect 92598 2248 92638 2288
rect 92680 2248 92720 2288
rect 96352 2248 96392 2288
rect 96434 2248 96474 2288
rect 96516 2248 96556 2288
rect 96598 2248 96638 2288
rect 96680 2248 96720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 7112 1492 7152 1532
rect 7194 1492 7234 1532
rect 7276 1492 7316 1532
rect 7358 1492 7398 1532
rect 7440 1492 7480 1532
rect 11112 1492 11152 1532
rect 11194 1492 11234 1532
rect 11276 1492 11316 1532
rect 11358 1492 11398 1532
rect 11440 1492 11480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 19112 1492 19152 1532
rect 19194 1492 19234 1532
rect 19276 1492 19316 1532
rect 19358 1492 19398 1532
rect 19440 1492 19480 1532
rect 23112 1492 23152 1532
rect 23194 1492 23234 1532
rect 23276 1492 23316 1532
rect 23358 1492 23398 1532
rect 23440 1492 23480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 31112 1492 31152 1532
rect 31194 1492 31234 1532
rect 31276 1492 31316 1532
rect 31358 1492 31398 1532
rect 31440 1492 31480 1532
rect 35112 1492 35152 1532
rect 35194 1492 35234 1532
rect 35276 1492 35316 1532
rect 35358 1492 35398 1532
rect 35440 1492 35480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 43112 1492 43152 1532
rect 43194 1492 43234 1532
rect 43276 1492 43316 1532
rect 43358 1492 43398 1532
rect 43440 1492 43480 1532
rect 47112 1492 47152 1532
rect 47194 1492 47234 1532
rect 47276 1492 47316 1532
rect 47358 1492 47398 1532
rect 47440 1492 47480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 55112 1492 55152 1532
rect 55194 1492 55234 1532
rect 55276 1492 55316 1532
rect 55358 1492 55398 1532
rect 55440 1492 55480 1532
rect 59112 1492 59152 1532
rect 59194 1492 59234 1532
rect 59276 1492 59316 1532
rect 59358 1492 59398 1532
rect 59440 1492 59480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 67112 1492 67152 1532
rect 67194 1492 67234 1532
rect 67276 1492 67316 1532
rect 67358 1492 67398 1532
rect 67440 1492 67480 1532
rect 71112 1492 71152 1532
rect 71194 1492 71234 1532
rect 71276 1492 71316 1532
rect 71358 1492 71398 1532
rect 71440 1492 71480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 79112 1492 79152 1532
rect 79194 1492 79234 1532
rect 79276 1492 79316 1532
rect 79358 1492 79398 1532
rect 79440 1492 79480 1532
rect 83112 1492 83152 1532
rect 83194 1492 83234 1532
rect 83276 1492 83316 1532
rect 83358 1492 83398 1532
rect 83440 1492 83480 1532
rect 87112 1492 87152 1532
rect 87194 1492 87234 1532
rect 87276 1492 87316 1532
rect 87358 1492 87398 1532
rect 87440 1492 87480 1532
rect 91112 1492 91152 1532
rect 91194 1492 91234 1532
rect 91276 1492 91316 1532
rect 91358 1492 91398 1532
rect 91440 1492 91480 1532
rect 95112 1492 95152 1532
rect 95194 1492 95234 1532
rect 95276 1492 95316 1532
rect 95358 1492 95398 1532
rect 95440 1492 95480 1532
rect 99112 1492 99152 1532
rect 99194 1492 99234 1532
rect 99276 1492 99316 1532
rect 99358 1492 99398 1532
rect 99440 1492 99480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 8352 736 8392 776
rect 8434 736 8474 776
rect 8516 736 8556 776
rect 8598 736 8638 776
rect 8680 736 8720 776
rect 12352 736 12392 776
rect 12434 736 12474 776
rect 12516 736 12556 776
rect 12598 736 12638 776
rect 12680 736 12720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 20352 736 20392 776
rect 20434 736 20474 776
rect 20516 736 20556 776
rect 20598 736 20638 776
rect 20680 736 20720 776
rect 24352 736 24392 776
rect 24434 736 24474 776
rect 24516 736 24556 776
rect 24598 736 24638 776
rect 24680 736 24720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 32352 736 32392 776
rect 32434 736 32474 776
rect 32516 736 32556 776
rect 32598 736 32638 776
rect 32680 736 32720 776
rect 36352 736 36392 776
rect 36434 736 36474 776
rect 36516 736 36556 776
rect 36598 736 36638 776
rect 36680 736 36720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 44352 736 44392 776
rect 44434 736 44474 776
rect 44516 736 44556 776
rect 44598 736 44638 776
rect 44680 736 44720 776
rect 48352 736 48392 776
rect 48434 736 48474 776
rect 48516 736 48556 776
rect 48598 736 48638 776
rect 48680 736 48720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 56352 736 56392 776
rect 56434 736 56474 776
rect 56516 736 56556 776
rect 56598 736 56638 776
rect 56680 736 56720 776
rect 60352 736 60392 776
rect 60434 736 60474 776
rect 60516 736 60556 776
rect 60598 736 60638 776
rect 60680 736 60720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 68352 736 68392 776
rect 68434 736 68474 776
rect 68516 736 68556 776
rect 68598 736 68638 776
rect 68680 736 68720 776
rect 72352 736 72392 776
rect 72434 736 72474 776
rect 72516 736 72556 776
rect 72598 736 72638 776
rect 72680 736 72720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
rect 80352 736 80392 776
rect 80434 736 80474 776
rect 80516 736 80556 776
rect 80598 736 80638 776
rect 80680 736 80720 776
rect 84352 736 84392 776
rect 84434 736 84474 776
rect 84516 736 84556 776
rect 84598 736 84638 776
rect 84680 736 84720 776
rect 88352 736 88392 776
rect 88434 736 88474 776
rect 88516 736 88556 776
rect 88598 736 88638 776
rect 88680 736 88720 776
rect 92352 736 92392 776
rect 92434 736 92474 776
rect 92516 736 92556 776
rect 92598 736 92638 776
rect 92680 736 92720 776
rect 96352 736 96392 776
rect 96434 736 96474 776
rect 96516 736 96556 776
rect 96598 736 96638 776
rect 96680 736 96720 776
<< metal3 >>
rect 4343 38536 4352 38576
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4720 38536 4729 38576
rect 8343 38536 8352 38576
rect 8392 38536 8434 38576
rect 8474 38536 8516 38576
rect 8556 38536 8598 38576
rect 8638 38536 8680 38576
rect 8720 38536 8729 38576
rect 12343 38536 12352 38576
rect 12392 38536 12434 38576
rect 12474 38536 12516 38576
rect 12556 38536 12598 38576
rect 12638 38536 12680 38576
rect 12720 38536 12729 38576
rect 16343 38536 16352 38576
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16720 38536 16729 38576
rect 20343 38536 20352 38576
rect 20392 38536 20434 38576
rect 20474 38536 20516 38576
rect 20556 38536 20598 38576
rect 20638 38536 20680 38576
rect 20720 38536 20729 38576
rect 24343 38536 24352 38576
rect 24392 38536 24434 38576
rect 24474 38536 24516 38576
rect 24556 38536 24598 38576
rect 24638 38536 24680 38576
rect 24720 38536 24729 38576
rect 28343 38536 28352 38576
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28720 38536 28729 38576
rect 32343 38536 32352 38576
rect 32392 38536 32434 38576
rect 32474 38536 32516 38576
rect 32556 38536 32598 38576
rect 32638 38536 32680 38576
rect 32720 38536 32729 38576
rect 36343 38536 36352 38576
rect 36392 38536 36434 38576
rect 36474 38536 36516 38576
rect 36556 38536 36598 38576
rect 36638 38536 36680 38576
rect 36720 38536 36729 38576
rect 40343 38536 40352 38576
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40720 38536 40729 38576
rect 44343 38536 44352 38576
rect 44392 38536 44434 38576
rect 44474 38536 44516 38576
rect 44556 38536 44598 38576
rect 44638 38536 44680 38576
rect 44720 38536 44729 38576
rect 48343 38536 48352 38576
rect 48392 38536 48434 38576
rect 48474 38536 48516 38576
rect 48556 38536 48598 38576
rect 48638 38536 48680 38576
rect 48720 38536 48729 38576
rect 52343 38536 52352 38576
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52720 38536 52729 38576
rect 56343 38536 56352 38576
rect 56392 38536 56434 38576
rect 56474 38536 56516 38576
rect 56556 38536 56598 38576
rect 56638 38536 56680 38576
rect 56720 38536 56729 38576
rect 60343 38536 60352 38576
rect 60392 38536 60434 38576
rect 60474 38536 60516 38576
rect 60556 38536 60598 38576
rect 60638 38536 60680 38576
rect 60720 38536 60729 38576
rect 64343 38536 64352 38576
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64720 38536 64729 38576
rect 68343 38536 68352 38576
rect 68392 38536 68434 38576
rect 68474 38536 68516 38576
rect 68556 38536 68598 38576
rect 68638 38536 68680 38576
rect 68720 38536 68729 38576
rect 72343 38536 72352 38576
rect 72392 38536 72434 38576
rect 72474 38536 72516 38576
rect 72556 38536 72598 38576
rect 72638 38536 72680 38576
rect 72720 38536 72729 38576
rect 76343 38536 76352 38576
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76720 38536 76729 38576
rect 80343 38536 80352 38576
rect 80392 38536 80434 38576
rect 80474 38536 80516 38576
rect 80556 38536 80598 38576
rect 80638 38536 80680 38576
rect 80720 38536 80729 38576
rect 84343 38536 84352 38576
rect 84392 38536 84434 38576
rect 84474 38536 84516 38576
rect 84556 38536 84598 38576
rect 84638 38536 84680 38576
rect 84720 38536 84729 38576
rect 88343 38536 88352 38576
rect 88392 38536 88434 38576
rect 88474 38536 88516 38576
rect 88556 38536 88598 38576
rect 88638 38536 88680 38576
rect 88720 38536 88729 38576
rect 92343 38536 92352 38576
rect 92392 38536 92434 38576
rect 92474 38536 92516 38576
rect 92556 38536 92598 38576
rect 92638 38536 92680 38576
rect 92720 38536 92729 38576
rect 96343 38536 96352 38576
rect 96392 38536 96434 38576
rect 96474 38536 96516 38576
rect 96556 38536 96598 38576
rect 96638 38536 96680 38576
rect 96720 38536 96729 38576
rect 3103 37780 3112 37820
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3480 37780 3489 37820
rect 7103 37780 7112 37820
rect 7152 37780 7194 37820
rect 7234 37780 7276 37820
rect 7316 37780 7358 37820
rect 7398 37780 7440 37820
rect 7480 37780 7489 37820
rect 11103 37780 11112 37820
rect 11152 37780 11194 37820
rect 11234 37780 11276 37820
rect 11316 37780 11358 37820
rect 11398 37780 11440 37820
rect 11480 37780 11489 37820
rect 15103 37780 15112 37820
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15480 37780 15489 37820
rect 19103 37780 19112 37820
rect 19152 37780 19194 37820
rect 19234 37780 19276 37820
rect 19316 37780 19358 37820
rect 19398 37780 19440 37820
rect 19480 37780 19489 37820
rect 23103 37780 23112 37820
rect 23152 37780 23194 37820
rect 23234 37780 23276 37820
rect 23316 37780 23358 37820
rect 23398 37780 23440 37820
rect 23480 37780 23489 37820
rect 27103 37780 27112 37820
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27480 37780 27489 37820
rect 31103 37780 31112 37820
rect 31152 37780 31194 37820
rect 31234 37780 31276 37820
rect 31316 37780 31358 37820
rect 31398 37780 31440 37820
rect 31480 37780 31489 37820
rect 35103 37780 35112 37820
rect 35152 37780 35194 37820
rect 35234 37780 35276 37820
rect 35316 37780 35358 37820
rect 35398 37780 35440 37820
rect 35480 37780 35489 37820
rect 39103 37780 39112 37820
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39480 37780 39489 37820
rect 43103 37780 43112 37820
rect 43152 37780 43194 37820
rect 43234 37780 43276 37820
rect 43316 37780 43358 37820
rect 43398 37780 43440 37820
rect 43480 37780 43489 37820
rect 47103 37780 47112 37820
rect 47152 37780 47194 37820
rect 47234 37780 47276 37820
rect 47316 37780 47358 37820
rect 47398 37780 47440 37820
rect 47480 37780 47489 37820
rect 51103 37780 51112 37820
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51480 37780 51489 37820
rect 55103 37780 55112 37820
rect 55152 37780 55194 37820
rect 55234 37780 55276 37820
rect 55316 37780 55358 37820
rect 55398 37780 55440 37820
rect 55480 37780 55489 37820
rect 59103 37780 59112 37820
rect 59152 37780 59194 37820
rect 59234 37780 59276 37820
rect 59316 37780 59358 37820
rect 59398 37780 59440 37820
rect 59480 37780 59489 37820
rect 63103 37780 63112 37820
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63480 37780 63489 37820
rect 67103 37780 67112 37820
rect 67152 37780 67194 37820
rect 67234 37780 67276 37820
rect 67316 37780 67358 37820
rect 67398 37780 67440 37820
rect 67480 37780 67489 37820
rect 71103 37780 71112 37820
rect 71152 37780 71194 37820
rect 71234 37780 71276 37820
rect 71316 37780 71358 37820
rect 71398 37780 71440 37820
rect 71480 37780 71489 37820
rect 75103 37780 75112 37820
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75480 37780 75489 37820
rect 79103 37780 79112 37820
rect 79152 37780 79194 37820
rect 79234 37780 79276 37820
rect 79316 37780 79358 37820
rect 79398 37780 79440 37820
rect 79480 37780 79489 37820
rect 83103 37780 83112 37820
rect 83152 37780 83194 37820
rect 83234 37780 83276 37820
rect 83316 37780 83358 37820
rect 83398 37780 83440 37820
rect 83480 37780 83489 37820
rect 87103 37780 87112 37820
rect 87152 37780 87194 37820
rect 87234 37780 87276 37820
rect 87316 37780 87358 37820
rect 87398 37780 87440 37820
rect 87480 37780 87489 37820
rect 91103 37780 91112 37820
rect 91152 37780 91194 37820
rect 91234 37780 91276 37820
rect 91316 37780 91358 37820
rect 91398 37780 91440 37820
rect 91480 37780 91489 37820
rect 95103 37780 95112 37820
rect 95152 37780 95194 37820
rect 95234 37780 95276 37820
rect 95316 37780 95358 37820
rect 95398 37780 95440 37820
rect 95480 37780 95489 37820
rect 99103 37780 99112 37820
rect 99152 37780 99194 37820
rect 99234 37780 99276 37820
rect 99316 37780 99358 37820
rect 99398 37780 99440 37820
rect 99480 37780 99489 37820
rect 0 37508 80 37588
rect 4343 37024 4352 37064
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4720 37024 4729 37064
rect 8343 37024 8352 37064
rect 8392 37024 8434 37064
rect 8474 37024 8516 37064
rect 8556 37024 8598 37064
rect 8638 37024 8680 37064
rect 8720 37024 8729 37064
rect 12343 37024 12352 37064
rect 12392 37024 12434 37064
rect 12474 37024 12516 37064
rect 12556 37024 12598 37064
rect 12638 37024 12680 37064
rect 12720 37024 12729 37064
rect 16343 37024 16352 37064
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16720 37024 16729 37064
rect 20343 37024 20352 37064
rect 20392 37024 20434 37064
rect 20474 37024 20516 37064
rect 20556 37024 20598 37064
rect 20638 37024 20680 37064
rect 20720 37024 20729 37064
rect 24343 37024 24352 37064
rect 24392 37024 24434 37064
rect 24474 37024 24516 37064
rect 24556 37024 24598 37064
rect 24638 37024 24680 37064
rect 24720 37024 24729 37064
rect 28343 37024 28352 37064
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28720 37024 28729 37064
rect 32343 37024 32352 37064
rect 32392 37024 32434 37064
rect 32474 37024 32516 37064
rect 32556 37024 32598 37064
rect 32638 37024 32680 37064
rect 32720 37024 32729 37064
rect 36343 37024 36352 37064
rect 36392 37024 36434 37064
rect 36474 37024 36516 37064
rect 36556 37024 36598 37064
rect 36638 37024 36680 37064
rect 36720 37024 36729 37064
rect 40343 37024 40352 37064
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40720 37024 40729 37064
rect 44343 37024 44352 37064
rect 44392 37024 44434 37064
rect 44474 37024 44516 37064
rect 44556 37024 44598 37064
rect 44638 37024 44680 37064
rect 44720 37024 44729 37064
rect 48343 37024 48352 37064
rect 48392 37024 48434 37064
rect 48474 37024 48516 37064
rect 48556 37024 48598 37064
rect 48638 37024 48680 37064
rect 48720 37024 48729 37064
rect 52343 37024 52352 37064
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52720 37024 52729 37064
rect 56343 37024 56352 37064
rect 56392 37024 56434 37064
rect 56474 37024 56516 37064
rect 56556 37024 56598 37064
rect 56638 37024 56680 37064
rect 56720 37024 56729 37064
rect 60343 37024 60352 37064
rect 60392 37024 60434 37064
rect 60474 37024 60516 37064
rect 60556 37024 60598 37064
rect 60638 37024 60680 37064
rect 60720 37024 60729 37064
rect 64343 37024 64352 37064
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64720 37024 64729 37064
rect 68343 37024 68352 37064
rect 68392 37024 68434 37064
rect 68474 37024 68516 37064
rect 68556 37024 68598 37064
rect 68638 37024 68680 37064
rect 68720 37024 68729 37064
rect 72343 37024 72352 37064
rect 72392 37024 72434 37064
rect 72474 37024 72516 37064
rect 72556 37024 72598 37064
rect 72638 37024 72680 37064
rect 72720 37024 72729 37064
rect 76343 37024 76352 37064
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76720 37024 76729 37064
rect 80343 37024 80352 37064
rect 80392 37024 80434 37064
rect 80474 37024 80516 37064
rect 80556 37024 80598 37064
rect 80638 37024 80680 37064
rect 80720 37024 80729 37064
rect 84343 37024 84352 37064
rect 84392 37024 84434 37064
rect 84474 37024 84516 37064
rect 84556 37024 84598 37064
rect 84638 37024 84680 37064
rect 84720 37024 84729 37064
rect 88343 37024 88352 37064
rect 88392 37024 88434 37064
rect 88474 37024 88516 37064
rect 88556 37024 88598 37064
rect 88638 37024 88680 37064
rect 88720 37024 88729 37064
rect 92343 37024 92352 37064
rect 92392 37024 92434 37064
rect 92474 37024 92516 37064
rect 92556 37024 92598 37064
rect 92638 37024 92680 37064
rect 92720 37024 92729 37064
rect 96343 37024 96352 37064
rect 96392 37024 96434 37064
rect 96474 37024 96516 37064
rect 96556 37024 96598 37064
rect 96638 37024 96680 37064
rect 96720 37024 96729 37064
rect 0 36668 80 36748
rect 3103 36268 3112 36308
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3480 36268 3489 36308
rect 7103 36268 7112 36308
rect 7152 36268 7194 36308
rect 7234 36268 7276 36308
rect 7316 36268 7358 36308
rect 7398 36268 7440 36308
rect 7480 36268 7489 36308
rect 11103 36268 11112 36308
rect 11152 36268 11194 36308
rect 11234 36268 11276 36308
rect 11316 36268 11358 36308
rect 11398 36268 11440 36308
rect 11480 36268 11489 36308
rect 15103 36268 15112 36308
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15480 36268 15489 36308
rect 19103 36268 19112 36308
rect 19152 36268 19194 36308
rect 19234 36268 19276 36308
rect 19316 36268 19358 36308
rect 19398 36268 19440 36308
rect 19480 36268 19489 36308
rect 23103 36268 23112 36308
rect 23152 36268 23194 36308
rect 23234 36268 23276 36308
rect 23316 36268 23358 36308
rect 23398 36268 23440 36308
rect 23480 36268 23489 36308
rect 27103 36268 27112 36308
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27480 36268 27489 36308
rect 31103 36268 31112 36308
rect 31152 36268 31194 36308
rect 31234 36268 31276 36308
rect 31316 36268 31358 36308
rect 31398 36268 31440 36308
rect 31480 36268 31489 36308
rect 35103 36268 35112 36308
rect 35152 36268 35194 36308
rect 35234 36268 35276 36308
rect 35316 36268 35358 36308
rect 35398 36268 35440 36308
rect 35480 36268 35489 36308
rect 39103 36268 39112 36308
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39480 36268 39489 36308
rect 43103 36268 43112 36308
rect 43152 36268 43194 36308
rect 43234 36268 43276 36308
rect 43316 36268 43358 36308
rect 43398 36268 43440 36308
rect 43480 36268 43489 36308
rect 47103 36268 47112 36308
rect 47152 36268 47194 36308
rect 47234 36268 47276 36308
rect 47316 36268 47358 36308
rect 47398 36268 47440 36308
rect 47480 36268 47489 36308
rect 51103 36268 51112 36308
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51480 36268 51489 36308
rect 55103 36268 55112 36308
rect 55152 36268 55194 36308
rect 55234 36268 55276 36308
rect 55316 36268 55358 36308
rect 55398 36268 55440 36308
rect 55480 36268 55489 36308
rect 59103 36268 59112 36308
rect 59152 36268 59194 36308
rect 59234 36268 59276 36308
rect 59316 36268 59358 36308
rect 59398 36268 59440 36308
rect 59480 36268 59489 36308
rect 63103 36268 63112 36308
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63480 36268 63489 36308
rect 67103 36268 67112 36308
rect 67152 36268 67194 36308
rect 67234 36268 67276 36308
rect 67316 36268 67358 36308
rect 67398 36268 67440 36308
rect 67480 36268 67489 36308
rect 71103 36268 71112 36308
rect 71152 36268 71194 36308
rect 71234 36268 71276 36308
rect 71316 36268 71358 36308
rect 71398 36268 71440 36308
rect 71480 36268 71489 36308
rect 75103 36268 75112 36308
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75480 36268 75489 36308
rect 79103 36268 79112 36308
rect 79152 36268 79194 36308
rect 79234 36268 79276 36308
rect 79316 36268 79358 36308
rect 79398 36268 79440 36308
rect 79480 36268 79489 36308
rect 83103 36268 83112 36308
rect 83152 36268 83194 36308
rect 83234 36268 83276 36308
rect 83316 36268 83358 36308
rect 83398 36268 83440 36308
rect 83480 36268 83489 36308
rect 87103 36268 87112 36308
rect 87152 36268 87194 36308
rect 87234 36268 87276 36308
rect 87316 36268 87358 36308
rect 87398 36268 87440 36308
rect 87480 36268 87489 36308
rect 91103 36268 91112 36308
rect 91152 36268 91194 36308
rect 91234 36268 91276 36308
rect 91316 36268 91358 36308
rect 91398 36268 91440 36308
rect 91480 36268 91489 36308
rect 95103 36268 95112 36308
rect 95152 36268 95194 36308
rect 95234 36268 95276 36308
rect 95316 36268 95358 36308
rect 95398 36268 95440 36308
rect 95480 36268 95489 36308
rect 99103 36268 99112 36308
rect 99152 36268 99194 36308
rect 99234 36268 99276 36308
rect 99316 36268 99358 36308
rect 99398 36268 99440 36308
rect 99480 36268 99489 36308
rect 0 35828 80 35908
rect 4343 35512 4352 35552
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4720 35512 4729 35552
rect 8343 35512 8352 35552
rect 8392 35512 8434 35552
rect 8474 35512 8516 35552
rect 8556 35512 8598 35552
rect 8638 35512 8680 35552
rect 8720 35512 8729 35552
rect 12343 35512 12352 35552
rect 12392 35512 12434 35552
rect 12474 35512 12516 35552
rect 12556 35512 12598 35552
rect 12638 35512 12680 35552
rect 12720 35512 12729 35552
rect 16343 35512 16352 35552
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16720 35512 16729 35552
rect 20343 35512 20352 35552
rect 20392 35512 20434 35552
rect 20474 35512 20516 35552
rect 20556 35512 20598 35552
rect 20638 35512 20680 35552
rect 20720 35512 20729 35552
rect 24343 35512 24352 35552
rect 24392 35512 24434 35552
rect 24474 35512 24516 35552
rect 24556 35512 24598 35552
rect 24638 35512 24680 35552
rect 24720 35512 24729 35552
rect 28343 35512 28352 35552
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28720 35512 28729 35552
rect 32343 35512 32352 35552
rect 32392 35512 32434 35552
rect 32474 35512 32516 35552
rect 32556 35512 32598 35552
rect 32638 35512 32680 35552
rect 32720 35512 32729 35552
rect 36343 35512 36352 35552
rect 36392 35512 36434 35552
rect 36474 35512 36516 35552
rect 36556 35512 36598 35552
rect 36638 35512 36680 35552
rect 36720 35512 36729 35552
rect 40343 35512 40352 35552
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40720 35512 40729 35552
rect 44343 35512 44352 35552
rect 44392 35512 44434 35552
rect 44474 35512 44516 35552
rect 44556 35512 44598 35552
rect 44638 35512 44680 35552
rect 44720 35512 44729 35552
rect 48343 35512 48352 35552
rect 48392 35512 48434 35552
rect 48474 35512 48516 35552
rect 48556 35512 48598 35552
rect 48638 35512 48680 35552
rect 48720 35512 48729 35552
rect 52343 35512 52352 35552
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52720 35512 52729 35552
rect 56343 35512 56352 35552
rect 56392 35512 56434 35552
rect 56474 35512 56516 35552
rect 56556 35512 56598 35552
rect 56638 35512 56680 35552
rect 56720 35512 56729 35552
rect 60343 35512 60352 35552
rect 60392 35512 60434 35552
rect 60474 35512 60516 35552
rect 60556 35512 60598 35552
rect 60638 35512 60680 35552
rect 60720 35512 60729 35552
rect 64343 35512 64352 35552
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64720 35512 64729 35552
rect 68343 35512 68352 35552
rect 68392 35512 68434 35552
rect 68474 35512 68516 35552
rect 68556 35512 68598 35552
rect 68638 35512 68680 35552
rect 68720 35512 68729 35552
rect 72343 35512 72352 35552
rect 72392 35512 72434 35552
rect 72474 35512 72516 35552
rect 72556 35512 72598 35552
rect 72638 35512 72680 35552
rect 72720 35512 72729 35552
rect 76343 35512 76352 35552
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76720 35512 76729 35552
rect 80343 35512 80352 35552
rect 80392 35512 80434 35552
rect 80474 35512 80516 35552
rect 80556 35512 80598 35552
rect 80638 35512 80680 35552
rect 80720 35512 80729 35552
rect 84343 35512 84352 35552
rect 84392 35512 84434 35552
rect 84474 35512 84516 35552
rect 84556 35512 84598 35552
rect 84638 35512 84680 35552
rect 84720 35512 84729 35552
rect 88343 35512 88352 35552
rect 88392 35512 88434 35552
rect 88474 35512 88516 35552
rect 88556 35512 88598 35552
rect 88638 35512 88680 35552
rect 88720 35512 88729 35552
rect 92343 35512 92352 35552
rect 92392 35512 92434 35552
rect 92474 35512 92516 35552
rect 92556 35512 92598 35552
rect 92638 35512 92680 35552
rect 92720 35512 92729 35552
rect 96343 35512 96352 35552
rect 96392 35512 96434 35552
rect 96474 35512 96516 35552
rect 96556 35512 96598 35552
rect 96638 35512 96680 35552
rect 96720 35512 96729 35552
rect 0 34988 80 35068
rect 3103 34756 3112 34796
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3480 34756 3489 34796
rect 7103 34756 7112 34796
rect 7152 34756 7194 34796
rect 7234 34756 7276 34796
rect 7316 34756 7358 34796
rect 7398 34756 7440 34796
rect 7480 34756 7489 34796
rect 11103 34756 11112 34796
rect 11152 34756 11194 34796
rect 11234 34756 11276 34796
rect 11316 34756 11358 34796
rect 11398 34756 11440 34796
rect 11480 34756 11489 34796
rect 15103 34756 15112 34796
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15480 34756 15489 34796
rect 19103 34756 19112 34796
rect 19152 34756 19194 34796
rect 19234 34756 19276 34796
rect 19316 34756 19358 34796
rect 19398 34756 19440 34796
rect 19480 34756 19489 34796
rect 23103 34756 23112 34796
rect 23152 34756 23194 34796
rect 23234 34756 23276 34796
rect 23316 34756 23358 34796
rect 23398 34756 23440 34796
rect 23480 34756 23489 34796
rect 27103 34756 27112 34796
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27480 34756 27489 34796
rect 31103 34756 31112 34796
rect 31152 34756 31194 34796
rect 31234 34756 31276 34796
rect 31316 34756 31358 34796
rect 31398 34756 31440 34796
rect 31480 34756 31489 34796
rect 35103 34756 35112 34796
rect 35152 34756 35194 34796
rect 35234 34756 35276 34796
rect 35316 34756 35358 34796
rect 35398 34756 35440 34796
rect 35480 34756 35489 34796
rect 39103 34756 39112 34796
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39480 34756 39489 34796
rect 43103 34756 43112 34796
rect 43152 34756 43194 34796
rect 43234 34756 43276 34796
rect 43316 34756 43358 34796
rect 43398 34756 43440 34796
rect 43480 34756 43489 34796
rect 47103 34756 47112 34796
rect 47152 34756 47194 34796
rect 47234 34756 47276 34796
rect 47316 34756 47358 34796
rect 47398 34756 47440 34796
rect 47480 34756 47489 34796
rect 51103 34756 51112 34796
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51480 34756 51489 34796
rect 55103 34756 55112 34796
rect 55152 34756 55194 34796
rect 55234 34756 55276 34796
rect 55316 34756 55358 34796
rect 55398 34756 55440 34796
rect 55480 34756 55489 34796
rect 59103 34756 59112 34796
rect 59152 34756 59194 34796
rect 59234 34756 59276 34796
rect 59316 34756 59358 34796
rect 59398 34756 59440 34796
rect 59480 34756 59489 34796
rect 63103 34756 63112 34796
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63480 34756 63489 34796
rect 67103 34756 67112 34796
rect 67152 34756 67194 34796
rect 67234 34756 67276 34796
rect 67316 34756 67358 34796
rect 67398 34756 67440 34796
rect 67480 34756 67489 34796
rect 71103 34756 71112 34796
rect 71152 34756 71194 34796
rect 71234 34756 71276 34796
rect 71316 34756 71358 34796
rect 71398 34756 71440 34796
rect 71480 34756 71489 34796
rect 75103 34756 75112 34796
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75480 34756 75489 34796
rect 79103 34756 79112 34796
rect 79152 34756 79194 34796
rect 79234 34756 79276 34796
rect 79316 34756 79358 34796
rect 79398 34756 79440 34796
rect 79480 34756 79489 34796
rect 83103 34756 83112 34796
rect 83152 34756 83194 34796
rect 83234 34756 83276 34796
rect 83316 34756 83358 34796
rect 83398 34756 83440 34796
rect 83480 34756 83489 34796
rect 87103 34756 87112 34796
rect 87152 34756 87194 34796
rect 87234 34756 87276 34796
rect 87316 34756 87358 34796
rect 87398 34756 87440 34796
rect 87480 34756 87489 34796
rect 91103 34756 91112 34796
rect 91152 34756 91194 34796
rect 91234 34756 91276 34796
rect 91316 34756 91358 34796
rect 91398 34756 91440 34796
rect 91480 34756 91489 34796
rect 95103 34756 95112 34796
rect 95152 34756 95194 34796
rect 95234 34756 95276 34796
rect 95316 34756 95358 34796
rect 95398 34756 95440 34796
rect 95480 34756 95489 34796
rect 99103 34756 99112 34796
rect 99152 34756 99194 34796
rect 99234 34756 99276 34796
rect 99316 34756 99358 34796
rect 99398 34756 99440 34796
rect 99480 34756 99489 34796
rect 0 34148 80 34228
rect 4343 34000 4352 34040
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4720 34000 4729 34040
rect 8343 34000 8352 34040
rect 8392 34000 8434 34040
rect 8474 34000 8516 34040
rect 8556 34000 8598 34040
rect 8638 34000 8680 34040
rect 8720 34000 8729 34040
rect 12343 34000 12352 34040
rect 12392 34000 12434 34040
rect 12474 34000 12516 34040
rect 12556 34000 12598 34040
rect 12638 34000 12680 34040
rect 12720 34000 12729 34040
rect 16343 34000 16352 34040
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16720 34000 16729 34040
rect 20343 34000 20352 34040
rect 20392 34000 20434 34040
rect 20474 34000 20516 34040
rect 20556 34000 20598 34040
rect 20638 34000 20680 34040
rect 20720 34000 20729 34040
rect 24343 34000 24352 34040
rect 24392 34000 24434 34040
rect 24474 34000 24516 34040
rect 24556 34000 24598 34040
rect 24638 34000 24680 34040
rect 24720 34000 24729 34040
rect 28343 34000 28352 34040
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28720 34000 28729 34040
rect 32343 34000 32352 34040
rect 32392 34000 32434 34040
rect 32474 34000 32516 34040
rect 32556 34000 32598 34040
rect 32638 34000 32680 34040
rect 32720 34000 32729 34040
rect 36343 34000 36352 34040
rect 36392 34000 36434 34040
rect 36474 34000 36516 34040
rect 36556 34000 36598 34040
rect 36638 34000 36680 34040
rect 36720 34000 36729 34040
rect 40343 34000 40352 34040
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40720 34000 40729 34040
rect 44343 34000 44352 34040
rect 44392 34000 44434 34040
rect 44474 34000 44516 34040
rect 44556 34000 44598 34040
rect 44638 34000 44680 34040
rect 44720 34000 44729 34040
rect 48343 34000 48352 34040
rect 48392 34000 48434 34040
rect 48474 34000 48516 34040
rect 48556 34000 48598 34040
rect 48638 34000 48680 34040
rect 48720 34000 48729 34040
rect 52343 34000 52352 34040
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52720 34000 52729 34040
rect 56343 34000 56352 34040
rect 56392 34000 56434 34040
rect 56474 34000 56516 34040
rect 56556 34000 56598 34040
rect 56638 34000 56680 34040
rect 56720 34000 56729 34040
rect 60343 34000 60352 34040
rect 60392 34000 60434 34040
rect 60474 34000 60516 34040
rect 60556 34000 60598 34040
rect 60638 34000 60680 34040
rect 60720 34000 60729 34040
rect 64343 34000 64352 34040
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64720 34000 64729 34040
rect 68343 34000 68352 34040
rect 68392 34000 68434 34040
rect 68474 34000 68516 34040
rect 68556 34000 68598 34040
rect 68638 34000 68680 34040
rect 68720 34000 68729 34040
rect 91267 33748 91276 33788
rect 91316 33748 91660 33788
rect 91700 33748 91709 33788
rect 95491 33748 95500 33788
rect 95540 33748 95549 33788
rect 95500 33704 95540 33748
rect 95299 33664 95308 33704
rect 95348 33664 96076 33704
rect 96116 33664 96460 33704
rect 96500 33664 96980 33704
rect 96940 33620 96980 33664
rect 74179 33580 74188 33620
rect 74228 33580 74476 33620
rect 74516 33580 74860 33620
rect 74900 33580 75340 33620
rect 75380 33580 75389 33620
rect 75811 33580 75820 33620
rect 75860 33580 76204 33620
rect 76244 33580 76253 33620
rect 77059 33580 77068 33620
rect 77108 33580 77452 33620
rect 77492 33580 77836 33620
rect 77876 33580 77885 33620
rect 78595 33580 78604 33620
rect 78644 33580 78988 33620
rect 79028 33580 79372 33620
rect 79412 33580 79756 33620
rect 79796 33580 79805 33620
rect 80323 33580 80332 33620
rect 80372 33580 81292 33620
rect 81332 33580 82444 33620
rect 82484 33580 83116 33620
rect 83156 33580 83165 33620
rect 85891 33580 85900 33620
rect 85940 33580 86284 33620
rect 86324 33580 86333 33620
rect 86659 33580 86668 33620
rect 86708 33580 87436 33620
rect 87476 33580 87820 33620
rect 87860 33580 87869 33620
rect 88579 33580 88588 33620
rect 88628 33580 88972 33620
rect 89012 33580 89356 33620
rect 89396 33580 89405 33620
rect 89539 33580 89548 33620
rect 89588 33580 90124 33620
rect 90164 33580 90508 33620
rect 90548 33580 90892 33620
rect 90932 33580 91180 33620
rect 91220 33580 91852 33620
rect 91892 33580 91901 33620
rect 93187 33580 93196 33620
rect 93236 33580 93388 33620
rect 93428 33580 93580 33620
rect 93620 33580 93629 33620
rect 94243 33580 94252 33620
rect 94292 33580 94636 33620
rect 94676 33580 94685 33620
rect 95683 33580 95692 33620
rect 95732 33580 96748 33620
rect 96788 33580 96797 33620
rect 96931 33580 96940 33620
rect 96980 33580 98380 33620
rect 98420 33580 98429 33620
rect 95692 33536 95732 33580
rect 80515 33496 80524 33536
rect 80564 33496 80908 33536
rect 80948 33496 81676 33536
rect 81716 33496 82060 33536
rect 82100 33496 82109 33536
rect 82243 33496 82252 33536
rect 82292 33496 82828 33536
rect 82868 33496 83212 33536
rect 83252 33496 83500 33536
rect 83540 33496 83549 33536
rect 92515 33496 92524 33536
rect 92564 33496 92812 33536
rect 92852 33496 93772 33536
rect 93812 33496 95732 33536
rect 87043 33452 87101 33453
rect 97228 33452 97268 33580
rect 86958 33412 87052 33452
rect 87092 33412 92620 33452
rect 92660 33412 92669 33452
rect 97219 33412 97228 33452
rect 97268 33412 97277 33452
rect 87043 33411 87101 33412
rect 0 33308 80 33388
rect 3103 33244 3112 33284
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3480 33244 3489 33284
rect 7103 33244 7112 33284
rect 7152 33244 7194 33284
rect 7234 33244 7276 33284
rect 7316 33244 7358 33284
rect 7398 33244 7440 33284
rect 7480 33244 7489 33284
rect 11103 33244 11112 33284
rect 11152 33244 11194 33284
rect 11234 33244 11276 33284
rect 11316 33244 11358 33284
rect 11398 33244 11440 33284
rect 11480 33244 11489 33284
rect 15103 33244 15112 33284
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15480 33244 15489 33284
rect 19103 33244 19112 33284
rect 19152 33244 19194 33284
rect 19234 33244 19276 33284
rect 19316 33244 19358 33284
rect 19398 33244 19440 33284
rect 19480 33244 19489 33284
rect 23103 33244 23112 33284
rect 23152 33244 23194 33284
rect 23234 33244 23276 33284
rect 23316 33244 23358 33284
rect 23398 33244 23440 33284
rect 23480 33244 23489 33284
rect 27103 33244 27112 33284
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27480 33244 27489 33284
rect 31103 33244 31112 33284
rect 31152 33244 31194 33284
rect 31234 33244 31276 33284
rect 31316 33244 31358 33284
rect 31398 33244 31440 33284
rect 31480 33244 31489 33284
rect 35103 33244 35112 33284
rect 35152 33244 35194 33284
rect 35234 33244 35276 33284
rect 35316 33244 35358 33284
rect 35398 33244 35440 33284
rect 35480 33244 35489 33284
rect 39103 33244 39112 33284
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39480 33244 39489 33284
rect 43103 33244 43112 33284
rect 43152 33244 43194 33284
rect 43234 33244 43276 33284
rect 43316 33244 43358 33284
rect 43398 33244 43440 33284
rect 43480 33244 43489 33284
rect 47103 33244 47112 33284
rect 47152 33244 47194 33284
rect 47234 33244 47276 33284
rect 47316 33244 47358 33284
rect 47398 33244 47440 33284
rect 47480 33244 47489 33284
rect 51103 33244 51112 33284
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51480 33244 51489 33284
rect 55103 33244 55112 33284
rect 55152 33244 55194 33284
rect 55234 33244 55276 33284
rect 55316 33244 55358 33284
rect 55398 33244 55440 33284
rect 55480 33244 55489 33284
rect 59103 33244 59112 33284
rect 59152 33244 59194 33284
rect 59234 33244 59276 33284
rect 59316 33244 59358 33284
rect 59398 33244 59440 33284
rect 59480 33244 59489 33284
rect 63103 33244 63112 33284
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63480 33244 63489 33284
rect 67103 33244 67112 33284
rect 67152 33244 67194 33284
rect 67234 33244 67276 33284
rect 67316 33244 67358 33284
rect 67398 33244 67440 33284
rect 67480 33244 67489 33284
rect 71779 33244 71788 33284
rect 71828 33244 74668 33284
rect 74708 33244 81100 33284
rect 81140 33244 81149 33284
rect 86275 33244 86284 33284
rect 86324 33244 86860 33284
rect 86900 33244 87916 33284
rect 87956 33244 88436 33284
rect 88963 33244 88972 33284
rect 89012 33244 89548 33284
rect 89588 33244 90316 33284
rect 90356 33244 90365 33284
rect 88396 33200 88436 33244
rect 75427 33160 75436 33200
rect 75476 33160 76300 33200
rect 76340 33160 76349 33200
rect 83107 33160 83116 33200
rect 83156 33160 84652 33200
rect 84692 33160 84701 33200
rect 86467 33160 86476 33200
rect 86516 33160 87052 33200
rect 87092 33160 87340 33200
rect 87380 33160 87628 33200
rect 87668 33160 88300 33200
rect 88340 33160 88349 33200
rect 88396 33160 89740 33200
rect 89780 33160 90700 33200
rect 90740 33160 90749 33200
rect 92323 33160 92332 33200
rect 92372 33160 93388 33200
rect 93428 33160 93676 33200
rect 93716 33160 94348 33200
rect 94388 33160 94828 33200
rect 94868 33160 94877 33200
rect 76195 33076 76204 33116
rect 76244 33076 76284 33116
rect 83587 33076 83596 33116
rect 83636 33076 83676 33116
rect 85123 33076 85132 33116
rect 85172 33076 85181 33116
rect 86851 33076 86860 33116
rect 86900 33076 87244 33116
rect 87284 33076 87293 33116
rect 88003 33076 88012 33116
rect 88052 33076 88396 33116
rect 88436 33076 88445 33116
rect 90883 33076 90892 33116
rect 90932 33076 91756 33116
rect 91796 33076 92812 33116
rect 92852 33076 93004 33116
rect 93044 33076 93053 33116
rect 94627 33076 94636 33116
rect 94676 33076 95212 33116
rect 95252 33076 95500 33116
rect 95540 33076 95692 33116
rect 95732 33076 95741 33116
rect 76204 33032 76244 33076
rect 83596 33032 83636 33076
rect 76003 32992 76012 33032
rect 76052 32992 76588 33032
rect 76628 32992 76637 33032
rect 76867 32992 76876 33032
rect 76916 32992 77452 33032
rect 77492 32992 77501 33032
rect 77827 32992 77836 33032
rect 77876 32992 78124 33032
rect 78164 32992 78412 33032
rect 78452 32992 79084 33032
rect 79124 32992 79133 33032
rect 83299 32992 83308 33032
rect 83348 32992 83884 33032
rect 83924 32992 84172 33032
rect 84212 32992 84460 33032
rect 84500 32992 84748 33032
rect 84788 32992 85036 33032
rect 85076 32992 85085 33032
rect 85132 32948 85172 33076
rect 85872 32992 85900 33032
rect 85940 32992 86668 33032
rect 86708 32992 86717 33032
rect 88099 32992 88108 33032
rect 88148 32992 88684 33032
rect 88724 32992 89452 33032
rect 89492 32992 89740 33032
rect 89780 32992 89932 33032
rect 89972 32992 89981 33032
rect 91171 32992 91180 33032
rect 91220 32992 91468 33032
rect 91508 32992 91517 33032
rect 91756 32992 92716 33032
rect 92756 32992 92765 33032
rect 93763 32992 93772 33032
rect 93812 32992 94924 33032
rect 94964 32992 94973 33032
rect 70723 32908 70732 32948
rect 70772 32908 72364 32948
rect 72404 32908 72652 32948
rect 72692 32908 73036 32948
rect 73076 32908 73228 32948
rect 73268 32908 73277 32948
rect 74371 32908 74380 32948
rect 74420 32908 74860 32948
rect 74900 32908 75148 32948
rect 75188 32908 75820 32948
rect 75860 32908 77260 32948
rect 77300 32908 78700 32948
rect 78740 32908 78749 32948
rect 78796 32908 79372 32948
rect 79412 32908 79421 32948
rect 79747 32908 79756 32948
rect 79796 32908 80044 32948
rect 80084 32908 80236 32948
rect 80276 32908 80285 32948
rect 80611 32908 80620 32948
rect 80660 32908 81100 32948
rect 81140 32908 81388 32948
rect 81428 32908 82252 32948
rect 82292 32908 82301 32948
rect 82636 32908 83596 32948
rect 83636 32908 83645 32948
rect 84835 32908 84844 32948
rect 84884 32908 85460 32948
rect 73603 32864 73661 32865
rect 78796 32864 78836 32908
rect 71587 32824 71596 32864
rect 71636 32824 72268 32864
rect 72308 32824 72317 32864
rect 73518 32824 73612 32864
rect 73652 32824 73661 32864
rect 73987 32824 73996 32864
rect 74036 32824 74188 32864
rect 74228 32824 74237 32864
rect 75436 32824 76204 32864
rect 76244 32824 76253 32864
rect 76579 32824 76588 32864
rect 76628 32824 76876 32864
rect 76916 32824 76925 32864
rect 76972 32824 77548 32864
rect 77588 32824 77597 32864
rect 77836 32824 78316 32864
rect 78356 32824 78365 32864
rect 78700 32824 78836 32864
rect 78979 32824 78988 32864
rect 79028 32824 79660 32864
rect 79700 32824 79709 32864
rect 80236 32824 81004 32864
rect 81044 32824 81053 32864
rect 81676 32824 82348 32864
rect 82388 32824 82397 32864
rect 73603 32823 73661 32824
rect 75436 32696 75476 32824
rect 76972 32780 77012 32824
rect 76932 32740 76972 32780
rect 77012 32740 77021 32780
rect 77836 32696 77876 32824
rect 78700 32780 78740 32824
rect 78660 32740 78700 32780
rect 78740 32740 78749 32780
rect 80236 32696 80276 32824
rect 81676 32780 81716 32824
rect 81475 32740 81484 32780
rect 81524 32740 81716 32780
rect 82636 32696 82676 32908
rect 85420 32864 85460 32908
rect 85996 32864 86036 32992
rect 86380 32908 86956 32948
rect 86996 32908 87005 32948
rect 87628 32908 88396 32948
rect 88436 32908 88445 32948
rect 89059 32908 89068 32948
rect 89108 32908 90028 32948
rect 90068 32908 90077 32948
rect 90124 32908 91084 32948
rect 91124 32908 91133 32948
rect 86380 32864 86420 32908
rect 83116 32824 83788 32864
rect 83828 32824 83837 32864
rect 84172 32824 85132 32864
rect 85172 32824 85181 32864
rect 85411 32824 85420 32864
rect 85460 32824 85708 32864
rect 85748 32824 85996 32864
rect 86036 32824 86045 32864
rect 86284 32824 86420 32864
rect 86668 32824 87244 32864
rect 87284 32824 87293 32864
rect 83116 32780 83156 32824
rect 84172 32780 84212 32824
rect 86284 32780 86324 32824
rect 83076 32740 83116 32780
rect 83156 32740 83165 32780
rect 84172 32740 84268 32780
rect 84308 32740 84317 32780
rect 85660 32740 85900 32780
rect 85940 32740 85949 32780
rect 86244 32740 86284 32780
rect 86324 32740 86333 32780
rect 85660 32696 85700 32740
rect 86668 32696 86708 32824
rect 87628 32696 87668 32908
rect 90124 32864 90164 32908
rect 87916 32824 88588 32864
rect 88628 32824 88637 32864
rect 88771 32824 88780 32864
rect 88820 32824 89644 32864
rect 89684 32824 89693 32864
rect 89932 32824 90164 32864
rect 90403 32824 90412 32864
rect 90452 32824 91372 32864
rect 91412 32824 91421 32864
rect 87916 32780 87956 32824
rect 87876 32740 87916 32780
rect 87956 32740 87965 32780
rect 89932 32696 89972 32824
rect 73891 32656 73900 32696
rect 73940 32656 74188 32696
rect 74228 32656 74237 32696
rect 74659 32656 74668 32696
rect 74708 32656 75052 32696
rect 75092 32656 75101 32696
rect 75427 32656 75436 32696
rect 75476 32656 75485 32696
rect 76291 32656 76300 32696
rect 76340 32656 76780 32696
rect 76820 32656 76829 32696
rect 77827 32656 77836 32696
rect 77876 32656 77885 32696
rect 79459 32656 79468 32696
rect 79508 32656 79948 32696
rect 79988 32656 79997 32696
rect 80227 32656 80236 32696
rect 80276 32656 80285 32696
rect 82627 32656 82636 32696
rect 82676 32656 82685 32696
rect 83875 32656 83884 32696
rect 83924 32656 84364 32696
rect 84404 32656 84413 32696
rect 85411 32656 85420 32696
rect 85460 32656 85700 32696
rect 86659 32656 86668 32696
rect 86708 32656 86717 32696
rect 87619 32656 87628 32696
rect 87668 32656 87677 32696
rect 89923 32656 89932 32696
rect 89972 32656 89981 32696
rect 90787 32656 90796 32696
rect 90836 32656 91660 32696
rect 91700 32656 91709 32696
rect 91756 32612 91796 32992
rect 91843 32908 91852 32948
rect 91892 32908 93100 32948
rect 93140 32908 93149 32948
rect 94147 32908 94156 32948
rect 94196 32908 95116 32948
rect 95156 32908 95165 32948
rect 92323 32824 92332 32864
rect 92372 32824 93292 32864
rect 93332 32824 93341 32864
rect 93772 32824 94252 32864
rect 94292 32824 94301 32864
rect 95011 32824 95020 32864
rect 95060 32824 95788 32864
rect 95828 32824 95837 32864
rect 96067 32824 96076 32864
rect 96116 32824 96364 32864
rect 96404 32824 96413 32864
rect 96931 32824 96940 32864
rect 96980 32824 97132 32864
rect 97172 32824 97516 32864
rect 97556 32824 97804 32864
rect 97844 32824 98092 32864
rect 98132 32824 99148 32864
rect 99188 32824 99197 32864
rect 93772 32780 93812 32824
rect 92611 32740 92620 32780
rect 92660 32740 93580 32780
rect 93620 32740 93629 32780
rect 93676 32740 93812 32780
rect 93859 32740 93868 32780
rect 93908 32740 94540 32780
rect 94580 32740 94589 32780
rect 95500 32740 95980 32780
rect 96020 32740 96029 32780
rect 93676 32696 93716 32740
rect 95500 32696 95540 32740
rect 92995 32656 93004 32696
rect 93044 32656 93716 32696
rect 95491 32656 95500 32696
rect 95540 32656 95549 32696
rect 97507 32656 97516 32696
rect 97556 32656 97996 32696
rect 98036 32656 98045 32696
rect 91459 32572 91468 32612
rect 91508 32572 91796 32612
rect 0 32468 80 32548
rect 4343 32488 4352 32528
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4720 32488 4729 32528
rect 8343 32488 8352 32528
rect 8392 32488 8434 32528
rect 8474 32488 8516 32528
rect 8556 32488 8598 32528
rect 8638 32488 8680 32528
rect 8720 32488 8729 32528
rect 12343 32488 12352 32528
rect 12392 32488 12434 32528
rect 12474 32488 12516 32528
rect 12556 32488 12598 32528
rect 12638 32488 12680 32528
rect 12720 32488 12729 32528
rect 16343 32488 16352 32528
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16720 32488 16729 32528
rect 20343 32488 20352 32528
rect 20392 32488 20434 32528
rect 20474 32488 20516 32528
rect 20556 32488 20598 32528
rect 20638 32488 20680 32528
rect 20720 32488 20729 32528
rect 24343 32488 24352 32528
rect 24392 32488 24434 32528
rect 24474 32488 24516 32528
rect 24556 32488 24598 32528
rect 24638 32488 24680 32528
rect 24720 32488 24729 32528
rect 28343 32488 28352 32528
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28720 32488 28729 32528
rect 32343 32488 32352 32528
rect 32392 32488 32434 32528
rect 32474 32488 32516 32528
rect 32556 32488 32598 32528
rect 32638 32488 32680 32528
rect 32720 32488 32729 32528
rect 36343 32488 36352 32528
rect 36392 32488 36434 32528
rect 36474 32488 36516 32528
rect 36556 32488 36598 32528
rect 36638 32488 36680 32528
rect 36720 32488 36729 32528
rect 40343 32488 40352 32528
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40720 32488 40729 32528
rect 44343 32488 44352 32528
rect 44392 32488 44434 32528
rect 44474 32488 44516 32528
rect 44556 32488 44598 32528
rect 44638 32488 44680 32528
rect 44720 32488 44729 32528
rect 48343 32488 48352 32528
rect 48392 32488 48434 32528
rect 48474 32488 48516 32528
rect 48556 32488 48598 32528
rect 48638 32488 48680 32528
rect 48720 32488 48729 32528
rect 52343 32488 52352 32528
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52720 32488 52729 32528
rect 56343 32488 56352 32528
rect 56392 32488 56434 32528
rect 56474 32488 56516 32528
rect 56556 32488 56598 32528
rect 56638 32488 56680 32528
rect 56720 32488 56729 32528
rect 60343 32488 60352 32528
rect 60392 32488 60434 32528
rect 60474 32488 60516 32528
rect 60556 32488 60598 32528
rect 60638 32488 60680 32528
rect 60720 32488 60729 32528
rect 64343 32488 64352 32528
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64720 32488 64729 32528
rect 68343 32488 68352 32528
rect 68392 32488 68434 32528
rect 68474 32488 68516 32528
rect 68556 32488 68598 32528
rect 68638 32488 68680 32528
rect 68720 32488 68729 32528
rect 72451 32488 72460 32528
rect 72500 32488 73132 32528
rect 73172 32488 73181 32528
rect 78019 32404 78028 32444
rect 78068 32404 78077 32444
rect 78028 32360 78068 32404
rect 71395 32320 71404 32360
rect 71444 32320 72415 32360
rect 72455 32320 72464 32360
rect 72835 32320 72844 32360
rect 72884 32320 73215 32360
rect 73255 32320 73264 32360
rect 77496 32320 77505 32360
rect 77545 32320 78068 32360
rect 79747 32320 79756 32360
rect 79796 32320 80332 32360
rect 80372 32320 80381 32360
rect 80696 32320 80705 32360
rect 80745 32320 81292 32360
rect 81332 32320 81341 32360
rect 82296 32320 82305 32360
rect 82345 32320 82828 32360
rect 82868 32320 82877 32360
rect 83496 32320 83505 32360
rect 83545 32320 84076 32360
rect 84116 32320 84125 32360
rect 85096 32320 85105 32360
rect 85145 32320 85612 32360
rect 85652 32320 85661 32360
rect 85896 32320 85905 32360
rect 85945 32320 86764 32360
rect 86804 32320 86813 32360
rect 87096 32320 87105 32360
rect 87145 32320 87532 32360
rect 87572 32320 87581 32360
rect 75896 32236 75905 32276
rect 75945 32236 76492 32276
rect 76532 32236 76541 32276
rect 78296 32236 78305 32276
rect 78345 32236 79180 32276
rect 79220 32236 79229 32276
rect 81096 32236 81105 32276
rect 81145 32236 81580 32276
rect 81620 32236 81629 32276
rect 91096 32236 91105 32276
rect 91145 32236 91852 32276
rect 91892 32236 91901 32276
rect 95896 32236 95905 32276
rect 95945 32236 96268 32276
rect 96308 32236 96317 32276
rect 96364 32236 97132 32276
rect 97172 32236 97181 32276
rect 70819 32152 70828 32192
rect 70868 32152 72815 32192
rect 72855 32152 72864 32192
rect 77059 32152 77068 32192
rect 77108 32152 77740 32192
rect 77780 32152 77789 32192
rect 96364 32108 96404 32236
rect 96696 32152 96705 32192
rect 96745 32152 97420 32192
rect 97460 32152 97469 32192
rect 98296 32152 98305 32192
rect 98345 32152 98956 32192
rect 98996 32152 99005 32192
rect 70531 32068 70540 32108
rect 70580 32068 70924 32108
rect 70964 32068 70973 32108
rect 71107 32068 71116 32108
rect 71156 32068 72705 32108
rect 72745 32068 72754 32108
rect 75096 32068 75105 32108
rect 75145 32068 75340 32108
rect 75380 32068 75389 32108
rect 76696 32068 76705 32108
rect 76745 32068 76972 32108
rect 77012 32068 77021 32108
rect 81896 32068 81905 32108
rect 81945 32068 82540 32108
rect 82580 32068 82589 32108
rect 84696 32068 84705 32108
rect 84745 32068 85324 32108
rect 85364 32068 85373 32108
rect 88296 32068 88305 32108
rect 88345 32068 89356 32108
rect 89396 32068 89405 32108
rect 89496 32068 89505 32108
rect 89545 32068 90220 32108
rect 90260 32068 90269 32108
rect 93496 32068 93505 32108
rect 93545 32068 93772 32108
rect 93812 32068 93821 32108
rect 94696 32068 94705 32108
rect 94745 32068 95404 32108
rect 95444 32068 95453 32108
rect 96296 32068 96305 32108
rect 96345 32068 96404 32108
rect 97096 32068 97105 32108
rect 97145 32068 97708 32108
rect 97748 32068 97757 32108
rect 97896 32068 97905 32108
rect 97945 32068 99244 32108
rect 99284 32068 99293 32108
rect 3103 31732 3112 31772
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3480 31732 3489 31772
rect 7103 31732 7112 31772
rect 7152 31732 7194 31772
rect 7234 31732 7276 31772
rect 7316 31732 7358 31772
rect 7398 31732 7440 31772
rect 7480 31732 7489 31772
rect 11103 31732 11112 31772
rect 11152 31732 11194 31772
rect 11234 31732 11276 31772
rect 11316 31732 11358 31772
rect 11398 31732 11440 31772
rect 11480 31732 11489 31772
rect 15103 31732 15112 31772
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15480 31732 15489 31772
rect 19103 31732 19112 31772
rect 19152 31732 19194 31772
rect 19234 31732 19276 31772
rect 19316 31732 19358 31772
rect 19398 31732 19440 31772
rect 19480 31732 19489 31772
rect 23103 31732 23112 31772
rect 23152 31732 23194 31772
rect 23234 31732 23276 31772
rect 23316 31732 23358 31772
rect 23398 31732 23440 31772
rect 23480 31732 23489 31772
rect 27103 31732 27112 31772
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27480 31732 27489 31772
rect 31103 31732 31112 31772
rect 31152 31732 31194 31772
rect 31234 31732 31276 31772
rect 31316 31732 31358 31772
rect 31398 31732 31440 31772
rect 31480 31732 31489 31772
rect 35103 31732 35112 31772
rect 35152 31732 35194 31772
rect 35234 31732 35276 31772
rect 35316 31732 35358 31772
rect 35398 31732 35440 31772
rect 35480 31732 35489 31772
rect 39103 31732 39112 31772
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39480 31732 39489 31772
rect 43103 31732 43112 31772
rect 43152 31732 43194 31772
rect 43234 31732 43276 31772
rect 43316 31732 43358 31772
rect 43398 31732 43440 31772
rect 43480 31732 43489 31772
rect 47103 31732 47112 31772
rect 47152 31732 47194 31772
rect 47234 31732 47276 31772
rect 47316 31732 47358 31772
rect 47398 31732 47440 31772
rect 47480 31732 47489 31772
rect 51103 31732 51112 31772
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51480 31732 51489 31772
rect 55103 31732 55112 31772
rect 55152 31732 55194 31772
rect 55234 31732 55276 31772
rect 55316 31732 55358 31772
rect 55398 31732 55440 31772
rect 55480 31732 55489 31772
rect 59103 31732 59112 31772
rect 59152 31732 59194 31772
rect 59234 31732 59276 31772
rect 59316 31732 59358 31772
rect 59398 31732 59440 31772
rect 59480 31732 59489 31772
rect 63103 31732 63112 31772
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63480 31732 63489 31772
rect 67103 31732 67112 31772
rect 67152 31732 67194 31772
rect 67234 31732 67276 31772
rect 67316 31732 67358 31772
rect 67398 31732 67440 31772
rect 67480 31732 67489 31772
rect 0 31628 80 31708
rect 4343 30976 4352 31016
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4720 30976 4729 31016
rect 8343 30976 8352 31016
rect 8392 30976 8434 31016
rect 8474 30976 8516 31016
rect 8556 30976 8598 31016
rect 8638 30976 8680 31016
rect 8720 30976 8729 31016
rect 12343 30976 12352 31016
rect 12392 30976 12434 31016
rect 12474 30976 12516 31016
rect 12556 30976 12598 31016
rect 12638 30976 12680 31016
rect 12720 30976 12729 31016
rect 16343 30976 16352 31016
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16720 30976 16729 31016
rect 20343 30976 20352 31016
rect 20392 30976 20434 31016
rect 20474 30976 20516 31016
rect 20556 30976 20598 31016
rect 20638 30976 20680 31016
rect 20720 30976 20729 31016
rect 24343 30976 24352 31016
rect 24392 30976 24434 31016
rect 24474 30976 24516 31016
rect 24556 30976 24598 31016
rect 24638 30976 24680 31016
rect 24720 30976 24729 31016
rect 28343 30976 28352 31016
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28720 30976 28729 31016
rect 32343 30976 32352 31016
rect 32392 30976 32434 31016
rect 32474 30976 32516 31016
rect 32556 30976 32598 31016
rect 32638 30976 32680 31016
rect 32720 30976 32729 31016
rect 36343 30976 36352 31016
rect 36392 30976 36434 31016
rect 36474 30976 36516 31016
rect 36556 30976 36598 31016
rect 36638 30976 36680 31016
rect 36720 30976 36729 31016
rect 40343 30976 40352 31016
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40720 30976 40729 31016
rect 44343 30976 44352 31016
rect 44392 30976 44434 31016
rect 44474 30976 44516 31016
rect 44556 30976 44598 31016
rect 44638 30976 44680 31016
rect 44720 30976 44729 31016
rect 48343 30976 48352 31016
rect 48392 30976 48434 31016
rect 48474 30976 48516 31016
rect 48556 30976 48598 31016
rect 48638 30976 48680 31016
rect 48720 30976 48729 31016
rect 52343 30976 52352 31016
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52720 30976 52729 31016
rect 56343 30976 56352 31016
rect 56392 30976 56434 31016
rect 56474 30976 56516 31016
rect 56556 30976 56598 31016
rect 56638 30976 56680 31016
rect 56720 30976 56729 31016
rect 60343 30976 60352 31016
rect 60392 30976 60434 31016
rect 60474 30976 60516 31016
rect 60556 30976 60598 31016
rect 60638 30976 60680 31016
rect 60720 30976 60729 31016
rect 64343 30976 64352 31016
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64720 30976 64729 31016
rect 68343 30976 68352 31016
rect 68392 30976 68434 31016
rect 68474 30976 68516 31016
rect 68556 30976 68598 31016
rect 68638 30976 68680 31016
rect 68720 30976 68729 31016
rect 0 30788 80 30868
rect 3103 30220 3112 30260
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3480 30220 3489 30260
rect 7103 30220 7112 30260
rect 7152 30220 7194 30260
rect 7234 30220 7276 30260
rect 7316 30220 7358 30260
rect 7398 30220 7440 30260
rect 7480 30220 7489 30260
rect 11103 30220 11112 30260
rect 11152 30220 11194 30260
rect 11234 30220 11276 30260
rect 11316 30220 11358 30260
rect 11398 30220 11440 30260
rect 11480 30220 11489 30260
rect 15103 30220 15112 30260
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15480 30220 15489 30260
rect 19103 30220 19112 30260
rect 19152 30220 19194 30260
rect 19234 30220 19276 30260
rect 19316 30220 19358 30260
rect 19398 30220 19440 30260
rect 19480 30220 19489 30260
rect 23103 30220 23112 30260
rect 23152 30220 23194 30260
rect 23234 30220 23276 30260
rect 23316 30220 23358 30260
rect 23398 30220 23440 30260
rect 23480 30220 23489 30260
rect 27103 30220 27112 30260
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27480 30220 27489 30260
rect 31103 30220 31112 30260
rect 31152 30220 31194 30260
rect 31234 30220 31276 30260
rect 31316 30220 31358 30260
rect 31398 30220 31440 30260
rect 31480 30220 31489 30260
rect 35103 30220 35112 30260
rect 35152 30220 35194 30260
rect 35234 30220 35276 30260
rect 35316 30220 35358 30260
rect 35398 30220 35440 30260
rect 35480 30220 35489 30260
rect 39103 30220 39112 30260
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39480 30220 39489 30260
rect 43103 30220 43112 30260
rect 43152 30220 43194 30260
rect 43234 30220 43276 30260
rect 43316 30220 43358 30260
rect 43398 30220 43440 30260
rect 43480 30220 43489 30260
rect 47103 30220 47112 30260
rect 47152 30220 47194 30260
rect 47234 30220 47276 30260
rect 47316 30220 47358 30260
rect 47398 30220 47440 30260
rect 47480 30220 47489 30260
rect 51103 30220 51112 30260
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51480 30220 51489 30260
rect 55103 30220 55112 30260
rect 55152 30220 55194 30260
rect 55234 30220 55276 30260
rect 55316 30220 55358 30260
rect 55398 30220 55440 30260
rect 55480 30220 55489 30260
rect 59103 30220 59112 30260
rect 59152 30220 59194 30260
rect 59234 30220 59276 30260
rect 59316 30220 59358 30260
rect 59398 30220 59440 30260
rect 59480 30220 59489 30260
rect 63103 30220 63112 30260
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63480 30220 63489 30260
rect 67103 30220 67112 30260
rect 67152 30220 67194 30260
rect 67234 30220 67276 30260
rect 67316 30220 67358 30260
rect 67398 30220 67440 30260
rect 67480 30220 67489 30260
rect 0 29948 80 30028
rect 4343 29464 4352 29504
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4720 29464 4729 29504
rect 8343 29464 8352 29504
rect 8392 29464 8434 29504
rect 8474 29464 8516 29504
rect 8556 29464 8598 29504
rect 8638 29464 8680 29504
rect 8720 29464 8729 29504
rect 12343 29464 12352 29504
rect 12392 29464 12434 29504
rect 12474 29464 12516 29504
rect 12556 29464 12598 29504
rect 12638 29464 12680 29504
rect 12720 29464 12729 29504
rect 16343 29464 16352 29504
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16720 29464 16729 29504
rect 20343 29464 20352 29504
rect 20392 29464 20434 29504
rect 20474 29464 20516 29504
rect 20556 29464 20598 29504
rect 20638 29464 20680 29504
rect 20720 29464 20729 29504
rect 24343 29464 24352 29504
rect 24392 29464 24434 29504
rect 24474 29464 24516 29504
rect 24556 29464 24598 29504
rect 24638 29464 24680 29504
rect 24720 29464 24729 29504
rect 28343 29464 28352 29504
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28720 29464 28729 29504
rect 32343 29464 32352 29504
rect 32392 29464 32434 29504
rect 32474 29464 32516 29504
rect 32556 29464 32598 29504
rect 32638 29464 32680 29504
rect 32720 29464 32729 29504
rect 36343 29464 36352 29504
rect 36392 29464 36434 29504
rect 36474 29464 36516 29504
rect 36556 29464 36598 29504
rect 36638 29464 36680 29504
rect 36720 29464 36729 29504
rect 40343 29464 40352 29504
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40720 29464 40729 29504
rect 44343 29464 44352 29504
rect 44392 29464 44434 29504
rect 44474 29464 44516 29504
rect 44556 29464 44598 29504
rect 44638 29464 44680 29504
rect 44720 29464 44729 29504
rect 48343 29464 48352 29504
rect 48392 29464 48434 29504
rect 48474 29464 48516 29504
rect 48556 29464 48598 29504
rect 48638 29464 48680 29504
rect 48720 29464 48729 29504
rect 52343 29464 52352 29504
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52720 29464 52729 29504
rect 56343 29464 56352 29504
rect 56392 29464 56434 29504
rect 56474 29464 56516 29504
rect 56556 29464 56598 29504
rect 56638 29464 56680 29504
rect 56720 29464 56729 29504
rect 60343 29464 60352 29504
rect 60392 29464 60434 29504
rect 60474 29464 60516 29504
rect 60556 29464 60598 29504
rect 60638 29464 60680 29504
rect 60720 29464 60729 29504
rect 64343 29464 64352 29504
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64720 29464 64729 29504
rect 68343 29464 68352 29504
rect 68392 29464 68434 29504
rect 68474 29464 68516 29504
rect 68556 29464 68598 29504
rect 68638 29464 68680 29504
rect 68720 29464 68729 29504
rect 0 29108 80 29188
rect 3103 28708 3112 28748
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3480 28708 3489 28748
rect 7103 28708 7112 28748
rect 7152 28708 7194 28748
rect 7234 28708 7276 28748
rect 7316 28708 7358 28748
rect 7398 28708 7440 28748
rect 7480 28708 7489 28748
rect 11103 28708 11112 28748
rect 11152 28708 11194 28748
rect 11234 28708 11276 28748
rect 11316 28708 11358 28748
rect 11398 28708 11440 28748
rect 11480 28708 11489 28748
rect 15103 28708 15112 28748
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15480 28708 15489 28748
rect 19103 28708 19112 28748
rect 19152 28708 19194 28748
rect 19234 28708 19276 28748
rect 19316 28708 19358 28748
rect 19398 28708 19440 28748
rect 19480 28708 19489 28748
rect 23103 28708 23112 28748
rect 23152 28708 23194 28748
rect 23234 28708 23276 28748
rect 23316 28708 23358 28748
rect 23398 28708 23440 28748
rect 23480 28708 23489 28748
rect 27103 28708 27112 28748
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27480 28708 27489 28748
rect 31103 28708 31112 28748
rect 31152 28708 31194 28748
rect 31234 28708 31276 28748
rect 31316 28708 31358 28748
rect 31398 28708 31440 28748
rect 31480 28708 31489 28748
rect 35103 28708 35112 28748
rect 35152 28708 35194 28748
rect 35234 28708 35276 28748
rect 35316 28708 35358 28748
rect 35398 28708 35440 28748
rect 35480 28708 35489 28748
rect 39103 28708 39112 28748
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39480 28708 39489 28748
rect 43103 28708 43112 28748
rect 43152 28708 43194 28748
rect 43234 28708 43276 28748
rect 43316 28708 43358 28748
rect 43398 28708 43440 28748
rect 43480 28708 43489 28748
rect 47103 28708 47112 28748
rect 47152 28708 47194 28748
rect 47234 28708 47276 28748
rect 47316 28708 47358 28748
rect 47398 28708 47440 28748
rect 47480 28708 47489 28748
rect 51103 28708 51112 28748
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51480 28708 51489 28748
rect 55103 28708 55112 28748
rect 55152 28708 55194 28748
rect 55234 28708 55276 28748
rect 55316 28708 55358 28748
rect 55398 28708 55440 28748
rect 55480 28708 55489 28748
rect 59103 28708 59112 28748
rect 59152 28708 59194 28748
rect 59234 28708 59276 28748
rect 59316 28708 59358 28748
rect 59398 28708 59440 28748
rect 59480 28708 59489 28748
rect 63103 28708 63112 28748
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63480 28708 63489 28748
rect 67103 28708 67112 28748
rect 67152 28708 67194 28748
rect 67234 28708 67276 28748
rect 67316 28708 67358 28748
rect 67398 28708 67440 28748
rect 67480 28708 67489 28748
rect 0 28268 80 28348
rect 4343 27952 4352 27992
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4720 27952 4729 27992
rect 8343 27952 8352 27992
rect 8392 27952 8434 27992
rect 8474 27952 8516 27992
rect 8556 27952 8598 27992
rect 8638 27952 8680 27992
rect 8720 27952 8729 27992
rect 12343 27952 12352 27992
rect 12392 27952 12434 27992
rect 12474 27952 12516 27992
rect 12556 27952 12598 27992
rect 12638 27952 12680 27992
rect 12720 27952 12729 27992
rect 16343 27952 16352 27992
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16720 27952 16729 27992
rect 20343 27952 20352 27992
rect 20392 27952 20434 27992
rect 20474 27952 20516 27992
rect 20556 27952 20598 27992
rect 20638 27952 20680 27992
rect 20720 27952 20729 27992
rect 24343 27952 24352 27992
rect 24392 27952 24434 27992
rect 24474 27952 24516 27992
rect 24556 27952 24598 27992
rect 24638 27952 24680 27992
rect 24720 27952 24729 27992
rect 28343 27952 28352 27992
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28720 27952 28729 27992
rect 32343 27952 32352 27992
rect 32392 27952 32434 27992
rect 32474 27952 32516 27992
rect 32556 27952 32598 27992
rect 32638 27952 32680 27992
rect 32720 27952 32729 27992
rect 36343 27952 36352 27992
rect 36392 27952 36434 27992
rect 36474 27952 36516 27992
rect 36556 27952 36598 27992
rect 36638 27952 36680 27992
rect 36720 27952 36729 27992
rect 40343 27952 40352 27992
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40720 27952 40729 27992
rect 44343 27952 44352 27992
rect 44392 27952 44434 27992
rect 44474 27952 44516 27992
rect 44556 27952 44598 27992
rect 44638 27952 44680 27992
rect 44720 27952 44729 27992
rect 48343 27952 48352 27992
rect 48392 27952 48434 27992
rect 48474 27952 48516 27992
rect 48556 27952 48598 27992
rect 48638 27952 48680 27992
rect 48720 27952 48729 27992
rect 52343 27952 52352 27992
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52720 27952 52729 27992
rect 56343 27952 56352 27992
rect 56392 27952 56434 27992
rect 56474 27952 56516 27992
rect 56556 27952 56598 27992
rect 56638 27952 56680 27992
rect 56720 27952 56729 27992
rect 60343 27952 60352 27992
rect 60392 27952 60434 27992
rect 60474 27952 60516 27992
rect 60556 27952 60598 27992
rect 60638 27952 60680 27992
rect 60720 27952 60729 27992
rect 64343 27952 64352 27992
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64720 27952 64729 27992
rect 68343 27952 68352 27992
rect 68392 27952 68434 27992
rect 68474 27952 68516 27992
rect 68556 27952 68598 27992
rect 68638 27952 68680 27992
rect 68720 27952 68729 27992
rect 69955 27616 69964 27656
rect 70004 27616 70924 27656
rect 70964 27616 70973 27656
rect 0 27428 80 27508
rect 3103 27196 3112 27236
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3480 27196 3489 27236
rect 7103 27196 7112 27236
rect 7152 27196 7194 27236
rect 7234 27196 7276 27236
rect 7316 27196 7358 27236
rect 7398 27196 7440 27236
rect 7480 27196 7489 27236
rect 11103 27196 11112 27236
rect 11152 27196 11194 27236
rect 11234 27196 11276 27236
rect 11316 27196 11358 27236
rect 11398 27196 11440 27236
rect 11480 27196 11489 27236
rect 15103 27196 15112 27236
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15480 27196 15489 27236
rect 19103 27196 19112 27236
rect 19152 27196 19194 27236
rect 19234 27196 19276 27236
rect 19316 27196 19358 27236
rect 19398 27196 19440 27236
rect 19480 27196 19489 27236
rect 23103 27196 23112 27236
rect 23152 27196 23194 27236
rect 23234 27196 23276 27236
rect 23316 27196 23358 27236
rect 23398 27196 23440 27236
rect 23480 27196 23489 27236
rect 27103 27196 27112 27236
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27480 27196 27489 27236
rect 31103 27196 31112 27236
rect 31152 27196 31194 27236
rect 31234 27196 31276 27236
rect 31316 27196 31358 27236
rect 31398 27196 31440 27236
rect 31480 27196 31489 27236
rect 35103 27196 35112 27236
rect 35152 27196 35194 27236
rect 35234 27196 35276 27236
rect 35316 27196 35358 27236
rect 35398 27196 35440 27236
rect 35480 27196 35489 27236
rect 39103 27196 39112 27236
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39480 27196 39489 27236
rect 43103 27196 43112 27236
rect 43152 27196 43194 27236
rect 43234 27196 43276 27236
rect 43316 27196 43358 27236
rect 43398 27196 43440 27236
rect 43480 27196 43489 27236
rect 47103 27196 47112 27236
rect 47152 27196 47194 27236
rect 47234 27196 47276 27236
rect 47316 27196 47358 27236
rect 47398 27196 47440 27236
rect 47480 27196 47489 27236
rect 51103 27196 51112 27236
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51480 27196 51489 27236
rect 55103 27196 55112 27236
rect 55152 27196 55194 27236
rect 55234 27196 55276 27236
rect 55316 27196 55358 27236
rect 55398 27196 55440 27236
rect 55480 27196 55489 27236
rect 59103 27196 59112 27236
rect 59152 27196 59194 27236
rect 59234 27196 59276 27236
rect 59316 27196 59358 27236
rect 59398 27196 59440 27236
rect 59480 27196 59489 27236
rect 63103 27196 63112 27236
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63480 27196 63489 27236
rect 67103 27196 67112 27236
rect 67152 27196 67194 27236
rect 67234 27196 67276 27236
rect 67316 27196 67358 27236
rect 67398 27196 67440 27236
rect 67480 27196 67489 27236
rect 71875 26816 71933 26817
rect 69763 26776 69772 26816
rect 69812 26776 70348 26816
rect 70388 26776 70732 26816
rect 70772 26776 71116 26816
rect 71156 26776 71884 26816
rect 71924 26776 71933 26816
rect 71875 26775 71933 26776
rect 69955 26692 69964 26732
rect 70004 26692 71884 26732
rect 71924 26692 71933 26732
rect 0 26588 80 26668
rect 71395 26608 71404 26648
rect 71444 26608 72305 26648
rect 72345 26608 72354 26648
rect 71299 26524 71308 26564
rect 71348 26524 72705 26564
rect 72745 26524 72754 26564
rect 96296 26524 96305 26564
rect 96345 26524 96556 26564
rect 96596 26524 96605 26564
rect 4343 26440 4352 26480
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4720 26440 4729 26480
rect 8343 26440 8352 26480
rect 8392 26440 8434 26480
rect 8474 26440 8516 26480
rect 8556 26440 8598 26480
rect 8638 26440 8680 26480
rect 8720 26440 8729 26480
rect 12343 26440 12352 26480
rect 12392 26440 12434 26480
rect 12474 26440 12516 26480
rect 12556 26440 12598 26480
rect 12638 26440 12680 26480
rect 12720 26440 12729 26480
rect 16343 26440 16352 26480
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16720 26440 16729 26480
rect 20343 26440 20352 26480
rect 20392 26440 20434 26480
rect 20474 26440 20516 26480
rect 20556 26440 20598 26480
rect 20638 26440 20680 26480
rect 20720 26440 20729 26480
rect 24343 26440 24352 26480
rect 24392 26440 24434 26480
rect 24474 26440 24516 26480
rect 24556 26440 24598 26480
rect 24638 26440 24680 26480
rect 24720 26440 24729 26480
rect 28343 26440 28352 26480
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28720 26440 28729 26480
rect 32343 26440 32352 26480
rect 32392 26440 32434 26480
rect 32474 26440 32516 26480
rect 32556 26440 32598 26480
rect 32638 26440 32680 26480
rect 32720 26440 32729 26480
rect 36343 26440 36352 26480
rect 36392 26440 36434 26480
rect 36474 26440 36516 26480
rect 36556 26440 36598 26480
rect 36638 26440 36680 26480
rect 36720 26440 36729 26480
rect 40343 26440 40352 26480
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40720 26440 40729 26480
rect 44343 26440 44352 26480
rect 44392 26440 44434 26480
rect 44474 26440 44516 26480
rect 44556 26440 44598 26480
rect 44638 26440 44680 26480
rect 44720 26440 44729 26480
rect 48343 26440 48352 26480
rect 48392 26440 48434 26480
rect 48474 26440 48516 26480
rect 48556 26440 48598 26480
rect 48638 26440 48680 26480
rect 48720 26440 48729 26480
rect 52343 26440 52352 26480
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52720 26440 52729 26480
rect 56343 26440 56352 26480
rect 56392 26440 56434 26480
rect 56474 26440 56516 26480
rect 56556 26440 56598 26480
rect 56638 26440 56680 26480
rect 56720 26440 56729 26480
rect 60343 26440 60352 26480
rect 60392 26440 60434 26480
rect 60474 26440 60516 26480
rect 60556 26440 60598 26480
rect 60638 26440 60680 26480
rect 60720 26440 60729 26480
rect 64343 26440 64352 26480
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64720 26440 64729 26480
rect 68343 26440 68352 26480
rect 68392 26440 68434 26480
rect 68474 26440 68516 26480
rect 68556 26440 68598 26480
rect 68638 26440 68680 26480
rect 68720 26440 68729 26480
rect 71395 26440 71404 26480
rect 71444 26440 72415 26480
rect 72455 26440 72464 26480
rect 72556 26440 73105 26480
rect 73145 26440 73154 26480
rect 75206 26440 75215 26480
rect 75255 26440 76204 26480
rect 76244 26440 76253 26480
rect 77206 26440 77215 26480
rect 77255 26440 78508 26480
rect 78548 26440 78557 26480
rect 72556 26396 72596 26440
rect 70531 26356 70540 26396
rect 70580 26356 72596 26396
rect 69283 26272 69292 26312
rect 69332 26272 70444 26312
rect 70484 26272 70493 26312
rect 71011 26272 71020 26312
rect 71060 26272 72844 26312
rect 72884 26272 72893 26312
rect 70819 26188 70828 26228
rect 70868 26188 73420 26228
rect 73460 26188 73469 26228
rect 70627 26104 70636 26144
rect 70676 26104 70924 26144
rect 70964 26104 70973 26144
rect 71107 26104 71116 26144
rect 71156 26104 73612 26144
rect 73652 26104 73661 26144
rect 76840 26104 98860 26144
rect 98900 26104 98909 26144
rect 71875 26020 71884 26060
rect 71924 26020 74668 26060
rect 74708 26020 74717 26060
rect 76840 25976 76880 26104
rect 71299 25936 71308 25976
rect 71348 25936 76880 25976
rect 0 25748 80 25828
rect 85699 25724 85757 25725
rect 3103 25684 3112 25724
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3480 25684 3489 25724
rect 7103 25684 7112 25724
rect 7152 25684 7194 25724
rect 7234 25684 7276 25724
rect 7316 25684 7358 25724
rect 7398 25684 7440 25724
rect 7480 25684 7489 25724
rect 11103 25684 11112 25724
rect 11152 25684 11194 25724
rect 11234 25684 11276 25724
rect 11316 25684 11358 25724
rect 11398 25684 11440 25724
rect 11480 25684 11489 25724
rect 15103 25684 15112 25724
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15480 25684 15489 25724
rect 19103 25684 19112 25724
rect 19152 25684 19194 25724
rect 19234 25684 19276 25724
rect 19316 25684 19358 25724
rect 19398 25684 19440 25724
rect 19480 25684 19489 25724
rect 23103 25684 23112 25724
rect 23152 25684 23194 25724
rect 23234 25684 23276 25724
rect 23316 25684 23358 25724
rect 23398 25684 23440 25724
rect 23480 25684 23489 25724
rect 27103 25684 27112 25724
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27480 25684 27489 25724
rect 31103 25684 31112 25724
rect 31152 25684 31194 25724
rect 31234 25684 31276 25724
rect 31316 25684 31358 25724
rect 31398 25684 31440 25724
rect 31480 25684 31489 25724
rect 35103 25684 35112 25724
rect 35152 25684 35194 25724
rect 35234 25684 35276 25724
rect 35316 25684 35358 25724
rect 35398 25684 35440 25724
rect 35480 25684 35489 25724
rect 39103 25684 39112 25724
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39480 25684 39489 25724
rect 43103 25684 43112 25724
rect 43152 25684 43194 25724
rect 43234 25684 43276 25724
rect 43316 25684 43358 25724
rect 43398 25684 43440 25724
rect 43480 25684 43489 25724
rect 47103 25684 47112 25724
rect 47152 25684 47194 25724
rect 47234 25684 47276 25724
rect 47316 25684 47358 25724
rect 47398 25684 47440 25724
rect 47480 25684 47489 25724
rect 51103 25684 51112 25724
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51480 25684 51489 25724
rect 55103 25684 55112 25724
rect 55152 25684 55194 25724
rect 55234 25684 55276 25724
rect 55316 25684 55358 25724
rect 55398 25684 55440 25724
rect 55480 25684 55489 25724
rect 59103 25684 59112 25724
rect 59152 25684 59194 25724
rect 59234 25684 59276 25724
rect 59316 25684 59358 25724
rect 59398 25684 59440 25724
rect 59480 25684 59489 25724
rect 63103 25684 63112 25724
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63480 25684 63489 25724
rect 67103 25684 67112 25724
rect 67152 25684 67194 25724
rect 67234 25684 67276 25724
rect 67316 25684 67358 25724
rect 67398 25684 67440 25724
rect 67480 25684 67489 25724
rect 73123 25684 73132 25724
rect 73172 25684 73804 25724
rect 73844 25684 85708 25724
rect 85748 25684 85757 25724
rect 85699 25683 85757 25684
rect 76483 25600 76492 25640
rect 76532 25600 76876 25640
rect 76916 25600 76925 25640
rect 72739 25516 72748 25556
rect 72788 25516 73228 25556
rect 73268 25516 73277 25556
rect 74851 25516 74860 25556
rect 74900 25516 75916 25556
rect 75956 25516 75965 25556
rect 76771 25516 76780 25556
rect 76820 25516 77164 25556
rect 77204 25516 77213 25556
rect 77635 25516 77644 25556
rect 77684 25516 77932 25556
rect 77972 25516 77981 25556
rect 78595 25516 78604 25556
rect 78644 25516 79756 25556
rect 79796 25516 79805 25556
rect 83683 25516 83692 25556
rect 83732 25516 83980 25556
rect 84020 25516 84029 25556
rect 86851 25516 86860 25556
rect 86900 25516 87532 25556
rect 87572 25516 87581 25556
rect 89635 25516 89644 25556
rect 89684 25516 89932 25556
rect 89972 25516 89981 25556
rect 95683 25516 95692 25556
rect 95732 25516 96076 25556
rect 96116 25516 96125 25556
rect 96451 25516 96460 25556
rect 96500 25516 97420 25556
rect 97460 25516 97469 25556
rect 75235 25432 75244 25472
rect 75284 25432 75532 25472
rect 75572 25432 75581 25472
rect 76003 25432 76012 25472
rect 76052 25432 76492 25472
rect 76532 25432 76541 25472
rect 86947 25432 86956 25472
rect 86996 25432 87380 25472
rect 86851 25388 86909 25389
rect 87340 25388 87380 25432
rect 70435 25348 70444 25388
rect 70484 25348 72940 25388
rect 72980 25348 72989 25388
rect 74467 25348 74476 25388
rect 74516 25348 74668 25388
rect 74708 25348 75052 25388
rect 75092 25348 77548 25388
rect 77588 25348 77597 25388
rect 81187 25348 81196 25388
rect 81236 25348 81580 25388
rect 81620 25348 81629 25388
rect 86851 25348 86860 25388
rect 86900 25348 87148 25388
rect 87188 25348 87197 25388
rect 87331 25348 87340 25388
rect 87380 25348 88876 25388
rect 88916 25348 89548 25388
rect 89588 25348 92332 25388
rect 92372 25348 95692 25388
rect 95732 25348 95741 25388
rect 86851 25347 86909 25348
rect 835 25264 844 25304
rect 884 25264 59240 25304
rect 70915 25264 70924 25304
rect 70964 25264 72652 25304
rect 72692 25264 73324 25304
rect 73364 25264 73373 25304
rect 75523 25264 75532 25304
rect 75572 25264 76012 25304
rect 76052 25264 76300 25304
rect 76340 25264 76588 25304
rect 76628 25264 76780 25304
rect 76820 25264 76829 25304
rect 77731 25264 77740 25304
rect 77780 25264 78028 25304
rect 78068 25264 78316 25304
rect 78356 25264 78892 25304
rect 78932 25264 79372 25304
rect 79412 25264 79852 25304
rect 79892 25264 80044 25304
rect 80084 25264 80093 25304
rect 83779 25264 83788 25304
rect 83828 25264 84076 25304
rect 84116 25264 84364 25304
rect 84404 25264 84652 25304
rect 84692 25264 84940 25304
rect 84980 25264 85132 25304
rect 85172 25264 85516 25304
rect 85556 25264 85900 25304
rect 85940 25264 85949 25304
rect 86563 25264 86572 25304
rect 86612 25264 86764 25304
rect 86804 25264 87628 25304
rect 87668 25264 87916 25304
rect 87956 25264 88204 25304
rect 88244 25264 88492 25304
rect 88532 25264 88684 25304
rect 88724 25264 88733 25304
rect 89731 25264 89740 25304
rect 89780 25264 90028 25304
rect 90068 25264 90316 25304
rect 90356 25264 90604 25304
rect 90644 25264 90892 25304
rect 90932 25264 91276 25304
rect 91316 25264 91948 25304
rect 91988 25264 91997 25304
rect 92515 25264 92524 25304
rect 92564 25264 92908 25304
rect 92948 25264 93676 25304
rect 93716 25264 93964 25304
rect 94004 25264 94156 25304
rect 94196 25264 94924 25304
rect 94964 25264 94973 25304
rect 96739 25264 96748 25304
rect 96788 25264 97036 25304
rect 97076 25264 97516 25304
rect 97556 25264 97804 25304
rect 97844 25264 97996 25304
rect 98036 25264 98045 25304
rect 59200 25220 59240 25264
rect 96748 25220 96788 25264
rect 59200 25180 71308 25220
rect 71348 25180 71357 25220
rect 80419 25180 80428 25220
rect 80468 25180 80716 25220
rect 80756 25180 80908 25220
rect 80948 25180 81100 25220
rect 81140 25180 81484 25220
rect 81524 25180 82252 25220
rect 82292 25180 82732 25220
rect 82772 25180 82781 25220
rect 95884 25180 96172 25220
rect 96212 25180 96460 25220
rect 96500 25180 96788 25220
rect 95884 25136 95924 25180
rect 73891 25096 73900 25136
rect 73940 25096 74284 25136
rect 74324 25096 74333 25136
rect 95875 25096 95884 25136
rect 95924 25096 95933 25136
rect 0 24968 80 24988
rect 0 24928 652 24968
rect 692 24928 701 24968
rect 4343 24928 4352 24968
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4720 24928 4729 24968
rect 8343 24928 8352 24968
rect 8392 24928 8434 24968
rect 8474 24928 8516 24968
rect 8556 24928 8598 24968
rect 8638 24928 8680 24968
rect 8720 24928 8729 24968
rect 12343 24928 12352 24968
rect 12392 24928 12434 24968
rect 12474 24928 12516 24968
rect 12556 24928 12598 24968
rect 12638 24928 12680 24968
rect 12720 24928 12729 24968
rect 16343 24928 16352 24968
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16720 24928 16729 24968
rect 20343 24928 20352 24968
rect 20392 24928 20434 24968
rect 20474 24928 20516 24968
rect 20556 24928 20598 24968
rect 20638 24928 20680 24968
rect 20720 24928 20729 24968
rect 24343 24928 24352 24968
rect 24392 24928 24434 24968
rect 24474 24928 24516 24968
rect 24556 24928 24598 24968
rect 24638 24928 24680 24968
rect 24720 24928 24729 24968
rect 28343 24928 28352 24968
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28720 24928 28729 24968
rect 32343 24928 32352 24968
rect 32392 24928 32434 24968
rect 32474 24928 32516 24968
rect 32556 24928 32598 24968
rect 32638 24928 32680 24968
rect 32720 24928 32729 24968
rect 36343 24928 36352 24968
rect 36392 24928 36434 24968
rect 36474 24928 36516 24968
rect 36556 24928 36598 24968
rect 36638 24928 36680 24968
rect 36720 24928 36729 24968
rect 40343 24928 40352 24968
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40720 24928 40729 24968
rect 44343 24928 44352 24968
rect 44392 24928 44434 24968
rect 44474 24928 44516 24968
rect 44556 24928 44598 24968
rect 44638 24928 44680 24968
rect 44720 24928 44729 24968
rect 48343 24928 48352 24968
rect 48392 24928 48434 24968
rect 48474 24928 48516 24968
rect 48556 24928 48598 24968
rect 48638 24928 48680 24968
rect 48720 24928 48729 24968
rect 52343 24928 52352 24968
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52720 24928 52729 24968
rect 56343 24928 56352 24968
rect 56392 24928 56434 24968
rect 56474 24928 56516 24968
rect 56556 24928 56598 24968
rect 56638 24928 56680 24968
rect 56720 24928 56729 24968
rect 60343 24928 60352 24968
rect 60392 24928 60434 24968
rect 60474 24928 60516 24968
rect 60556 24928 60598 24968
rect 60638 24928 60680 24968
rect 60720 24928 60729 24968
rect 64343 24928 64352 24968
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64720 24928 64729 24968
rect 68343 24928 68352 24968
rect 68392 24928 68434 24968
rect 68474 24928 68516 24968
rect 68556 24928 68598 24968
rect 68638 24928 68680 24968
rect 68720 24928 68729 24968
rect 73315 24928 73324 24968
rect 73364 24928 73996 24968
rect 74036 24928 74045 24968
rect 76867 24928 76876 24968
rect 76916 24928 77068 24968
rect 77108 24928 77117 24968
rect 0 24908 80 24928
rect 73507 24760 73516 24800
rect 73556 24760 74380 24800
rect 74420 24760 74429 24800
rect 81379 24760 81388 24800
rect 81428 24760 81964 24800
rect 82004 24760 82013 24800
rect 95395 24760 95404 24800
rect 95444 24760 95980 24800
rect 96020 24760 96364 24800
rect 96404 24760 96748 24800
rect 96788 24760 97132 24800
rect 97172 24760 97516 24800
rect 97556 24760 97565 24800
rect 71779 24676 71788 24716
rect 71828 24676 73996 24716
rect 74036 24676 74188 24716
rect 74228 24676 75724 24716
rect 75764 24676 75773 24716
rect 73219 24632 73277 24633
rect 835 24592 844 24632
rect 884 24592 71020 24632
rect 71060 24592 71069 24632
rect 73134 24592 73228 24632
rect 73268 24592 73277 24632
rect 73219 24591 73277 24592
rect 73603 24508 73612 24548
rect 73652 24508 74284 24548
rect 74324 24508 74668 24548
rect 74708 24508 75244 24548
rect 75284 24508 76012 24548
rect 76052 24508 76396 24548
rect 76436 24508 76876 24548
rect 76916 24508 76925 24548
rect 77251 24508 77260 24548
rect 77300 24508 77836 24548
rect 77876 24508 78220 24548
rect 78260 24508 78604 24548
rect 78644 24508 78988 24548
rect 79028 24508 79372 24548
rect 79412 24508 79756 24548
rect 79796 24508 80140 24548
rect 80180 24508 80189 24548
rect 83299 24508 83308 24548
rect 83348 24508 83692 24548
rect 83732 24508 84268 24548
rect 84308 24508 84652 24548
rect 84692 24508 85036 24548
rect 85076 24508 85324 24548
rect 85364 24508 85373 24548
rect 86083 24508 86092 24548
rect 86132 24508 86476 24548
rect 86516 24508 86764 24548
rect 86804 24508 86956 24548
rect 86996 24508 87340 24548
rect 87380 24508 87820 24548
rect 87860 24508 88108 24548
rect 88148 24508 88492 24548
rect 88532 24508 88541 24548
rect 89059 24508 89068 24548
rect 89108 24508 89260 24548
rect 89300 24508 89740 24548
rect 89780 24508 90124 24548
rect 90164 24508 90508 24548
rect 90548 24508 90988 24548
rect 91028 24508 91660 24548
rect 91700 24508 91709 24548
rect 92323 24508 92332 24548
rect 92372 24508 92524 24548
rect 92564 24508 93100 24548
rect 93140 24508 93484 24548
rect 93524 24508 93772 24548
rect 93812 24508 94156 24548
rect 94196 24508 94540 24548
rect 94580 24508 94589 24548
rect 97507 24508 97516 24548
rect 97556 24508 97900 24548
rect 97940 24508 98284 24548
rect 98324 24508 98333 24548
rect 74371 24340 74380 24380
rect 74420 24340 74764 24380
rect 74804 24340 80620 24380
rect 80660 24340 83596 24380
rect 83636 24340 84076 24380
rect 84116 24340 84125 24380
rect 3103 24172 3112 24212
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3480 24172 3489 24212
rect 7103 24172 7112 24212
rect 7152 24172 7194 24212
rect 7234 24172 7276 24212
rect 7316 24172 7358 24212
rect 7398 24172 7440 24212
rect 7480 24172 7489 24212
rect 11103 24172 11112 24212
rect 11152 24172 11194 24212
rect 11234 24172 11276 24212
rect 11316 24172 11358 24212
rect 11398 24172 11440 24212
rect 11480 24172 11489 24212
rect 15103 24172 15112 24212
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15480 24172 15489 24212
rect 19103 24172 19112 24212
rect 19152 24172 19194 24212
rect 19234 24172 19276 24212
rect 19316 24172 19358 24212
rect 19398 24172 19440 24212
rect 19480 24172 19489 24212
rect 23103 24172 23112 24212
rect 23152 24172 23194 24212
rect 23234 24172 23276 24212
rect 23316 24172 23358 24212
rect 23398 24172 23440 24212
rect 23480 24172 23489 24212
rect 27103 24172 27112 24212
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27480 24172 27489 24212
rect 31103 24172 31112 24212
rect 31152 24172 31194 24212
rect 31234 24172 31276 24212
rect 31316 24172 31358 24212
rect 31398 24172 31440 24212
rect 31480 24172 31489 24212
rect 35103 24172 35112 24212
rect 35152 24172 35194 24212
rect 35234 24172 35276 24212
rect 35316 24172 35358 24212
rect 35398 24172 35440 24212
rect 35480 24172 35489 24212
rect 39103 24172 39112 24212
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39480 24172 39489 24212
rect 43103 24172 43112 24212
rect 43152 24172 43194 24212
rect 43234 24172 43276 24212
rect 43316 24172 43358 24212
rect 43398 24172 43440 24212
rect 43480 24172 43489 24212
rect 47103 24172 47112 24212
rect 47152 24172 47194 24212
rect 47234 24172 47276 24212
rect 47316 24172 47358 24212
rect 47398 24172 47440 24212
rect 47480 24172 47489 24212
rect 51103 24172 51112 24212
rect 51152 24172 51194 24212
rect 51234 24172 51276 24212
rect 51316 24172 51358 24212
rect 51398 24172 51440 24212
rect 51480 24172 51489 24212
rect 55103 24172 55112 24212
rect 55152 24172 55194 24212
rect 55234 24172 55276 24212
rect 55316 24172 55358 24212
rect 55398 24172 55440 24212
rect 55480 24172 55489 24212
rect 59103 24172 59112 24212
rect 59152 24172 59194 24212
rect 59234 24172 59276 24212
rect 59316 24172 59358 24212
rect 59398 24172 59440 24212
rect 59480 24172 59489 24212
rect 63103 24172 63112 24212
rect 63152 24172 63194 24212
rect 63234 24172 63276 24212
rect 63316 24172 63358 24212
rect 63398 24172 63440 24212
rect 63480 24172 63489 24212
rect 67103 24172 67112 24212
rect 67152 24172 67194 24212
rect 67234 24172 67276 24212
rect 67316 24172 67358 24212
rect 67398 24172 67440 24212
rect 67480 24172 67489 24212
rect 71103 24172 71112 24212
rect 71152 24172 71194 24212
rect 71234 24172 71276 24212
rect 71316 24172 71358 24212
rect 71398 24172 71440 24212
rect 71480 24172 71489 24212
rect 75103 24172 75112 24212
rect 75152 24172 75194 24212
rect 75234 24172 75276 24212
rect 75316 24172 75358 24212
rect 75398 24172 75440 24212
rect 75480 24172 75489 24212
rect 79103 24172 79112 24212
rect 79152 24172 79194 24212
rect 79234 24172 79276 24212
rect 79316 24172 79358 24212
rect 79398 24172 79440 24212
rect 79480 24172 79489 24212
rect 83103 24172 83112 24212
rect 83152 24172 83194 24212
rect 83234 24172 83276 24212
rect 83316 24172 83358 24212
rect 83398 24172 83440 24212
rect 83480 24172 83489 24212
rect 87103 24172 87112 24212
rect 87152 24172 87194 24212
rect 87234 24172 87276 24212
rect 87316 24172 87358 24212
rect 87398 24172 87440 24212
rect 87480 24172 87489 24212
rect 91103 24172 91112 24212
rect 91152 24172 91194 24212
rect 91234 24172 91276 24212
rect 91316 24172 91358 24212
rect 91398 24172 91440 24212
rect 91480 24172 91489 24212
rect 95103 24172 95112 24212
rect 95152 24172 95194 24212
rect 95234 24172 95276 24212
rect 95316 24172 95358 24212
rect 95398 24172 95440 24212
rect 95480 24172 95489 24212
rect 99103 24172 99112 24212
rect 99152 24172 99194 24212
rect 99234 24172 99276 24212
rect 99316 24172 99358 24212
rect 99398 24172 99440 24212
rect 99480 24172 99489 24212
rect 0 24128 80 24148
rect 0 24088 652 24128
rect 692 24088 701 24128
rect 0 24068 80 24088
rect 80323 23836 80332 23876
rect 80372 23836 80812 23876
rect 80852 23836 81388 23876
rect 81428 23836 81676 23876
rect 81716 23836 82156 23876
rect 82196 23836 82444 23876
rect 82484 23836 82493 23876
rect 84931 23836 84940 23876
rect 84980 23836 85708 23876
rect 85748 23836 85757 23876
rect 835 23752 844 23792
rect 884 23752 2092 23792
rect 2132 23752 2141 23792
rect 4343 23416 4352 23456
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4720 23416 4729 23456
rect 8343 23416 8352 23456
rect 8392 23416 8434 23456
rect 8474 23416 8516 23456
rect 8556 23416 8598 23456
rect 8638 23416 8680 23456
rect 8720 23416 8729 23456
rect 12343 23416 12352 23456
rect 12392 23416 12434 23456
rect 12474 23416 12516 23456
rect 12556 23416 12598 23456
rect 12638 23416 12680 23456
rect 12720 23416 12729 23456
rect 16343 23416 16352 23456
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16720 23416 16729 23456
rect 20343 23416 20352 23456
rect 20392 23416 20434 23456
rect 20474 23416 20516 23456
rect 20556 23416 20598 23456
rect 20638 23416 20680 23456
rect 20720 23416 20729 23456
rect 24343 23416 24352 23456
rect 24392 23416 24434 23456
rect 24474 23416 24516 23456
rect 24556 23416 24598 23456
rect 24638 23416 24680 23456
rect 24720 23416 24729 23456
rect 28343 23416 28352 23456
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28720 23416 28729 23456
rect 32343 23416 32352 23456
rect 32392 23416 32434 23456
rect 32474 23416 32516 23456
rect 32556 23416 32598 23456
rect 32638 23416 32680 23456
rect 32720 23416 32729 23456
rect 36343 23416 36352 23456
rect 36392 23416 36434 23456
rect 36474 23416 36516 23456
rect 36556 23416 36598 23456
rect 36638 23416 36680 23456
rect 36720 23416 36729 23456
rect 40343 23416 40352 23456
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40720 23416 40729 23456
rect 44343 23416 44352 23456
rect 44392 23416 44434 23456
rect 44474 23416 44516 23456
rect 44556 23416 44598 23456
rect 44638 23416 44680 23456
rect 44720 23416 44729 23456
rect 48343 23416 48352 23456
rect 48392 23416 48434 23456
rect 48474 23416 48516 23456
rect 48556 23416 48598 23456
rect 48638 23416 48680 23456
rect 48720 23416 48729 23456
rect 52343 23416 52352 23456
rect 52392 23416 52434 23456
rect 52474 23416 52516 23456
rect 52556 23416 52598 23456
rect 52638 23416 52680 23456
rect 52720 23416 52729 23456
rect 56343 23416 56352 23456
rect 56392 23416 56434 23456
rect 56474 23416 56516 23456
rect 56556 23416 56598 23456
rect 56638 23416 56680 23456
rect 56720 23416 56729 23456
rect 60343 23416 60352 23456
rect 60392 23416 60434 23456
rect 60474 23416 60516 23456
rect 60556 23416 60598 23456
rect 60638 23416 60680 23456
rect 60720 23416 60729 23456
rect 64343 23416 64352 23456
rect 64392 23416 64434 23456
rect 64474 23416 64516 23456
rect 64556 23416 64598 23456
rect 64638 23416 64680 23456
rect 64720 23416 64729 23456
rect 68343 23416 68352 23456
rect 68392 23416 68434 23456
rect 68474 23416 68516 23456
rect 68556 23416 68598 23456
rect 68638 23416 68680 23456
rect 68720 23416 68729 23456
rect 72343 23416 72352 23456
rect 72392 23416 72434 23456
rect 72474 23416 72516 23456
rect 72556 23416 72598 23456
rect 72638 23416 72680 23456
rect 72720 23416 72729 23456
rect 76343 23416 76352 23456
rect 76392 23416 76434 23456
rect 76474 23416 76516 23456
rect 76556 23416 76598 23456
rect 76638 23416 76680 23456
rect 76720 23416 76729 23456
rect 80343 23416 80352 23456
rect 80392 23416 80434 23456
rect 80474 23416 80516 23456
rect 80556 23416 80598 23456
rect 80638 23416 80680 23456
rect 80720 23416 80729 23456
rect 84343 23416 84352 23456
rect 84392 23416 84434 23456
rect 84474 23416 84516 23456
rect 84556 23416 84598 23456
rect 84638 23416 84680 23456
rect 84720 23416 84729 23456
rect 88343 23416 88352 23456
rect 88392 23416 88434 23456
rect 88474 23416 88516 23456
rect 88556 23416 88598 23456
rect 88638 23416 88680 23456
rect 88720 23416 88729 23456
rect 92343 23416 92352 23456
rect 92392 23416 92434 23456
rect 92474 23416 92516 23456
rect 92556 23416 92598 23456
rect 92638 23416 92680 23456
rect 92720 23416 92729 23456
rect 96343 23416 96352 23456
rect 96392 23416 96434 23456
rect 96474 23416 96516 23456
rect 96556 23416 96598 23456
rect 96638 23416 96680 23456
rect 96720 23416 96729 23456
rect 0 23288 80 23308
rect 0 23248 652 23288
rect 692 23248 701 23288
rect 2083 23248 2092 23288
rect 2132 23248 69292 23288
rect 69332 23248 69341 23288
rect 0 23228 80 23248
rect 835 23080 844 23120
rect 884 23080 1996 23120
rect 2036 23080 2045 23120
rect 3103 22660 3112 22700
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3480 22660 3489 22700
rect 7103 22660 7112 22700
rect 7152 22660 7194 22700
rect 7234 22660 7276 22700
rect 7316 22660 7358 22700
rect 7398 22660 7440 22700
rect 7480 22660 7489 22700
rect 11103 22660 11112 22700
rect 11152 22660 11194 22700
rect 11234 22660 11276 22700
rect 11316 22660 11358 22700
rect 11398 22660 11440 22700
rect 11480 22660 11489 22700
rect 15103 22660 15112 22700
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15480 22660 15489 22700
rect 19103 22660 19112 22700
rect 19152 22660 19194 22700
rect 19234 22660 19276 22700
rect 19316 22660 19358 22700
rect 19398 22660 19440 22700
rect 19480 22660 19489 22700
rect 23103 22660 23112 22700
rect 23152 22660 23194 22700
rect 23234 22660 23276 22700
rect 23316 22660 23358 22700
rect 23398 22660 23440 22700
rect 23480 22660 23489 22700
rect 27103 22660 27112 22700
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27480 22660 27489 22700
rect 31103 22660 31112 22700
rect 31152 22660 31194 22700
rect 31234 22660 31276 22700
rect 31316 22660 31358 22700
rect 31398 22660 31440 22700
rect 31480 22660 31489 22700
rect 35103 22660 35112 22700
rect 35152 22660 35194 22700
rect 35234 22660 35276 22700
rect 35316 22660 35358 22700
rect 35398 22660 35440 22700
rect 35480 22660 35489 22700
rect 39103 22660 39112 22700
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39480 22660 39489 22700
rect 43103 22660 43112 22700
rect 43152 22660 43194 22700
rect 43234 22660 43276 22700
rect 43316 22660 43358 22700
rect 43398 22660 43440 22700
rect 43480 22660 43489 22700
rect 47103 22660 47112 22700
rect 47152 22660 47194 22700
rect 47234 22660 47276 22700
rect 47316 22660 47358 22700
rect 47398 22660 47440 22700
rect 47480 22660 47489 22700
rect 51103 22660 51112 22700
rect 51152 22660 51194 22700
rect 51234 22660 51276 22700
rect 51316 22660 51358 22700
rect 51398 22660 51440 22700
rect 51480 22660 51489 22700
rect 55103 22660 55112 22700
rect 55152 22660 55194 22700
rect 55234 22660 55276 22700
rect 55316 22660 55358 22700
rect 55398 22660 55440 22700
rect 55480 22660 55489 22700
rect 59103 22660 59112 22700
rect 59152 22660 59194 22700
rect 59234 22660 59276 22700
rect 59316 22660 59358 22700
rect 59398 22660 59440 22700
rect 59480 22660 59489 22700
rect 63103 22660 63112 22700
rect 63152 22660 63194 22700
rect 63234 22660 63276 22700
rect 63316 22660 63358 22700
rect 63398 22660 63440 22700
rect 63480 22660 63489 22700
rect 67103 22660 67112 22700
rect 67152 22660 67194 22700
rect 67234 22660 67276 22700
rect 67316 22660 67358 22700
rect 67398 22660 67440 22700
rect 67480 22660 67489 22700
rect 71103 22660 71112 22700
rect 71152 22660 71194 22700
rect 71234 22660 71276 22700
rect 71316 22660 71358 22700
rect 71398 22660 71440 22700
rect 71480 22660 71489 22700
rect 75103 22660 75112 22700
rect 75152 22660 75194 22700
rect 75234 22660 75276 22700
rect 75316 22660 75358 22700
rect 75398 22660 75440 22700
rect 75480 22660 75489 22700
rect 79103 22660 79112 22700
rect 79152 22660 79194 22700
rect 79234 22660 79276 22700
rect 79316 22660 79358 22700
rect 79398 22660 79440 22700
rect 79480 22660 79489 22700
rect 83103 22660 83112 22700
rect 83152 22660 83194 22700
rect 83234 22660 83276 22700
rect 83316 22660 83358 22700
rect 83398 22660 83440 22700
rect 83480 22660 83489 22700
rect 87103 22660 87112 22700
rect 87152 22660 87194 22700
rect 87234 22660 87276 22700
rect 87316 22660 87358 22700
rect 87398 22660 87440 22700
rect 87480 22660 87489 22700
rect 91103 22660 91112 22700
rect 91152 22660 91194 22700
rect 91234 22660 91276 22700
rect 91316 22660 91358 22700
rect 91398 22660 91440 22700
rect 91480 22660 91489 22700
rect 95103 22660 95112 22700
rect 95152 22660 95194 22700
rect 95234 22660 95276 22700
rect 95316 22660 95358 22700
rect 95398 22660 95440 22700
rect 95480 22660 95489 22700
rect 99103 22660 99112 22700
rect 99152 22660 99194 22700
rect 99234 22660 99276 22700
rect 99316 22660 99358 22700
rect 99398 22660 99440 22700
rect 99480 22660 99489 22700
rect 0 22448 80 22468
rect 0 22408 556 22448
rect 596 22408 605 22448
rect 0 22388 80 22408
rect 4343 21904 4352 21944
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4720 21904 4729 21944
rect 8343 21904 8352 21944
rect 8392 21904 8434 21944
rect 8474 21904 8516 21944
rect 8556 21904 8598 21944
rect 8638 21904 8680 21944
rect 8720 21904 8729 21944
rect 12343 21904 12352 21944
rect 12392 21904 12434 21944
rect 12474 21904 12516 21944
rect 12556 21904 12598 21944
rect 12638 21904 12680 21944
rect 12720 21904 12729 21944
rect 16343 21904 16352 21944
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16720 21904 16729 21944
rect 20343 21904 20352 21944
rect 20392 21904 20434 21944
rect 20474 21904 20516 21944
rect 20556 21904 20598 21944
rect 20638 21904 20680 21944
rect 20720 21904 20729 21944
rect 24343 21904 24352 21944
rect 24392 21904 24434 21944
rect 24474 21904 24516 21944
rect 24556 21904 24598 21944
rect 24638 21904 24680 21944
rect 24720 21904 24729 21944
rect 28343 21904 28352 21944
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28720 21904 28729 21944
rect 32343 21904 32352 21944
rect 32392 21904 32434 21944
rect 32474 21904 32516 21944
rect 32556 21904 32598 21944
rect 32638 21904 32680 21944
rect 32720 21904 32729 21944
rect 36343 21904 36352 21944
rect 36392 21904 36434 21944
rect 36474 21904 36516 21944
rect 36556 21904 36598 21944
rect 36638 21904 36680 21944
rect 36720 21904 36729 21944
rect 40343 21904 40352 21944
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40720 21904 40729 21944
rect 44343 21904 44352 21944
rect 44392 21904 44434 21944
rect 44474 21904 44516 21944
rect 44556 21904 44598 21944
rect 44638 21904 44680 21944
rect 44720 21904 44729 21944
rect 48343 21904 48352 21944
rect 48392 21904 48434 21944
rect 48474 21904 48516 21944
rect 48556 21904 48598 21944
rect 48638 21904 48680 21944
rect 48720 21904 48729 21944
rect 52343 21904 52352 21944
rect 52392 21904 52434 21944
rect 52474 21904 52516 21944
rect 52556 21904 52598 21944
rect 52638 21904 52680 21944
rect 52720 21904 52729 21944
rect 56343 21904 56352 21944
rect 56392 21904 56434 21944
rect 56474 21904 56516 21944
rect 56556 21904 56598 21944
rect 56638 21904 56680 21944
rect 56720 21904 56729 21944
rect 60343 21904 60352 21944
rect 60392 21904 60434 21944
rect 60474 21904 60516 21944
rect 60556 21904 60598 21944
rect 60638 21904 60680 21944
rect 60720 21904 60729 21944
rect 64343 21904 64352 21944
rect 64392 21904 64434 21944
rect 64474 21904 64516 21944
rect 64556 21904 64598 21944
rect 64638 21904 64680 21944
rect 64720 21904 64729 21944
rect 68343 21904 68352 21944
rect 68392 21904 68434 21944
rect 68474 21904 68516 21944
rect 68556 21904 68598 21944
rect 68638 21904 68680 21944
rect 68720 21904 68729 21944
rect 72343 21904 72352 21944
rect 72392 21904 72434 21944
rect 72474 21904 72516 21944
rect 72556 21904 72598 21944
rect 72638 21904 72680 21944
rect 72720 21904 72729 21944
rect 76343 21904 76352 21944
rect 76392 21904 76434 21944
rect 76474 21904 76516 21944
rect 76556 21904 76598 21944
rect 76638 21904 76680 21944
rect 76720 21904 76729 21944
rect 80343 21904 80352 21944
rect 80392 21904 80434 21944
rect 80474 21904 80516 21944
rect 80556 21904 80598 21944
rect 80638 21904 80680 21944
rect 80720 21904 80729 21944
rect 84343 21904 84352 21944
rect 84392 21904 84434 21944
rect 84474 21904 84516 21944
rect 84556 21904 84598 21944
rect 84638 21904 84680 21944
rect 84720 21904 84729 21944
rect 88343 21904 88352 21944
rect 88392 21904 88434 21944
rect 88474 21904 88516 21944
rect 88556 21904 88598 21944
rect 88638 21904 88680 21944
rect 88720 21904 88729 21944
rect 92343 21904 92352 21944
rect 92392 21904 92434 21944
rect 92474 21904 92516 21944
rect 92556 21904 92598 21944
rect 92638 21904 92680 21944
rect 92720 21904 92729 21944
rect 96343 21904 96352 21944
rect 96392 21904 96434 21944
rect 96474 21904 96516 21944
rect 96556 21904 96598 21944
rect 96638 21904 96680 21944
rect 96720 21904 96729 21944
rect 0 21608 80 21628
rect 0 21568 652 21608
rect 692 21568 701 21608
rect 0 21548 80 21568
rect 3103 21148 3112 21188
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3480 21148 3489 21188
rect 7103 21148 7112 21188
rect 7152 21148 7194 21188
rect 7234 21148 7276 21188
rect 7316 21148 7358 21188
rect 7398 21148 7440 21188
rect 7480 21148 7489 21188
rect 11103 21148 11112 21188
rect 11152 21148 11194 21188
rect 11234 21148 11276 21188
rect 11316 21148 11358 21188
rect 11398 21148 11440 21188
rect 11480 21148 11489 21188
rect 15103 21148 15112 21188
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15480 21148 15489 21188
rect 19103 21148 19112 21188
rect 19152 21148 19194 21188
rect 19234 21148 19276 21188
rect 19316 21148 19358 21188
rect 19398 21148 19440 21188
rect 19480 21148 19489 21188
rect 23103 21148 23112 21188
rect 23152 21148 23194 21188
rect 23234 21148 23276 21188
rect 23316 21148 23358 21188
rect 23398 21148 23440 21188
rect 23480 21148 23489 21188
rect 27103 21148 27112 21188
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27480 21148 27489 21188
rect 31103 21148 31112 21188
rect 31152 21148 31194 21188
rect 31234 21148 31276 21188
rect 31316 21148 31358 21188
rect 31398 21148 31440 21188
rect 31480 21148 31489 21188
rect 35103 21148 35112 21188
rect 35152 21148 35194 21188
rect 35234 21148 35276 21188
rect 35316 21148 35358 21188
rect 35398 21148 35440 21188
rect 35480 21148 35489 21188
rect 39103 21148 39112 21188
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39480 21148 39489 21188
rect 43103 21148 43112 21188
rect 43152 21148 43194 21188
rect 43234 21148 43276 21188
rect 43316 21148 43358 21188
rect 43398 21148 43440 21188
rect 43480 21148 43489 21188
rect 47103 21148 47112 21188
rect 47152 21148 47194 21188
rect 47234 21148 47276 21188
rect 47316 21148 47358 21188
rect 47398 21148 47440 21188
rect 47480 21148 47489 21188
rect 51103 21148 51112 21188
rect 51152 21148 51194 21188
rect 51234 21148 51276 21188
rect 51316 21148 51358 21188
rect 51398 21148 51440 21188
rect 51480 21148 51489 21188
rect 55103 21148 55112 21188
rect 55152 21148 55194 21188
rect 55234 21148 55276 21188
rect 55316 21148 55358 21188
rect 55398 21148 55440 21188
rect 55480 21148 55489 21188
rect 59103 21148 59112 21188
rect 59152 21148 59194 21188
rect 59234 21148 59276 21188
rect 59316 21148 59358 21188
rect 59398 21148 59440 21188
rect 59480 21148 59489 21188
rect 63103 21148 63112 21188
rect 63152 21148 63194 21188
rect 63234 21148 63276 21188
rect 63316 21148 63358 21188
rect 63398 21148 63440 21188
rect 63480 21148 63489 21188
rect 67103 21148 67112 21188
rect 67152 21148 67194 21188
rect 67234 21148 67276 21188
rect 67316 21148 67358 21188
rect 67398 21148 67440 21188
rect 67480 21148 67489 21188
rect 71103 21148 71112 21188
rect 71152 21148 71194 21188
rect 71234 21148 71276 21188
rect 71316 21148 71358 21188
rect 71398 21148 71440 21188
rect 71480 21148 71489 21188
rect 75103 21148 75112 21188
rect 75152 21148 75194 21188
rect 75234 21148 75276 21188
rect 75316 21148 75358 21188
rect 75398 21148 75440 21188
rect 75480 21148 75489 21188
rect 79103 21148 79112 21188
rect 79152 21148 79194 21188
rect 79234 21148 79276 21188
rect 79316 21148 79358 21188
rect 79398 21148 79440 21188
rect 79480 21148 79489 21188
rect 83103 21148 83112 21188
rect 83152 21148 83194 21188
rect 83234 21148 83276 21188
rect 83316 21148 83358 21188
rect 83398 21148 83440 21188
rect 83480 21148 83489 21188
rect 87103 21148 87112 21188
rect 87152 21148 87194 21188
rect 87234 21148 87276 21188
rect 87316 21148 87358 21188
rect 87398 21148 87440 21188
rect 87480 21148 87489 21188
rect 91103 21148 91112 21188
rect 91152 21148 91194 21188
rect 91234 21148 91276 21188
rect 91316 21148 91358 21188
rect 91398 21148 91440 21188
rect 91480 21148 91489 21188
rect 95103 21148 95112 21188
rect 95152 21148 95194 21188
rect 95234 21148 95276 21188
rect 95316 21148 95358 21188
rect 95398 21148 95440 21188
rect 95480 21148 95489 21188
rect 99103 21148 99112 21188
rect 99152 21148 99194 21188
rect 99234 21148 99276 21188
rect 99316 21148 99358 21188
rect 99398 21148 99440 21188
rect 99480 21148 99489 21188
rect 0 20768 80 20788
rect 0 20728 652 20768
rect 692 20728 701 20768
rect 0 20708 80 20728
rect 4343 20392 4352 20432
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4720 20392 4729 20432
rect 8343 20392 8352 20432
rect 8392 20392 8434 20432
rect 8474 20392 8516 20432
rect 8556 20392 8598 20432
rect 8638 20392 8680 20432
rect 8720 20392 8729 20432
rect 12343 20392 12352 20432
rect 12392 20392 12434 20432
rect 12474 20392 12516 20432
rect 12556 20392 12598 20432
rect 12638 20392 12680 20432
rect 12720 20392 12729 20432
rect 16343 20392 16352 20432
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16720 20392 16729 20432
rect 20343 20392 20352 20432
rect 20392 20392 20434 20432
rect 20474 20392 20516 20432
rect 20556 20392 20598 20432
rect 20638 20392 20680 20432
rect 20720 20392 20729 20432
rect 24343 20392 24352 20432
rect 24392 20392 24434 20432
rect 24474 20392 24516 20432
rect 24556 20392 24598 20432
rect 24638 20392 24680 20432
rect 24720 20392 24729 20432
rect 28343 20392 28352 20432
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28720 20392 28729 20432
rect 32343 20392 32352 20432
rect 32392 20392 32434 20432
rect 32474 20392 32516 20432
rect 32556 20392 32598 20432
rect 32638 20392 32680 20432
rect 32720 20392 32729 20432
rect 36343 20392 36352 20432
rect 36392 20392 36434 20432
rect 36474 20392 36516 20432
rect 36556 20392 36598 20432
rect 36638 20392 36680 20432
rect 36720 20392 36729 20432
rect 40343 20392 40352 20432
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40720 20392 40729 20432
rect 44343 20392 44352 20432
rect 44392 20392 44434 20432
rect 44474 20392 44516 20432
rect 44556 20392 44598 20432
rect 44638 20392 44680 20432
rect 44720 20392 44729 20432
rect 48343 20392 48352 20432
rect 48392 20392 48434 20432
rect 48474 20392 48516 20432
rect 48556 20392 48598 20432
rect 48638 20392 48680 20432
rect 48720 20392 48729 20432
rect 52343 20392 52352 20432
rect 52392 20392 52434 20432
rect 52474 20392 52516 20432
rect 52556 20392 52598 20432
rect 52638 20392 52680 20432
rect 52720 20392 52729 20432
rect 56343 20392 56352 20432
rect 56392 20392 56434 20432
rect 56474 20392 56516 20432
rect 56556 20392 56598 20432
rect 56638 20392 56680 20432
rect 56720 20392 56729 20432
rect 60343 20392 60352 20432
rect 60392 20392 60434 20432
rect 60474 20392 60516 20432
rect 60556 20392 60598 20432
rect 60638 20392 60680 20432
rect 60720 20392 60729 20432
rect 64343 20392 64352 20432
rect 64392 20392 64434 20432
rect 64474 20392 64516 20432
rect 64556 20392 64598 20432
rect 64638 20392 64680 20432
rect 64720 20392 64729 20432
rect 68343 20392 68352 20432
rect 68392 20392 68434 20432
rect 68474 20392 68516 20432
rect 68556 20392 68598 20432
rect 68638 20392 68680 20432
rect 68720 20392 68729 20432
rect 72343 20392 72352 20432
rect 72392 20392 72434 20432
rect 72474 20392 72516 20432
rect 72556 20392 72598 20432
rect 72638 20392 72680 20432
rect 72720 20392 72729 20432
rect 76343 20392 76352 20432
rect 76392 20392 76434 20432
rect 76474 20392 76516 20432
rect 76556 20392 76598 20432
rect 76638 20392 76680 20432
rect 76720 20392 76729 20432
rect 80343 20392 80352 20432
rect 80392 20392 80434 20432
rect 80474 20392 80516 20432
rect 80556 20392 80598 20432
rect 80638 20392 80680 20432
rect 80720 20392 80729 20432
rect 84343 20392 84352 20432
rect 84392 20392 84434 20432
rect 84474 20392 84516 20432
rect 84556 20392 84598 20432
rect 84638 20392 84680 20432
rect 84720 20392 84729 20432
rect 88343 20392 88352 20432
rect 88392 20392 88434 20432
rect 88474 20392 88516 20432
rect 88556 20392 88598 20432
rect 88638 20392 88680 20432
rect 88720 20392 88729 20432
rect 92343 20392 92352 20432
rect 92392 20392 92434 20432
rect 92474 20392 92516 20432
rect 92556 20392 92598 20432
rect 92638 20392 92680 20432
rect 92720 20392 92729 20432
rect 96343 20392 96352 20432
rect 96392 20392 96434 20432
rect 96474 20392 96516 20432
rect 96556 20392 96598 20432
rect 96638 20392 96680 20432
rect 96720 20392 96729 20432
rect 0 19928 80 19948
rect 0 19888 652 19928
rect 692 19888 701 19928
rect 0 19868 80 19888
rect 3103 19636 3112 19676
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3480 19636 3489 19676
rect 7103 19636 7112 19676
rect 7152 19636 7194 19676
rect 7234 19636 7276 19676
rect 7316 19636 7358 19676
rect 7398 19636 7440 19676
rect 7480 19636 7489 19676
rect 11103 19636 11112 19676
rect 11152 19636 11194 19676
rect 11234 19636 11276 19676
rect 11316 19636 11358 19676
rect 11398 19636 11440 19676
rect 11480 19636 11489 19676
rect 15103 19636 15112 19676
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15480 19636 15489 19676
rect 19103 19636 19112 19676
rect 19152 19636 19194 19676
rect 19234 19636 19276 19676
rect 19316 19636 19358 19676
rect 19398 19636 19440 19676
rect 19480 19636 19489 19676
rect 23103 19636 23112 19676
rect 23152 19636 23194 19676
rect 23234 19636 23276 19676
rect 23316 19636 23358 19676
rect 23398 19636 23440 19676
rect 23480 19636 23489 19676
rect 27103 19636 27112 19676
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27480 19636 27489 19676
rect 31103 19636 31112 19676
rect 31152 19636 31194 19676
rect 31234 19636 31276 19676
rect 31316 19636 31358 19676
rect 31398 19636 31440 19676
rect 31480 19636 31489 19676
rect 35103 19636 35112 19676
rect 35152 19636 35194 19676
rect 35234 19636 35276 19676
rect 35316 19636 35358 19676
rect 35398 19636 35440 19676
rect 35480 19636 35489 19676
rect 39103 19636 39112 19676
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39480 19636 39489 19676
rect 43103 19636 43112 19676
rect 43152 19636 43194 19676
rect 43234 19636 43276 19676
rect 43316 19636 43358 19676
rect 43398 19636 43440 19676
rect 43480 19636 43489 19676
rect 47103 19636 47112 19676
rect 47152 19636 47194 19676
rect 47234 19636 47276 19676
rect 47316 19636 47358 19676
rect 47398 19636 47440 19676
rect 47480 19636 47489 19676
rect 51103 19636 51112 19676
rect 51152 19636 51194 19676
rect 51234 19636 51276 19676
rect 51316 19636 51358 19676
rect 51398 19636 51440 19676
rect 51480 19636 51489 19676
rect 55103 19636 55112 19676
rect 55152 19636 55194 19676
rect 55234 19636 55276 19676
rect 55316 19636 55358 19676
rect 55398 19636 55440 19676
rect 55480 19636 55489 19676
rect 59103 19636 59112 19676
rect 59152 19636 59194 19676
rect 59234 19636 59276 19676
rect 59316 19636 59358 19676
rect 59398 19636 59440 19676
rect 59480 19636 59489 19676
rect 63103 19636 63112 19676
rect 63152 19636 63194 19676
rect 63234 19636 63276 19676
rect 63316 19636 63358 19676
rect 63398 19636 63440 19676
rect 63480 19636 63489 19676
rect 67103 19636 67112 19676
rect 67152 19636 67194 19676
rect 67234 19636 67276 19676
rect 67316 19636 67358 19676
rect 67398 19636 67440 19676
rect 67480 19636 67489 19676
rect 71103 19636 71112 19676
rect 71152 19636 71194 19676
rect 71234 19636 71276 19676
rect 71316 19636 71358 19676
rect 71398 19636 71440 19676
rect 71480 19636 71489 19676
rect 75103 19636 75112 19676
rect 75152 19636 75194 19676
rect 75234 19636 75276 19676
rect 75316 19636 75358 19676
rect 75398 19636 75440 19676
rect 75480 19636 75489 19676
rect 79103 19636 79112 19676
rect 79152 19636 79194 19676
rect 79234 19636 79276 19676
rect 79316 19636 79358 19676
rect 79398 19636 79440 19676
rect 79480 19636 79489 19676
rect 83103 19636 83112 19676
rect 83152 19636 83194 19676
rect 83234 19636 83276 19676
rect 83316 19636 83358 19676
rect 83398 19636 83440 19676
rect 83480 19636 83489 19676
rect 87103 19636 87112 19676
rect 87152 19636 87194 19676
rect 87234 19636 87276 19676
rect 87316 19636 87358 19676
rect 87398 19636 87440 19676
rect 87480 19636 87489 19676
rect 91103 19636 91112 19676
rect 91152 19636 91194 19676
rect 91234 19636 91276 19676
rect 91316 19636 91358 19676
rect 91398 19636 91440 19676
rect 91480 19636 91489 19676
rect 95103 19636 95112 19676
rect 95152 19636 95194 19676
rect 95234 19636 95276 19676
rect 95316 19636 95358 19676
rect 95398 19636 95440 19676
rect 95480 19636 95489 19676
rect 99103 19636 99112 19676
rect 99152 19636 99194 19676
rect 99234 19636 99276 19676
rect 99316 19636 99358 19676
rect 99398 19636 99440 19676
rect 99480 19636 99489 19676
rect 0 19088 80 19108
rect 0 19048 652 19088
rect 692 19048 701 19088
rect 0 19028 80 19048
rect 4343 18880 4352 18920
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4720 18880 4729 18920
rect 8343 18880 8352 18920
rect 8392 18880 8434 18920
rect 8474 18880 8516 18920
rect 8556 18880 8598 18920
rect 8638 18880 8680 18920
rect 8720 18880 8729 18920
rect 12343 18880 12352 18920
rect 12392 18880 12434 18920
rect 12474 18880 12516 18920
rect 12556 18880 12598 18920
rect 12638 18880 12680 18920
rect 12720 18880 12729 18920
rect 16343 18880 16352 18920
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16720 18880 16729 18920
rect 20343 18880 20352 18920
rect 20392 18880 20434 18920
rect 20474 18880 20516 18920
rect 20556 18880 20598 18920
rect 20638 18880 20680 18920
rect 20720 18880 20729 18920
rect 24343 18880 24352 18920
rect 24392 18880 24434 18920
rect 24474 18880 24516 18920
rect 24556 18880 24598 18920
rect 24638 18880 24680 18920
rect 24720 18880 24729 18920
rect 28343 18880 28352 18920
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28720 18880 28729 18920
rect 32343 18880 32352 18920
rect 32392 18880 32434 18920
rect 32474 18880 32516 18920
rect 32556 18880 32598 18920
rect 32638 18880 32680 18920
rect 32720 18880 32729 18920
rect 36343 18880 36352 18920
rect 36392 18880 36434 18920
rect 36474 18880 36516 18920
rect 36556 18880 36598 18920
rect 36638 18880 36680 18920
rect 36720 18880 36729 18920
rect 40343 18880 40352 18920
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40720 18880 40729 18920
rect 44343 18880 44352 18920
rect 44392 18880 44434 18920
rect 44474 18880 44516 18920
rect 44556 18880 44598 18920
rect 44638 18880 44680 18920
rect 44720 18880 44729 18920
rect 48343 18880 48352 18920
rect 48392 18880 48434 18920
rect 48474 18880 48516 18920
rect 48556 18880 48598 18920
rect 48638 18880 48680 18920
rect 48720 18880 48729 18920
rect 52343 18880 52352 18920
rect 52392 18880 52434 18920
rect 52474 18880 52516 18920
rect 52556 18880 52598 18920
rect 52638 18880 52680 18920
rect 52720 18880 52729 18920
rect 56343 18880 56352 18920
rect 56392 18880 56434 18920
rect 56474 18880 56516 18920
rect 56556 18880 56598 18920
rect 56638 18880 56680 18920
rect 56720 18880 56729 18920
rect 60343 18880 60352 18920
rect 60392 18880 60434 18920
rect 60474 18880 60516 18920
rect 60556 18880 60598 18920
rect 60638 18880 60680 18920
rect 60720 18880 60729 18920
rect 64343 18880 64352 18920
rect 64392 18880 64434 18920
rect 64474 18880 64516 18920
rect 64556 18880 64598 18920
rect 64638 18880 64680 18920
rect 64720 18880 64729 18920
rect 68343 18880 68352 18920
rect 68392 18880 68434 18920
rect 68474 18880 68516 18920
rect 68556 18880 68598 18920
rect 68638 18880 68680 18920
rect 68720 18880 68729 18920
rect 72343 18880 72352 18920
rect 72392 18880 72434 18920
rect 72474 18880 72516 18920
rect 72556 18880 72598 18920
rect 72638 18880 72680 18920
rect 72720 18880 72729 18920
rect 76343 18880 76352 18920
rect 76392 18880 76434 18920
rect 76474 18880 76516 18920
rect 76556 18880 76598 18920
rect 76638 18880 76680 18920
rect 76720 18880 76729 18920
rect 80343 18880 80352 18920
rect 80392 18880 80434 18920
rect 80474 18880 80516 18920
rect 80556 18880 80598 18920
rect 80638 18880 80680 18920
rect 80720 18880 80729 18920
rect 84343 18880 84352 18920
rect 84392 18880 84434 18920
rect 84474 18880 84516 18920
rect 84556 18880 84598 18920
rect 84638 18880 84680 18920
rect 84720 18880 84729 18920
rect 88343 18880 88352 18920
rect 88392 18880 88434 18920
rect 88474 18880 88516 18920
rect 88556 18880 88598 18920
rect 88638 18880 88680 18920
rect 88720 18880 88729 18920
rect 92343 18880 92352 18920
rect 92392 18880 92434 18920
rect 92474 18880 92516 18920
rect 92556 18880 92598 18920
rect 92638 18880 92680 18920
rect 92720 18880 92729 18920
rect 96343 18880 96352 18920
rect 96392 18880 96434 18920
rect 96474 18880 96516 18920
rect 96556 18880 96598 18920
rect 96638 18880 96680 18920
rect 96720 18880 96729 18920
rect 0 18248 80 18268
rect 0 18208 652 18248
rect 692 18208 701 18248
rect 0 18188 80 18208
rect 3103 18124 3112 18164
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3480 18124 3489 18164
rect 7103 18124 7112 18164
rect 7152 18124 7194 18164
rect 7234 18124 7276 18164
rect 7316 18124 7358 18164
rect 7398 18124 7440 18164
rect 7480 18124 7489 18164
rect 11103 18124 11112 18164
rect 11152 18124 11194 18164
rect 11234 18124 11276 18164
rect 11316 18124 11358 18164
rect 11398 18124 11440 18164
rect 11480 18124 11489 18164
rect 15103 18124 15112 18164
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15480 18124 15489 18164
rect 19103 18124 19112 18164
rect 19152 18124 19194 18164
rect 19234 18124 19276 18164
rect 19316 18124 19358 18164
rect 19398 18124 19440 18164
rect 19480 18124 19489 18164
rect 23103 18124 23112 18164
rect 23152 18124 23194 18164
rect 23234 18124 23276 18164
rect 23316 18124 23358 18164
rect 23398 18124 23440 18164
rect 23480 18124 23489 18164
rect 27103 18124 27112 18164
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27480 18124 27489 18164
rect 31103 18124 31112 18164
rect 31152 18124 31194 18164
rect 31234 18124 31276 18164
rect 31316 18124 31358 18164
rect 31398 18124 31440 18164
rect 31480 18124 31489 18164
rect 35103 18124 35112 18164
rect 35152 18124 35194 18164
rect 35234 18124 35276 18164
rect 35316 18124 35358 18164
rect 35398 18124 35440 18164
rect 35480 18124 35489 18164
rect 39103 18124 39112 18164
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39480 18124 39489 18164
rect 43103 18124 43112 18164
rect 43152 18124 43194 18164
rect 43234 18124 43276 18164
rect 43316 18124 43358 18164
rect 43398 18124 43440 18164
rect 43480 18124 43489 18164
rect 47103 18124 47112 18164
rect 47152 18124 47194 18164
rect 47234 18124 47276 18164
rect 47316 18124 47358 18164
rect 47398 18124 47440 18164
rect 47480 18124 47489 18164
rect 51103 18124 51112 18164
rect 51152 18124 51194 18164
rect 51234 18124 51276 18164
rect 51316 18124 51358 18164
rect 51398 18124 51440 18164
rect 51480 18124 51489 18164
rect 55103 18124 55112 18164
rect 55152 18124 55194 18164
rect 55234 18124 55276 18164
rect 55316 18124 55358 18164
rect 55398 18124 55440 18164
rect 55480 18124 55489 18164
rect 59103 18124 59112 18164
rect 59152 18124 59194 18164
rect 59234 18124 59276 18164
rect 59316 18124 59358 18164
rect 59398 18124 59440 18164
rect 59480 18124 59489 18164
rect 63103 18124 63112 18164
rect 63152 18124 63194 18164
rect 63234 18124 63276 18164
rect 63316 18124 63358 18164
rect 63398 18124 63440 18164
rect 63480 18124 63489 18164
rect 67103 18124 67112 18164
rect 67152 18124 67194 18164
rect 67234 18124 67276 18164
rect 67316 18124 67358 18164
rect 67398 18124 67440 18164
rect 67480 18124 67489 18164
rect 71103 18124 71112 18164
rect 71152 18124 71194 18164
rect 71234 18124 71276 18164
rect 71316 18124 71358 18164
rect 71398 18124 71440 18164
rect 71480 18124 71489 18164
rect 75103 18124 75112 18164
rect 75152 18124 75194 18164
rect 75234 18124 75276 18164
rect 75316 18124 75358 18164
rect 75398 18124 75440 18164
rect 75480 18124 75489 18164
rect 79103 18124 79112 18164
rect 79152 18124 79194 18164
rect 79234 18124 79276 18164
rect 79316 18124 79358 18164
rect 79398 18124 79440 18164
rect 79480 18124 79489 18164
rect 83103 18124 83112 18164
rect 83152 18124 83194 18164
rect 83234 18124 83276 18164
rect 83316 18124 83358 18164
rect 83398 18124 83440 18164
rect 83480 18124 83489 18164
rect 87103 18124 87112 18164
rect 87152 18124 87194 18164
rect 87234 18124 87276 18164
rect 87316 18124 87358 18164
rect 87398 18124 87440 18164
rect 87480 18124 87489 18164
rect 91103 18124 91112 18164
rect 91152 18124 91194 18164
rect 91234 18124 91276 18164
rect 91316 18124 91358 18164
rect 91398 18124 91440 18164
rect 91480 18124 91489 18164
rect 95103 18124 95112 18164
rect 95152 18124 95194 18164
rect 95234 18124 95276 18164
rect 95316 18124 95358 18164
rect 95398 18124 95440 18164
rect 95480 18124 95489 18164
rect 99103 18124 99112 18164
rect 99152 18124 99194 18164
rect 99234 18124 99276 18164
rect 99316 18124 99358 18164
rect 99398 18124 99440 18164
rect 99480 18124 99489 18164
rect 0 17408 80 17428
rect 0 17368 652 17408
rect 692 17368 701 17408
rect 4343 17368 4352 17408
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4720 17368 4729 17408
rect 8343 17368 8352 17408
rect 8392 17368 8434 17408
rect 8474 17368 8516 17408
rect 8556 17368 8598 17408
rect 8638 17368 8680 17408
rect 8720 17368 8729 17408
rect 12343 17368 12352 17408
rect 12392 17368 12434 17408
rect 12474 17368 12516 17408
rect 12556 17368 12598 17408
rect 12638 17368 12680 17408
rect 12720 17368 12729 17408
rect 16343 17368 16352 17408
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16720 17368 16729 17408
rect 20343 17368 20352 17408
rect 20392 17368 20434 17408
rect 20474 17368 20516 17408
rect 20556 17368 20598 17408
rect 20638 17368 20680 17408
rect 20720 17368 20729 17408
rect 24343 17368 24352 17408
rect 24392 17368 24434 17408
rect 24474 17368 24516 17408
rect 24556 17368 24598 17408
rect 24638 17368 24680 17408
rect 24720 17368 24729 17408
rect 28343 17368 28352 17408
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28720 17368 28729 17408
rect 32343 17368 32352 17408
rect 32392 17368 32434 17408
rect 32474 17368 32516 17408
rect 32556 17368 32598 17408
rect 32638 17368 32680 17408
rect 32720 17368 32729 17408
rect 36343 17368 36352 17408
rect 36392 17368 36434 17408
rect 36474 17368 36516 17408
rect 36556 17368 36598 17408
rect 36638 17368 36680 17408
rect 36720 17368 36729 17408
rect 40343 17368 40352 17408
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40720 17368 40729 17408
rect 44343 17368 44352 17408
rect 44392 17368 44434 17408
rect 44474 17368 44516 17408
rect 44556 17368 44598 17408
rect 44638 17368 44680 17408
rect 44720 17368 44729 17408
rect 48343 17368 48352 17408
rect 48392 17368 48434 17408
rect 48474 17368 48516 17408
rect 48556 17368 48598 17408
rect 48638 17368 48680 17408
rect 48720 17368 48729 17408
rect 52343 17368 52352 17408
rect 52392 17368 52434 17408
rect 52474 17368 52516 17408
rect 52556 17368 52598 17408
rect 52638 17368 52680 17408
rect 52720 17368 52729 17408
rect 56343 17368 56352 17408
rect 56392 17368 56434 17408
rect 56474 17368 56516 17408
rect 56556 17368 56598 17408
rect 56638 17368 56680 17408
rect 56720 17368 56729 17408
rect 60343 17368 60352 17408
rect 60392 17368 60434 17408
rect 60474 17368 60516 17408
rect 60556 17368 60598 17408
rect 60638 17368 60680 17408
rect 60720 17368 60729 17408
rect 64343 17368 64352 17408
rect 64392 17368 64434 17408
rect 64474 17368 64516 17408
rect 64556 17368 64598 17408
rect 64638 17368 64680 17408
rect 64720 17368 64729 17408
rect 68343 17368 68352 17408
rect 68392 17368 68434 17408
rect 68474 17368 68516 17408
rect 68556 17368 68598 17408
rect 68638 17368 68680 17408
rect 68720 17368 68729 17408
rect 72343 17368 72352 17408
rect 72392 17368 72434 17408
rect 72474 17368 72516 17408
rect 72556 17368 72598 17408
rect 72638 17368 72680 17408
rect 72720 17368 72729 17408
rect 76343 17368 76352 17408
rect 76392 17368 76434 17408
rect 76474 17368 76516 17408
rect 76556 17368 76598 17408
rect 76638 17368 76680 17408
rect 76720 17368 76729 17408
rect 80343 17368 80352 17408
rect 80392 17368 80434 17408
rect 80474 17368 80516 17408
rect 80556 17368 80598 17408
rect 80638 17368 80680 17408
rect 80720 17368 80729 17408
rect 84343 17368 84352 17408
rect 84392 17368 84434 17408
rect 84474 17368 84516 17408
rect 84556 17368 84598 17408
rect 84638 17368 84680 17408
rect 84720 17368 84729 17408
rect 88343 17368 88352 17408
rect 88392 17368 88434 17408
rect 88474 17368 88516 17408
rect 88556 17368 88598 17408
rect 88638 17368 88680 17408
rect 88720 17368 88729 17408
rect 92343 17368 92352 17408
rect 92392 17368 92434 17408
rect 92474 17368 92516 17408
rect 92556 17368 92598 17408
rect 92638 17368 92680 17408
rect 92720 17368 92729 17408
rect 96343 17368 96352 17408
rect 96392 17368 96434 17408
rect 96474 17368 96516 17408
rect 96556 17368 96598 17408
rect 96638 17368 96680 17408
rect 96720 17368 96729 17408
rect 0 17348 80 17368
rect 3103 16612 3112 16652
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3480 16612 3489 16652
rect 7103 16612 7112 16652
rect 7152 16612 7194 16652
rect 7234 16612 7276 16652
rect 7316 16612 7358 16652
rect 7398 16612 7440 16652
rect 7480 16612 7489 16652
rect 11103 16612 11112 16652
rect 11152 16612 11194 16652
rect 11234 16612 11276 16652
rect 11316 16612 11358 16652
rect 11398 16612 11440 16652
rect 11480 16612 11489 16652
rect 15103 16612 15112 16652
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15480 16612 15489 16652
rect 19103 16612 19112 16652
rect 19152 16612 19194 16652
rect 19234 16612 19276 16652
rect 19316 16612 19358 16652
rect 19398 16612 19440 16652
rect 19480 16612 19489 16652
rect 23103 16612 23112 16652
rect 23152 16612 23194 16652
rect 23234 16612 23276 16652
rect 23316 16612 23358 16652
rect 23398 16612 23440 16652
rect 23480 16612 23489 16652
rect 27103 16612 27112 16652
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27480 16612 27489 16652
rect 31103 16612 31112 16652
rect 31152 16612 31194 16652
rect 31234 16612 31276 16652
rect 31316 16612 31358 16652
rect 31398 16612 31440 16652
rect 31480 16612 31489 16652
rect 35103 16612 35112 16652
rect 35152 16612 35194 16652
rect 35234 16612 35276 16652
rect 35316 16612 35358 16652
rect 35398 16612 35440 16652
rect 35480 16612 35489 16652
rect 39103 16612 39112 16652
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39480 16612 39489 16652
rect 43103 16612 43112 16652
rect 43152 16612 43194 16652
rect 43234 16612 43276 16652
rect 43316 16612 43358 16652
rect 43398 16612 43440 16652
rect 43480 16612 43489 16652
rect 47103 16612 47112 16652
rect 47152 16612 47194 16652
rect 47234 16612 47276 16652
rect 47316 16612 47358 16652
rect 47398 16612 47440 16652
rect 47480 16612 47489 16652
rect 51103 16612 51112 16652
rect 51152 16612 51194 16652
rect 51234 16612 51276 16652
rect 51316 16612 51358 16652
rect 51398 16612 51440 16652
rect 51480 16612 51489 16652
rect 55103 16612 55112 16652
rect 55152 16612 55194 16652
rect 55234 16612 55276 16652
rect 55316 16612 55358 16652
rect 55398 16612 55440 16652
rect 55480 16612 55489 16652
rect 59103 16612 59112 16652
rect 59152 16612 59194 16652
rect 59234 16612 59276 16652
rect 59316 16612 59358 16652
rect 59398 16612 59440 16652
rect 59480 16612 59489 16652
rect 63103 16612 63112 16652
rect 63152 16612 63194 16652
rect 63234 16612 63276 16652
rect 63316 16612 63358 16652
rect 63398 16612 63440 16652
rect 63480 16612 63489 16652
rect 67103 16612 67112 16652
rect 67152 16612 67194 16652
rect 67234 16612 67276 16652
rect 67316 16612 67358 16652
rect 67398 16612 67440 16652
rect 67480 16612 67489 16652
rect 71103 16612 71112 16652
rect 71152 16612 71194 16652
rect 71234 16612 71276 16652
rect 71316 16612 71358 16652
rect 71398 16612 71440 16652
rect 71480 16612 71489 16652
rect 75103 16612 75112 16652
rect 75152 16612 75194 16652
rect 75234 16612 75276 16652
rect 75316 16612 75358 16652
rect 75398 16612 75440 16652
rect 75480 16612 75489 16652
rect 79103 16612 79112 16652
rect 79152 16612 79194 16652
rect 79234 16612 79276 16652
rect 79316 16612 79358 16652
rect 79398 16612 79440 16652
rect 79480 16612 79489 16652
rect 83103 16612 83112 16652
rect 83152 16612 83194 16652
rect 83234 16612 83276 16652
rect 83316 16612 83358 16652
rect 83398 16612 83440 16652
rect 83480 16612 83489 16652
rect 87103 16612 87112 16652
rect 87152 16612 87194 16652
rect 87234 16612 87276 16652
rect 87316 16612 87358 16652
rect 87398 16612 87440 16652
rect 87480 16612 87489 16652
rect 91103 16612 91112 16652
rect 91152 16612 91194 16652
rect 91234 16612 91276 16652
rect 91316 16612 91358 16652
rect 91398 16612 91440 16652
rect 91480 16612 91489 16652
rect 95103 16612 95112 16652
rect 95152 16612 95194 16652
rect 95234 16612 95276 16652
rect 95316 16612 95358 16652
rect 95398 16612 95440 16652
rect 95480 16612 95489 16652
rect 99103 16612 99112 16652
rect 99152 16612 99194 16652
rect 99234 16612 99276 16652
rect 99316 16612 99358 16652
rect 99398 16612 99440 16652
rect 99480 16612 99489 16652
rect 0 16568 80 16588
rect 0 16528 652 16568
rect 692 16528 701 16568
rect 0 16508 80 16528
rect 86179 16400 86237 16401
rect 71779 16360 71788 16400
rect 71828 16360 73940 16400
rect 83107 16360 83116 16400
rect 83156 16360 83404 16400
rect 83444 16360 83788 16400
rect 83828 16360 83837 16400
rect 86094 16360 86188 16400
rect 86228 16360 86764 16400
rect 86804 16360 92468 16400
rect 73900 16316 73940 16360
rect 86179 16359 86237 16360
rect 92428 16316 92468 16360
rect 73891 16276 73900 16316
rect 73940 16276 74476 16316
rect 74516 16276 77164 16316
rect 77204 16276 80428 16316
rect 80468 16276 80477 16316
rect 80611 16276 80620 16316
rect 80660 16276 81772 16316
rect 81812 16276 83308 16316
rect 83348 16276 84652 16316
rect 84692 16276 84701 16316
rect 86371 16276 86380 16316
rect 86420 16276 86572 16316
rect 86612 16276 88204 16316
rect 88244 16276 89356 16316
rect 89396 16276 90220 16316
rect 90260 16276 90604 16316
rect 90644 16276 90653 16316
rect 92419 16276 92428 16316
rect 92468 16276 95596 16316
rect 95636 16276 95645 16316
rect 73123 16192 73132 16232
rect 73172 16192 74284 16232
rect 74324 16192 86476 16232
rect 86516 16192 86525 16232
rect 76771 16024 76780 16064
rect 76820 16024 77356 16064
rect 77396 16024 77405 16064
rect 81571 16024 81580 16064
rect 81620 16024 81772 16064
rect 81812 16024 82252 16064
rect 82292 16024 82301 16064
rect 4343 15856 4352 15896
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4720 15856 4729 15896
rect 8343 15856 8352 15896
rect 8392 15856 8434 15896
rect 8474 15856 8516 15896
rect 8556 15856 8598 15896
rect 8638 15856 8680 15896
rect 8720 15856 8729 15896
rect 12343 15856 12352 15896
rect 12392 15856 12434 15896
rect 12474 15856 12516 15896
rect 12556 15856 12598 15896
rect 12638 15856 12680 15896
rect 12720 15856 12729 15896
rect 16343 15856 16352 15896
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16720 15856 16729 15896
rect 20343 15856 20352 15896
rect 20392 15856 20434 15896
rect 20474 15856 20516 15896
rect 20556 15856 20598 15896
rect 20638 15856 20680 15896
rect 20720 15856 20729 15896
rect 24343 15856 24352 15896
rect 24392 15856 24434 15896
rect 24474 15856 24516 15896
rect 24556 15856 24598 15896
rect 24638 15856 24680 15896
rect 24720 15856 24729 15896
rect 28343 15856 28352 15896
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28720 15856 28729 15896
rect 32343 15856 32352 15896
rect 32392 15856 32434 15896
rect 32474 15856 32516 15896
rect 32556 15856 32598 15896
rect 32638 15856 32680 15896
rect 32720 15856 32729 15896
rect 36343 15856 36352 15896
rect 36392 15856 36434 15896
rect 36474 15856 36516 15896
rect 36556 15856 36598 15896
rect 36638 15856 36680 15896
rect 36720 15856 36729 15896
rect 40343 15856 40352 15896
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40720 15856 40729 15896
rect 44343 15856 44352 15896
rect 44392 15856 44434 15896
rect 44474 15856 44516 15896
rect 44556 15856 44598 15896
rect 44638 15856 44680 15896
rect 44720 15856 44729 15896
rect 48343 15856 48352 15896
rect 48392 15856 48434 15896
rect 48474 15856 48516 15896
rect 48556 15856 48598 15896
rect 48638 15856 48680 15896
rect 48720 15856 48729 15896
rect 52343 15856 52352 15896
rect 52392 15856 52434 15896
rect 52474 15856 52516 15896
rect 52556 15856 52598 15896
rect 52638 15856 52680 15896
rect 52720 15856 52729 15896
rect 56343 15856 56352 15896
rect 56392 15856 56434 15896
rect 56474 15856 56516 15896
rect 56556 15856 56598 15896
rect 56638 15856 56680 15896
rect 56720 15856 56729 15896
rect 60343 15856 60352 15896
rect 60392 15856 60434 15896
rect 60474 15856 60516 15896
rect 60556 15856 60598 15896
rect 60638 15856 60680 15896
rect 60720 15856 60729 15896
rect 64343 15856 64352 15896
rect 64392 15856 64434 15896
rect 64474 15856 64516 15896
rect 64556 15856 64598 15896
rect 64638 15856 64680 15896
rect 64720 15856 64729 15896
rect 68343 15856 68352 15896
rect 68392 15856 68434 15896
rect 68474 15856 68516 15896
rect 68556 15856 68598 15896
rect 68638 15856 68680 15896
rect 68720 15856 68729 15896
rect 72343 15856 72352 15896
rect 72392 15856 72434 15896
rect 72474 15856 72516 15896
rect 72556 15856 72598 15896
rect 72638 15856 72680 15896
rect 72720 15856 72729 15896
rect 76343 15856 76352 15896
rect 76392 15856 76434 15896
rect 76474 15856 76516 15896
rect 76556 15856 76598 15896
rect 76638 15856 76680 15896
rect 76720 15856 76729 15896
rect 80343 15856 80352 15896
rect 80392 15856 80434 15896
rect 80474 15856 80516 15896
rect 80556 15856 80598 15896
rect 80638 15856 80680 15896
rect 80720 15856 80729 15896
rect 84343 15856 84352 15896
rect 84392 15856 84434 15896
rect 84474 15856 84516 15896
rect 84556 15856 84598 15896
rect 84638 15856 84680 15896
rect 84720 15856 84729 15896
rect 88343 15856 88352 15896
rect 88392 15856 88434 15896
rect 88474 15856 88516 15896
rect 88556 15856 88598 15896
rect 88638 15856 88680 15896
rect 88720 15856 88729 15896
rect 92343 15856 92352 15896
rect 92392 15856 92434 15896
rect 92474 15856 92516 15896
rect 92556 15856 92598 15896
rect 92638 15856 92680 15896
rect 92720 15856 92729 15896
rect 96343 15856 96352 15896
rect 96392 15856 96434 15896
rect 96474 15856 96516 15896
rect 96556 15856 96598 15896
rect 96638 15856 96680 15896
rect 96720 15856 96729 15896
rect 0 15728 80 15748
rect 0 15688 652 15728
rect 692 15688 701 15728
rect 0 15668 80 15688
rect 95491 15520 95500 15560
rect 95540 15520 96076 15560
rect 96116 15520 96556 15560
rect 96596 15520 96844 15560
rect 96884 15520 98036 15560
rect 97996 15476 98036 15520
rect 73699 15436 73708 15476
rect 73748 15436 74092 15476
rect 74132 15436 74476 15476
rect 74516 15436 74860 15476
rect 74900 15436 74909 15476
rect 80227 15436 80236 15476
rect 80276 15436 80716 15476
rect 80756 15436 81100 15476
rect 81140 15436 81388 15476
rect 81428 15436 82540 15476
rect 82580 15436 82589 15476
rect 83011 15436 83020 15476
rect 83060 15436 83404 15476
rect 83444 15436 83884 15476
rect 83924 15436 84172 15476
rect 84212 15436 84221 15476
rect 84547 15436 84556 15476
rect 84596 15436 85036 15476
rect 85076 15436 85420 15476
rect 85460 15436 85804 15476
rect 85844 15436 85853 15476
rect 86179 15436 86188 15476
rect 86228 15436 86380 15476
rect 86420 15436 86572 15476
rect 86612 15436 87052 15476
rect 87092 15436 87436 15476
rect 87476 15436 87485 15476
rect 88291 15436 88300 15476
rect 88340 15436 88684 15476
rect 88724 15436 88733 15476
rect 89059 15436 89068 15476
rect 89108 15436 89452 15476
rect 89492 15436 89836 15476
rect 89876 15436 91084 15476
rect 91124 15436 91948 15476
rect 91988 15436 91997 15476
rect 93859 15436 93868 15476
rect 93908 15436 94252 15476
rect 94292 15436 94636 15476
rect 94676 15436 94924 15476
rect 94964 15436 94973 15476
rect 95971 15436 95980 15476
rect 96020 15436 97228 15476
rect 97268 15436 97708 15476
rect 97748 15436 97757 15476
rect 97987 15436 97996 15476
rect 98036 15436 98380 15476
rect 98420 15436 98429 15476
rect 74860 15308 74900 15436
rect 78787 15352 78796 15392
rect 78836 15352 79180 15392
rect 79220 15352 79372 15392
rect 79412 15352 79660 15392
rect 79700 15352 79709 15392
rect 90883 15308 90941 15309
rect 73891 15268 73900 15308
rect 73940 15268 74380 15308
rect 74420 15268 74429 15308
rect 74860 15268 75340 15308
rect 75380 15268 75820 15308
rect 75860 15268 76204 15308
rect 76244 15268 76588 15308
rect 76628 15268 76637 15308
rect 83971 15268 83980 15308
rect 84020 15268 84268 15308
rect 84308 15268 84317 15308
rect 90798 15268 90892 15308
rect 90932 15268 90941 15308
rect 92227 15268 92236 15308
rect 92276 15268 92716 15308
rect 92756 15268 93388 15308
rect 93428 15268 95020 15308
rect 95060 15268 95069 15308
rect 90883 15267 90941 15268
rect 76963 15184 76972 15224
rect 77012 15184 77356 15224
rect 77396 15184 77740 15224
rect 77780 15184 78124 15224
rect 78164 15184 79756 15224
rect 79796 15184 79805 15224
rect 90499 15184 90508 15224
rect 90548 15184 91084 15224
rect 91124 15184 91564 15224
rect 91604 15184 91756 15224
rect 91796 15184 91805 15224
rect 79756 15140 79796 15184
rect 3103 15100 3112 15140
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3480 15100 3489 15140
rect 7103 15100 7112 15140
rect 7152 15100 7194 15140
rect 7234 15100 7276 15140
rect 7316 15100 7358 15140
rect 7398 15100 7440 15140
rect 7480 15100 7489 15140
rect 11103 15100 11112 15140
rect 11152 15100 11194 15140
rect 11234 15100 11276 15140
rect 11316 15100 11358 15140
rect 11398 15100 11440 15140
rect 11480 15100 11489 15140
rect 15103 15100 15112 15140
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15480 15100 15489 15140
rect 19103 15100 19112 15140
rect 19152 15100 19194 15140
rect 19234 15100 19276 15140
rect 19316 15100 19358 15140
rect 19398 15100 19440 15140
rect 19480 15100 19489 15140
rect 23103 15100 23112 15140
rect 23152 15100 23194 15140
rect 23234 15100 23276 15140
rect 23316 15100 23358 15140
rect 23398 15100 23440 15140
rect 23480 15100 23489 15140
rect 27103 15100 27112 15140
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27480 15100 27489 15140
rect 31103 15100 31112 15140
rect 31152 15100 31194 15140
rect 31234 15100 31276 15140
rect 31316 15100 31358 15140
rect 31398 15100 31440 15140
rect 31480 15100 31489 15140
rect 35103 15100 35112 15140
rect 35152 15100 35194 15140
rect 35234 15100 35276 15140
rect 35316 15100 35358 15140
rect 35398 15100 35440 15140
rect 35480 15100 35489 15140
rect 39103 15100 39112 15140
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39480 15100 39489 15140
rect 43103 15100 43112 15140
rect 43152 15100 43194 15140
rect 43234 15100 43276 15140
rect 43316 15100 43358 15140
rect 43398 15100 43440 15140
rect 43480 15100 43489 15140
rect 47103 15100 47112 15140
rect 47152 15100 47194 15140
rect 47234 15100 47276 15140
rect 47316 15100 47358 15140
rect 47398 15100 47440 15140
rect 47480 15100 47489 15140
rect 51103 15100 51112 15140
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51480 15100 51489 15140
rect 55103 15100 55112 15140
rect 55152 15100 55194 15140
rect 55234 15100 55276 15140
rect 55316 15100 55358 15140
rect 55398 15100 55440 15140
rect 55480 15100 55489 15140
rect 59103 15100 59112 15140
rect 59152 15100 59194 15140
rect 59234 15100 59276 15140
rect 59316 15100 59358 15140
rect 59398 15100 59440 15140
rect 59480 15100 59489 15140
rect 63103 15100 63112 15140
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63480 15100 63489 15140
rect 67103 15100 67112 15140
rect 67152 15100 67194 15140
rect 67234 15100 67276 15140
rect 67316 15100 67358 15140
rect 67398 15100 67440 15140
rect 67480 15100 67489 15140
rect 76867 15100 76876 15140
rect 76916 15100 77836 15140
rect 77876 15100 78604 15140
rect 78644 15100 78653 15140
rect 79756 15100 80428 15140
rect 80468 15100 80477 15140
rect 92419 15100 92428 15140
rect 92468 15100 92812 15140
rect 92852 15100 94156 15140
rect 94196 15100 94205 15140
rect 97027 15100 97036 15140
rect 97076 15100 97516 15140
rect 97556 15100 97565 15140
rect 835 14932 844 14972
rect 884 14932 1420 14972
rect 1460 14932 1469 14972
rect 0 14888 80 14908
rect 0 14848 652 14888
rect 692 14848 701 14888
rect 0 14828 80 14848
rect 1987 14764 1996 14804
rect 2036 14764 70636 14804
rect 70676 14764 70685 14804
rect 71299 14680 71308 14720
rect 71348 14680 72748 14720
rect 72788 14680 73036 14720
rect 73076 14680 73516 14720
rect 73556 14680 73900 14720
rect 73940 14680 73949 14720
rect 74179 14680 74188 14720
rect 74228 14680 74860 14720
rect 74900 14680 75244 14720
rect 75284 14680 75820 14720
rect 75860 14680 76108 14720
rect 76148 14680 76157 14720
rect 94147 14680 94156 14720
rect 94196 14680 94636 14720
rect 94676 14680 94685 14720
rect 72835 14512 72844 14552
rect 72884 14512 73100 14552
rect 92803 14512 92812 14552
rect 92852 14512 93100 14552
rect 93140 14512 93149 14552
rect 97123 14512 97132 14552
rect 97172 14512 97804 14552
rect 97844 14512 97853 14552
rect 73060 14468 73100 14512
rect 73060 14428 74188 14468
rect 74228 14428 74237 14468
rect 4343 14344 4352 14384
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4720 14344 4729 14384
rect 8343 14344 8352 14384
rect 8392 14344 8434 14384
rect 8474 14344 8516 14384
rect 8556 14344 8598 14384
rect 8638 14344 8680 14384
rect 8720 14344 8729 14384
rect 12343 14344 12352 14384
rect 12392 14344 12434 14384
rect 12474 14344 12516 14384
rect 12556 14344 12598 14384
rect 12638 14344 12680 14384
rect 12720 14344 12729 14384
rect 16343 14344 16352 14384
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16720 14344 16729 14384
rect 20343 14344 20352 14384
rect 20392 14344 20434 14384
rect 20474 14344 20516 14384
rect 20556 14344 20598 14384
rect 20638 14344 20680 14384
rect 20720 14344 20729 14384
rect 24343 14344 24352 14384
rect 24392 14344 24434 14384
rect 24474 14344 24516 14384
rect 24556 14344 24598 14384
rect 24638 14344 24680 14384
rect 24720 14344 24729 14384
rect 28343 14344 28352 14384
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28720 14344 28729 14384
rect 32343 14344 32352 14384
rect 32392 14344 32434 14384
rect 32474 14344 32516 14384
rect 32556 14344 32598 14384
rect 32638 14344 32680 14384
rect 32720 14344 32729 14384
rect 36343 14344 36352 14384
rect 36392 14344 36434 14384
rect 36474 14344 36516 14384
rect 36556 14344 36598 14384
rect 36638 14344 36680 14384
rect 36720 14344 36729 14384
rect 40343 14344 40352 14384
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40720 14344 40729 14384
rect 44343 14344 44352 14384
rect 44392 14344 44434 14384
rect 44474 14344 44516 14384
rect 44556 14344 44598 14384
rect 44638 14344 44680 14384
rect 44720 14344 44729 14384
rect 48343 14344 48352 14384
rect 48392 14344 48434 14384
rect 48474 14344 48516 14384
rect 48556 14344 48598 14384
rect 48638 14344 48680 14384
rect 48720 14344 48729 14384
rect 52343 14344 52352 14384
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52720 14344 52729 14384
rect 56343 14344 56352 14384
rect 56392 14344 56434 14384
rect 56474 14344 56516 14384
rect 56556 14344 56598 14384
rect 56638 14344 56680 14384
rect 56720 14344 56729 14384
rect 60343 14344 60352 14384
rect 60392 14344 60434 14384
rect 60474 14344 60516 14384
rect 60556 14344 60598 14384
rect 60638 14344 60680 14384
rect 60720 14344 60729 14384
rect 64343 14344 64352 14384
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64720 14344 64729 14384
rect 68343 14344 68352 14384
rect 68392 14344 68434 14384
rect 68474 14344 68516 14384
rect 68556 14344 68598 14384
rect 68638 14344 68680 14384
rect 68720 14344 68729 14384
rect 0 14048 80 14068
rect 0 14008 652 14048
rect 692 14008 701 14048
rect 70531 14008 70540 14048
rect 70580 14008 70828 14048
rect 70868 14008 73132 14048
rect 73172 14008 73181 14048
rect 0 13988 80 14008
rect 1219 13924 1228 13964
rect 1268 13924 1804 13964
rect 1844 13924 1853 13964
rect 70723 13924 70732 13964
rect 70772 13924 71308 13964
rect 71348 13924 71357 13964
rect 71395 13840 71404 13880
rect 71444 13840 73516 13880
rect 73556 13840 73565 13880
rect 79075 13840 79084 13880
rect 79124 13840 79756 13880
rect 79796 13840 79805 13880
rect 70627 13756 70636 13796
rect 70676 13756 73132 13796
rect 73172 13756 73181 13796
rect 71011 13672 71020 13712
rect 71060 13672 72652 13712
rect 72692 13672 72701 13712
rect 80515 13672 80524 13712
rect 80564 13672 80573 13712
rect 96556 13672 98380 13712
rect 98420 13672 98764 13712
rect 98804 13672 98813 13712
rect 3103 13588 3112 13628
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3480 13588 3489 13628
rect 7103 13588 7112 13628
rect 7152 13588 7194 13628
rect 7234 13588 7276 13628
rect 7316 13588 7358 13628
rect 7398 13588 7440 13628
rect 7480 13588 7489 13628
rect 11103 13588 11112 13628
rect 11152 13588 11194 13628
rect 11234 13588 11276 13628
rect 11316 13588 11358 13628
rect 11398 13588 11440 13628
rect 11480 13588 11489 13628
rect 15103 13588 15112 13628
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15480 13588 15489 13628
rect 19103 13588 19112 13628
rect 19152 13588 19194 13628
rect 19234 13588 19276 13628
rect 19316 13588 19358 13628
rect 19398 13588 19440 13628
rect 19480 13588 19489 13628
rect 23103 13588 23112 13628
rect 23152 13588 23194 13628
rect 23234 13588 23276 13628
rect 23316 13588 23358 13628
rect 23398 13588 23440 13628
rect 23480 13588 23489 13628
rect 27103 13588 27112 13628
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27480 13588 27489 13628
rect 31103 13588 31112 13628
rect 31152 13588 31194 13628
rect 31234 13588 31276 13628
rect 31316 13588 31358 13628
rect 31398 13588 31440 13628
rect 31480 13588 31489 13628
rect 35103 13588 35112 13628
rect 35152 13588 35194 13628
rect 35234 13588 35276 13628
rect 35316 13588 35358 13628
rect 35398 13588 35440 13628
rect 35480 13588 35489 13628
rect 39103 13588 39112 13628
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39480 13588 39489 13628
rect 43103 13588 43112 13628
rect 43152 13588 43194 13628
rect 43234 13588 43276 13628
rect 43316 13588 43358 13628
rect 43398 13588 43440 13628
rect 43480 13588 43489 13628
rect 47103 13588 47112 13628
rect 47152 13588 47194 13628
rect 47234 13588 47276 13628
rect 47316 13588 47358 13628
rect 47398 13588 47440 13628
rect 47480 13588 47489 13628
rect 51103 13588 51112 13628
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51480 13588 51489 13628
rect 55103 13588 55112 13628
rect 55152 13588 55194 13628
rect 55234 13588 55276 13628
rect 55316 13588 55358 13628
rect 55398 13588 55440 13628
rect 55480 13588 55489 13628
rect 59103 13588 59112 13628
rect 59152 13588 59194 13628
rect 59234 13588 59276 13628
rect 59316 13588 59358 13628
rect 59398 13588 59440 13628
rect 59480 13588 59489 13628
rect 63103 13588 63112 13628
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63480 13588 63489 13628
rect 67103 13588 67112 13628
rect 67152 13588 67194 13628
rect 67234 13588 67276 13628
rect 67316 13588 67358 13628
rect 67398 13588 67440 13628
rect 67480 13588 67489 13628
rect 70051 13588 70060 13628
rect 70100 13588 73100 13628
rect 74275 13588 74284 13628
rect 74324 13588 74668 13628
rect 74708 13588 74717 13628
rect 73060 13544 73100 13588
rect 70924 13504 72844 13544
rect 72884 13504 72893 13544
rect 73060 13504 73228 13544
rect 73268 13504 73277 13544
rect 70924 13460 70964 13504
rect 80524 13460 80564 13672
rect 82051 13588 82060 13628
rect 82100 13588 82109 13628
rect 70915 13420 70924 13460
rect 70964 13420 70973 13460
rect 71299 13420 71308 13460
rect 71348 13420 72415 13460
rect 72455 13420 72464 13460
rect 72556 13420 73100 13460
rect 79896 13420 79905 13460
rect 79945 13420 80564 13460
rect 82060 13460 82100 13588
rect 90883 13460 90941 13461
rect 82060 13420 82305 13460
rect 82345 13420 82354 13460
rect 90406 13420 90415 13460
rect 90455 13420 90892 13460
rect 90932 13420 90941 13460
rect 72451 13376 72509 13377
rect 72556 13376 72596 13420
rect 835 13336 844 13376
rect 884 13336 1612 13376
rect 1652 13336 1661 13376
rect 71203 13336 71212 13376
rect 71252 13336 72305 13376
rect 72345 13336 72354 13376
rect 72451 13336 72460 13376
rect 72500 13336 72596 13376
rect 73060 13376 73100 13420
rect 90883 13419 90941 13420
rect 96556 13376 96596 13672
rect 97896 13420 97905 13460
rect 97945 13420 98668 13460
rect 98708 13420 98717 13460
rect 73060 13336 96596 13376
rect 96696 13336 96705 13376
rect 96745 13336 96940 13376
rect 96980 13336 96989 13376
rect 72451 13335 72509 13336
rect 71875 13292 71933 13293
rect 71107 13252 71116 13292
rect 71156 13252 71884 13292
rect 71924 13252 71933 13292
rect 71875 13251 71933 13252
rect 0 13208 80 13228
rect 0 13168 652 13208
rect 692 13168 701 13208
rect 69859 13168 69868 13208
rect 69908 13168 70348 13208
rect 70388 13168 70732 13208
rect 70772 13168 70781 13208
rect 0 13148 80 13168
rect 4343 12832 4352 12872
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4720 12832 4729 12872
rect 8343 12832 8352 12872
rect 8392 12832 8434 12872
rect 8474 12832 8516 12872
rect 8556 12832 8598 12872
rect 8638 12832 8680 12872
rect 8720 12832 8729 12872
rect 12343 12832 12352 12872
rect 12392 12832 12434 12872
rect 12474 12832 12516 12872
rect 12556 12832 12598 12872
rect 12638 12832 12680 12872
rect 12720 12832 12729 12872
rect 16343 12832 16352 12872
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16720 12832 16729 12872
rect 20343 12832 20352 12872
rect 20392 12832 20434 12872
rect 20474 12832 20516 12872
rect 20556 12832 20598 12872
rect 20638 12832 20680 12872
rect 20720 12832 20729 12872
rect 24343 12832 24352 12872
rect 24392 12832 24434 12872
rect 24474 12832 24516 12872
rect 24556 12832 24598 12872
rect 24638 12832 24680 12872
rect 24720 12832 24729 12872
rect 28343 12832 28352 12872
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28720 12832 28729 12872
rect 32343 12832 32352 12872
rect 32392 12832 32434 12872
rect 32474 12832 32516 12872
rect 32556 12832 32598 12872
rect 32638 12832 32680 12872
rect 32720 12832 32729 12872
rect 36343 12832 36352 12872
rect 36392 12832 36434 12872
rect 36474 12832 36516 12872
rect 36556 12832 36598 12872
rect 36638 12832 36680 12872
rect 36720 12832 36729 12872
rect 40343 12832 40352 12872
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40720 12832 40729 12872
rect 44343 12832 44352 12872
rect 44392 12832 44434 12872
rect 44474 12832 44516 12872
rect 44556 12832 44598 12872
rect 44638 12832 44680 12872
rect 44720 12832 44729 12872
rect 48343 12832 48352 12872
rect 48392 12832 48434 12872
rect 48474 12832 48516 12872
rect 48556 12832 48598 12872
rect 48638 12832 48680 12872
rect 48720 12832 48729 12872
rect 52343 12832 52352 12872
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52720 12832 52729 12872
rect 56343 12832 56352 12872
rect 56392 12832 56434 12872
rect 56474 12832 56516 12872
rect 56556 12832 56598 12872
rect 56638 12832 56680 12872
rect 56720 12832 56729 12872
rect 60343 12832 60352 12872
rect 60392 12832 60434 12872
rect 60474 12832 60516 12872
rect 60556 12832 60598 12872
rect 60638 12832 60680 12872
rect 60720 12832 60729 12872
rect 64343 12832 64352 12872
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64720 12832 64729 12872
rect 68343 12832 68352 12872
rect 68392 12832 68434 12872
rect 68474 12832 68516 12872
rect 68556 12832 68598 12872
rect 68638 12832 68680 12872
rect 68720 12832 68729 12872
rect 0 12368 80 12388
rect 0 12328 652 12368
rect 692 12328 701 12368
rect 0 12308 80 12328
rect 3103 12076 3112 12116
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3480 12076 3489 12116
rect 7103 12076 7112 12116
rect 7152 12076 7194 12116
rect 7234 12076 7276 12116
rect 7316 12076 7358 12116
rect 7398 12076 7440 12116
rect 7480 12076 7489 12116
rect 11103 12076 11112 12116
rect 11152 12076 11194 12116
rect 11234 12076 11276 12116
rect 11316 12076 11358 12116
rect 11398 12076 11440 12116
rect 11480 12076 11489 12116
rect 15103 12076 15112 12116
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15480 12076 15489 12116
rect 19103 12076 19112 12116
rect 19152 12076 19194 12116
rect 19234 12076 19276 12116
rect 19316 12076 19358 12116
rect 19398 12076 19440 12116
rect 19480 12076 19489 12116
rect 23103 12076 23112 12116
rect 23152 12076 23194 12116
rect 23234 12076 23276 12116
rect 23316 12076 23358 12116
rect 23398 12076 23440 12116
rect 23480 12076 23489 12116
rect 27103 12076 27112 12116
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27480 12076 27489 12116
rect 31103 12076 31112 12116
rect 31152 12076 31194 12116
rect 31234 12076 31276 12116
rect 31316 12076 31358 12116
rect 31398 12076 31440 12116
rect 31480 12076 31489 12116
rect 35103 12076 35112 12116
rect 35152 12076 35194 12116
rect 35234 12076 35276 12116
rect 35316 12076 35358 12116
rect 35398 12076 35440 12116
rect 35480 12076 35489 12116
rect 39103 12076 39112 12116
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39480 12076 39489 12116
rect 43103 12076 43112 12116
rect 43152 12076 43194 12116
rect 43234 12076 43276 12116
rect 43316 12076 43358 12116
rect 43398 12076 43440 12116
rect 43480 12076 43489 12116
rect 47103 12076 47112 12116
rect 47152 12076 47194 12116
rect 47234 12076 47276 12116
rect 47316 12076 47358 12116
rect 47398 12076 47440 12116
rect 47480 12076 47489 12116
rect 51103 12076 51112 12116
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51480 12076 51489 12116
rect 55103 12076 55112 12116
rect 55152 12076 55194 12116
rect 55234 12076 55276 12116
rect 55316 12076 55358 12116
rect 55398 12076 55440 12116
rect 55480 12076 55489 12116
rect 59103 12076 59112 12116
rect 59152 12076 59194 12116
rect 59234 12076 59276 12116
rect 59316 12076 59358 12116
rect 59398 12076 59440 12116
rect 59480 12076 59489 12116
rect 63103 12076 63112 12116
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63480 12076 63489 12116
rect 67103 12076 67112 12116
rect 67152 12076 67194 12116
rect 67234 12076 67276 12116
rect 67316 12076 67358 12116
rect 67398 12076 67440 12116
rect 67480 12076 67489 12116
rect 0 11528 80 11548
rect 0 11488 652 11528
rect 692 11488 701 11528
rect 0 11468 80 11488
rect 4343 11320 4352 11360
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4720 11320 4729 11360
rect 8343 11320 8352 11360
rect 8392 11320 8434 11360
rect 8474 11320 8516 11360
rect 8556 11320 8598 11360
rect 8638 11320 8680 11360
rect 8720 11320 8729 11360
rect 12343 11320 12352 11360
rect 12392 11320 12434 11360
rect 12474 11320 12516 11360
rect 12556 11320 12598 11360
rect 12638 11320 12680 11360
rect 12720 11320 12729 11360
rect 16343 11320 16352 11360
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16720 11320 16729 11360
rect 20343 11320 20352 11360
rect 20392 11320 20434 11360
rect 20474 11320 20516 11360
rect 20556 11320 20598 11360
rect 20638 11320 20680 11360
rect 20720 11320 20729 11360
rect 24343 11320 24352 11360
rect 24392 11320 24434 11360
rect 24474 11320 24516 11360
rect 24556 11320 24598 11360
rect 24638 11320 24680 11360
rect 24720 11320 24729 11360
rect 28343 11320 28352 11360
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28720 11320 28729 11360
rect 32343 11320 32352 11360
rect 32392 11320 32434 11360
rect 32474 11320 32516 11360
rect 32556 11320 32598 11360
rect 32638 11320 32680 11360
rect 32720 11320 32729 11360
rect 36343 11320 36352 11360
rect 36392 11320 36434 11360
rect 36474 11320 36516 11360
rect 36556 11320 36598 11360
rect 36638 11320 36680 11360
rect 36720 11320 36729 11360
rect 40343 11320 40352 11360
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40720 11320 40729 11360
rect 44343 11320 44352 11360
rect 44392 11320 44434 11360
rect 44474 11320 44516 11360
rect 44556 11320 44598 11360
rect 44638 11320 44680 11360
rect 44720 11320 44729 11360
rect 48343 11320 48352 11360
rect 48392 11320 48434 11360
rect 48474 11320 48516 11360
rect 48556 11320 48598 11360
rect 48638 11320 48680 11360
rect 48720 11320 48729 11360
rect 52343 11320 52352 11360
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52720 11320 52729 11360
rect 56343 11320 56352 11360
rect 56392 11320 56434 11360
rect 56474 11320 56516 11360
rect 56556 11320 56598 11360
rect 56638 11320 56680 11360
rect 56720 11320 56729 11360
rect 60343 11320 60352 11360
rect 60392 11320 60434 11360
rect 60474 11320 60516 11360
rect 60556 11320 60598 11360
rect 60638 11320 60680 11360
rect 60720 11320 60729 11360
rect 64343 11320 64352 11360
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64720 11320 64729 11360
rect 68343 11320 68352 11360
rect 68392 11320 68434 11360
rect 68474 11320 68516 11360
rect 68556 11320 68598 11360
rect 68638 11320 68680 11360
rect 68720 11320 68729 11360
rect 643 10732 652 10772
rect 692 10732 701 10772
rect 0 10688 80 10708
rect 652 10688 692 10732
rect 0 10648 692 10688
rect 0 10628 80 10648
rect 3103 10564 3112 10604
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3480 10564 3489 10604
rect 7103 10564 7112 10604
rect 7152 10564 7194 10604
rect 7234 10564 7276 10604
rect 7316 10564 7358 10604
rect 7398 10564 7440 10604
rect 7480 10564 7489 10604
rect 11103 10564 11112 10604
rect 11152 10564 11194 10604
rect 11234 10564 11276 10604
rect 11316 10564 11358 10604
rect 11398 10564 11440 10604
rect 11480 10564 11489 10604
rect 15103 10564 15112 10604
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15480 10564 15489 10604
rect 19103 10564 19112 10604
rect 19152 10564 19194 10604
rect 19234 10564 19276 10604
rect 19316 10564 19358 10604
rect 19398 10564 19440 10604
rect 19480 10564 19489 10604
rect 23103 10564 23112 10604
rect 23152 10564 23194 10604
rect 23234 10564 23276 10604
rect 23316 10564 23358 10604
rect 23398 10564 23440 10604
rect 23480 10564 23489 10604
rect 27103 10564 27112 10604
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27480 10564 27489 10604
rect 31103 10564 31112 10604
rect 31152 10564 31194 10604
rect 31234 10564 31276 10604
rect 31316 10564 31358 10604
rect 31398 10564 31440 10604
rect 31480 10564 31489 10604
rect 35103 10564 35112 10604
rect 35152 10564 35194 10604
rect 35234 10564 35276 10604
rect 35316 10564 35358 10604
rect 35398 10564 35440 10604
rect 35480 10564 35489 10604
rect 39103 10564 39112 10604
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39480 10564 39489 10604
rect 43103 10564 43112 10604
rect 43152 10564 43194 10604
rect 43234 10564 43276 10604
rect 43316 10564 43358 10604
rect 43398 10564 43440 10604
rect 43480 10564 43489 10604
rect 47103 10564 47112 10604
rect 47152 10564 47194 10604
rect 47234 10564 47276 10604
rect 47316 10564 47358 10604
rect 47398 10564 47440 10604
rect 47480 10564 47489 10604
rect 51103 10564 51112 10604
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51480 10564 51489 10604
rect 55103 10564 55112 10604
rect 55152 10564 55194 10604
rect 55234 10564 55276 10604
rect 55316 10564 55358 10604
rect 55398 10564 55440 10604
rect 55480 10564 55489 10604
rect 59103 10564 59112 10604
rect 59152 10564 59194 10604
rect 59234 10564 59276 10604
rect 59316 10564 59358 10604
rect 59398 10564 59440 10604
rect 59480 10564 59489 10604
rect 63103 10564 63112 10604
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63480 10564 63489 10604
rect 67103 10564 67112 10604
rect 67152 10564 67194 10604
rect 67234 10564 67276 10604
rect 67316 10564 67358 10604
rect 67398 10564 67440 10604
rect 67480 10564 67489 10604
rect 835 10480 844 10520
rect 884 10480 1420 10520
rect 1460 10480 1469 10520
rect 1219 10228 1228 10268
rect 1268 10228 1612 10268
rect 1652 10228 1661 10268
rect 0 9848 80 9868
rect 0 9808 652 9848
rect 692 9808 701 9848
rect 4343 9808 4352 9848
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4720 9808 4729 9848
rect 8343 9808 8352 9848
rect 8392 9808 8434 9848
rect 8474 9808 8516 9848
rect 8556 9808 8598 9848
rect 8638 9808 8680 9848
rect 8720 9808 8729 9848
rect 12343 9808 12352 9848
rect 12392 9808 12434 9848
rect 12474 9808 12516 9848
rect 12556 9808 12598 9848
rect 12638 9808 12680 9848
rect 12720 9808 12729 9848
rect 16343 9808 16352 9848
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16720 9808 16729 9848
rect 20343 9808 20352 9848
rect 20392 9808 20434 9848
rect 20474 9808 20516 9848
rect 20556 9808 20598 9848
rect 20638 9808 20680 9848
rect 20720 9808 20729 9848
rect 24343 9808 24352 9848
rect 24392 9808 24434 9848
rect 24474 9808 24516 9848
rect 24556 9808 24598 9848
rect 24638 9808 24680 9848
rect 24720 9808 24729 9848
rect 28343 9808 28352 9848
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28720 9808 28729 9848
rect 32343 9808 32352 9848
rect 32392 9808 32434 9848
rect 32474 9808 32516 9848
rect 32556 9808 32598 9848
rect 32638 9808 32680 9848
rect 32720 9808 32729 9848
rect 36343 9808 36352 9848
rect 36392 9808 36434 9848
rect 36474 9808 36516 9848
rect 36556 9808 36598 9848
rect 36638 9808 36680 9848
rect 36720 9808 36729 9848
rect 40343 9808 40352 9848
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40720 9808 40729 9848
rect 44343 9808 44352 9848
rect 44392 9808 44434 9848
rect 44474 9808 44516 9848
rect 44556 9808 44598 9848
rect 44638 9808 44680 9848
rect 44720 9808 44729 9848
rect 48343 9808 48352 9848
rect 48392 9808 48434 9848
rect 48474 9808 48516 9848
rect 48556 9808 48598 9848
rect 48638 9808 48680 9848
rect 48720 9808 48729 9848
rect 52343 9808 52352 9848
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52720 9808 52729 9848
rect 56343 9808 56352 9848
rect 56392 9808 56434 9848
rect 56474 9808 56516 9848
rect 56556 9808 56598 9848
rect 56638 9808 56680 9848
rect 56720 9808 56729 9848
rect 60343 9808 60352 9848
rect 60392 9808 60434 9848
rect 60474 9808 60516 9848
rect 60556 9808 60598 9848
rect 60638 9808 60680 9848
rect 60720 9808 60729 9848
rect 64343 9808 64352 9848
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64720 9808 64729 9848
rect 68343 9808 68352 9848
rect 68392 9808 68434 9848
rect 68474 9808 68516 9848
rect 68556 9808 68598 9848
rect 68638 9808 68680 9848
rect 68720 9808 68729 9848
rect 0 9788 80 9808
rect 3103 9052 3112 9092
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3480 9052 3489 9092
rect 7103 9052 7112 9092
rect 7152 9052 7194 9092
rect 7234 9052 7276 9092
rect 7316 9052 7358 9092
rect 7398 9052 7440 9092
rect 7480 9052 7489 9092
rect 11103 9052 11112 9092
rect 11152 9052 11194 9092
rect 11234 9052 11276 9092
rect 11316 9052 11358 9092
rect 11398 9052 11440 9092
rect 11480 9052 11489 9092
rect 15103 9052 15112 9092
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15480 9052 15489 9092
rect 19103 9052 19112 9092
rect 19152 9052 19194 9092
rect 19234 9052 19276 9092
rect 19316 9052 19358 9092
rect 19398 9052 19440 9092
rect 19480 9052 19489 9092
rect 23103 9052 23112 9092
rect 23152 9052 23194 9092
rect 23234 9052 23276 9092
rect 23316 9052 23358 9092
rect 23398 9052 23440 9092
rect 23480 9052 23489 9092
rect 27103 9052 27112 9092
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27480 9052 27489 9092
rect 31103 9052 31112 9092
rect 31152 9052 31194 9092
rect 31234 9052 31276 9092
rect 31316 9052 31358 9092
rect 31398 9052 31440 9092
rect 31480 9052 31489 9092
rect 35103 9052 35112 9092
rect 35152 9052 35194 9092
rect 35234 9052 35276 9092
rect 35316 9052 35358 9092
rect 35398 9052 35440 9092
rect 35480 9052 35489 9092
rect 39103 9052 39112 9092
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39480 9052 39489 9092
rect 43103 9052 43112 9092
rect 43152 9052 43194 9092
rect 43234 9052 43276 9092
rect 43316 9052 43358 9092
rect 43398 9052 43440 9092
rect 43480 9052 43489 9092
rect 47103 9052 47112 9092
rect 47152 9052 47194 9092
rect 47234 9052 47276 9092
rect 47316 9052 47358 9092
rect 47398 9052 47440 9092
rect 47480 9052 47489 9092
rect 51103 9052 51112 9092
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51480 9052 51489 9092
rect 55103 9052 55112 9092
rect 55152 9052 55194 9092
rect 55234 9052 55276 9092
rect 55316 9052 55358 9092
rect 55398 9052 55440 9092
rect 55480 9052 55489 9092
rect 59103 9052 59112 9092
rect 59152 9052 59194 9092
rect 59234 9052 59276 9092
rect 59316 9052 59358 9092
rect 59398 9052 59440 9092
rect 59480 9052 59489 9092
rect 63103 9052 63112 9092
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63480 9052 63489 9092
rect 67103 9052 67112 9092
rect 67152 9052 67194 9092
rect 67234 9052 67276 9092
rect 67316 9052 67358 9092
rect 67398 9052 67440 9092
rect 67480 9052 67489 9092
rect 0 9008 80 9028
rect 0 8968 652 9008
rect 692 8968 701 9008
rect 0 8948 80 8968
rect 739 8800 748 8840
rect 788 8800 1516 8840
rect 1556 8800 1565 8840
rect 4343 8296 4352 8336
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4720 8296 4729 8336
rect 8343 8296 8352 8336
rect 8392 8296 8434 8336
rect 8474 8296 8516 8336
rect 8556 8296 8598 8336
rect 8638 8296 8680 8336
rect 8720 8296 8729 8336
rect 12343 8296 12352 8336
rect 12392 8296 12434 8336
rect 12474 8296 12516 8336
rect 12556 8296 12598 8336
rect 12638 8296 12680 8336
rect 12720 8296 12729 8336
rect 16343 8296 16352 8336
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16720 8296 16729 8336
rect 20343 8296 20352 8336
rect 20392 8296 20434 8336
rect 20474 8296 20516 8336
rect 20556 8296 20598 8336
rect 20638 8296 20680 8336
rect 20720 8296 20729 8336
rect 24343 8296 24352 8336
rect 24392 8296 24434 8336
rect 24474 8296 24516 8336
rect 24556 8296 24598 8336
rect 24638 8296 24680 8336
rect 24720 8296 24729 8336
rect 28343 8296 28352 8336
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28720 8296 28729 8336
rect 32343 8296 32352 8336
rect 32392 8296 32434 8336
rect 32474 8296 32516 8336
rect 32556 8296 32598 8336
rect 32638 8296 32680 8336
rect 32720 8296 32729 8336
rect 36343 8296 36352 8336
rect 36392 8296 36434 8336
rect 36474 8296 36516 8336
rect 36556 8296 36598 8336
rect 36638 8296 36680 8336
rect 36720 8296 36729 8336
rect 40343 8296 40352 8336
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40720 8296 40729 8336
rect 44343 8296 44352 8336
rect 44392 8296 44434 8336
rect 44474 8296 44516 8336
rect 44556 8296 44598 8336
rect 44638 8296 44680 8336
rect 44720 8296 44729 8336
rect 48343 8296 48352 8336
rect 48392 8296 48434 8336
rect 48474 8296 48516 8336
rect 48556 8296 48598 8336
rect 48638 8296 48680 8336
rect 48720 8296 48729 8336
rect 52343 8296 52352 8336
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52720 8296 52729 8336
rect 56343 8296 56352 8336
rect 56392 8296 56434 8336
rect 56474 8296 56516 8336
rect 56556 8296 56598 8336
rect 56638 8296 56680 8336
rect 56720 8296 56729 8336
rect 60343 8296 60352 8336
rect 60392 8296 60434 8336
rect 60474 8296 60516 8336
rect 60556 8296 60598 8336
rect 60638 8296 60680 8336
rect 60720 8296 60729 8336
rect 64343 8296 64352 8336
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64720 8296 64729 8336
rect 68343 8296 68352 8336
rect 68392 8296 68434 8336
rect 68474 8296 68516 8336
rect 68556 8296 68598 8336
rect 68638 8296 68680 8336
rect 68720 8296 68729 8336
rect 0 8168 80 8188
rect 0 8128 652 8168
rect 692 8128 701 8168
rect 0 8108 80 8128
rect 71011 7876 71020 7916
rect 71060 7876 72705 7916
rect 72745 7876 72754 7916
rect 93763 7832 93821 7833
rect 71395 7792 71404 7832
rect 71444 7792 72305 7832
rect 72345 7792 72354 7832
rect 72406 7792 72415 7832
rect 72455 7792 72500 7832
rect 84406 7792 84415 7832
rect 84455 7792 85324 7832
rect 85364 7792 85373 7832
rect 93763 7792 93772 7832
rect 93812 7792 93905 7832
rect 93945 7792 93954 7832
rect 72460 7748 72500 7792
rect 93763 7791 93821 7792
rect 71491 7708 71500 7748
rect 71540 7708 72500 7748
rect 89606 7708 89615 7748
rect 89655 7708 90508 7748
rect 90548 7708 90557 7748
rect 90979 7708 90988 7748
rect 91028 7708 91215 7748
rect 91255 7708 91264 7748
rect 75606 7624 75615 7664
rect 75655 7624 76204 7664
rect 76244 7624 76253 7664
rect 78406 7624 78415 7664
rect 78455 7624 79276 7664
rect 79316 7624 79325 7664
rect 83606 7624 83615 7664
rect 83655 7624 84172 7664
rect 84212 7624 84221 7664
rect 90806 7624 90815 7664
rect 90855 7624 91756 7664
rect 91796 7624 91805 7664
rect 97496 7624 97505 7664
rect 97545 7624 97708 7664
rect 97748 7624 97757 7664
rect 3103 7540 3112 7580
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3480 7540 3489 7580
rect 7103 7540 7112 7580
rect 7152 7540 7194 7580
rect 7234 7540 7276 7580
rect 7316 7540 7358 7580
rect 7398 7540 7440 7580
rect 7480 7540 7489 7580
rect 11103 7540 11112 7580
rect 11152 7540 11194 7580
rect 11234 7540 11276 7580
rect 11316 7540 11358 7580
rect 11398 7540 11440 7580
rect 11480 7540 11489 7580
rect 15103 7540 15112 7580
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15480 7540 15489 7580
rect 19103 7540 19112 7580
rect 19152 7540 19194 7580
rect 19234 7540 19276 7580
rect 19316 7540 19358 7580
rect 19398 7540 19440 7580
rect 19480 7540 19489 7580
rect 23103 7540 23112 7580
rect 23152 7540 23194 7580
rect 23234 7540 23276 7580
rect 23316 7540 23358 7580
rect 23398 7540 23440 7580
rect 23480 7540 23489 7580
rect 27103 7540 27112 7580
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27480 7540 27489 7580
rect 31103 7540 31112 7580
rect 31152 7540 31194 7580
rect 31234 7540 31276 7580
rect 31316 7540 31358 7580
rect 31398 7540 31440 7580
rect 31480 7540 31489 7580
rect 35103 7540 35112 7580
rect 35152 7540 35194 7580
rect 35234 7540 35276 7580
rect 35316 7540 35358 7580
rect 35398 7540 35440 7580
rect 35480 7540 35489 7580
rect 39103 7540 39112 7580
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39480 7540 39489 7580
rect 43103 7540 43112 7580
rect 43152 7540 43194 7580
rect 43234 7540 43276 7580
rect 43316 7540 43358 7580
rect 43398 7540 43440 7580
rect 43480 7540 43489 7580
rect 47103 7540 47112 7580
rect 47152 7540 47194 7580
rect 47234 7540 47276 7580
rect 47316 7540 47358 7580
rect 47398 7540 47440 7580
rect 47480 7540 47489 7580
rect 51103 7540 51112 7580
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51480 7540 51489 7580
rect 55103 7540 55112 7580
rect 55152 7540 55194 7580
rect 55234 7540 55276 7580
rect 55316 7540 55358 7580
rect 55398 7540 55440 7580
rect 55480 7540 55489 7580
rect 59103 7540 59112 7580
rect 59152 7540 59194 7580
rect 59234 7540 59276 7580
rect 59316 7540 59358 7580
rect 59398 7540 59440 7580
rect 59480 7540 59489 7580
rect 63103 7540 63112 7580
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63480 7540 63489 7580
rect 67103 7540 67112 7580
rect 67152 7540 67194 7580
rect 67234 7540 67276 7580
rect 67316 7540 67358 7580
rect 67398 7540 67440 7580
rect 67480 7540 67489 7580
rect 74668 7540 80372 7580
rect 82051 7540 82060 7580
rect 82100 7540 82828 7580
rect 82868 7540 82877 7580
rect 87811 7540 87820 7580
rect 87860 7540 88780 7580
rect 88820 7540 88829 7580
rect 93763 7540 93772 7580
rect 93812 7540 94924 7580
rect 94964 7540 94973 7580
rect 72547 7456 72556 7496
rect 72596 7456 73132 7496
rect 73172 7456 73181 7496
rect 74668 7412 74708 7540
rect 80332 7496 80372 7540
rect 86659 7496 86717 7497
rect 75235 7456 75244 7496
rect 75284 7456 75916 7496
rect 75956 7456 75965 7496
rect 77635 7456 77644 7496
rect 77684 7456 78124 7496
rect 78164 7456 78173 7496
rect 80323 7456 80332 7496
rect 80372 7456 80381 7496
rect 81187 7456 81196 7496
rect 81236 7456 82348 7496
rect 82388 7456 82397 7496
rect 82915 7456 82924 7496
rect 82964 7456 83980 7496
rect 84020 7456 84029 7496
rect 84835 7456 84844 7496
rect 84884 7456 85516 7496
rect 85556 7456 85565 7496
rect 86574 7456 86668 7496
rect 86708 7456 86717 7496
rect 86851 7456 86860 7496
rect 86900 7456 87724 7496
rect 87764 7456 87773 7496
rect 88387 7456 88396 7496
rect 88436 7456 89644 7496
rect 89684 7456 89693 7496
rect 90019 7456 90028 7496
rect 90068 7456 91316 7496
rect 92419 7456 92428 7496
rect 92468 7456 93484 7496
rect 93524 7456 93533 7496
rect 98083 7456 98092 7496
rect 98132 7456 99244 7496
rect 99284 7456 99293 7496
rect 86659 7455 86717 7456
rect 91276 7412 91316 7456
rect 835 7372 844 7412
rect 884 7372 1516 7412
rect 1556 7372 1565 7412
rect 71779 7372 71788 7412
rect 71828 7372 74668 7412
rect 74708 7372 74717 7412
rect 74851 7372 74860 7412
rect 74900 7372 75148 7412
rect 75188 7372 75197 7412
rect 76483 7372 76492 7412
rect 76532 7372 76780 7412
rect 76820 7372 76829 7412
rect 77251 7372 77260 7412
rect 77300 7372 77836 7412
rect 77876 7372 77885 7412
rect 78019 7372 78028 7412
rect 78068 7372 78412 7412
rect 78452 7372 78461 7412
rect 78787 7372 78796 7412
rect 78836 7372 79468 7412
rect 79508 7372 79517 7412
rect 80035 7372 80044 7412
rect 80084 7372 81100 7412
rect 81140 7372 81149 7412
rect 81667 7372 81676 7412
rect 81716 7372 82540 7412
rect 82580 7372 82589 7412
rect 84067 7372 84076 7412
rect 84116 7372 84460 7412
rect 84500 7372 84509 7412
rect 85219 7372 85228 7412
rect 85268 7372 85804 7412
rect 85844 7372 85853 7412
rect 86467 7372 86476 7412
rect 86516 7372 87436 7412
rect 87476 7372 87485 7412
rect 88003 7372 88012 7412
rect 88052 7372 88972 7412
rect 89012 7372 89021 7412
rect 89251 7372 89260 7412
rect 89300 7372 90220 7412
rect 90260 7372 90269 7412
rect 90595 7372 90604 7412
rect 90644 7372 90740 7412
rect 91267 7372 91276 7412
rect 91316 7372 91325 7412
rect 92803 7372 92812 7412
rect 92852 7372 93772 7412
rect 93812 7372 93821 7412
rect 95587 7372 95596 7412
rect 95636 7372 96460 7412
rect 96500 7372 96509 7412
rect 96835 7372 96844 7412
rect 96884 7372 97804 7412
rect 97844 7372 97853 7412
rect 98275 7372 98284 7412
rect 98324 7372 98476 7412
rect 98516 7372 98525 7412
rect 0 7328 80 7348
rect 90700 7328 90740 7372
rect 0 7288 652 7328
rect 692 7288 701 7328
rect 74275 7288 74284 7328
rect 74324 7288 75532 7328
rect 75572 7288 76628 7328
rect 76867 7288 76876 7328
rect 76916 7288 77644 7328
rect 77684 7288 77693 7328
rect 79171 7288 79180 7328
rect 79220 7288 80524 7328
rect 80564 7288 80573 7328
rect 82435 7288 82444 7328
rect 82484 7288 83596 7328
rect 83636 7288 83645 7328
rect 85699 7288 85708 7328
rect 85748 7288 86860 7328
rect 86900 7288 86909 7328
rect 87235 7288 87244 7328
rect 87284 7288 88396 7328
rect 88436 7288 88445 7328
rect 88867 7288 88876 7328
rect 88916 7288 90028 7328
rect 90068 7288 90077 7328
rect 90700 7288 91564 7328
rect 91604 7288 91613 7328
rect 91843 7288 91852 7328
rect 91892 7288 93004 7328
rect 93044 7288 93196 7328
rect 93236 7288 93245 7328
rect 93571 7288 93580 7328
rect 93620 7288 93868 7328
rect 93908 7288 94540 7328
rect 94580 7288 94589 7328
rect 94819 7288 94828 7328
rect 94868 7288 95980 7328
rect 96020 7288 96029 7328
rect 96259 7288 96268 7328
rect 96308 7288 96317 7328
rect 97219 7288 97228 7328
rect 97268 7288 98092 7328
rect 98132 7288 98141 7328
rect 0 7268 80 7288
rect 76588 7244 76628 7288
rect 74467 7204 74476 7244
rect 74516 7204 74860 7244
rect 74900 7204 74909 7244
rect 76099 7204 76108 7244
rect 76148 7204 76492 7244
rect 76532 7204 76541 7244
rect 76588 7204 77356 7244
rect 77396 7204 78796 7244
rect 78836 7204 78845 7244
rect 79747 7204 79756 7244
rect 79796 7204 80140 7244
rect 80180 7204 81580 7244
rect 81620 7204 83212 7244
rect 83252 7204 84844 7244
rect 84884 7204 84893 7244
rect 86275 7204 86284 7244
rect 86324 7204 86476 7244
rect 86516 7204 88204 7244
rect 88244 7204 89260 7244
rect 89300 7204 90796 7244
rect 90836 7204 90845 7244
rect 90979 7204 90988 7244
rect 91028 7204 91180 7244
rect 91220 7204 91229 7244
rect 91651 7204 91660 7244
rect 91700 7204 92908 7244
rect 92948 7204 92957 7244
rect 94435 7204 94444 7244
rect 94484 7204 95596 7244
rect 95636 7204 95645 7244
rect 96163 7204 96172 7244
rect 96212 7204 96221 7244
rect 96172 7160 96212 7204
rect 71107 7120 71116 7160
rect 71156 7120 72076 7160
rect 72116 7120 72364 7160
rect 72404 7120 72940 7160
rect 72980 7120 73612 7160
rect 73652 7120 73661 7160
rect 75715 7120 75724 7160
rect 75764 7120 76300 7160
rect 76340 7120 76588 7160
rect 76628 7120 76876 7160
rect 76916 7120 77548 7160
rect 77588 7120 77597 7160
rect 77923 7120 77932 7160
rect 77972 7120 78220 7160
rect 78260 7120 78508 7160
rect 78548 7120 79180 7160
rect 79220 7120 79229 7160
rect 80899 7120 80908 7160
rect 80948 7120 80957 7160
rect 81187 7120 81196 7160
rect 81236 7120 82060 7160
rect 82100 7120 82252 7160
rect 82292 7120 82301 7160
rect 82627 7120 82636 7160
rect 82676 7120 82924 7160
rect 82964 7120 83692 7160
rect 83732 7120 83884 7160
rect 83924 7120 83933 7160
rect 85027 7120 85036 7160
rect 85076 7120 85612 7160
rect 85652 7120 85900 7160
rect 85940 7120 86956 7160
rect 86996 7120 87148 7160
rect 87188 7120 87197 7160
rect 87331 7120 87340 7160
rect 87380 7120 87532 7160
rect 87572 7120 87820 7160
rect 87860 7120 88492 7160
rect 88532 7120 88684 7160
rect 88724 7120 88733 7160
rect 88867 7120 88876 7160
rect 88916 7120 89068 7160
rect 89108 7120 89740 7160
rect 89780 7120 89932 7160
rect 89972 7120 89981 7160
rect 90307 7120 90316 7160
rect 90356 7120 90604 7160
rect 90644 7120 91276 7160
rect 91316 7120 91468 7160
rect 91508 7120 91517 7160
rect 93283 7120 93292 7160
rect 93332 7120 94484 7160
rect 94531 7120 94540 7160
rect 94580 7120 94732 7160
rect 94772 7120 94781 7160
rect 95299 7120 95308 7160
rect 95348 7120 96212 7160
rect 96268 7160 96308 7288
rect 96547 7204 96556 7244
rect 96596 7204 97324 7244
rect 97364 7204 97373 7244
rect 96268 7120 97228 7160
rect 97268 7120 97277 7160
rect 97603 7120 97612 7160
rect 97652 7120 98900 7160
rect 73228 7076 73268 7120
rect 73219 7036 73228 7076
rect 73268 7036 73308 7076
rect 80908 6992 80948 7120
rect 90316 7076 90356 7120
rect 94444 7076 94484 7120
rect 98860 7076 98900 7120
rect 86179 7036 86188 7076
rect 86228 7036 87244 7076
rect 87284 7036 87293 7076
rect 89443 7036 89452 7076
rect 89492 7036 90356 7076
rect 92323 7036 92332 7076
rect 92372 7036 92524 7076
rect 92564 7036 94252 7076
rect 94292 7036 94301 7076
rect 94435 7036 94444 7076
rect 94484 7036 94493 7076
rect 96259 7036 96268 7076
rect 96308 7036 96556 7076
rect 96596 7036 96605 7076
rect 98851 7036 98860 7076
rect 98900 7036 98909 7076
rect 74083 6952 74092 6992
rect 74132 6952 74956 6992
rect 74996 6952 75244 6992
rect 75284 6952 76012 6992
rect 76052 6952 76492 6992
rect 76532 6952 76541 6992
rect 78979 6952 78988 6992
rect 79028 6952 79564 6992
rect 79604 6952 79756 6992
rect 79796 6952 80620 6992
rect 80660 6952 80812 6992
rect 80852 6952 80861 6992
rect 80908 6952 81964 6992
rect 82004 6952 82013 6992
rect 84259 6952 84268 6992
rect 84308 6952 84556 6992
rect 84596 6952 85228 6992
rect 85268 6952 85277 6992
rect 92035 6952 92044 6992
rect 92084 6952 93292 6992
rect 93332 6952 93341 6992
rect 96643 6952 96652 6992
rect 96692 6952 97612 6992
rect 97652 6952 97661 6992
rect 98179 6952 98188 6992
rect 98228 6952 98956 6992
rect 98996 6952 99005 6992
rect 79651 6868 79660 6908
rect 79700 6868 80908 6908
rect 80948 6868 80957 6908
rect 86659 6868 86668 6908
rect 86708 6868 92716 6908
rect 92756 6868 92765 6908
rect 94243 6868 94252 6908
rect 94292 6868 95212 6908
rect 95252 6868 96844 6908
rect 96884 6868 96893 6908
rect 4343 6784 4352 6824
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4720 6784 4729 6824
rect 8343 6784 8352 6824
rect 8392 6784 8434 6824
rect 8474 6784 8516 6824
rect 8556 6784 8598 6824
rect 8638 6784 8680 6824
rect 8720 6784 8729 6824
rect 12343 6784 12352 6824
rect 12392 6784 12434 6824
rect 12474 6784 12516 6824
rect 12556 6784 12598 6824
rect 12638 6784 12680 6824
rect 12720 6784 12729 6824
rect 16343 6784 16352 6824
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16720 6784 16729 6824
rect 20343 6784 20352 6824
rect 20392 6784 20434 6824
rect 20474 6784 20516 6824
rect 20556 6784 20598 6824
rect 20638 6784 20680 6824
rect 20720 6784 20729 6824
rect 24343 6784 24352 6824
rect 24392 6784 24434 6824
rect 24474 6784 24516 6824
rect 24556 6784 24598 6824
rect 24638 6784 24680 6824
rect 24720 6784 24729 6824
rect 28343 6784 28352 6824
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28720 6784 28729 6824
rect 32343 6784 32352 6824
rect 32392 6784 32434 6824
rect 32474 6784 32516 6824
rect 32556 6784 32598 6824
rect 32638 6784 32680 6824
rect 32720 6784 32729 6824
rect 36343 6784 36352 6824
rect 36392 6784 36434 6824
rect 36474 6784 36516 6824
rect 36556 6784 36598 6824
rect 36638 6784 36680 6824
rect 36720 6784 36729 6824
rect 40343 6784 40352 6824
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40720 6784 40729 6824
rect 44343 6784 44352 6824
rect 44392 6784 44434 6824
rect 44474 6784 44516 6824
rect 44556 6784 44598 6824
rect 44638 6784 44680 6824
rect 44720 6784 44729 6824
rect 48343 6784 48352 6824
rect 48392 6784 48434 6824
rect 48474 6784 48516 6824
rect 48556 6784 48598 6824
rect 48638 6784 48680 6824
rect 48720 6784 48729 6824
rect 52343 6784 52352 6824
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52720 6784 52729 6824
rect 56343 6784 56352 6824
rect 56392 6784 56434 6824
rect 56474 6784 56516 6824
rect 56556 6784 56598 6824
rect 56638 6784 56680 6824
rect 56720 6784 56729 6824
rect 60343 6784 60352 6824
rect 60392 6784 60434 6824
rect 60474 6784 60516 6824
rect 60556 6784 60598 6824
rect 60638 6784 60680 6824
rect 60720 6784 60729 6824
rect 64343 6784 64352 6824
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64720 6784 64729 6824
rect 68343 6784 68352 6824
rect 68392 6784 68434 6824
rect 68474 6784 68516 6824
rect 68556 6784 68598 6824
rect 68638 6784 68680 6824
rect 68720 6784 68729 6824
rect 97027 6784 97036 6824
rect 97076 6784 97228 6824
rect 97268 6784 97277 6824
rect 93763 6656 93821 6657
rect 835 6616 844 6656
rect 884 6616 1708 6656
rect 1748 6616 1757 6656
rect 80419 6616 80428 6656
rect 80468 6616 80908 6656
rect 80948 6616 80957 6656
rect 93678 6616 93772 6656
rect 93812 6616 93821 6656
rect 93763 6615 93821 6616
rect 0 6488 80 6508
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 93955 6448 93964 6488
rect 94004 6448 94156 6488
rect 94196 6448 94540 6488
rect 94580 6448 94924 6488
rect 94964 6448 95692 6488
rect 95732 6448 95741 6488
rect 0 6428 80 6448
rect 73987 6364 73996 6404
rect 74036 6364 74380 6404
rect 74420 6364 74860 6404
rect 74900 6364 74909 6404
rect 76867 6364 76876 6404
rect 76916 6364 77260 6404
rect 77300 6364 77644 6404
rect 77684 6364 78124 6404
rect 78164 6364 78173 6404
rect 78499 6364 78508 6404
rect 78548 6364 78892 6404
rect 78932 6364 79276 6404
rect 79316 6364 79756 6404
rect 79796 6364 79805 6404
rect 80131 6364 80140 6404
rect 80180 6364 80524 6404
rect 80564 6364 81004 6404
rect 81044 6364 81196 6404
rect 81236 6364 81245 6404
rect 81763 6364 81772 6404
rect 81812 6364 82060 6404
rect 82100 6364 82540 6404
rect 82580 6364 82589 6404
rect 83395 6364 83404 6404
rect 83444 6364 83692 6404
rect 83732 6364 84076 6404
rect 84116 6364 84460 6404
rect 84500 6364 84509 6404
rect 84835 6364 84844 6404
rect 84884 6364 85324 6404
rect 85364 6364 85373 6404
rect 86083 6364 86092 6404
rect 86132 6364 86476 6404
rect 86516 6364 86860 6404
rect 86900 6364 87340 6404
rect 87380 6364 87389 6404
rect 87907 6364 87916 6404
rect 87956 6364 88108 6404
rect 88148 6364 88492 6404
rect 88532 6364 88876 6404
rect 88916 6364 88925 6404
rect 89251 6364 89260 6404
rect 89300 6364 89740 6404
rect 89780 6364 90124 6404
rect 90164 6364 90508 6404
rect 90548 6364 90557 6404
rect 90979 6364 90988 6404
rect 91028 6364 91276 6404
rect 91316 6364 91756 6404
rect 91796 6364 91805 6404
rect 92131 6364 92140 6404
rect 92180 6364 92524 6404
rect 92564 6364 92908 6404
rect 92948 6364 93388 6404
rect 93428 6364 93437 6404
rect 95395 6364 95404 6404
rect 95444 6364 95788 6404
rect 95828 6364 96172 6404
rect 96212 6364 96221 6404
rect 97219 6364 97228 6404
rect 97268 6364 97708 6404
rect 97748 6364 98092 6404
rect 98132 6364 98141 6404
rect 3103 6028 3112 6068
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3480 6028 3489 6068
rect 7103 6028 7112 6068
rect 7152 6028 7194 6068
rect 7234 6028 7276 6068
rect 7316 6028 7358 6068
rect 7398 6028 7440 6068
rect 7480 6028 7489 6068
rect 11103 6028 11112 6068
rect 11152 6028 11194 6068
rect 11234 6028 11276 6068
rect 11316 6028 11358 6068
rect 11398 6028 11440 6068
rect 11480 6028 11489 6068
rect 15103 6028 15112 6068
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15480 6028 15489 6068
rect 19103 6028 19112 6068
rect 19152 6028 19194 6068
rect 19234 6028 19276 6068
rect 19316 6028 19358 6068
rect 19398 6028 19440 6068
rect 19480 6028 19489 6068
rect 23103 6028 23112 6068
rect 23152 6028 23194 6068
rect 23234 6028 23276 6068
rect 23316 6028 23358 6068
rect 23398 6028 23440 6068
rect 23480 6028 23489 6068
rect 27103 6028 27112 6068
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27480 6028 27489 6068
rect 31103 6028 31112 6068
rect 31152 6028 31194 6068
rect 31234 6028 31276 6068
rect 31316 6028 31358 6068
rect 31398 6028 31440 6068
rect 31480 6028 31489 6068
rect 35103 6028 35112 6068
rect 35152 6028 35194 6068
rect 35234 6028 35276 6068
rect 35316 6028 35358 6068
rect 35398 6028 35440 6068
rect 35480 6028 35489 6068
rect 39103 6028 39112 6068
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39480 6028 39489 6068
rect 43103 6028 43112 6068
rect 43152 6028 43194 6068
rect 43234 6028 43276 6068
rect 43316 6028 43358 6068
rect 43398 6028 43440 6068
rect 43480 6028 43489 6068
rect 47103 6028 47112 6068
rect 47152 6028 47194 6068
rect 47234 6028 47276 6068
rect 47316 6028 47358 6068
rect 47398 6028 47440 6068
rect 47480 6028 47489 6068
rect 51103 6028 51112 6068
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51480 6028 51489 6068
rect 55103 6028 55112 6068
rect 55152 6028 55194 6068
rect 55234 6028 55276 6068
rect 55316 6028 55358 6068
rect 55398 6028 55440 6068
rect 55480 6028 55489 6068
rect 59103 6028 59112 6068
rect 59152 6028 59194 6068
rect 59234 6028 59276 6068
rect 59316 6028 59358 6068
rect 59398 6028 59440 6068
rect 59480 6028 59489 6068
rect 63103 6028 63112 6068
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63480 6028 63489 6068
rect 67103 6028 67112 6068
rect 67152 6028 67194 6068
rect 67234 6028 67276 6068
rect 67316 6028 67358 6068
rect 67398 6028 67440 6068
rect 67480 6028 67489 6068
rect 0 5648 80 5668
rect 0 5608 652 5648
rect 692 5608 701 5648
rect 0 5588 80 5608
rect 4343 5272 4352 5312
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4720 5272 4729 5312
rect 8343 5272 8352 5312
rect 8392 5272 8434 5312
rect 8474 5272 8516 5312
rect 8556 5272 8598 5312
rect 8638 5272 8680 5312
rect 8720 5272 8729 5312
rect 12343 5272 12352 5312
rect 12392 5272 12434 5312
rect 12474 5272 12516 5312
rect 12556 5272 12598 5312
rect 12638 5272 12680 5312
rect 12720 5272 12729 5312
rect 16343 5272 16352 5312
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16720 5272 16729 5312
rect 20343 5272 20352 5312
rect 20392 5272 20434 5312
rect 20474 5272 20516 5312
rect 20556 5272 20598 5312
rect 20638 5272 20680 5312
rect 20720 5272 20729 5312
rect 24343 5272 24352 5312
rect 24392 5272 24434 5312
rect 24474 5272 24516 5312
rect 24556 5272 24598 5312
rect 24638 5272 24680 5312
rect 24720 5272 24729 5312
rect 28343 5272 28352 5312
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28720 5272 28729 5312
rect 32343 5272 32352 5312
rect 32392 5272 32434 5312
rect 32474 5272 32516 5312
rect 32556 5272 32598 5312
rect 32638 5272 32680 5312
rect 32720 5272 32729 5312
rect 36343 5272 36352 5312
rect 36392 5272 36434 5312
rect 36474 5272 36516 5312
rect 36556 5272 36598 5312
rect 36638 5272 36680 5312
rect 36720 5272 36729 5312
rect 40343 5272 40352 5312
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40720 5272 40729 5312
rect 44343 5272 44352 5312
rect 44392 5272 44434 5312
rect 44474 5272 44516 5312
rect 44556 5272 44598 5312
rect 44638 5272 44680 5312
rect 44720 5272 44729 5312
rect 48343 5272 48352 5312
rect 48392 5272 48434 5312
rect 48474 5272 48516 5312
rect 48556 5272 48598 5312
rect 48638 5272 48680 5312
rect 48720 5272 48729 5312
rect 52343 5272 52352 5312
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52720 5272 52729 5312
rect 56343 5272 56352 5312
rect 56392 5272 56434 5312
rect 56474 5272 56516 5312
rect 56556 5272 56598 5312
rect 56638 5272 56680 5312
rect 56720 5272 56729 5312
rect 60343 5272 60352 5312
rect 60392 5272 60434 5312
rect 60474 5272 60516 5312
rect 60556 5272 60598 5312
rect 60638 5272 60680 5312
rect 60720 5272 60729 5312
rect 64343 5272 64352 5312
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64720 5272 64729 5312
rect 68343 5272 68352 5312
rect 68392 5272 68434 5312
rect 68474 5272 68516 5312
rect 68556 5272 68598 5312
rect 68638 5272 68680 5312
rect 68720 5272 68729 5312
rect 72343 5272 72352 5312
rect 72392 5272 72434 5312
rect 72474 5272 72516 5312
rect 72556 5272 72598 5312
rect 72638 5272 72680 5312
rect 72720 5272 72729 5312
rect 76343 5272 76352 5312
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76720 5272 76729 5312
rect 80343 5272 80352 5312
rect 80392 5272 80434 5312
rect 80474 5272 80516 5312
rect 80556 5272 80598 5312
rect 80638 5272 80680 5312
rect 80720 5272 80729 5312
rect 84343 5272 84352 5312
rect 84392 5272 84434 5312
rect 84474 5272 84516 5312
rect 84556 5272 84598 5312
rect 84638 5272 84680 5312
rect 84720 5272 84729 5312
rect 88343 5272 88352 5312
rect 88392 5272 88434 5312
rect 88474 5272 88516 5312
rect 88556 5272 88598 5312
rect 88638 5272 88680 5312
rect 88720 5272 88729 5312
rect 92343 5272 92352 5312
rect 92392 5272 92434 5312
rect 92474 5272 92516 5312
rect 92556 5272 92598 5312
rect 92638 5272 92680 5312
rect 92720 5272 92729 5312
rect 96343 5272 96352 5312
rect 96392 5272 96434 5312
rect 96474 5272 96516 5312
rect 96556 5272 96598 5312
rect 96638 5272 96680 5312
rect 96720 5272 96729 5312
rect 1027 4852 1036 4892
rect 1076 4852 1420 4892
rect 1460 4852 1804 4892
rect 1844 4852 2188 4892
rect 2228 4852 2237 4892
rect 0 4808 80 4828
rect 0 4768 652 4808
rect 692 4768 701 4808
rect 0 4748 80 4768
rect 739 4684 748 4724
rect 788 4684 1996 4724
rect 2036 4684 2045 4724
rect 3103 4516 3112 4556
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3480 4516 3489 4556
rect 7103 4516 7112 4556
rect 7152 4516 7194 4556
rect 7234 4516 7276 4556
rect 7316 4516 7358 4556
rect 7398 4516 7440 4556
rect 7480 4516 7489 4556
rect 11103 4516 11112 4556
rect 11152 4516 11194 4556
rect 11234 4516 11276 4556
rect 11316 4516 11358 4556
rect 11398 4516 11440 4556
rect 11480 4516 11489 4556
rect 15103 4516 15112 4556
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15480 4516 15489 4556
rect 19103 4516 19112 4556
rect 19152 4516 19194 4556
rect 19234 4516 19276 4556
rect 19316 4516 19358 4556
rect 19398 4516 19440 4556
rect 19480 4516 19489 4556
rect 23103 4516 23112 4556
rect 23152 4516 23194 4556
rect 23234 4516 23276 4556
rect 23316 4516 23358 4556
rect 23398 4516 23440 4556
rect 23480 4516 23489 4556
rect 27103 4516 27112 4556
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27480 4516 27489 4556
rect 31103 4516 31112 4556
rect 31152 4516 31194 4556
rect 31234 4516 31276 4556
rect 31316 4516 31358 4556
rect 31398 4516 31440 4556
rect 31480 4516 31489 4556
rect 35103 4516 35112 4556
rect 35152 4516 35194 4556
rect 35234 4516 35276 4556
rect 35316 4516 35358 4556
rect 35398 4516 35440 4556
rect 35480 4516 35489 4556
rect 39103 4516 39112 4556
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39480 4516 39489 4556
rect 43103 4516 43112 4556
rect 43152 4516 43194 4556
rect 43234 4516 43276 4556
rect 43316 4516 43358 4556
rect 43398 4516 43440 4556
rect 43480 4516 43489 4556
rect 47103 4516 47112 4556
rect 47152 4516 47194 4556
rect 47234 4516 47276 4556
rect 47316 4516 47358 4556
rect 47398 4516 47440 4556
rect 47480 4516 47489 4556
rect 51103 4516 51112 4556
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51480 4516 51489 4556
rect 55103 4516 55112 4556
rect 55152 4516 55194 4556
rect 55234 4516 55276 4556
rect 55316 4516 55358 4556
rect 55398 4516 55440 4556
rect 55480 4516 55489 4556
rect 59103 4516 59112 4556
rect 59152 4516 59194 4556
rect 59234 4516 59276 4556
rect 59316 4516 59358 4556
rect 59398 4516 59440 4556
rect 59480 4516 59489 4556
rect 63103 4516 63112 4556
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63480 4516 63489 4556
rect 67103 4516 67112 4556
rect 67152 4516 67194 4556
rect 67234 4516 67276 4556
rect 67316 4516 67358 4556
rect 67398 4516 67440 4556
rect 67480 4516 67489 4556
rect 71103 4516 71112 4556
rect 71152 4516 71194 4556
rect 71234 4516 71276 4556
rect 71316 4516 71358 4556
rect 71398 4516 71440 4556
rect 71480 4516 71489 4556
rect 75103 4516 75112 4556
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75480 4516 75489 4556
rect 79103 4516 79112 4556
rect 79152 4516 79194 4556
rect 79234 4516 79276 4556
rect 79316 4516 79358 4556
rect 79398 4516 79440 4556
rect 79480 4516 79489 4556
rect 83103 4516 83112 4556
rect 83152 4516 83194 4556
rect 83234 4516 83276 4556
rect 83316 4516 83358 4556
rect 83398 4516 83440 4556
rect 83480 4516 83489 4556
rect 87103 4516 87112 4556
rect 87152 4516 87194 4556
rect 87234 4516 87276 4556
rect 87316 4516 87358 4556
rect 87398 4516 87440 4556
rect 87480 4516 87489 4556
rect 91103 4516 91112 4556
rect 91152 4516 91194 4556
rect 91234 4516 91276 4556
rect 91316 4516 91358 4556
rect 91398 4516 91440 4556
rect 91480 4516 91489 4556
rect 95103 4516 95112 4556
rect 95152 4516 95194 4556
rect 95234 4516 95276 4556
rect 95316 4516 95358 4556
rect 95398 4516 95440 4556
rect 95480 4516 95489 4556
rect 99103 4516 99112 4556
rect 99152 4516 99194 4556
rect 99234 4516 99276 4556
rect 99316 4516 99358 4556
rect 99398 4516 99440 4556
rect 99480 4516 99489 4556
rect 835 4180 844 4220
rect 884 4180 1612 4220
rect 1652 4180 1661 4220
rect 0 3968 80 3988
rect 0 3928 1036 3968
rect 1076 3928 1085 3968
rect 0 3908 80 3928
rect 4343 3760 4352 3800
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4720 3760 4729 3800
rect 8343 3760 8352 3800
rect 8392 3760 8434 3800
rect 8474 3760 8516 3800
rect 8556 3760 8598 3800
rect 8638 3760 8680 3800
rect 8720 3760 8729 3800
rect 12343 3760 12352 3800
rect 12392 3760 12434 3800
rect 12474 3760 12516 3800
rect 12556 3760 12598 3800
rect 12638 3760 12680 3800
rect 12720 3760 12729 3800
rect 16343 3760 16352 3800
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16720 3760 16729 3800
rect 20343 3760 20352 3800
rect 20392 3760 20434 3800
rect 20474 3760 20516 3800
rect 20556 3760 20598 3800
rect 20638 3760 20680 3800
rect 20720 3760 20729 3800
rect 24343 3760 24352 3800
rect 24392 3760 24434 3800
rect 24474 3760 24516 3800
rect 24556 3760 24598 3800
rect 24638 3760 24680 3800
rect 24720 3760 24729 3800
rect 28343 3760 28352 3800
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28720 3760 28729 3800
rect 32343 3760 32352 3800
rect 32392 3760 32434 3800
rect 32474 3760 32516 3800
rect 32556 3760 32598 3800
rect 32638 3760 32680 3800
rect 32720 3760 32729 3800
rect 36343 3760 36352 3800
rect 36392 3760 36434 3800
rect 36474 3760 36516 3800
rect 36556 3760 36598 3800
rect 36638 3760 36680 3800
rect 36720 3760 36729 3800
rect 40343 3760 40352 3800
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40720 3760 40729 3800
rect 44343 3760 44352 3800
rect 44392 3760 44434 3800
rect 44474 3760 44516 3800
rect 44556 3760 44598 3800
rect 44638 3760 44680 3800
rect 44720 3760 44729 3800
rect 48343 3760 48352 3800
rect 48392 3760 48434 3800
rect 48474 3760 48516 3800
rect 48556 3760 48598 3800
rect 48638 3760 48680 3800
rect 48720 3760 48729 3800
rect 52343 3760 52352 3800
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52720 3760 52729 3800
rect 56343 3760 56352 3800
rect 56392 3760 56434 3800
rect 56474 3760 56516 3800
rect 56556 3760 56598 3800
rect 56638 3760 56680 3800
rect 56720 3760 56729 3800
rect 60343 3760 60352 3800
rect 60392 3760 60434 3800
rect 60474 3760 60516 3800
rect 60556 3760 60598 3800
rect 60638 3760 60680 3800
rect 60720 3760 60729 3800
rect 64343 3760 64352 3800
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64720 3760 64729 3800
rect 68343 3760 68352 3800
rect 68392 3760 68434 3800
rect 68474 3760 68516 3800
rect 68556 3760 68598 3800
rect 68638 3760 68680 3800
rect 68720 3760 68729 3800
rect 72343 3760 72352 3800
rect 72392 3760 72434 3800
rect 72474 3760 72516 3800
rect 72556 3760 72598 3800
rect 72638 3760 72680 3800
rect 72720 3760 72729 3800
rect 76343 3760 76352 3800
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76720 3760 76729 3800
rect 80343 3760 80352 3800
rect 80392 3760 80434 3800
rect 80474 3760 80516 3800
rect 80556 3760 80598 3800
rect 80638 3760 80680 3800
rect 80720 3760 80729 3800
rect 84343 3760 84352 3800
rect 84392 3760 84434 3800
rect 84474 3760 84516 3800
rect 84556 3760 84598 3800
rect 84638 3760 84680 3800
rect 84720 3760 84729 3800
rect 88343 3760 88352 3800
rect 88392 3760 88434 3800
rect 88474 3760 88516 3800
rect 88556 3760 88598 3800
rect 88638 3760 88680 3800
rect 88720 3760 88729 3800
rect 92343 3760 92352 3800
rect 92392 3760 92434 3800
rect 92474 3760 92516 3800
rect 92556 3760 92598 3800
rect 92638 3760 92680 3800
rect 92720 3760 92729 3800
rect 96343 3760 96352 3800
rect 96392 3760 96434 3800
rect 96474 3760 96516 3800
rect 96556 3760 96598 3800
rect 96638 3760 96680 3800
rect 96720 3760 96729 3800
rect 643 3172 652 3212
rect 692 3172 701 3212
rect 0 3128 80 3148
rect 652 3128 692 3172
rect 0 3088 692 3128
rect 0 3068 80 3088
rect 3103 3004 3112 3044
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3480 3004 3489 3044
rect 7103 3004 7112 3044
rect 7152 3004 7194 3044
rect 7234 3004 7276 3044
rect 7316 3004 7358 3044
rect 7398 3004 7440 3044
rect 7480 3004 7489 3044
rect 11103 3004 11112 3044
rect 11152 3004 11194 3044
rect 11234 3004 11276 3044
rect 11316 3004 11358 3044
rect 11398 3004 11440 3044
rect 11480 3004 11489 3044
rect 15103 3004 15112 3044
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15480 3004 15489 3044
rect 19103 3004 19112 3044
rect 19152 3004 19194 3044
rect 19234 3004 19276 3044
rect 19316 3004 19358 3044
rect 19398 3004 19440 3044
rect 19480 3004 19489 3044
rect 23103 3004 23112 3044
rect 23152 3004 23194 3044
rect 23234 3004 23276 3044
rect 23316 3004 23358 3044
rect 23398 3004 23440 3044
rect 23480 3004 23489 3044
rect 27103 3004 27112 3044
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27480 3004 27489 3044
rect 31103 3004 31112 3044
rect 31152 3004 31194 3044
rect 31234 3004 31276 3044
rect 31316 3004 31358 3044
rect 31398 3004 31440 3044
rect 31480 3004 31489 3044
rect 35103 3004 35112 3044
rect 35152 3004 35194 3044
rect 35234 3004 35276 3044
rect 35316 3004 35358 3044
rect 35398 3004 35440 3044
rect 35480 3004 35489 3044
rect 39103 3004 39112 3044
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39480 3004 39489 3044
rect 43103 3004 43112 3044
rect 43152 3004 43194 3044
rect 43234 3004 43276 3044
rect 43316 3004 43358 3044
rect 43398 3004 43440 3044
rect 43480 3004 43489 3044
rect 47103 3004 47112 3044
rect 47152 3004 47194 3044
rect 47234 3004 47276 3044
rect 47316 3004 47358 3044
rect 47398 3004 47440 3044
rect 47480 3004 47489 3044
rect 51103 3004 51112 3044
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51480 3004 51489 3044
rect 55103 3004 55112 3044
rect 55152 3004 55194 3044
rect 55234 3004 55276 3044
rect 55316 3004 55358 3044
rect 55398 3004 55440 3044
rect 55480 3004 55489 3044
rect 59103 3004 59112 3044
rect 59152 3004 59194 3044
rect 59234 3004 59276 3044
rect 59316 3004 59358 3044
rect 59398 3004 59440 3044
rect 59480 3004 59489 3044
rect 63103 3004 63112 3044
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63480 3004 63489 3044
rect 67103 3004 67112 3044
rect 67152 3004 67194 3044
rect 67234 3004 67276 3044
rect 67316 3004 67358 3044
rect 67398 3004 67440 3044
rect 67480 3004 67489 3044
rect 71103 3004 71112 3044
rect 71152 3004 71194 3044
rect 71234 3004 71276 3044
rect 71316 3004 71358 3044
rect 71398 3004 71440 3044
rect 71480 3004 71489 3044
rect 75103 3004 75112 3044
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75480 3004 75489 3044
rect 79103 3004 79112 3044
rect 79152 3004 79194 3044
rect 79234 3004 79276 3044
rect 79316 3004 79358 3044
rect 79398 3004 79440 3044
rect 79480 3004 79489 3044
rect 83103 3004 83112 3044
rect 83152 3004 83194 3044
rect 83234 3004 83276 3044
rect 83316 3004 83358 3044
rect 83398 3004 83440 3044
rect 83480 3004 83489 3044
rect 87103 3004 87112 3044
rect 87152 3004 87194 3044
rect 87234 3004 87276 3044
rect 87316 3004 87358 3044
rect 87398 3004 87440 3044
rect 87480 3004 87489 3044
rect 91103 3004 91112 3044
rect 91152 3004 91194 3044
rect 91234 3004 91276 3044
rect 91316 3004 91358 3044
rect 91398 3004 91440 3044
rect 91480 3004 91489 3044
rect 95103 3004 95112 3044
rect 95152 3004 95194 3044
rect 95234 3004 95276 3044
rect 95316 3004 95358 3044
rect 95398 3004 95440 3044
rect 95480 3004 95489 3044
rect 99103 3004 99112 3044
rect 99152 3004 99194 3044
rect 99234 3004 99276 3044
rect 99316 3004 99358 3044
rect 99398 3004 99440 3044
rect 99480 3004 99489 3044
rect 0 2288 80 2308
rect 0 2248 652 2288
rect 692 2248 701 2288
rect 4343 2248 4352 2288
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4720 2248 4729 2288
rect 8343 2248 8352 2288
rect 8392 2248 8434 2288
rect 8474 2248 8516 2288
rect 8556 2248 8598 2288
rect 8638 2248 8680 2288
rect 8720 2248 8729 2288
rect 12343 2248 12352 2288
rect 12392 2248 12434 2288
rect 12474 2248 12516 2288
rect 12556 2248 12598 2288
rect 12638 2248 12680 2288
rect 12720 2248 12729 2288
rect 16343 2248 16352 2288
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16720 2248 16729 2288
rect 20343 2248 20352 2288
rect 20392 2248 20434 2288
rect 20474 2248 20516 2288
rect 20556 2248 20598 2288
rect 20638 2248 20680 2288
rect 20720 2248 20729 2288
rect 24343 2248 24352 2288
rect 24392 2248 24434 2288
rect 24474 2248 24516 2288
rect 24556 2248 24598 2288
rect 24638 2248 24680 2288
rect 24720 2248 24729 2288
rect 28343 2248 28352 2288
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28720 2248 28729 2288
rect 32343 2248 32352 2288
rect 32392 2248 32434 2288
rect 32474 2248 32516 2288
rect 32556 2248 32598 2288
rect 32638 2248 32680 2288
rect 32720 2248 32729 2288
rect 36343 2248 36352 2288
rect 36392 2248 36434 2288
rect 36474 2248 36516 2288
rect 36556 2248 36598 2288
rect 36638 2248 36680 2288
rect 36720 2248 36729 2288
rect 40343 2248 40352 2288
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40720 2248 40729 2288
rect 44343 2248 44352 2288
rect 44392 2248 44434 2288
rect 44474 2248 44516 2288
rect 44556 2248 44598 2288
rect 44638 2248 44680 2288
rect 44720 2248 44729 2288
rect 48343 2248 48352 2288
rect 48392 2248 48434 2288
rect 48474 2248 48516 2288
rect 48556 2248 48598 2288
rect 48638 2248 48680 2288
rect 48720 2248 48729 2288
rect 52343 2248 52352 2288
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52720 2248 52729 2288
rect 56343 2248 56352 2288
rect 56392 2248 56434 2288
rect 56474 2248 56516 2288
rect 56556 2248 56598 2288
rect 56638 2248 56680 2288
rect 56720 2248 56729 2288
rect 60343 2248 60352 2288
rect 60392 2248 60434 2288
rect 60474 2248 60516 2288
rect 60556 2248 60598 2288
rect 60638 2248 60680 2288
rect 60720 2248 60729 2288
rect 64343 2248 64352 2288
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64720 2248 64729 2288
rect 68343 2248 68352 2288
rect 68392 2248 68434 2288
rect 68474 2248 68516 2288
rect 68556 2248 68598 2288
rect 68638 2248 68680 2288
rect 68720 2248 68729 2288
rect 72343 2248 72352 2288
rect 72392 2248 72434 2288
rect 72474 2248 72516 2288
rect 72556 2248 72598 2288
rect 72638 2248 72680 2288
rect 72720 2248 72729 2288
rect 76343 2248 76352 2288
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76720 2248 76729 2288
rect 80343 2248 80352 2288
rect 80392 2248 80434 2288
rect 80474 2248 80516 2288
rect 80556 2248 80598 2288
rect 80638 2248 80680 2288
rect 80720 2248 80729 2288
rect 84343 2248 84352 2288
rect 84392 2248 84434 2288
rect 84474 2248 84516 2288
rect 84556 2248 84598 2288
rect 84638 2248 84680 2288
rect 84720 2248 84729 2288
rect 88343 2248 88352 2288
rect 88392 2248 88434 2288
rect 88474 2248 88516 2288
rect 88556 2248 88598 2288
rect 88638 2248 88680 2288
rect 88720 2248 88729 2288
rect 92343 2248 92352 2288
rect 92392 2248 92434 2288
rect 92474 2248 92516 2288
rect 92556 2248 92598 2288
rect 92638 2248 92680 2288
rect 92720 2248 92729 2288
rect 96343 2248 96352 2288
rect 96392 2248 96434 2288
rect 96474 2248 96516 2288
rect 96556 2248 96598 2288
rect 96638 2248 96680 2288
rect 96720 2248 96729 2288
rect 0 2228 80 2248
rect 3103 1492 3112 1532
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3480 1492 3489 1532
rect 7103 1492 7112 1532
rect 7152 1492 7194 1532
rect 7234 1492 7276 1532
rect 7316 1492 7358 1532
rect 7398 1492 7440 1532
rect 7480 1492 7489 1532
rect 11103 1492 11112 1532
rect 11152 1492 11194 1532
rect 11234 1492 11276 1532
rect 11316 1492 11358 1532
rect 11398 1492 11440 1532
rect 11480 1492 11489 1532
rect 15103 1492 15112 1532
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15480 1492 15489 1532
rect 19103 1492 19112 1532
rect 19152 1492 19194 1532
rect 19234 1492 19276 1532
rect 19316 1492 19358 1532
rect 19398 1492 19440 1532
rect 19480 1492 19489 1532
rect 23103 1492 23112 1532
rect 23152 1492 23194 1532
rect 23234 1492 23276 1532
rect 23316 1492 23358 1532
rect 23398 1492 23440 1532
rect 23480 1492 23489 1532
rect 27103 1492 27112 1532
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27480 1492 27489 1532
rect 31103 1492 31112 1532
rect 31152 1492 31194 1532
rect 31234 1492 31276 1532
rect 31316 1492 31358 1532
rect 31398 1492 31440 1532
rect 31480 1492 31489 1532
rect 35103 1492 35112 1532
rect 35152 1492 35194 1532
rect 35234 1492 35276 1532
rect 35316 1492 35358 1532
rect 35398 1492 35440 1532
rect 35480 1492 35489 1532
rect 39103 1492 39112 1532
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39480 1492 39489 1532
rect 43103 1492 43112 1532
rect 43152 1492 43194 1532
rect 43234 1492 43276 1532
rect 43316 1492 43358 1532
rect 43398 1492 43440 1532
rect 43480 1492 43489 1532
rect 47103 1492 47112 1532
rect 47152 1492 47194 1532
rect 47234 1492 47276 1532
rect 47316 1492 47358 1532
rect 47398 1492 47440 1532
rect 47480 1492 47489 1532
rect 51103 1492 51112 1532
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51480 1492 51489 1532
rect 55103 1492 55112 1532
rect 55152 1492 55194 1532
rect 55234 1492 55276 1532
rect 55316 1492 55358 1532
rect 55398 1492 55440 1532
rect 55480 1492 55489 1532
rect 59103 1492 59112 1532
rect 59152 1492 59194 1532
rect 59234 1492 59276 1532
rect 59316 1492 59358 1532
rect 59398 1492 59440 1532
rect 59480 1492 59489 1532
rect 63103 1492 63112 1532
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63480 1492 63489 1532
rect 67103 1492 67112 1532
rect 67152 1492 67194 1532
rect 67234 1492 67276 1532
rect 67316 1492 67358 1532
rect 67398 1492 67440 1532
rect 67480 1492 67489 1532
rect 71103 1492 71112 1532
rect 71152 1492 71194 1532
rect 71234 1492 71276 1532
rect 71316 1492 71358 1532
rect 71398 1492 71440 1532
rect 71480 1492 71489 1532
rect 75103 1492 75112 1532
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75480 1492 75489 1532
rect 79103 1492 79112 1532
rect 79152 1492 79194 1532
rect 79234 1492 79276 1532
rect 79316 1492 79358 1532
rect 79398 1492 79440 1532
rect 79480 1492 79489 1532
rect 83103 1492 83112 1532
rect 83152 1492 83194 1532
rect 83234 1492 83276 1532
rect 83316 1492 83358 1532
rect 83398 1492 83440 1532
rect 83480 1492 83489 1532
rect 87103 1492 87112 1532
rect 87152 1492 87194 1532
rect 87234 1492 87276 1532
rect 87316 1492 87358 1532
rect 87398 1492 87440 1532
rect 87480 1492 87489 1532
rect 91103 1492 91112 1532
rect 91152 1492 91194 1532
rect 91234 1492 91276 1532
rect 91316 1492 91358 1532
rect 91398 1492 91440 1532
rect 91480 1492 91489 1532
rect 95103 1492 95112 1532
rect 95152 1492 95194 1532
rect 95234 1492 95276 1532
rect 95316 1492 95358 1532
rect 95398 1492 95440 1532
rect 95480 1492 95489 1532
rect 99103 1492 99112 1532
rect 99152 1492 99194 1532
rect 99234 1492 99276 1532
rect 99316 1492 99358 1532
rect 99398 1492 99440 1532
rect 99480 1492 99489 1532
rect 4343 736 4352 776
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4720 736 4729 776
rect 8343 736 8352 776
rect 8392 736 8434 776
rect 8474 736 8516 776
rect 8556 736 8598 776
rect 8638 736 8680 776
rect 8720 736 8729 776
rect 12343 736 12352 776
rect 12392 736 12434 776
rect 12474 736 12516 776
rect 12556 736 12598 776
rect 12638 736 12680 776
rect 12720 736 12729 776
rect 16343 736 16352 776
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16720 736 16729 776
rect 20343 736 20352 776
rect 20392 736 20434 776
rect 20474 736 20516 776
rect 20556 736 20598 776
rect 20638 736 20680 776
rect 20720 736 20729 776
rect 24343 736 24352 776
rect 24392 736 24434 776
rect 24474 736 24516 776
rect 24556 736 24598 776
rect 24638 736 24680 776
rect 24720 736 24729 776
rect 28343 736 28352 776
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28720 736 28729 776
rect 32343 736 32352 776
rect 32392 736 32434 776
rect 32474 736 32516 776
rect 32556 736 32598 776
rect 32638 736 32680 776
rect 32720 736 32729 776
rect 36343 736 36352 776
rect 36392 736 36434 776
rect 36474 736 36516 776
rect 36556 736 36598 776
rect 36638 736 36680 776
rect 36720 736 36729 776
rect 40343 736 40352 776
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40720 736 40729 776
rect 44343 736 44352 776
rect 44392 736 44434 776
rect 44474 736 44516 776
rect 44556 736 44598 776
rect 44638 736 44680 776
rect 44720 736 44729 776
rect 48343 736 48352 776
rect 48392 736 48434 776
rect 48474 736 48516 776
rect 48556 736 48598 776
rect 48638 736 48680 776
rect 48720 736 48729 776
rect 52343 736 52352 776
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52720 736 52729 776
rect 56343 736 56352 776
rect 56392 736 56434 776
rect 56474 736 56516 776
rect 56556 736 56598 776
rect 56638 736 56680 776
rect 56720 736 56729 776
rect 60343 736 60352 776
rect 60392 736 60434 776
rect 60474 736 60516 776
rect 60556 736 60598 776
rect 60638 736 60680 776
rect 60720 736 60729 776
rect 64343 736 64352 776
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64720 736 64729 776
rect 68343 736 68352 776
rect 68392 736 68434 776
rect 68474 736 68516 776
rect 68556 736 68598 776
rect 68638 736 68680 776
rect 68720 736 68729 776
rect 72343 736 72352 776
rect 72392 736 72434 776
rect 72474 736 72516 776
rect 72556 736 72598 776
rect 72638 736 72680 776
rect 72720 736 72729 776
rect 76343 736 76352 776
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76720 736 76729 776
rect 80343 736 80352 776
rect 80392 736 80434 776
rect 80474 736 80516 776
rect 80556 736 80598 776
rect 80638 736 80680 776
rect 80720 736 80729 776
rect 84343 736 84352 776
rect 84392 736 84434 776
rect 84474 736 84516 776
rect 84556 736 84598 776
rect 84638 736 84680 776
rect 84720 736 84729 776
rect 88343 736 88352 776
rect 88392 736 88434 776
rect 88474 736 88516 776
rect 88556 736 88598 776
rect 88638 736 88680 776
rect 88720 736 88729 776
rect 92343 736 92352 776
rect 92392 736 92434 776
rect 92474 736 92516 776
rect 92556 736 92598 776
rect 92638 736 92680 776
rect 92720 736 92729 776
rect 96343 736 96352 776
rect 96392 736 96434 776
rect 96474 736 96516 776
rect 96556 736 96598 776
rect 96638 736 96680 776
rect 96720 736 96729 776
<< via3 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 8352 38536 8392 38576
rect 8434 38536 8474 38576
rect 8516 38536 8556 38576
rect 8598 38536 8638 38576
rect 8680 38536 8720 38576
rect 12352 38536 12392 38576
rect 12434 38536 12474 38576
rect 12516 38536 12556 38576
rect 12598 38536 12638 38576
rect 12680 38536 12720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 20352 38536 20392 38576
rect 20434 38536 20474 38576
rect 20516 38536 20556 38576
rect 20598 38536 20638 38576
rect 20680 38536 20720 38576
rect 24352 38536 24392 38576
rect 24434 38536 24474 38576
rect 24516 38536 24556 38576
rect 24598 38536 24638 38576
rect 24680 38536 24720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 32352 38536 32392 38576
rect 32434 38536 32474 38576
rect 32516 38536 32556 38576
rect 32598 38536 32638 38576
rect 32680 38536 32720 38576
rect 36352 38536 36392 38576
rect 36434 38536 36474 38576
rect 36516 38536 36556 38576
rect 36598 38536 36638 38576
rect 36680 38536 36720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 44352 38536 44392 38576
rect 44434 38536 44474 38576
rect 44516 38536 44556 38576
rect 44598 38536 44638 38576
rect 44680 38536 44720 38576
rect 48352 38536 48392 38576
rect 48434 38536 48474 38576
rect 48516 38536 48556 38576
rect 48598 38536 48638 38576
rect 48680 38536 48720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 56352 38536 56392 38576
rect 56434 38536 56474 38576
rect 56516 38536 56556 38576
rect 56598 38536 56638 38576
rect 56680 38536 56720 38576
rect 60352 38536 60392 38576
rect 60434 38536 60474 38576
rect 60516 38536 60556 38576
rect 60598 38536 60638 38576
rect 60680 38536 60720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 68352 38536 68392 38576
rect 68434 38536 68474 38576
rect 68516 38536 68556 38576
rect 68598 38536 68638 38576
rect 68680 38536 68720 38576
rect 72352 38536 72392 38576
rect 72434 38536 72474 38576
rect 72516 38536 72556 38576
rect 72598 38536 72638 38576
rect 72680 38536 72720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 80352 38536 80392 38576
rect 80434 38536 80474 38576
rect 80516 38536 80556 38576
rect 80598 38536 80638 38576
rect 80680 38536 80720 38576
rect 84352 38536 84392 38576
rect 84434 38536 84474 38576
rect 84516 38536 84556 38576
rect 84598 38536 84638 38576
rect 84680 38536 84720 38576
rect 88352 38536 88392 38576
rect 88434 38536 88474 38576
rect 88516 38536 88556 38576
rect 88598 38536 88638 38576
rect 88680 38536 88720 38576
rect 92352 38536 92392 38576
rect 92434 38536 92474 38576
rect 92516 38536 92556 38576
rect 92598 38536 92638 38576
rect 92680 38536 92720 38576
rect 96352 38536 96392 38576
rect 96434 38536 96474 38576
rect 96516 38536 96556 38576
rect 96598 38536 96638 38576
rect 96680 38536 96720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 7112 37780 7152 37820
rect 7194 37780 7234 37820
rect 7276 37780 7316 37820
rect 7358 37780 7398 37820
rect 7440 37780 7480 37820
rect 11112 37780 11152 37820
rect 11194 37780 11234 37820
rect 11276 37780 11316 37820
rect 11358 37780 11398 37820
rect 11440 37780 11480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 19112 37780 19152 37820
rect 19194 37780 19234 37820
rect 19276 37780 19316 37820
rect 19358 37780 19398 37820
rect 19440 37780 19480 37820
rect 23112 37780 23152 37820
rect 23194 37780 23234 37820
rect 23276 37780 23316 37820
rect 23358 37780 23398 37820
rect 23440 37780 23480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 31112 37780 31152 37820
rect 31194 37780 31234 37820
rect 31276 37780 31316 37820
rect 31358 37780 31398 37820
rect 31440 37780 31480 37820
rect 35112 37780 35152 37820
rect 35194 37780 35234 37820
rect 35276 37780 35316 37820
rect 35358 37780 35398 37820
rect 35440 37780 35480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 43112 37780 43152 37820
rect 43194 37780 43234 37820
rect 43276 37780 43316 37820
rect 43358 37780 43398 37820
rect 43440 37780 43480 37820
rect 47112 37780 47152 37820
rect 47194 37780 47234 37820
rect 47276 37780 47316 37820
rect 47358 37780 47398 37820
rect 47440 37780 47480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 55112 37780 55152 37820
rect 55194 37780 55234 37820
rect 55276 37780 55316 37820
rect 55358 37780 55398 37820
rect 55440 37780 55480 37820
rect 59112 37780 59152 37820
rect 59194 37780 59234 37820
rect 59276 37780 59316 37820
rect 59358 37780 59398 37820
rect 59440 37780 59480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 67112 37780 67152 37820
rect 67194 37780 67234 37820
rect 67276 37780 67316 37820
rect 67358 37780 67398 37820
rect 67440 37780 67480 37820
rect 71112 37780 71152 37820
rect 71194 37780 71234 37820
rect 71276 37780 71316 37820
rect 71358 37780 71398 37820
rect 71440 37780 71480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 79112 37780 79152 37820
rect 79194 37780 79234 37820
rect 79276 37780 79316 37820
rect 79358 37780 79398 37820
rect 79440 37780 79480 37820
rect 83112 37780 83152 37820
rect 83194 37780 83234 37820
rect 83276 37780 83316 37820
rect 83358 37780 83398 37820
rect 83440 37780 83480 37820
rect 87112 37780 87152 37820
rect 87194 37780 87234 37820
rect 87276 37780 87316 37820
rect 87358 37780 87398 37820
rect 87440 37780 87480 37820
rect 91112 37780 91152 37820
rect 91194 37780 91234 37820
rect 91276 37780 91316 37820
rect 91358 37780 91398 37820
rect 91440 37780 91480 37820
rect 95112 37780 95152 37820
rect 95194 37780 95234 37820
rect 95276 37780 95316 37820
rect 95358 37780 95398 37820
rect 95440 37780 95480 37820
rect 99112 37780 99152 37820
rect 99194 37780 99234 37820
rect 99276 37780 99316 37820
rect 99358 37780 99398 37820
rect 99440 37780 99480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 8352 37024 8392 37064
rect 8434 37024 8474 37064
rect 8516 37024 8556 37064
rect 8598 37024 8638 37064
rect 8680 37024 8720 37064
rect 12352 37024 12392 37064
rect 12434 37024 12474 37064
rect 12516 37024 12556 37064
rect 12598 37024 12638 37064
rect 12680 37024 12720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 20352 37024 20392 37064
rect 20434 37024 20474 37064
rect 20516 37024 20556 37064
rect 20598 37024 20638 37064
rect 20680 37024 20720 37064
rect 24352 37024 24392 37064
rect 24434 37024 24474 37064
rect 24516 37024 24556 37064
rect 24598 37024 24638 37064
rect 24680 37024 24720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 32352 37024 32392 37064
rect 32434 37024 32474 37064
rect 32516 37024 32556 37064
rect 32598 37024 32638 37064
rect 32680 37024 32720 37064
rect 36352 37024 36392 37064
rect 36434 37024 36474 37064
rect 36516 37024 36556 37064
rect 36598 37024 36638 37064
rect 36680 37024 36720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 44352 37024 44392 37064
rect 44434 37024 44474 37064
rect 44516 37024 44556 37064
rect 44598 37024 44638 37064
rect 44680 37024 44720 37064
rect 48352 37024 48392 37064
rect 48434 37024 48474 37064
rect 48516 37024 48556 37064
rect 48598 37024 48638 37064
rect 48680 37024 48720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 56352 37024 56392 37064
rect 56434 37024 56474 37064
rect 56516 37024 56556 37064
rect 56598 37024 56638 37064
rect 56680 37024 56720 37064
rect 60352 37024 60392 37064
rect 60434 37024 60474 37064
rect 60516 37024 60556 37064
rect 60598 37024 60638 37064
rect 60680 37024 60720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 68352 37024 68392 37064
rect 68434 37024 68474 37064
rect 68516 37024 68556 37064
rect 68598 37024 68638 37064
rect 68680 37024 68720 37064
rect 72352 37024 72392 37064
rect 72434 37024 72474 37064
rect 72516 37024 72556 37064
rect 72598 37024 72638 37064
rect 72680 37024 72720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 80352 37024 80392 37064
rect 80434 37024 80474 37064
rect 80516 37024 80556 37064
rect 80598 37024 80638 37064
rect 80680 37024 80720 37064
rect 84352 37024 84392 37064
rect 84434 37024 84474 37064
rect 84516 37024 84556 37064
rect 84598 37024 84638 37064
rect 84680 37024 84720 37064
rect 88352 37024 88392 37064
rect 88434 37024 88474 37064
rect 88516 37024 88556 37064
rect 88598 37024 88638 37064
rect 88680 37024 88720 37064
rect 92352 37024 92392 37064
rect 92434 37024 92474 37064
rect 92516 37024 92556 37064
rect 92598 37024 92638 37064
rect 92680 37024 92720 37064
rect 96352 37024 96392 37064
rect 96434 37024 96474 37064
rect 96516 37024 96556 37064
rect 96598 37024 96638 37064
rect 96680 37024 96720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 7112 36268 7152 36308
rect 7194 36268 7234 36308
rect 7276 36268 7316 36308
rect 7358 36268 7398 36308
rect 7440 36268 7480 36308
rect 11112 36268 11152 36308
rect 11194 36268 11234 36308
rect 11276 36268 11316 36308
rect 11358 36268 11398 36308
rect 11440 36268 11480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 19112 36268 19152 36308
rect 19194 36268 19234 36308
rect 19276 36268 19316 36308
rect 19358 36268 19398 36308
rect 19440 36268 19480 36308
rect 23112 36268 23152 36308
rect 23194 36268 23234 36308
rect 23276 36268 23316 36308
rect 23358 36268 23398 36308
rect 23440 36268 23480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 31112 36268 31152 36308
rect 31194 36268 31234 36308
rect 31276 36268 31316 36308
rect 31358 36268 31398 36308
rect 31440 36268 31480 36308
rect 35112 36268 35152 36308
rect 35194 36268 35234 36308
rect 35276 36268 35316 36308
rect 35358 36268 35398 36308
rect 35440 36268 35480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 43112 36268 43152 36308
rect 43194 36268 43234 36308
rect 43276 36268 43316 36308
rect 43358 36268 43398 36308
rect 43440 36268 43480 36308
rect 47112 36268 47152 36308
rect 47194 36268 47234 36308
rect 47276 36268 47316 36308
rect 47358 36268 47398 36308
rect 47440 36268 47480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 55112 36268 55152 36308
rect 55194 36268 55234 36308
rect 55276 36268 55316 36308
rect 55358 36268 55398 36308
rect 55440 36268 55480 36308
rect 59112 36268 59152 36308
rect 59194 36268 59234 36308
rect 59276 36268 59316 36308
rect 59358 36268 59398 36308
rect 59440 36268 59480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 67112 36268 67152 36308
rect 67194 36268 67234 36308
rect 67276 36268 67316 36308
rect 67358 36268 67398 36308
rect 67440 36268 67480 36308
rect 71112 36268 71152 36308
rect 71194 36268 71234 36308
rect 71276 36268 71316 36308
rect 71358 36268 71398 36308
rect 71440 36268 71480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 79112 36268 79152 36308
rect 79194 36268 79234 36308
rect 79276 36268 79316 36308
rect 79358 36268 79398 36308
rect 79440 36268 79480 36308
rect 83112 36268 83152 36308
rect 83194 36268 83234 36308
rect 83276 36268 83316 36308
rect 83358 36268 83398 36308
rect 83440 36268 83480 36308
rect 87112 36268 87152 36308
rect 87194 36268 87234 36308
rect 87276 36268 87316 36308
rect 87358 36268 87398 36308
rect 87440 36268 87480 36308
rect 91112 36268 91152 36308
rect 91194 36268 91234 36308
rect 91276 36268 91316 36308
rect 91358 36268 91398 36308
rect 91440 36268 91480 36308
rect 95112 36268 95152 36308
rect 95194 36268 95234 36308
rect 95276 36268 95316 36308
rect 95358 36268 95398 36308
rect 95440 36268 95480 36308
rect 99112 36268 99152 36308
rect 99194 36268 99234 36308
rect 99276 36268 99316 36308
rect 99358 36268 99398 36308
rect 99440 36268 99480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 8352 35512 8392 35552
rect 8434 35512 8474 35552
rect 8516 35512 8556 35552
rect 8598 35512 8638 35552
rect 8680 35512 8720 35552
rect 12352 35512 12392 35552
rect 12434 35512 12474 35552
rect 12516 35512 12556 35552
rect 12598 35512 12638 35552
rect 12680 35512 12720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 20352 35512 20392 35552
rect 20434 35512 20474 35552
rect 20516 35512 20556 35552
rect 20598 35512 20638 35552
rect 20680 35512 20720 35552
rect 24352 35512 24392 35552
rect 24434 35512 24474 35552
rect 24516 35512 24556 35552
rect 24598 35512 24638 35552
rect 24680 35512 24720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 32352 35512 32392 35552
rect 32434 35512 32474 35552
rect 32516 35512 32556 35552
rect 32598 35512 32638 35552
rect 32680 35512 32720 35552
rect 36352 35512 36392 35552
rect 36434 35512 36474 35552
rect 36516 35512 36556 35552
rect 36598 35512 36638 35552
rect 36680 35512 36720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 44352 35512 44392 35552
rect 44434 35512 44474 35552
rect 44516 35512 44556 35552
rect 44598 35512 44638 35552
rect 44680 35512 44720 35552
rect 48352 35512 48392 35552
rect 48434 35512 48474 35552
rect 48516 35512 48556 35552
rect 48598 35512 48638 35552
rect 48680 35512 48720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 56352 35512 56392 35552
rect 56434 35512 56474 35552
rect 56516 35512 56556 35552
rect 56598 35512 56638 35552
rect 56680 35512 56720 35552
rect 60352 35512 60392 35552
rect 60434 35512 60474 35552
rect 60516 35512 60556 35552
rect 60598 35512 60638 35552
rect 60680 35512 60720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 68352 35512 68392 35552
rect 68434 35512 68474 35552
rect 68516 35512 68556 35552
rect 68598 35512 68638 35552
rect 68680 35512 68720 35552
rect 72352 35512 72392 35552
rect 72434 35512 72474 35552
rect 72516 35512 72556 35552
rect 72598 35512 72638 35552
rect 72680 35512 72720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 80352 35512 80392 35552
rect 80434 35512 80474 35552
rect 80516 35512 80556 35552
rect 80598 35512 80638 35552
rect 80680 35512 80720 35552
rect 84352 35512 84392 35552
rect 84434 35512 84474 35552
rect 84516 35512 84556 35552
rect 84598 35512 84638 35552
rect 84680 35512 84720 35552
rect 88352 35512 88392 35552
rect 88434 35512 88474 35552
rect 88516 35512 88556 35552
rect 88598 35512 88638 35552
rect 88680 35512 88720 35552
rect 92352 35512 92392 35552
rect 92434 35512 92474 35552
rect 92516 35512 92556 35552
rect 92598 35512 92638 35552
rect 92680 35512 92720 35552
rect 96352 35512 96392 35552
rect 96434 35512 96474 35552
rect 96516 35512 96556 35552
rect 96598 35512 96638 35552
rect 96680 35512 96720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 7112 34756 7152 34796
rect 7194 34756 7234 34796
rect 7276 34756 7316 34796
rect 7358 34756 7398 34796
rect 7440 34756 7480 34796
rect 11112 34756 11152 34796
rect 11194 34756 11234 34796
rect 11276 34756 11316 34796
rect 11358 34756 11398 34796
rect 11440 34756 11480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 19112 34756 19152 34796
rect 19194 34756 19234 34796
rect 19276 34756 19316 34796
rect 19358 34756 19398 34796
rect 19440 34756 19480 34796
rect 23112 34756 23152 34796
rect 23194 34756 23234 34796
rect 23276 34756 23316 34796
rect 23358 34756 23398 34796
rect 23440 34756 23480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 31112 34756 31152 34796
rect 31194 34756 31234 34796
rect 31276 34756 31316 34796
rect 31358 34756 31398 34796
rect 31440 34756 31480 34796
rect 35112 34756 35152 34796
rect 35194 34756 35234 34796
rect 35276 34756 35316 34796
rect 35358 34756 35398 34796
rect 35440 34756 35480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 43112 34756 43152 34796
rect 43194 34756 43234 34796
rect 43276 34756 43316 34796
rect 43358 34756 43398 34796
rect 43440 34756 43480 34796
rect 47112 34756 47152 34796
rect 47194 34756 47234 34796
rect 47276 34756 47316 34796
rect 47358 34756 47398 34796
rect 47440 34756 47480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 55112 34756 55152 34796
rect 55194 34756 55234 34796
rect 55276 34756 55316 34796
rect 55358 34756 55398 34796
rect 55440 34756 55480 34796
rect 59112 34756 59152 34796
rect 59194 34756 59234 34796
rect 59276 34756 59316 34796
rect 59358 34756 59398 34796
rect 59440 34756 59480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 67112 34756 67152 34796
rect 67194 34756 67234 34796
rect 67276 34756 67316 34796
rect 67358 34756 67398 34796
rect 67440 34756 67480 34796
rect 71112 34756 71152 34796
rect 71194 34756 71234 34796
rect 71276 34756 71316 34796
rect 71358 34756 71398 34796
rect 71440 34756 71480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 79112 34756 79152 34796
rect 79194 34756 79234 34796
rect 79276 34756 79316 34796
rect 79358 34756 79398 34796
rect 79440 34756 79480 34796
rect 83112 34756 83152 34796
rect 83194 34756 83234 34796
rect 83276 34756 83316 34796
rect 83358 34756 83398 34796
rect 83440 34756 83480 34796
rect 87112 34756 87152 34796
rect 87194 34756 87234 34796
rect 87276 34756 87316 34796
rect 87358 34756 87398 34796
rect 87440 34756 87480 34796
rect 91112 34756 91152 34796
rect 91194 34756 91234 34796
rect 91276 34756 91316 34796
rect 91358 34756 91398 34796
rect 91440 34756 91480 34796
rect 95112 34756 95152 34796
rect 95194 34756 95234 34796
rect 95276 34756 95316 34796
rect 95358 34756 95398 34796
rect 95440 34756 95480 34796
rect 99112 34756 99152 34796
rect 99194 34756 99234 34796
rect 99276 34756 99316 34796
rect 99358 34756 99398 34796
rect 99440 34756 99480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 8352 34000 8392 34040
rect 8434 34000 8474 34040
rect 8516 34000 8556 34040
rect 8598 34000 8638 34040
rect 8680 34000 8720 34040
rect 12352 34000 12392 34040
rect 12434 34000 12474 34040
rect 12516 34000 12556 34040
rect 12598 34000 12638 34040
rect 12680 34000 12720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 20352 34000 20392 34040
rect 20434 34000 20474 34040
rect 20516 34000 20556 34040
rect 20598 34000 20638 34040
rect 20680 34000 20720 34040
rect 24352 34000 24392 34040
rect 24434 34000 24474 34040
rect 24516 34000 24556 34040
rect 24598 34000 24638 34040
rect 24680 34000 24720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 32352 34000 32392 34040
rect 32434 34000 32474 34040
rect 32516 34000 32556 34040
rect 32598 34000 32638 34040
rect 32680 34000 32720 34040
rect 36352 34000 36392 34040
rect 36434 34000 36474 34040
rect 36516 34000 36556 34040
rect 36598 34000 36638 34040
rect 36680 34000 36720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 44352 34000 44392 34040
rect 44434 34000 44474 34040
rect 44516 34000 44556 34040
rect 44598 34000 44638 34040
rect 44680 34000 44720 34040
rect 48352 34000 48392 34040
rect 48434 34000 48474 34040
rect 48516 34000 48556 34040
rect 48598 34000 48638 34040
rect 48680 34000 48720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 56352 34000 56392 34040
rect 56434 34000 56474 34040
rect 56516 34000 56556 34040
rect 56598 34000 56638 34040
rect 56680 34000 56720 34040
rect 60352 34000 60392 34040
rect 60434 34000 60474 34040
rect 60516 34000 60556 34040
rect 60598 34000 60638 34040
rect 60680 34000 60720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 68352 34000 68392 34040
rect 68434 34000 68474 34040
rect 68516 34000 68556 34040
rect 68598 34000 68638 34040
rect 68680 34000 68720 34040
rect 87052 33412 87092 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 7112 33244 7152 33284
rect 7194 33244 7234 33284
rect 7276 33244 7316 33284
rect 7358 33244 7398 33284
rect 7440 33244 7480 33284
rect 11112 33244 11152 33284
rect 11194 33244 11234 33284
rect 11276 33244 11316 33284
rect 11358 33244 11398 33284
rect 11440 33244 11480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 19112 33244 19152 33284
rect 19194 33244 19234 33284
rect 19276 33244 19316 33284
rect 19358 33244 19398 33284
rect 19440 33244 19480 33284
rect 23112 33244 23152 33284
rect 23194 33244 23234 33284
rect 23276 33244 23316 33284
rect 23358 33244 23398 33284
rect 23440 33244 23480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 31112 33244 31152 33284
rect 31194 33244 31234 33284
rect 31276 33244 31316 33284
rect 31358 33244 31398 33284
rect 31440 33244 31480 33284
rect 35112 33244 35152 33284
rect 35194 33244 35234 33284
rect 35276 33244 35316 33284
rect 35358 33244 35398 33284
rect 35440 33244 35480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 43112 33244 43152 33284
rect 43194 33244 43234 33284
rect 43276 33244 43316 33284
rect 43358 33244 43398 33284
rect 43440 33244 43480 33284
rect 47112 33244 47152 33284
rect 47194 33244 47234 33284
rect 47276 33244 47316 33284
rect 47358 33244 47398 33284
rect 47440 33244 47480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 55112 33244 55152 33284
rect 55194 33244 55234 33284
rect 55276 33244 55316 33284
rect 55358 33244 55398 33284
rect 55440 33244 55480 33284
rect 59112 33244 59152 33284
rect 59194 33244 59234 33284
rect 59276 33244 59316 33284
rect 59358 33244 59398 33284
rect 59440 33244 59480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 67112 33244 67152 33284
rect 67194 33244 67234 33284
rect 67276 33244 67316 33284
rect 67358 33244 67398 33284
rect 67440 33244 67480 33284
rect 73612 32824 73652 32864
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 8352 32488 8392 32528
rect 8434 32488 8474 32528
rect 8516 32488 8556 32528
rect 8598 32488 8638 32528
rect 8680 32488 8720 32528
rect 12352 32488 12392 32528
rect 12434 32488 12474 32528
rect 12516 32488 12556 32528
rect 12598 32488 12638 32528
rect 12680 32488 12720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 20352 32488 20392 32528
rect 20434 32488 20474 32528
rect 20516 32488 20556 32528
rect 20598 32488 20638 32528
rect 20680 32488 20720 32528
rect 24352 32488 24392 32528
rect 24434 32488 24474 32528
rect 24516 32488 24556 32528
rect 24598 32488 24638 32528
rect 24680 32488 24720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 32352 32488 32392 32528
rect 32434 32488 32474 32528
rect 32516 32488 32556 32528
rect 32598 32488 32638 32528
rect 32680 32488 32720 32528
rect 36352 32488 36392 32528
rect 36434 32488 36474 32528
rect 36516 32488 36556 32528
rect 36598 32488 36638 32528
rect 36680 32488 36720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 44352 32488 44392 32528
rect 44434 32488 44474 32528
rect 44516 32488 44556 32528
rect 44598 32488 44638 32528
rect 44680 32488 44720 32528
rect 48352 32488 48392 32528
rect 48434 32488 48474 32528
rect 48516 32488 48556 32528
rect 48598 32488 48638 32528
rect 48680 32488 48720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 56352 32488 56392 32528
rect 56434 32488 56474 32528
rect 56516 32488 56556 32528
rect 56598 32488 56638 32528
rect 56680 32488 56720 32528
rect 60352 32488 60392 32528
rect 60434 32488 60474 32528
rect 60516 32488 60556 32528
rect 60598 32488 60638 32528
rect 60680 32488 60720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 68352 32488 68392 32528
rect 68434 32488 68474 32528
rect 68516 32488 68556 32528
rect 68598 32488 68638 32528
rect 68680 32488 68720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 7112 31732 7152 31772
rect 7194 31732 7234 31772
rect 7276 31732 7316 31772
rect 7358 31732 7398 31772
rect 7440 31732 7480 31772
rect 11112 31732 11152 31772
rect 11194 31732 11234 31772
rect 11276 31732 11316 31772
rect 11358 31732 11398 31772
rect 11440 31732 11480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 19112 31732 19152 31772
rect 19194 31732 19234 31772
rect 19276 31732 19316 31772
rect 19358 31732 19398 31772
rect 19440 31732 19480 31772
rect 23112 31732 23152 31772
rect 23194 31732 23234 31772
rect 23276 31732 23316 31772
rect 23358 31732 23398 31772
rect 23440 31732 23480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 31112 31732 31152 31772
rect 31194 31732 31234 31772
rect 31276 31732 31316 31772
rect 31358 31732 31398 31772
rect 31440 31732 31480 31772
rect 35112 31732 35152 31772
rect 35194 31732 35234 31772
rect 35276 31732 35316 31772
rect 35358 31732 35398 31772
rect 35440 31732 35480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 43112 31732 43152 31772
rect 43194 31732 43234 31772
rect 43276 31732 43316 31772
rect 43358 31732 43398 31772
rect 43440 31732 43480 31772
rect 47112 31732 47152 31772
rect 47194 31732 47234 31772
rect 47276 31732 47316 31772
rect 47358 31732 47398 31772
rect 47440 31732 47480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 55112 31732 55152 31772
rect 55194 31732 55234 31772
rect 55276 31732 55316 31772
rect 55358 31732 55398 31772
rect 55440 31732 55480 31772
rect 59112 31732 59152 31772
rect 59194 31732 59234 31772
rect 59276 31732 59316 31772
rect 59358 31732 59398 31772
rect 59440 31732 59480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 67112 31732 67152 31772
rect 67194 31732 67234 31772
rect 67276 31732 67316 31772
rect 67358 31732 67398 31772
rect 67440 31732 67480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 8352 30976 8392 31016
rect 8434 30976 8474 31016
rect 8516 30976 8556 31016
rect 8598 30976 8638 31016
rect 8680 30976 8720 31016
rect 12352 30976 12392 31016
rect 12434 30976 12474 31016
rect 12516 30976 12556 31016
rect 12598 30976 12638 31016
rect 12680 30976 12720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 20352 30976 20392 31016
rect 20434 30976 20474 31016
rect 20516 30976 20556 31016
rect 20598 30976 20638 31016
rect 20680 30976 20720 31016
rect 24352 30976 24392 31016
rect 24434 30976 24474 31016
rect 24516 30976 24556 31016
rect 24598 30976 24638 31016
rect 24680 30976 24720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 32352 30976 32392 31016
rect 32434 30976 32474 31016
rect 32516 30976 32556 31016
rect 32598 30976 32638 31016
rect 32680 30976 32720 31016
rect 36352 30976 36392 31016
rect 36434 30976 36474 31016
rect 36516 30976 36556 31016
rect 36598 30976 36638 31016
rect 36680 30976 36720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 44352 30976 44392 31016
rect 44434 30976 44474 31016
rect 44516 30976 44556 31016
rect 44598 30976 44638 31016
rect 44680 30976 44720 31016
rect 48352 30976 48392 31016
rect 48434 30976 48474 31016
rect 48516 30976 48556 31016
rect 48598 30976 48638 31016
rect 48680 30976 48720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 56352 30976 56392 31016
rect 56434 30976 56474 31016
rect 56516 30976 56556 31016
rect 56598 30976 56638 31016
rect 56680 30976 56720 31016
rect 60352 30976 60392 31016
rect 60434 30976 60474 31016
rect 60516 30976 60556 31016
rect 60598 30976 60638 31016
rect 60680 30976 60720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 68352 30976 68392 31016
rect 68434 30976 68474 31016
rect 68516 30976 68556 31016
rect 68598 30976 68638 31016
rect 68680 30976 68720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 7112 30220 7152 30260
rect 7194 30220 7234 30260
rect 7276 30220 7316 30260
rect 7358 30220 7398 30260
rect 7440 30220 7480 30260
rect 11112 30220 11152 30260
rect 11194 30220 11234 30260
rect 11276 30220 11316 30260
rect 11358 30220 11398 30260
rect 11440 30220 11480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 19112 30220 19152 30260
rect 19194 30220 19234 30260
rect 19276 30220 19316 30260
rect 19358 30220 19398 30260
rect 19440 30220 19480 30260
rect 23112 30220 23152 30260
rect 23194 30220 23234 30260
rect 23276 30220 23316 30260
rect 23358 30220 23398 30260
rect 23440 30220 23480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 31112 30220 31152 30260
rect 31194 30220 31234 30260
rect 31276 30220 31316 30260
rect 31358 30220 31398 30260
rect 31440 30220 31480 30260
rect 35112 30220 35152 30260
rect 35194 30220 35234 30260
rect 35276 30220 35316 30260
rect 35358 30220 35398 30260
rect 35440 30220 35480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 43112 30220 43152 30260
rect 43194 30220 43234 30260
rect 43276 30220 43316 30260
rect 43358 30220 43398 30260
rect 43440 30220 43480 30260
rect 47112 30220 47152 30260
rect 47194 30220 47234 30260
rect 47276 30220 47316 30260
rect 47358 30220 47398 30260
rect 47440 30220 47480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 55112 30220 55152 30260
rect 55194 30220 55234 30260
rect 55276 30220 55316 30260
rect 55358 30220 55398 30260
rect 55440 30220 55480 30260
rect 59112 30220 59152 30260
rect 59194 30220 59234 30260
rect 59276 30220 59316 30260
rect 59358 30220 59398 30260
rect 59440 30220 59480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 67112 30220 67152 30260
rect 67194 30220 67234 30260
rect 67276 30220 67316 30260
rect 67358 30220 67398 30260
rect 67440 30220 67480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 8352 29464 8392 29504
rect 8434 29464 8474 29504
rect 8516 29464 8556 29504
rect 8598 29464 8638 29504
rect 8680 29464 8720 29504
rect 12352 29464 12392 29504
rect 12434 29464 12474 29504
rect 12516 29464 12556 29504
rect 12598 29464 12638 29504
rect 12680 29464 12720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 20352 29464 20392 29504
rect 20434 29464 20474 29504
rect 20516 29464 20556 29504
rect 20598 29464 20638 29504
rect 20680 29464 20720 29504
rect 24352 29464 24392 29504
rect 24434 29464 24474 29504
rect 24516 29464 24556 29504
rect 24598 29464 24638 29504
rect 24680 29464 24720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 32352 29464 32392 29504
rect 32434 29464 32474 29504
rect 32516 29464 32556 29504
rect 32598 29464 32638 29504
rect 32680 29464 32720 29504
rect 36352 29464 36392 29504
rect 36434 29464 36474 29504
rect 36516 29464 36556 29504
rect 36598 29464 36638 29504
rect 36680 29464 36720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 44352 29464 44392 29504
rect 44434 29464 44474 29504
rect 44516 29464 44556 29504
rect 44598 29464 44638 29504
rect 44680 29464 44720 29504
rect 48352 29464 48392 29504
rect 48434 29464 48474 29504
rect 48516 29464 48556 29504
rect 48598 29464 48638 29504
rect 48680 29464 48720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 56352 29464 56392 29504
rect 56434 29464 56474 29504
rect 56516 29464 56556 29504
rect 56598 29464 56638 29504
rect 56680 29464 56720 29504
rect 60352 29464 60392 29504
rect 60434 29464 60474 29504
rect 60516 29464 60556 29504
rect 60598 29464 60638 29504
rect 60680 29464 60720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 68352 29464 68392 29504
rect 68434 29464 68474 29504
rect 68516 29464 68556 29504
rect 68598 29464 68638 29504
rect 68680 29464 68720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 7112 28708 7152 28748
rect 7194 28708 7234 28748
rect 7276 28708 7316 28748
rect 7358 28708 7398 28748
rect 7440 28708 7480 28748
rect 11112 28708 11152 28748
rect 11194 28708 11234 28748
rect 11276 28708 11316 28748
rect 11358 28708 11398 28748
rect 11440 28708 11480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 19112 28708 19152 28748
rect 19194 28708 19234 28748
rect 19276 28708 19316 28748
rect 19358 28708 19398 28748
rect 19440 28708 19480 28748
rect 23112 28708 23152 28748
rect 23194 28708 23234 28748
rect 23276 28708 23316 28748
rect 23358 28708 23398 28748
rect 23440 28708 23480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 31112 28708 31152 28748
rect 31194 28708 31234 28748
rect 31276 28708 31316 28748
rect 31358 28708 31398 28748
rect 31440 28708 31480 28748
rect 35112 28708 35152 28748
rect 35194 28708 35234 28748
rect 35276 28708 35316 28748
rect 35358 28708 35398 28748
rect 35440 28708 35480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 43112 28708 43152 28748
rect 43194 28708 43234 28748
rect 43276 28708 43316 28748
rect 43358 28708 43398 28748
rect 43440 28708 43480 28748
rect 47112 28708 47152 28748
rect 47194 28708 47234 28748
rect 47276 28708 47316 28748
rect 47358 28708 47398 28748
rect 47440 28708 47480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 55112 28708 55152 28748
rect 55194 28708 55234 28748
rect 55276 28708 55316 28748
rect 55358 28708 55398 28748
rect 55440 28708 55480 28748
rect 59112 28708 59152 28748
rect 59194 28708 59234 28748
rect 59276 28708 59316 28748
rect 59358 28708 59398 28748
rect 59440 28708 59480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 67112 28708 67152 28748
rect 67194 28708 67234 28748
rect 67276 28708 67316 28748
rect 67358 28708 67398 28748
rect 67440 28708 67480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 8352 27952 8392 27992
rect 8434 27952 8474 27992
rect 8516 27952 8556 27992
rect 8598 27952 8638 27992
rect 8680 27952 8720 27992
rect 12352 27952 12392 27992
rect 12434 27952 12474 27992
rect 12516 27952 12556 27992
rect 12598 27952 12638 27992
rect 12680 27952 12720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 20352 27952 20392 27992
rect 20434 27952 20474 27992
rect 20516 27952 20556 27992
rect 20598 27952 20638 27992
rect 20680 27952 20720 27992
rect 24352 27952 24392 27992
rect 24434 27952 24474 27992
rect 24516 27952 24556 27992
rect 24598 27952 24638 27992
rect 24680 27952 24720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 32352 27952 32392 27992
rect 32434 27952 32474 27992
rect 32516 27952 32556 27992
rect 32598 27952 32638 27992
rect 32680 27952 32720 27992
rect 36352 27952 36392 27992
rect 36434 27952 36474 27992
rect 36516 27952 36556 27992
rect 36598 27952 36638 27992
rect 36680 27952 36720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 44352 27952 44392 27992
rect 44434 27952 44474 27992
rect 44516 27952 44556 27992
rect 44598 27952 44638 27992
rect 44680 27952 44720 27992
rect 48352 27952 48392 27992
rect 48434 27952 48474 27992
rect 48516 27952 48556 27992
rect 48598 27952 48638 27992
rect 48680 27952 48720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 56352 27952 56392 27992
rect 56434 27952 56474 27992
rect 56516 27952 56556 27992
rect 56598 27952 56638 27992
rect 56680 27952 56720 27992
rect 60352 27952 60392 27992
rect 60434 27952 60474 27992
rect 60516 27952 60556 27992
rect 60598 27952 60638 27992
rect 60680 27952 60720 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 68352 27952 68392 27992
rect 68434 27952 68474 27992
rect 68516 27952 68556 27992
rect 68598 27952 68638 27992
rect 68680 27952 68720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 7112 27196 7152 27236
rect 7194 27196 7234 27236
rect 7276 27196 7316 27236
rect 7358 27196 7398 27236
rect 7440 27196 7480 27236
rect 11112 27196 11152 27236
rect 11194 27196 11234 27236
rect 11276 27196 11316 27236
rect 11358 27196 11398 27236
rect 11440 27196 11480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 19112 27196 19152 27236
rect 19194 27196 19234 27236
rect 19276 27196 19316 27236
rect 19358 27196 19398 27236
rect 19440 27196 19480 27236
rect 23112 27196 23152 27236
rect 23194 27196 23234 27236
rect 23276 27196 23316 27236
rect 23358 27196 23398 27236
rect 23440 27196 23480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 31112 27196 31152 27236
rect 31194 27196 31234 27236
rect 31276 27196 31316 27236
rect 31358 27196 31398 27236
rect 31440 27196 31480 27236
rect 35112 27196 35152 27236
rect 35194 27196 35234 27236
rect 35276 27196 35316 27236
rect 35358 27196 35398 27236
rect 35440 27196 35480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 43112 27196 43152 27236
rect 43194 27196 43234 27236
rect 43276 27196 43316 27236
rect 43358 27196 43398 27236
rect 43440 27196 43480 27236
rect 47112 27196 47152 27236
rect 47194 27196 47234 27236
rect 47276 27196 47316 27236
rect 47358 27196 47398 27236
rect 47440 27196 47480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 55112 27196 55152 27236
rect 55194 27196 55234 27236
rect 55276 27196 55316 27236
rect 55358 27196 55398 27236
rect 55440 27196 55480 27236
rect 59112 27196 59152 27236
rect 59194 27196 59234 27236
rect 59276 27196 59316 27236
rect 59358 27196 59398 27236
rect 59440 27196 59480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 67112 27196 67152 27236
rect 67194 27196 67234 27236
rect 67276 27196 67316 27236
rect 67358 27196 67398 27236
rect 67440 27196 67480 27236
rect 71884 26776 71924 26816
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 8352 26440 8392 26480
rect 8434 26440 8474 26480
rect 8516 26440 8556 26480
rect 8598 26440 8638 26480
rect 8680 26440 8720 26480
rect 12352 26440 12392 26480
rect 12434 26440 12474 26480
rect 12516 26440 12556 26480
rect 12598 26440 12638 26480
rect 12680 26440 12720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 20352 26440 20392 26480
rect 20434 26440 20474 26480
rect 20516 26440 20556 26480
rect 20598 26440 20638 26480
rect 20680 26440 20720 26480
rect 24352 26440 24392 26480
rect 24434 26440 24474 26480
rect 24516 26440 24556 26480
rect 24598 26440 24638 26480
rect 24680 26440 24720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 32352 26440 32392 26480
rect 32434 26440 32474 26480
rect 32516 26440 32556 26480
rect 32598 26440 32638 26480
rect 32680 26440 32720 26480
rect 36352 26440 36392 26480
rect 36434 26440 36474 26480
rect 36516 26440 36556 26480
rect 36598 26440 36638 26480
rect 36680 26440 36720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 44352 26440 44392 26480
rect 44434 26440 44474 26480
rect 44516 26440 44556 26480
rect 44598 26440 44638 26480
rect 44680 26440 44720 26480
rect 48352 26440 48392 26480
rect 48434 26440 48474 26480
rect 48516 26440 48556 26480
rect 48598 26440 48638 26480
rect 48680 26440 48720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 56352 26440 56392 26480
rect 56434 26440 56474 26480
rect 56516 26440 56556 26480
rect 56598 26440 56638 26480
rect 56680 26440 56720 26480
rect 60352 26440 60392 26480
rect 60434 26440 60474 26480
rect 60516 26440 60556 26480
rect 60598 26440 60638 26480
rect 60680 26440 60720 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 68352 26440 68392 26480
rect 68434 26440 68474 26480
rect 68516 26440 68556 26480
rect 68598 26440 68638 26480
rect 68680 26440 68720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 7112 25684 7152 25724
rect 7194 25684 7234 25724
rect 7276 25684 7316 25724
rect 7358 25684 7398 25724
rect 7440 25684 7480 25724
rect 11112 25684 11152 25724
rect 11194 25684 11234 25724
rect 11276 25684 11316 25724
rect 11358 25684 11398 25724
rect 11440 25684 11480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 19112 25684 19152 25724
rect 19194 25684 19234 25724
rect 19276 25684 19316 25724
rect 19358 25684 19398 25724
rect 19440 25684 19480 25724
rect 23112 25684 23152 25724
rect 23194 25684 23234 25724
rect 23276 25684 23316 25724
rect 23358 25684 23398 25724
rect 23440 25684 23480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 31112 25684 31152 25724
rect 31194 25684 31234 25724
rect 31276 25684 31316 25724
rect 31358 25684 31398 25724
rect 31440 25684 31480 25724
rect 35112 25684 35152 25724
rect 35194 25684 35234 25724
rect 35276 25684 35316 25724
rect 35358 25684 35398 25724
rect 35440 25684 35480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 43112 25684 43152 25724
rect 43194 25684 43234 25724
rect 43276 25684 43316 25724
rect 43358 25684 43398 25724
rect 43440 25684 43480 25724
rect 47112 25684 47152 25724
rect 47194 25684 47234 25724
rect 47276 25684 47316 25724
rect 47358 25684 47398 25724
rect 47440 25684 47480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 55112 25684 55152 25724
rect 55194 25684 55234 25724
rect 55276 25684 55316 25724
rect 55358 25684 55398 25724
rect 55440 25684 55480 25724
rect 59112 25684 59152 25724
rect 59194 25684 59234 25724
rect 59276 25684 59316 25724
rect 59358 25684 59398 25724
rect 59440 25684 59480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 67112 25684 67152 25724
rect 67194 25684 67234 25724
rect 67276 25684 67316 25724
rect 67358 25684 67398 25724
rect 67440 25684 67480 25724
rect 85708 25684 85748 25724
rect 86860 25348 86900 25388
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 8352 24928 8392 24968
rect 8434 24928 8474 24968
rect 8516 24928 8556 24968
rect 8598 24928 8638 24968
rect 8680 24928 8720 24968
rect 12352 24928 12392 24968
rect 12434 24928 12474 24968
rect 12516 24928 12556 24968
rect 12598 24928 12638 24968
rect 12680 24928 12720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 20352 24928 20392 24968
rect 20434 24928 20474 24968
rect 20516 24928 20556 24968
rect 20598 24928 20638 24968
rect 20680 24928 20720 24968
rect 24352 24928 24392 24968
rect 24434 24928 24474 24968
rect 24516 24928 24556 24968
rect 24598 24928 24638 24968
rect 24680 24928 24720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 32352 24928 32392 24968
rect 32434 24928 32474 24968
rect 32516 24928 32556 24968
rect 32598 24928 32638 24968
rect 32680 24928 32720 24968
rect 36352 24928 36392 24968
rect 36434 24928 36474 24968
rect 36516 24928 36556 24968
rect 36598 24928 36638 24968
rect 36680 24928 36720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 44352 24928 44392 24968
rect 44434 24928 44474 24968
rect 44516 24928 44556 24968
rect 44598 24928 44638 24968
rect 44680 24928 44720 24968
rect 48352 24928 48392 24968
rect 48434 24928 48474 24968
rect 48516 24928 48556 24968
rect 48598 24928 48638 24968
rect 48680 24928 48720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 56352 24928 56392 24968
rect 56434 24928 56474 24968
rect 56516 24928 56556 24968
rect 56598 24928 56638 24968
rect 56680 24928 56720 24968
rect 60352 24928 60392 24968
rect 60434 24928 60474 24968
rect 60516 24928 60556 24968
rect 60598 24928 60638 24968
rect 60680 24928 60720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 68352 24928 68392 24968
rect 68434 24928 68474 24968
rect 68516 24928 68556 24968
rect 68598 24928 68638 24968
rect 68680 24928 68720 24968
rect 73228 24592 73268 24632
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 7112 24172 7152 24212
rect 7194 24172 7234 24212
rect 7276 24172 7316 24212
rect 7358 24172 7398 24212
rect 7440 24172 7480 24212
rect 11112 24172 11152 24212
rect 11194 24172 11234 24212
rect 11276 24172 11316 24212
rect 11358 24172 11398 24212
rect 11440 24172 11480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 19112 24172 19152 24212
rect 19194 24172 19234 24212
rect 19276 24172 19316 24212
rect 19358 24172 19398 24212
rect 19440 24172 19480 24212
rect 23112 24172 23152 24212
rect 23194 24172 23234 24212
rect 23276 24172 23316 24212
rect 23358 24172 23398 24212
rect 23440 24172 23480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 31112 24172 31152 24212
rect 31194 24172 31234 24212
rect 31276 24172 31316 24212
rect 31358 24172 31398 24212
rect 31440 24172 31480 24212
rect 35112 24172 35152 24212
rect 35194 24172 35234 24212
rect 35276 24172 35316 24212
rect 35358 24172 35398 24212
rect 35440 24172 35480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 43112 24172 43152 24212
rect 43194 24172 43234 24212
rect 43276 24172 43316 24212
rect 43358 24172 43398 24212
rect 43440 24172 43480 24212
rect 47112 24172 47152 24212
rect 47194 24172 47234 24212
rect 47276 24172 47316 24212
rect 47358 24172 47398 24212
rect 47440 24172 47480 24212
rect 51112 24172 51152 24212
rect 51194 24172 51234 24212
rect 51276 24172 51316 24212
rect 51358 24172 51398 24212
rect 51440 24172 51480 24212
rect 55112 24172 55152 24212
rect 55194 24172 55234 24212
rect 55276 24172 55316 24212
rect 55358 24172 55398 24212
rect 55440 24172 55480 24212
rect 59112 24172 59152 24212
rect 59194 24172 59234 24212
rect 59276 24172 59316 24212
rect 59358 24172 59398 24212
rect 59440 24172 59480 24212
rect 63112 24172 63152 24212
rect 63194 24172 63234 24212
rect 63276 24172 63316 24212
rect 63358 24172 63398 24212
rect 63440 24172 63480 24212
rect 67112 24172 67152 24212
rect 67194 24172 67234 24212
rect 67276 24172 67316 24212
rect 67358 24172 67398 24212
rect 67440 24172 67480 24212
rect 71112 24172 71152 24212
rect 71194 24172 71234 24212
rect 71276 24172 71316 24212
rect 71358 24172 71398 24212
rect 71440 24172 71480 24212
rect 75112 24172 75152 24212
rect 75194 24172 75234 24212
rect 75276 24172 75316 24212
rect 75358 24172 75398 24212
rect 75440 24172 75480 24212
rect 79112 24172 79152 24212
rect 79194 24172 79234 24212
rect 79276 24172 79316 24212
rect 79358 24172 79398 24212
rect 79440 24172 79480 24212
rect 83112 24172 83152 24212
rect 83194 24172 83234 24212
rect 83276 24172 83316 24212
rect 83358 24172 83398 24212
rect 83440 24172 83480 24212
rect 87112 24172 87152 24212
rect 87194 24172 87234 24212
rect 87276 24172 87316 24212
rect 87358 24172 87398 24212
rect 87440 24172 87480 24212
rect 91112 24172 91152 24212
rect 91194 24172 91234 24212
rect 91276 24172 91316 24212
rect 91358 24172 91398 24212
rect 91440 24172 91480 24212
rect 95112 24172 95152 24212
rect 95194 24172 95234 24212
rect 95276 24172 95316 24212
rect 95358 24172 95398 24212
rect 95440 24172 95480 24212
rect 99112 24172 99152 24212
rect 99194 24172 99234 24212
rect 99276 24172 99316 24212
rect 99358 24172 99398 24212
rect 99440 24172 99480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 8352 23416 8392 23456
rect 8434 23416 8474 23456
rect 8516 23416 8556 23456
rect 8598 23416 8638 23456
rect 8680 23416 8720 23456
rect 12352 23416 12392 23456
rect 12434 23416 12474 23456
rect 12516 23416 12556 23456
rect 12598 23416 12638 23456
rect 12680 23416 12720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 20352 23416 20392 23456
rect 20434 23416 20474 23456
rect 20516 23416 20556 23456
rect 20598 23416 20638 23456
rect 20680 23416 20720 23456
rect 24352 23416 24392 23456
rect 24434 23416 24474 23456
rect 24516 23416 24556 23456
rect 24598 23416 24638 23456
rect 24680 23416 24720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 32352 23416 32392 23456
rect 32434 23416 32474 23456
rect 32516 23416 32556 23456
rect 32598 23416 32638 23456
rect 32680 23416 32720 23456
rect 36352 23416 36392 23456
rect 36434 23416 36474 23456
rect 36516 23416 36556 23456
rect 36598 23416 36638 23456
rect 36680 23416 36720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 44352 23416 44392 23456
rect 44434 23416 44474 23456
rect 44516 23416 44556 23456
rect 44598 23416 44638 23456
rect 44680 23416 44720 23456
rect 48352 23416 48392 23456
rect 48434 23416 48474 23456
rect 48516 23416 48556 23456
rect 48598 23416 48638 23456
rect 48680 23416 48720 23456
rect 52352 23416 52392 23456
rect 52434 23416 52474 23456
rect 52516 23416 52556 23456
rect 52598 23416 52638 23456
rect 52680 23416 52720 23456
rect 56352 23416 56392 23456
rect 56434 23416 56474 23456
rect 56516 23416 56556 23456
rect 56598 23416 56638 23456
rect 56680 23416 56720 23456
rect 60352 23416 60392 23456
rect 60434 23416 60474 23456
rect 60516 23416 60556 23456
rect 60598 23416 60638 23456
rect 60680 23416 60720 23456
rect 64352 23416 64392 23456
rect 64434 23416 64474 23456
rect 64516 23416 64556 23456
rect 64598 23416 64638 23456
rect 64680 23416 64720 23456
rect 68352 23416 68392 23456
rect 68434 23416 68474 23456
rect 68516 23416 68556 23456
rect 68598 23416 68638 23456
rect 68680 23416 68720 23456
rect 72352 23416 72392 23456
rect 72434 23416 72474 23456
rect 72516 23416 72556 23456
rect 72598 23416 72638 23456
rect 72680 23416 72720 23456
rect 76352 23416 76392 23456
rect 76434 23416 76474 23456
rect 76516 23416 76556 23456
rect 76598 23416 76638 23456
rect 76680 23416 76720 23456
rect 80352 23416 80392 23456
rect 80434 23416 80474 23456
rect 80516 23416 80556 23456
rect 80598 23416 80638 23456
rect 80680 23416 80720 23456
rect 84352 23416 84392 23456
rect 84434 23416 84474 23456
rect 84516 23416 84556 23456
rect 84598 23416 84638 23456
rect 84680 23416 84720 23456
rect 88352 23416 88392 23456
rect 88434 23416 88474 23456
rect 88516 23416 88556 23456
rect 88598 23416 88638 23456
rect 88680 23416 88720 23456
rect 92352 23416 92392 23456
rect 92434 23416 92474 23456
rect 92516 23416 92556 23456
rect 92598 23416 92638 23456
rect 92680 23416 92720 23456
rect 96352 23416 96392 23456
rect 96434 23416 96474 23456
rect 96516 23416 96556 23456
rect 96598 23416 96638 23456
rect 96680 23416 96720 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 7112 22660 7152 22700
rect 7194 22660 7234 22700
rect 7276 22660 7316 22700
rect 7358 22660 7398 22700
rect 7440 22660 7480 22700
rect 11112 22660 11152 22700
rect 11194 22660 11234 22700
rect 11276 22660 11316 22700
rect 11358 22660 11398 22700
rect 11440 22660 11480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 19112 22660 19152 22700
rect 19194 22660 19234 22700
rect 19276 22660 19316 22700
rect 19358 22660 19398 22700
rect 19440 22660 19480 22700
rect 23112 22660 23152 22700
rect 23194 22660 23234 22700
rect 23276 22660 23316 22700
rect 23358 22660 23398 22700
rect 23440 22660 23480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 31112 22660 31152 22700
rect 31194 22660 31234 22700
rect 31276 22660 31316 22700
rect 31358 22660 31398 22700
rect 31440 22660 31480 22700
rect 35112 22660 35152 22700
rect 35194 22660 35234 22700
rect 35276 22660 35316 22700
rect 35358 22660 35398 22700
rect 35440 22660 35480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 43112 22660 43152 22700
rect 43194 22660 43234 22700
rect 43276 22660 43316 22700
rect 43358 22660 43398 22700
rect 43440 22660 43480 22700
rect 47112 22660 47152 22700
rect 47194 22660 47234 22700
rect 47276 22660 47316 22700
rect 47358 22660 47398 22700
rect 47440 22660 47480 22700
rect 51112 22660 51152 22700
rect 51194 22660 51234 22700
rect 51276 22660 51316 22700
rect 51358 22660 51398 22700
rect 51440 22660 51480 22700
rect 55112 22660 55152 22700
rect 55194 22660 55234 22700
rect 55276 22660 55316 22700
rect 55358 22660 55398 22700
rect 55440 22660 55480 22700
rect 59112 22660 59152 22700
rect 59194 22660 59234 22700
rect 59276 22660 59316 22700
rect 59358 22660 59398 22700
rect 59440 22660 59480 22700
rect 63112 22660 63152 22700
rect 63194 22660 63234 22700
rect 63276 22660 63316 22700
rect 63358 22660 63398 22700
rect 63440 22660 63480 22700
rect 67112 22660 67152 22700
rect 67194 22660 67234 22700
rect 67276 22660 67316 22700
rect 67358 22660 67398 22700
rect 67440 22660 67480 22700
rect 71112 22660 71152 22700
rect 71194 22660 71234 22700
rect 71276 22660 71316 22700
rect 71358 22660 71398 22700
rect 71440 22660 71480 22700
rect 75112 22660 75152 22700
rect 75194 22660 75234 22700
rect 75276 22660 75316 22700
rect 75358 22660 75398 22700
rect 75440 22660 75480 22700
rect 79112 22660 79152 22700
rect 79194 22660 79234 22700
rect 79276 22660 79316 22700
rect 79358 22660 79398 22700
rect 79440 22660 79480 22700
rect 83112 22660 83152 22700
rect 83194 22660 83234 22700
rect 83276 22660 83316 22700
rect 83358 22660 83398 22700
rect 83440 22660 83480 22700
rect 87112 22660 87152 22700
rect 87194 22660 87234 22700
rect 87276 22660 87316 22700
rect 87358 22660 87398 22700
rect 87440 22660 87480 22700
rect 91112 22660 91152 22700
rect 91194 22660 91234 22700
rect 91276 22660 91316 22700
rect 91358 22660 91398 22700
rect 91440 22660 91480 22700
rect 95112 22660 95152 22700
rect 95194 22660 95234 22700
rect 95276 22660 95316 22700
rect 95358 22660 95398 22700
rect 95440 22660 95480 22700
rect 99112 22660 99152 22700
rect 99194 22660 99234 22700
rect 99276 22660 99316 22700
rect 99358 22660 99398 22700
rect 99440 22660 99480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 8352 21904 8392 21944
rect 8434 21904 8474 21944
rect 8516 21904 8556 21944
rect 8598 21904 8638 21944
rect 8680 21904 8720 21944
rect 12352 21904 12392 21944
rect 12434 21904 12474 21944
rect 12516 21904 12556 21944
rect 12598 21904 12638 21944
rect 12680 21904 12720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 20352 21904 20392 21944
rect 20434 21904 20474 21944
rect 20516 21904 20556 21944
rect 20598 21904 20638 21944
rect 20680 21904 20720 21944
rect 24352 21904 24392 21944
rect 24434 21904 24474 21944
rect 24516 21904 24556 21944
rect 24598 21904 24638 21944
rect 24680 21904 24720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 32352 21904 32392 21944
rect 32434 21904 32474 21944
rect 32516 21904 32556 21944
rect 32598 21904 32638 21944
rect 32680 21904 32720 21944
rect 36352 21904 36392 21944
rect 36434 21904 36474 21944
rect 36516 21904 36556 21944
rect 36598 21904 36638 21944
rect 36680 21904 36720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 44352 21904 44392 21944
rect 44434 21904 44474 21944
rect 44516 21904 44556 21944
rect 44598 21904 44638 21944
rect 44680 21904 44720 21944
rect 48352 21904 48392 21944
rect 48434 21904 48474 21944
rect 48516 21904 48556 21944
rect 48598 21904 48638 21944
rect 48680 21904 48720 21944
rect 52352 21904 52392 21944
rect 52434 21904 52474 21944
rect 52516 21904 52556 21944
rect 52598 21904 52638 21944
rect 52680 21904 52720 21944
rect 56352 21904 56392 21944
rect 56434 21904 56474 21944
rect 56516 21904 56556 21944
rect 56598 21904 56638 21944
rect 56680 21904 56720 21944
rect 60352 21904 60392 21944
rect 60434 21904 60474 21944
rect 60516 21904 60556 21944
rect 60598 21904 60638 21944
rect 60680 21904 60720 21944
rect 64352 21904 64392 21944
rect 64434 21904 64474 21944
rect 64516 21904 64556 21944
rect 64598 21904 64638 21944
rect 64680 21904 64720 21944
rect 68352 21904 68392 21944
rect 68434 21904 68474 21944
rect 68516 21904 68556 21944
rect 68598 21904 68638 21944
rect 68680 21904 68720 21944
rect 72352 21904 72392 21944
rect 72434 21904 72474 21944
rect 72516 21904 72556 21944
rect 72598 21904 72638 21944
rect 72680 21904 72720 21944
rect 76352 21904 76392 21944
rect 76434 21904 76474 21944
rect 76516 21904 76556 21944
rect 76598 21904 76638 21944
rect 76680 21904 76720 21944
rect 80352 21904 80392 21944
rect 80434 21904 80474 21944
rect 80516 21904 80556 21944
rect 80598 21904 80638 21944
rect 80680 21904 80720 21944
rect 84352 21904 84392 21944
rect 84434 21904 84474 21944
rect 84516 21904 84556 21944
rect 84598 21904 84638 21944
rect 84680 21904 84720 21944
rect 88352 21904 88392 21944
rect 88434 21904 88474 21944
rect 88516 21904 88556 21944
rect 88598 21904 88638 21944
rect 88680 21904 88720 21944
rect 92352 21904 92392 21944
rect 92434 21904 92474 21944
rect 92516 21904 92556 21944
rect 92598 21904 92638 21944
rect 92680 21904 92720 21944
rect 96352 21904 96392 21944
rect 96434 21904 96474 21944
rect 96516 21904 96556 21944
rect 96598 21904 96638 21944
rect 96680 21904 96720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 7112 21148 7152 21188
rect 7194 21148 7234 21188
rect 7276 21148 7316 21188
rect 7358 21148 7398 21188
rect 7440 21148 7480 21188
rect 11112 21148 11152 21188
rect 11194 21148 11234 21188
rect 11276 21148 11316 21188
rect 11358 21148 11398 21188
rect 11440 21148 11480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 19112 21148 19152 21188
rect 19194 21148 19234 21188
rect 19276 21148 19316 21188
rect 19358 21148 19398 21188
rect 19440 21148 19480 21188
rect 23112 21148 23152 21188
rect 23194 21148 23234 21188
rect 23276 21148 23316 21188
rect 23358 21148 23398 21188
rect 23440 21148 23480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 31112 21148 31152 21188
rect 31194 21148 31234 21188
rect 31276 21148 31316 21188
rect 31358 21148 31398 21188
rect 31440 21148 31480 21188
rect 35112 21148 35152 21188
rect 35194 21148 35234 21188
rect 35276 21148 35316 21188
rect 35358 21148 35398 21188
rect 35440 21148 35480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 43112 21148 43152 21188
rect 43194 21148 43234 21188
rect 43276 21148 43316 21188
rect 43358 21148 43398 21188
rect 43440 21148 43480 21188
rect 47112 21148 47152 21188
rect 47194 21148 47234 21188
rect 47276 21148 47316 21188
rect 47358 21148 47398 21188
rect 47440 21148 47480 21188
rect 51112 21148 51152 21188
rect 51194 21148 51234 21188
rect 51276 21148 51316 21188
rect 51358 21148 51398 21188
rect 51440 21148 51480 21188
rect 55112 21148 55152 21188
rect 55194 21148 55234 21188
rect 55276 21148 55316 21188
rect 55358 21148 55398 21188
rect 55440 21148 55480 21188
rect 59112 21148 59152 21188
rect 59194 21148 59234 21188
rect 59276 21148 59316 21188
rect 59358 21148 59398 21188
rect 59440 21148 59480 21188
rect 63112 21148 63152 21188
rect 63194 21148 63234 21188
rect 63276 21148 63316 21188
rect 63358 21148 63398 21188
rect 63440 21148 63480 21188
rect 67112 21148 67152 21188
rect 67194 21148 67234 21188
rect 67276 21148 67316 21188
rect 67358 21148 67398 21188
rect 67440 21148 67480 21188
rect 71112 21148 71152 21188
rect 71194 21148 71234 21188
rect 71276 21148 71316 21188
rect 71358 21148 71398 21188
rect 71440 21148 71480 21188
rect 75112 21148 75152 21188
rect 75194 21148 75234 21188
rect 75276 21148 75316 21188
rect 75358 21148 75398 21188
rect 75440 21148 75480 21188
rect 79112 21148 79152 21188
rect 79194 21148 79234 21188
rect 79276 21148 79316 21188
rect 79358 21148 79398 21188
rect 79440 21148 79480 21188
rect 83112 21148 83152 21188
rect 83194 21148 83234 21188
rect 83276 21148 83316 21188
rect 83358 21148 83398 21188
rect 83440 21148 83480 21188
rect 87112 21148 87152 21188
rect 87194 21148 87234 21188
rect 87276 21148 87316 21188
rect 87358 21148 87398 21188
rect 87440 21148 87480 21188
rect 91112 21148 91152 21188
rect 91194 21148 91234 21188
rect 91276 21148 91316 21188
rect 91358 21148 91398 21188
rect 91440 21148 91480 21188
rect 95112 21148 95152 21188
rect 95194 21148 95234 21188
rect 95276 21148 95316 21188
rect 95358 21148 95398 21188
rect 95440 21148 95480 21188
rect 99112 21148 99152 21188
rect 99194 21148 99234 21188
rect 99276 21148 99316 21188
rect 99358 21148 99398 21188
rect 99440 21148 99480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 8352 20392 8392 20432
rect 8434 20392 8474 20432
rect 8516 20392 8556 20432
rect 8598 20392 8638 20432
rect 8680 20392 8720 20432
rect 12352 20392 12392 20432
rect 12434 20392 12474 20432
rect 12516 20392 12556 20432
rect 12598 20392 12638 20432
rect 12680 20392 12720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 20352 20392 20392 20432
rect 20434 20392 20474 20432
rect 20516 20392 20556 20432
rect 20598 20392 20638 20432
rect 20680 20392 20720 20432
rect 24352 20392 24392 20432
rect 24434 20392 24474 20432
rect 24516 20392 24556 20432
rect 24598 20392 24638 20432
rect 24680 20392 24720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 32352 20392 32392 20432
rect 32434 20392 32474 20432
rect 32516 20392 32556 20432
rect 32598 20392 32638 20432
rect 32680 20392 32720 20432
rect 36352 20392 36392 20432
rect 36434 20392 36474 20432
rect 36516 20392 36556 20432
rect 36598 20392 36638 20432
rect 36680 20392 36720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 44352 20392 44392 20432
rect 44434 20392 44474 20432
rect 44516 20392 44556 20432
rect 44598 20392 44638 20432
rect 44680 20392 44720 20432
rect 48352 20392 48392 20432
rect 48434 20392 48474 20432
rect 48516 20392 48556 20432
rect 48598 20392 48638 20432
rect 48680 20392 48720 20432
rect 52352 20392 52392 20432
rect 52434 20392 52474 20432
rect 52516 20392 52556 20432
rect 52598 20392 52638 20432
rect 52680 20392 52720 20432
rect 56352 20392 56392 20432
rect 56434 20392 56474 20432
rect 56516 20392 56556 20432
rect 56598 20392 56638 20432
rect 56680 20392 56720 20432
rect 60352 20392 60392 20432
rect 60434 20392 60474 20432
rect 60516 20392 60556 20432
rect 60598 20392 60638 20432
rect 60680 20392 60720 20432
rect 64352 20392 64392 20432
rect 64434 20392 64474 20432
rect 64516 20392 64556 20432
rect 64598 20392 64638 20432
rect 64680 20392 64720 20432
rect 68352 20392 68392 20432
rect 68434 20392 68474 20432
rect 68516 20392 68556 20432
rect 68598 20392 68638 20432
rect 68680 20392 68720 20432
rect 72352 20392 72392 20432
rect 72434 20392 72474 20432
rect 72516 20392 72556 20432
rect 72598 20392 72638 20432
rect 72680 20392 72720 20432
rect 76352 20392 76392 20432
rect 76434 20392 76474 20432
rect 76516 20392 76556 20432
rect 76598 20392 76638 20432
rect 76680 20392 76720 20432
rect 80352 20392 80392 20432
rect 80434 20392 80474 20432
rect 80516 20392 80556 20432
rect 80598 20392 80638 20432
rect 80680 20392 80720 20432
rect 84352 20392 84392 20432
rect 84434 20392 84474 20432
rect 84516 20392 84556 20432
rect 84598 20392 84638 20432
rect 84680 20392 84720 20432
rect 88352 20392 88392 20432
rect 88434 20392 88474 20432
rect 88516 20392 88556 20432
rect 88598 20392 88638 20432
rect 88680 20392 88720 20432
rect 92352 20392 92392 20432
rect 92434 20392 92474 20432
rect 92516 20392 92556 20432
rect 92598 20392 92638 20432
rect 92680 20392 92720 20432
rect 96352 20392 96392 20432
rect 96434 20392 96474 20432
rect 96516 20392 96556 20432
rect 96598 20392 96638 20432
rect 96680 20392 96720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 7112 19636 7152 19676
rect 7194 19636 7234 19676
rect 7276 19636 7316 19676
rect 7358 19636 7398 19676
rect 7440 19636 7480 19676
rect 11112 19636 11152 19676
rect 11194 19636 11234 19676
rect 11276 19636 11316 19676
rect 11358 19636 11398 19676
rect 11440 19636 11480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 19112 19636 19152 19676
rect 19194 19636 19234 19676
rect 19276 19636 19316 19676
rect 19358 19636 19398 19676
rect 19440 19636 19480 19676
rect 23112 19636 23152 19676
rect 23194 19636 23234 19676
rect 23276 19636 23316 19676
rect 23358 19636 23398 19676
rect 23440 19636 23480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 31112 19636 31152 19676
rect 31194 19636 31234 19676
rect 31276 19636 31316 19676
rect 31358 19636 31398 19676
rect 31440 19636 31480 19676
rect 35112 19636 35152 19676
rect 35194 19636 35234 19676
rect 35276 19636 35316 19676
rect 35358 19636 35398 19676
rect 35440 19636 35480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 43112 19636 43152 19676
rect 43194 19636 43234 19676
rect 43276 19636 43316 19676
rect 43358 19636 43398 19676
rect 43440 19636 43480 19676
rect 47112 19636 47152 19676
rect 47194 19636 47234 19676
rect 47276 19636 47316 19676
rect 47358 19636 47398 19676
rect 47440 19636 47480 19676
rect 51112 19636 51152 19676
rect 51194 19636 51234 19676
rect 51276 19636 51316 19676
rect 51358 19636 51398 19676
rect 51440 19636 51480 19676
rect 55112 19636 55152 19676
rect 55194 19636 55234 19676
rect 55276 19636 55316 19676
rect 55358 19636 55398 19676
rect 55440 19636 55480 19676
rect 59112 19636 59152 19676
rect 59194 19636 59234 19676
rect 59276 19636 59316 19676
rect 59358 19636 59398 19676
rect 59440 19636 59480 19676
rect 63112 19636 63152 19676
rect 63194 19636 63234 19676
rect 63276 19636 63316 19676
rect 63358 19636 63398 19676
rect 63440 19636 63480 19676
rect 67112 19636 67152 19676
rect 67194 19636 67234 19676
rect 67276 19636 67316 19676
rect 67358 19636 67398 19676
rect 67440 19636 67480 19676
rect 71112 19636 71152 19676
rect 71194 19636 71234 19676
rect 71276 19636 71316 19676
rect 71358 19636 71398 19676
rect 71440 19636 71480 19676
rect 75112 19636 75152 19676
rect 75194 19636 75234 19676
rect 75276 19636 75316 19676
rect 75358 19636 75398 19676
rect 75440 19636 75480 19676
rect 79112 19636 79152 19676
rect 79194 19636 79234 19676
rect 79276 19636 79316 19676
rect 79358 19636 79398 19676
rect 79440 19636 79480 19676
rect 83112 19636 83152 19676
rect 83194 19636 83234 19676
rect 83276 19636 83316 19676
rect 83358 19636 83398 19676
rect 83440 19636 83480 19676
rect 87112 19636 87152 19676
rect 87194 19636 87234 19676
rect 87276 19636 87316 19676
rect 87358 19636 87398 19676
rect 87440 19636 87480 19676
rect 91112 19636 91152 19676
rect 91194 19636 91234 19676
rect 91276 19636 91316 19676
rect 91358 19636 91398 19676
rect 91440 19636 91480 19676
rect 95112 19636 95152 19676
rect 95194 19636 95234 19676
rect 95276 19636 95316 19676
rect 95358 19636 95398 19676
rect 95440 19636 95480 19676
rect 99112 19636 99152 19676
rect 99194 19636 99234 19676
rect 99276 19636 99316 19676
rect 99358 19636 99398 19676
rect 99440 19636 99480 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 8352 18880 8392 18920
rect 8434 18880 8474 18920
rect 8516 18880 8556 18920
rect 8598 18880 8638 18920
rect 8680 18880 8720 18920
rect 12352 18880 12392 18920
rect 12434 18880 12474 18920
rect 12516 18880 12556 18920
rect 12598 18880 12638 18920
rect 12680 18880 12720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 20352 18880 20392 18920
rect 20434 18880 20474 18920
rect 20516 18880 20556 18920
rect 20598 18880 20638 18920
rect 20680 18880 20720 18920
rect 24352 18880 24392 18920
rect 24434 18880 24474 18920
rect 24516 18880 24556 18920
rect 24598 18880 24638 18920
rect 24680 18880 24720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 32352 18880 32392 18920
rect 32434 18880 32474 18920
rect 32516 18880 32556 18920
rect 32598 18880 32638 18920
rect 32680 18880 32720 18920
rect 36352 18880 36392 18920
rect 36434 18880 36474 18920
rect 36516 18880 36556 18920
rect 36598 18880 36638 18920
rect 36680 18880 36720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 44352 18880 44392 18920
rect 44434 18880 44474 18920
rect 44516 18880 44556 18920
rect 44598 18880 44638 18920
rect 44680 18880 44720 18920
rect 48352 18880 48392 18920
rect 48434 18880 48474 18920
rect 48516 18880 48556 18920
rect 48598 18880 48638 18920
rect 48680 18880 48720 18920
rect 52352 18880 52392 18920
rect 52434 18880 52474 18920
rect 52516 18880 52556 18920
rect 52598 18880 52638 18920
rect 52680 18880 52720 18920
rect 56352 18880 56392 18920
rect 56434 18880 56474 18920
rect 56516 18880 56556 18920
rect 56598 18880 56638 18920
rect 56680 18880 56720 18920
rect 60352 18880 60392 18920
rect 60434 18880 60474 18920
rect 60516 18880 60556 18920
rect 60598 18880 60638 18920
rect 60680 18880 60720 18920
rect 64352 18880 64392 18920
rect 64434 18880 64474 18920
rect 64516 18880 64556 18920
rect 64598 18880 64638 18920
rect 64680 18880 64720 18920
rect 68352 18880 68392 18920
rect 68434 18880 68474 18920
rect 68516 18880 68556 18920
rect 68598 18880 68638 18920
rect 68680 18880 68720 18920
rect 72352 18880 72392 18920
rect 72434 18880 72474 18920
rect 72516 18880 72556 18920
rect 72598 18880 72638 18920
rect 72680 18880 72720 18920
rect 76352 18880 76392 18920
rect 76434 18880 76474 18920
rect 76516 18880 76556 18920
rect 76598 18880 76638 18920
rect 76680 18880 76720 18920
rect 80352 18880 80392 18920
rect 80434 18880 80474 18920
rect 80516 18880 80556 18920
rect 80598 18880 80638 18920
rect 80680 18880 80720 18920
rect 84352 18880 84392 18920
rect 84434 18880 84474 18920
rect 84516 18880 84556 18920
rect 84598 18880 84638 18920
rect 84680 18880 84720 18920
rect 88352 18880 88392 18920
rect 88434 18880 88474 18920
rect 88516 18880 88556 18920
rect 88598 18880 88638 18920
rect 88680 18880 88720 18920
rect 92352 18880 92392 18920
rect 92434 18880 92474 18920
rect 92516 18880 92556 18920
rect 92598 18880 92638 18920
rect 92680 18880 92720 18920
rect 96352 18880 96392 18920
rect 96434 18880 96474 18920
rect 96516 18880 96556 18920
rect 96598 18880 96638 18920
rect 96680 18880 96720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 7112 18124 7152 18164
rect 7194 18124 7234 18164
rect 7276 18124 7316 18164
rect 7358 18124 7398 18164
rect 7440 18124 7480 18164
rect 11112 18124 11152 18164
rect 11194 18124 11234 18164
rect 11276 18124 11316 18164
rect 11358 18124 11398 18164
rect 11440 18124 11480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 19112 18124 19152 18164
rect 19194 18124 19234 18164
rect 19276 18124 19316 18164
rect 19358 18124 19398 18164
rect 19440 18124 19480 18164
rect 23112 18124 23152 18164
rect 23194 18124 23234 18164
rect 23276 18124 23316 18164
rect 23358 18124 23398 18164
rect 23440 18124 23480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 31112 18124 31152 18164
rect 31194 18124 31234 18164
rect 31276 18124 31316 18164
rect 31358 18124 31398 18164
rect 31440 18124 31480 18164
rect 35112 18124 35152 18164
rect 35194 18124 35234 18164
rect 35276 18124 35316 18164
rect 35358 18124 35398 18164
rect 35440 18124 35480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 43112 18124 43152 18164
rect 43194 18124 43234 18164
rect 43276 18124 43316 18164
rect 43358 18124 43398 18164
rect 43440 18124 43480 18164
rect 47112 18124 47152 18164
rect 47194 18124 47234 18164
rect 47276 18124 47316 18164
rect 47358 18124 47398 18164
rect 47440 18124 47480 18164
rect 51112 18124 51152 18164
rect 51194 18124 51234 18164
rect 51276 18124 51316 18164
rect 51358 18124 51398 18164
rect 51440 18124 51480 18164
rect 55112 18124 55152 18164
rect 55194 18124 55234 18164
rect 55276 18124 55316 18164
rect 55358 18124 55398 18164
rect 55440 18124 55480 18164
rect 59112 18124 59152 18164
rect 59194 18124 59234 18164
rect 59276 18124 59316 18164
rect 59358 18124 59398 18164
rect 59440 18124 59480 18164
rect 63112 18124 63152 18164
rect 63194 18124 63234 18164
rect 63276 18124 63316 18164
rect 63358 18124 63398 18164
rect 63440 18124 63480 18164
rect 67112 18124 67152 18164
rect 67194 18124 67234 18164
rect 67276 18124 67316 18164
rect 67358 18124 67398 18164
rect 67440 18124 67480 18164
rect 71112 18124 71152 18164
rect 71194 18124 71234 18164
rect 71276 18124 71316 18164
rect 71358 18124 71398 18164
rect 71440 18124 71480 18164
rect 75112 18124 75152 18164
rect 75194 18124 75234 18164
rect 75276 18124 75316 18164
rect 75358 18124 75398 18164
rect 75440 18124 75480 18164
rect 79112 18124 79152 18164
rect 79194 18124 79234 18164
rect 79276 18124 79316 18164
rect 79358 18124 79398 18164
rect 79440 18124 79480 18164
rect 83112 18124 83152 18164
rect 83194 18124 83234 18164
rect 83276 18124 83316 18164
rect 83358 18124 83398 18164
rect 83440 18124 83480 18164
rect 87112 18124 87152 18164
rect 87194 18124 87234 18164
rect 87276 18124 87316 18164
rect 87358 18124 87398 18164
rect 87440 18124 87480 18164
rect 91112 18124 91152 18164
rect 91194 18124 91234 18164
rect 91276 18124 91316 18164
rect 91358 18124 91398 18164
rect 91440 18124 91480 18164
rect 95112 18124 95152 18164
rect 95194 18124 95234 18164
rect 95276 18124 95316 18164
rect 95358 18124 95398 18164
rect 95440 18124 95480 18164
rect 99112 18124 99152 18164
rect 99194 18124 99234 18164
rect 99276 18124 99316 18164
rect 99358 18124 99398 18164
rect 99440 18124 99480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 8352 17368 8392 17408
rect 8434 17368 8474 17408
rect 8516 17368 8556 17408
rect 8598 17368 8638 17408
rect 8680 17368 8720 17408
rect 12352 17368 12392 17408
rect 12434 17368 12474 17408
rect 12516 17368 12556 17408
rect 12598 17368 12638 17408
rect 12680 17368 12720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 20352 17368 20392 17408
rect 20434 17368 20474 17408
rect 20516 17368 20556 17408
rect 20598 17368 20638 17408
rect 20680 17368 20720 17408
rect 24352 17368 24392 17408
rect 24434 17368 24474 17408
rect 24516 17368 24556 17408
rect 24598 17368 24638 17408
rect 24680 17368 24720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 32352 17368 32392 17408
rect 32434 17368 32474 17408
rect 32516 17368 32556 17408
rect 32598 17368 32638 17408
rect 32680 17368 32720 17408
rect 36352 17368 36392 17408
rect 36434 17368 36474 17408
rect 36516 17368 36556 17408
rect 36598 17368 36638 17408
rect 36680 17368 36720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 44352 17368 44392 17408
rect 44434 17368 44474 17408
rect 44516 17368 44556 17408
rect 44598 17368 44638 17408
rect 44680 17368 44720 17408
rect 48352 17368 48392 17408
rect 48434 17368 48474 17408
rect 48516 17368 48556 17408
rect 48598 17368 48638 17408
rect 48680 17368 48720 17408
rect 52352 17368 52392 17408
rect 52434 17368 52474 17408
rect 52516 17368 52556 17408
rect 52598 17368 52638 17408
rect 52680 17368 52720 17408
rect 56352 17368 56392 17408
rect 56434 17368 56474 17408
rect 56516 17368 56556 17408
rect 56598 17368 56638 17408
rect 56680 17368 56720 17408
rect 60352 17368 60392 17408
rect 60434 17368 60474 17408
rect 60516 17368 60556 17408
rect 60598 17368 60638 17408
rect 60680 17368 60720 17408
rect 64352 17368 64392 17408
rect 64434 17368 64474 17408
rect 64516 17368 64556 17408
rect 64598 17368 64638 17408
rect 64680 17368 64720 17408
rect 68352 17368 68392 17408
rect 68434 17368 68474 17408
rect 68516 17368 68556 17408
rect 68598 17368 68638 17408
rect 68680 17368 68720 17408
rect 72352 17368 72392 17408
rect 72434 17368 72474 17408
rect 72516 17368 72556 17408
rect 72598 17368 72638 17408
rect 72680 17368 72720 17408
rect 76352 17368 76392 17408
rect 76434 17368 76474 17408
rect 76516 17368 76556 17408
rect 76598 17368 76638 17408
rect 76680 17368 76720 17408
rect 80352 17368 80392 17408
rect 80434 17368 80474 17408
rect 80516 17368 80556 17408
rect 80598 17368 80638 17408
rect 80680 17368 80720 17408
rect 84352 17368 84392 17408
rect 84434 17368 84474 17408
rect 84516 17368 84556 17408
rect 84598 17368 84638 17408
rect 84680 17368 84720 17408
rect 88352 17368 88392 17408
rect 88434 17368 88474 17408
rect 88516 17368 88556 17408
rect 88598 17368 88638 17408
rect 88680 17368 88720 17408
rect 92352 17368 92392 17408
rect 92434 17368 92474 17408
rect 92516 17368 92556 17408
rect 92598 17368 92638 17408
rect 92680 17368 92720 17408
rect 96352 17368 96392 17408
rect 96434 17368 96474 17408
rect 96516 17368 96556 17408
rect 96598 17368 96638 17408
rect 96680 17368 96720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 7112 16612 7152 16652
rect 7194 16612 7234 16652
rect 7276 16612 7316 16652
rect 7358 16612 7398 16652
rect 7440 16612 7480 16652
rect 11112 16612 11152 16652
rect 11194 16612 11234 16652
rect 11276 16612 11316 16652
rect 11358 16612 11398 16652
rect 11440 16612 11480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 19112 16612 19152 16652
rect 19194 16612 19234 16652
rect 19276 16612 19316 16652
rect 19358 16612 19398 16652
rect 19440 16612 19480 16652
rect 23112 16612 23152 16652
rect 23194 16612 23234 16652
rect 23276 16612 23316 16652
rect 23358 16612 23398 16652
rect 23440 16612 23480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 31112 16612 31152 16652
rect 31194 16612 31234 16652
rect 31276 16612 31316 16652
rect 31358 16612 31398 16652
rect 31440 16612 31480 16652
rect 35112 16612 35152 16652
rect 35194 16612 35234 16652
rect 35276 16612 35316 16652
rect 35358 16612 35398 16652
rect 35440 16612 35480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 43112 16612 43152 16652
rect 43194 16612 43234 16652
rect 43276 16612 43316 16652
rect 43358 16612 43398 16652
rect 43440 16612 43480 16652
rect 47112 16612 47152 16652
rect 47194 16612 47234 16652
rect 47276 16612 47316 16652
rect 47358 16612 47398 16652
rect 47440 16612 47480 16652
rect 51112 16612 51152 16652
rect 51194 16612 51234 16652
rect 51276 16612 51316 16652
rect 51358 16612 51398 16652
rect 51440 16612 51480 16652
rect 55112 16612 55152 16652
rect 55194 16612 55234 16652
rect 55276 16612 55316 16652
rect 55358 16612 55398 16652
rect 55440 16612 55480 16652
rect 59112 16612 59152 16652
rect 59194 16612 59234 16652
rect 59276 16612 59316 16652
rect 59358 16612 59398 16652
rect 59440 16612 59480 16652
rect 63112 16612 63152 16652
rect 63194 16612 63234 16652
rect 63276 16612 63316 16652
rect 63358 16612 63398 16652
rect 63440 16612 63480 16652
rect 67112 16612 67152 16652
rect 67194 16612 67234 16652
rect 67276 16612 67316 16652
rect 67358 16612 67398 16652
rect 67440 16612 67480 16652
rect 71112 16612 71152 16652
rect 71194 16612 71234 16652
rect 71276 16612 71316 16652
rect 71358 16612 71398 16652
rect 71440 16612 71480 16652
rect 75112 16612 75152 16652
rect 75194 16612 75234 16652
rect 75276 16612 75316 16652
rect 75358 16612 75398 16652
rect 75440 16612 75480 16652
rect 79112 16612 79152 16652
rect 79194 16612 79234 16652
rect 79276 16612 79316 16652
rect 79358 16612 79398 16652
rect 79440 16612 79480 16652
rect 83112 16612 83152 16652
rect 83194 16612 83234 16652
rect 83276 16612 83316 16652
rect 83358 16612 83398 16652
rect 83440 16612 83480 16652
rect 87112 16612 87152 16652
rect 87194 16612 87234 16652
rect 87276 16612 87316 16652
rect 87358 16612 87398 16652
rect 87440 16612 87480 16652
rect 91112 16612 91152 16652
rect 91194 16612 91234 16652
rect 91276 16612 91316 16652
rect 91358 16612 91398 16652
rect 91440 16612 91480 16652
rect 95112 16612 95152 16652
rect 95194 16612 95234 16652
rect 95276 16612 95316 16652
rect 95358 16612 95398 16652
rect 95440 16612 95480 16652
rect 99112 16612 99152 16652
rect 99194 16612 99234 16652
rect 99276 16612 99316 16652
rect 99358 16612 99398 16652
rect 99440 16612 99480 16652
rect 86188 16360 86228 16400
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 8352 15856 8392 15896
rect 8434 15856 8474 15896
rect 8516 15856 8556 15896
rect 8598 15856 8638 15896
rect 8680 15856 8720 15896
rect 12352 15856 12392 15896
rect 12434 15856 12474 15896
rect 12516 15856 12556 15896
rect 12598 15856 12638 15896
rect 12680 15856 12720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 20352 15856 20392 15896
rect 20434 15856 20474 15896
rect 20516 15856 20556 15896
rect 20598 15856 20638 15896
rect 20680 15856 20720 15896
rect 24352 15856 24392 15896
rect 24434 15856 24474 15896
rect 24516 15856 24556 15896
rect 24598 15856 24638 15896
rect 24680 15856 24720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 32352 15856 32392 15896
rect 32434 15856 32474 15896
rect 32516 15856 32556 15896
rect 32598 15856 32638 15896
rect 32680 15856 32720 15896
rect 36352 15856 36392 15896
rect 36434 15856 36474 15896
rect 36516 15856 36556 15896
rect 36598 15856 36638 15896
rect 36680 15856 36720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 44352 15856 44392 15896
rect 44434 15856 44474 15896
rect 44516 15856 44556 15896
rect 44598 15856 44638 15896
rect 44680 15856 44720 15896
rect 48352 15856 48392 15896
rect 48434 15856 48474 15896
rect 48516 15856 48556 15896
rect 48598 15856 48638 15896
rect 48680 15856 48720 15896
rect 52352 15856 52392 15896
rect 52434 15856 52474 15896
rect 52516 15856 52556 15896
rect 52598 15856 52638 15896
rect 52680 15856 52720 15896
rect 56352 15856 56392 15896
rect 56434 15856 56474 15896
rect 56516 15856 56556 15896
rect 56598 15856 56638 15896
rect 56680 15856 56720 15896
rect 60352 15856 60392 15896
rect 60434 15856 60474 15896
rect 60516 15856 60556 15896
rect 60598 15856 60638 15896
rect 60680 15856 60720 15896
rect 64352 15856 64392 15896
rect 64434 15856 64474 15896
rect 64516 15856 64556 15896
rect 64598 15856 64638 15896
rect 64680 15856 64720 15896
rect 68352 15856 68392 15896
rect 68434 15856 68474 15896
rect 68516 15856 68556 15896
rect 68598 15856 68638 15896
rect 68680 15856 68720 15896
rect 72352 15856 72392 15896
rect 72434 15856 72474 15896
rect 72516 15856 72556 15896
rect 72598 15856 72638 15896
rect 72680 15856 72720 15896
rect 76352 15856 76392 15896
rect 76434 15856 76474 15896
rect 76516 15856 76556 15896
rect 76598 15856 76638 15896
rect 76680 15856 76720 15896
rect 80352 15856 80392 15896
rect 80434 15856 80474 15896
rect 80516 15856 80556 15896
rect 80598 15856 80638 15896
rect 80680 15856 80720 15896
rect 84352 15856 84392 15896
rect 84434 15856 84474 15896
rect 84516 15856 84556 15896
rect 84598 15856 84638 15896
rect 84680 15856 84720 15896
rect 88352 15856 88392 15896
rect 88434 15856 88474 15896
rect 88516 15856 88556 15896
rect 88598 15856 88638 15896
rect 88680 15856 88720 15896
rect 92352 15856 92392 15896
rect 92434 15856 92474 15896
rect 92516 15856 92556 15896
rect 92598 15856 92638 15896
rect 92680 15856 92720 15896
rect 96352 15856 96392 15896
rect 96434 15856 96474 15896
rect 96516 15856 96556 15896
rect 96598 15856 96638 15896
rect 96680 15856 96720 15896
rect 90892 15268 90932 15308
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 7112 15100 7152 15140
rect 7194 15100 7234 15140
rect 7276 15100 7316 15140
rect 7358 15100 7398 15140
rect 7440 15100 7480 15140
rect 11112 15100 11152 15140
rect 11194 15100 11234 15140
rect 11276 15100 11316 15140
rect 11358 15100 11398 15140
rect 11440 15100 11480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 19112 15100 19152 15140
rect 19194 15100 19234 15140
rect 19276 15100 19316 15140
rect 19358 15100 19398 15140
rect 19440 15100 19480 15140
rect 23112 15100 23152 15140
rect 23194 15100 23234 15140
rect 23276 15100 23316 15140
rect 23358 15100 23398 15140
rect 23440 15100 23480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 31112 15100 31152 15140
rect 31194 15100 31234 15140
rect 31276 15100 31316 15140
rect 31358 15100 31398 15140
rect 31440 15100 31480 15140
rect 35112 15100 35152 15140
rect 35194 15100 35234 15140
rect 35276 15100 35316 15140
rect 35358 15100 35398 15140
rect 35440 15100 35480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 43112 15100 43152 15140
rect 43194 15100 43234 15140
rect 43276 15100 43316 15140
rect 43358 15100 43398 15140
rect 43440 15100 43480 15140
rect 47112 15100 47152 15140
rect 47194 15100 47234 15140
rect 47276 15100 47316 15140
rect 47358 15100 47398 15140
rect 47440 15100 47480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 55112 15100 55152 15140
rect 55194 15100 55234 15140
rect 55276 15100 55316 15140
rect 55358 15100 55398 15140
rect 55440 15100 55480 15140
rect 59112 15100 59152 15140
rect 59194 15100 59234 15140
rect 59276 15100 59316 15140
rect 59358 15100 59398 15140
rect 59440 15100 59480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 67112 15100 67152 15140
rect 67194 15100 67234 15140
rect 67276 15100 67316 15140
rect 67358 15100 67398 15140
rect 67440 15100 67480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 8352 14344 8392 14384
rect 8434 14344 8474 14384
rect 8516 14344 8556 14384
rect 8598 14344 8638 14384
rect 8680 14344 8720 14384
rect 12352 14344 12392 14384
rect 12434 14344 12474 14384
rect 12516 14344 12556 14384
rect 12598 14344 12638 14384
rect 12680 14344 12720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 20352 14344 20392 14384
rect 20434 14344 20474 14384
rect 20516 14344 20556 14384
rect 20598 14344 20638 14384
rect 20680 14344 20720 14384
rect 24352 14344 24392 14384
rect 24434 14344 24474 14384
rect 24516 14344 24556 14384
rect 24598 14344 24638 14384
rect 24680 14344 24720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 32352 14344 32392 14384
rect 32434 14344 32474 14384
rect 32516 14344 32556 14384
rect 32598 14344 32638 14384
rect 32680 14344 32720 14384
rect 36352 14344 36392 14384
rect 36434 14344 36474 14384
rect 36516 14344 36556 14384
rect 36598 14344 36638 14384
rect 36680 14344 36720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 44352 14344 44392 14384
rect 44434 14344 44474 14384
rect 44516 14344 44556 14384
rect 44598 14344 44638 14384
rect 44680 14344 44720 14384
rect 48352 14344 48392 14384
rect 48434 14344 48474 14384
rect 48516 14344 48556 14384
rect 48598 14344 48638 14384
rect 48680 14344 48720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 56352 14344 56392 14384
rect 56434 14344 56474 14384
rect 56516 14344 56556 14384
rect 56598 14344 56638 14384
rect 56680 14344 56720 14384
rect 60352 14344 60392 14384
rect 60434 14344 60474 14384
rect 60516 14344 60556 14384
rect 60598 14344 60638 14384
rect 60680 14344 60720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 68352 14344 68392 14384
rect 68434 14344 68474 14384
rect 68516 14344 68556 14384
rect 68598 14344 68638 14384
rect 68680 14344 68720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 7112 13588 7152 13628
rect 7194 13588 7234 13628
rect 7276 13588 7316 13628
rect 7358 13588 7398 13628
rect 7440 13588 7480 13628
rect 11112 13588 11152 13628
rect 11194 13588 11234 13628
rect 11276 13588 11316 13628
rect 11358 13588 11398 13628
rect 11440 13588 11480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 19112 13588 19152 13628
rect 19194 13588 19234 13628
rect 19276 13588 19316 13628
rect 19358 13588 19398 13628
rect 19440 13588 19480 13628
rect 23112 13588 23152 13628
rect 23194 13588 23234 13628
rect 23276 13588 23316 13628
rect 23358 13588 23398 13628
rect 23440 13588 23480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 31112 13588 31152 13628
rect 31194 13588 31234 13628
rect 31276 13588 31316 13628
rect 31358 13588 31398 13628
rect 31440 13588 31480 13628
rect 35112 13588 35152 13628
rect 35194 13588 35234 13628
rect 35276 13588 35316 13628
rect 35358 13588 35398 13628
rect 35440 13588 35480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 43112 13588 43152 13628
rect 43194 13588 43234 13628
rect 43276 13588 43316 13628
rect 43358 13588 43398 13628
rect 43440 13588 43480 13628
rect 47112 13588 47152 13628
rect 47194 13588 47234 13628
rect 47276 13588 47316 13628
rect 47358 13588 47398 13628
rect 47440 13588 47480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 55112 13588 55152 13628
rect 55194 13588 55234 13628
rect 55276 13588 55316 13628
rect 55358 13588 55398 13628
rect 55440 13588 55480 13628
rect 59112 13588 59152 13628
rect 59194 13588 59234 13628
rect 59276 13588 59316 13628
rect 59358 13588 59398 13628
rect 59440 13588 59480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 67112 13588 67152 13628
rect 67194 13588 67234 13628
rect 67276 13588 67316 13628
rect 67358 13588 67398 13628
rect 67440 13588 67480 13628
rect 90892 13420 90932 13460
rect 72460 13336 72500 13376
rect 71884 13252 71924 13292
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 8352 12832 8392 12872
rect 8434 12832 8474 12872
rect 8516 12832 8556 12872
rect 8598 12832 8638 12872
rect 8680 12832 8720 12872
rect 12352 12832 12392 12872
rect 12434 12832 12474 12872
rect 12516 12832 12556 12872
rect 12598 12832 12638 12872
rect 12680 12832 12720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 20352 12832 20392 12872
rect 20434 12832 20474 12872
rect 20516 12832 20556 12872
rect 20598 12832 20638 12872
rect 20680 12832 20720 12872
rect 24352 12832 24392 12872
rect 24434 12832 24474 12872
rect 24516 12832 24556 12872
rect 24598 12832 24638 12872
rect 24680 12832 24720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 32352 12832 32392 12872
rect 32434 12832 32474 12872
rect 32516 12832 32556 12872
rect 32598 12832 32638 12872
rect 32680 12832 32720 12872
rect 36352 12832 36392 12872
rect 36434 12832 36474 12872
rect 36516 12832 36556 12872
rect 36598 12832 36638 12872
rect 36680 12832 36720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 44352 12832 44392 12872
rect 44434 12832 44474 12872
rect 44516 12832 44556 12872
rect 44598 12832 44638 12872
rect 44680 12832 44720 12872
rect 48352 12832 48392 12872
rect 48434 12832 48474 12872
rect 48516 12832 48556 12872
rect 48598 12832 48638 12872
rect 48680 12832 48720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 56352 12832 56392 12872
rect 56434 12832 56474 12872
rect 56516 12832 56556 12872
rect 56598 12832 56638 12872
rect 56680 12832 56720 12872
rect 60352 12832 60392 12872
rect 60434 12832 60474 12872
rect 60516 12832 60556 12872
rect 60598 12832 60638 12872
rect 60680 12832 60720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 68352 12832 68392 12872
rect 68434 12832 68474 12872
rect 68516 12832 68556 12872
rect 68598 12832 68638 12872
rect 68680 12832 68720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 7112 12076 7152 12116
rect 7194 12076 7234 12116
rect 7276 12076 7316 12116
rect 7358 12076 7398 12116
rect 7440 12076 7480 12116
rect 11112 12076 11152 12116
rect 11194 12076 11234 12116
rect 11276 12076 11316 12116
rect 11358 12076 11398 12116
rect 11440 12076 11480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 19112 12076 19152 12116
rect 19194 12076 19234 12116
rect 19276 12076 19316 12116
rect 19358 12076 19398 12116
rect 19440 12076 19480 12116
rect 23112 12076 23152 12116
rect 23194 12076 23234 12116
rect 23276 12076 23316 12116
rect 23358 12076 23398 12116
rect 23440 12076 23480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 31112 12076 31152 12116
rect 31194 12076 31234 12116
rect 31276 12076 31316 12116
rect 31358 12076 31398 12116
rect 31440 12076 31480 12116
rect 35112 12076 35152 12116
rect 35194 12076 35234 12116
rect 35276 12076 35316 12116
rect 35358 12076 35398 12116
rect 35440 12076 35480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 43112 12076 43152 12116
rect 43194 12076 43234 12116
rect 43276 12076 43316 12116
rect 43358 12076 43398 12116
rect 43440 12076 43480 12116
rect 47112 12076 47152 12116
rect 47194 12076 47234 12116
rect 47276 12076 47316 12116
rect 47358 12076 47398 12116
rect 47440 12076 47480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 55112 12076 55152 12116
rect 55194 12076 55234 12116
rect 55276 12076 55316 12116
rect 55358 12076 55398 12116
rect 55440 12076 55480 12116
rect 59112 12076 59152 12116
rect 59194 12076 59234 12116
rect 59276 12076 59316 12116
rect 59358 12076 59398 12116
rect 59440 12076 59480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 67112 12076 67152 12116
rect 67194 12076 67234 12116
rect 67276 12076 67316 12116
rect 67358 12076 67398 12116
rect 67440 12076 67480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 8352 11320 8392 11360
rect 8434 11320 8474 11360
rect 8516 11320 8556 11360
rect 8598 11320 8638 11360
rect 8680 11320 8720 11360
rect 12352 11320 12392 11360
rect 12434 11320 12474 11360
rect 12516 11320 12556 11360
rect 12598 11320 12638 11360
rect 12680 11320 12720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 20352 11320 20392 11360
rect 20434 11320 20474 11360
rect 20516 11320 20556 11360
rect 20598 11320 20638 11360
rect 20680 11320 20720 11360
rect 24352 11320 24392 11360
rect 24434 11320 24474 11360
rect 24516 11320 24556 11360
rect 24598 11320 24638 11360
rect 24680 11320 24720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 32352 11320 32392 11360
rect 32434 11320 32474 11360
rect 32516 11320 32556 11360
rect 32598 11320 32638 11360
rect 32680 11320 32720 11360
rect 36352 11320 36392 11360
rect 36434 11320 36474 11360
rect 36516 11320 36556 11360
rect 36598 11320 36638 11360
rect 36680 11320 36720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 44352 11320 44392 11360
rect 44434 11320 44474 11360
rect 44516 11320 44556 11360
rect 44598 11320 44638 11360
rect 44680 11320 44720 11360
rect 48352 11320 48392 11360
rect 48434 11320 48474 11360
rect 48516 11320 48556 11360
rect 48598 11320 48638 11360
rect 48680 11320 48720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 56352 11320 56392 11360
rect 56434 11320 56474 11360
rect 56516 11320 56556 11360
rect 56598 11320 56638 11360
rect 56680 11320 56720 11360
rect 60352 11320 60392 11360
rect 60434 11320 60474 11360
rect 60516 11320 60556 11360
rect 60598 11320 60638 11360
rect 60680 11320 60720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 68352 11320 68392 11360
rect 68434 11320 68474 11360
rect 68516 11320 68556 11360
rect 68598 11320 68638 11360
rect 68680 11320 68720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 7112 10564 7152 10604
rect 7194 10564 7234 10604
rect 7276 10564 7316 10604
rect 7358 10564 7398 10604
rect 7440 10564 7480 10604
rect 11112 10564 11152 10604
rect 11194 10564 11234 10604
rect 11276 10564 11316 10604
rect 11358 10564 11398 10604
rect 11440 10564 11480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 19112 10564 19152 10604
rect 19194 10564 19234 10604
rect 19276 10564 19316 10604
rect 19358 10564 19398 10604
rect 19440 10564 19480 10604
rect 23112 10564 23152 10604
rect 23194 10564 23234 10604
rect 23276 10564 23316 10604
rect 23358 10564 23398 10604
rect 23440 10564 23480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 31112 10564 31152 10604
rect 31194 10564 31234 10604
rect 31276 10564 31316 10604
rect 31358 10564 31398 10604
rect 31440 10564 31480 10604
rect 35112 10564 35152 10604
rect 35194 10564 35234 10604
rect 35276 10564 35316 10604
rect 35358 10564 35398 10604
rect 35440 10564 35480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 43112 10564 43152 10604
rect 43194 10564 43234 10604
rect 43276 10564 43316 10604
rect 43358 10564 43398 10604
rect 43440 10564 43480 10604
rect 47112 10564 47152 10604
rect 47194 10564 47234 10604
rect 47276 10564 47316 10604
rect 47358 10564 47398 10604
rect 47440 10564 47480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 55112 10564 55152 10604
rect 55194 10564 55234 10604
rect 55276 10564 55316 10604
rect 55358 10564 55398 10604
rect 55440 10564 55480 10604
rect 59112 10564 59152 10604
rect 59194 10564 59234 10604
rect 59276 10564 59316 10604
rect 59358 10564 59398 10604
rect 59440 10564 59480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 67112 10564 67152 10604
rect 67194 10564 67234 10604
rect 67276 10564 67316 10604
rect 67358 10564 67398 10604
rect 67440 10564 67480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 8352 9808 8392 9848
rect 8434 9808 8474 9848
rect 8516 9808 8556 9848
rect 8598 9808 8638 9848
rect 8680 9808 8720 9848
rect 12352 9808 12392 9848
rect 12434 9808 12474 9848
rect 12516 9808 12556 9848
rect 12598 9808 12638 9848
rect 12680 9808 12720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 20352 9808 20392 9848
rect 20434 9808 20474 9848
rect 20516 9808 20556 9848
rect 20598 9808 20638 9848
rect 20680 9808 20720 9848
rect 24352 9808 24392 9848
rect 24434 9808 24474 9848
rect 24516 9808 24556 9848
rect 24598 9808 24638 9848
rect 24680 9808 24720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 32352 9808 32392 9848
rect 32434 9808 32474 9848
rect 32516 9808 32556 9848
rect 32598 9808 32638 9848
rect 32680 9808 32720 9848
rect 36352 9808 36392 9848
rect 36434 9808 36474 9848
rect 36516 9808 36556 9848
rect 36598 9808 36638 9848
rect 36680 9808 36720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 44352 9808 44392 9848
rect 44434 9808 44474 9848
rect 44516 9808 44556 9848
rect 44598 9808 44638 9848
rect 44680 9808 44720 9848
rect 48352 9808 48392 9848
rect 48434 9808 48474 9848
rect 48516 9808 48556 9848
rect 48598 9808 48638 9848
rect 48680 9808 48720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 56352 9808 56392 9848
rect 56434 9808 56474 9848
rect 56516 9808 56556 9848
rect 56598 9808 56638 9848
rect 56680 9808 56720 9848
rect 60352 9808 60392 9848
rect 60434 9808 60474 9848
rect 60516 9808 60556 9848
rect 60598 9808 60638 9848
rect 60680 9808 60720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 68352 9808 68392 9848
rect 68434 9808 68474 9848
rect 68516 9808 68556 9848
rect 68598 9808 68638 9848
rect 68680 9808 68720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 7112 9052 7152 9092
rect 7194 9052 7234 9092
rect 7276 9052 7316 9092
rect 7358 9052 7398 9092
rect 7440 9052 7480 9092
rect 11112 9052 11152 9092
rect 11194 9052 11234 9092
rect 11276 9052 11316 9092
rect 11358 9052 11398 9092
rect 11440 9052 11480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 19112 9052 19152 9092
rect 19194 9052 19234 9092
rect 19276 9052 19316 9092
rect 19358 9052 19398 9092
rect 19440 9052 19480 9092
rect 23112 9052 23152 9092
rect 23194 9052 23234 9092
rect 23276 9052 23316 9092
rect 23358 9052 23398 9092
rect 23440 9052 23480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 31112 9052 31152 9092
rect 31194 9052 31234 9092
rect 31276 9052 31316 9092
rect 31358 9052 31398 9092
rect 31440 9052 31480 9092
rect 35112 9052 35152 9092
rect 35194 9052 35234 9092
rect 35276 9052 35316 9092
rect 35358 9052 35398 9092
rect 35440 9052 35480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 43112 9052 43152 9092
rect 43194 9052 43234 9092
rect 43276 9052 43316 9092
rect 43358 9052 43398 9092
rect 43440 9052 43480 9092
rect 47112 9052 47152 9092
rect 47194 9052 47234 9092
rect 47276 9052 47316 9092
rect 47358 9052 47398 9092
rect 47440 9052 47480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 55112 9052 55152 9092
rect 55194 9052 55234 9092
rect 55276 9052 55316 9092
rect 55358 9052 55398 9092
rect 55440 9052 55480 9092
rect 59112 9052 59152 9092
rect 59194 9052 59234 9092
rect 59276 9052 59316 9092
rect 59358 9052 59398 9092
rect 59440 9052 59480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 67112 9052 67152 9092
rect 67194 9052 67234 9092
rect 67276 9052 67316 9092
rect 67358 9052 67398 9092
rect 67440 9052 67480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 8352 8296 8392 8336
rect 8434 8296 8474 8336
rect 8516 8296 8556 8336
rect 8598 8296 8638 8336
rect 8680 8296 8720 8336
rect 12352 8296 12392 8336
rect 12434 8296 12474 8336
rect 12516 8296 12556 8336
rect 12598 8296 12638 8336
rect 12680 8296 12720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 20352 8296 20392 8336
rect 20434 8296 20474 8336
rect 20516 8296 20556 8336
rect 20598 8296 20638 8336
rect 20680 8296 20720 8336
rect 24352 8296 24392 8336
rect 24434 8296 24474 8336
rect 24516 8296 24556 8336
rect 24598 8296 24638 8336
rect 24680 8296 24720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 32352 8296 32392 8336
rect 32434 8296 32474 8336
rect 32516 8296 32556 8336
rect 32598 8296 32638 8336
rect 32680 8296 32720 8336
rect 36352 8296 36392 8336
rect 36434 8296 36474 8336
rect 36516 8296 36556 8336
rect 36598 8296 36638 8336
rect 36680 8296 36720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 44352 8296 44392 8336
rect 44434 8296 44474 8336
rect 44516 8296 44556 8336
rect 44598 8296 44638 8336
rect 44680 8296 44720 8336
rect 48352 8296 48392 8336
rect 48434 8296 48474 8336
rect 48516 8296 48556 8336
rect 48598 8296 48638 8336
rect 48680 8296 48720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 56352 8296 56392 8336
rect 56434 8296 56474 8336
rect 56516 8296 56556 8336
rect 56598 8296 56638 8336
rect 56680 8296 56720 8336
rect 60352 8296 60392 8336
rect 60434 8296 60474 8336
rect 60516 8296 60556 8336
rect 60598 8296 60638 8336
rect 60680 8296 60720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 68352 8296 68392 8336
rect 68434 8296 68474 8336
rect 68516 8296 68556 8336
rect 68598 8296 68638 8336
rect 68680 8296 68720 8336
rect 93772 7792 93812 7832
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 7112 7540 7152 7580
rect 7194 7540 7234 7580
rect 7276 7540 7316 7580
rect 7358 7540 7398 7580
rect 7440 7540 7480 7580
rect 11112 7540 11152 7580
rect 11194 7540 11234 7580
rect 11276 7540 11316 7580
rect 11358 7540 11398 7580
rect 11440 7540 11480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 19112 7540 19152 7580
rect 19194 7540 19234 7580
rect 19276 7540 19316 7580
rect 19358 7540 19398 7580
rect 19440 7540 19480 7580
rect 23112 7540 23152 7580
rect 23194 7540 23234 7580
rect 23276 7540 23316 7580
rect 23358 7540 23398 7580
rect 23440 7540 23480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 31112 7540 31152 7580
rect 31194 7540 31234 7580
rect 31276 7540 31316 7580
rect 31358 7540 31398 7580
rect 31440 7540 31480 7580
rect 35112 7540 35152 7580
rect 35194 7540 35234 7580
rect 35276 7540 35316 7580
rect 35358 7540 35398 7580
rect 35440 7540 35480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 43112 7540 43152 7580
rect 43194 7540 43234 7580
rect 43276 7540 43316 7580
rect 43358 7540 43398 7580
rect 43440 7540 43480 7580
rect 47112 7540 47152 7580
rect 47194 7540 47234 7580
rect 47276 7540 47316 7580
rect 47358 7540 47398 7580
rect 47440 7540 47480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 55112 7540 55152 7580
rect 55194 7540 55234 7580
rect 55276 7540 55316 7580
rect 55358 7540 55398 7580
rect 55440 7540 55480 7580
rect 59112 7540 59152 7580
rect 59194 7540 59234 7580
rect 59276 7540 59316 7580
rect 59358 7540 59398 7580
rect 59440 7540 59480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 67112 7540 67152 7580
rect 67194 7540 67234 7580
rect 67276 7540 67316 7580
rect 67358 7540 67398 7580
rect 67440 7540 67480 7580
rect 86668 7456 86708 7496
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 8352 6784 8392 6824
rect 8434 6784 8474 6824
rect 8516 6784 8556 6824
rect 8598 6784 8638 6824
rect 8680 6784 8720 6824
rect 12352 6784 12392 6824
rect 12434 6784 12474 6824
rect 12516 6784 12556 6824
rect 12598 6784 12638 6824
rect 12680 6784 12720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 20352 6784 20392 6824
rect 20434 6784 20474 6824
rect 20516 6784 20556 6824
rect 20598 6784 20638 6824
rect 20680 6784 20720 6824
rect 24352 6784 24392 6824
rect 24434 6784 24474 6824
rect 24516 6784 24556 6824
rect 24598 6784 24638 6824
rect 24680 6784 24720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 32352 6784 32392 6824
rect 32434 6784 32474 6824
rect 32516 6784 32556 6824
rect 32598 6784 32638 6824
rect 32680 6784 32720 6824
rect 36352 6784 36392 6824
rect 36434 6784 36474 6824
rect 36516 6784 36556 6824
rect 36598 6784 36638 6824
rect 36680 6784 36720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 44352 6784 44392 6824
rect 44434 6784 44474 6824
rect 44516 6784 44556 6824
rect 44598 6784 44638 6824
rect 44680 6784 44720 6824
rect 48352 6784 48392 6824
rect 48434 6784 48474 6824
rect 48516 6784 48556 6824
rect 48598 6784 48638 6824
rect 48680 6784 48720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 56352 6784 56392 6824
rect 56434 6784 56474 6824
rect 56516 6784 56556 6824
rect 56598 6784 56638 6824
rect 56680 6784 56720 6824
rect 60352 6784 60392 6824
rect 60434 6784 60474 6824
rect 60516 6784 60556 6824
rect 60598 6784 60638 6824
rect 60680 6784 60720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 68352 6784 68392 6824
rect 68434 6784 68474 6824
rect 68516 6784 68556 6824
rect 68598 6784 68638 6824
rect 68680 6784 68720 6824
rect 93772 6616 93812 6656
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 7112 6028 7152 6068
rect 7194 6028 7234 6068
rect 7276 6028 7316 6068
rect 7358 6028 7398 6068
rect 7440 6028 7480 6068
rect 11112 6028 11152 6068
rect 11194 6028 11234 6068
rect 11276 6028 11316 6068
rect 11358 6028 11398 6068
rect 11440 6028 11480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 19112 6028 19152 6068
rect 19194 6028 19234 6068
rect 19276 6028 19316 6068
rect 19358 6028 19398 6068
rect 19440 6028 19480 6068
rect 23112 6028 23152 6068
rect 23194 6028 23234 6068
rect 23276 6028 23316 6068
rect 23358 6028 23398 6068
rect 23440 6028 23480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 31112 6028 31152 6068
rect 31194 6028 31234 6068
rect 31276 6028 31316 6068
rect 31358 6028 31398 6068
rect 31440 6028 31480 6068
rect 35112 6028 35152 6068
rect 35194 6028 35234 6068
rect 35276 6028 35316 6068
rect 35358 6028 35398 6068
rect 35440 6028 35480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 43112 6028 43152 6068
rect 43194 6028 43234 6068
rect 43276 6028 43316 6068
rect 43358 6028 43398 6068
rect 43440 6028 43480 6068
rect 47112 6028 47152 6068
rect 47194 6028 47234 6068
rect 47276 6028 47316 6068
rect 47358 6028 47398 6068
rect 47440 6028 47480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 55112 6028 55152 6068
rect 55194 6028 55234 6068
rect 55276 6028 55316 6068
rect 55358 6028 55398 6068
rect 55440 6028 55480 6068
rect 59112 6028 59152 6068
rect 59194 6028 59234 6068
rect 59276 6028 59316 6068
rect 59358 6028 59398 6068
rect 59440 6028 59480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 67112 6028 67152 6068
rect 67194 6028 67234 6068
rect 67276 6028 67316 6068
rect 67358 6028 67398 6068
rect 67440 6028 67480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 8352 5272 8392 5312
rect 8434 5272 8474 5312
rect 8516 5272 8556 5312
rect 8598 5272 8638 5312
rect 8680 5272 8720 5312
rect 12352 5272 12392 5312
rect 12434 5272 12474 5312
rect 12516 5272 12556 5312
rect 12598 5272 12638 5312
rect 12680 5272 12720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 20352 5272 20392 5312
rect 20434 5272 20474 5312
rect 20516 5272 20556 5312
rect 20598 5272 20638 5312
rect 20680 5272 20720 5312
rect 24352 5272 24392 5312
rect 24434 5272 24474 5312
rect 24516 5272 24556 5312
rect 24598 5272 24638 5312
rect 24680 5272 24720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 32352 5272 32392 5312
rect 32434 5272 32474 5312
rect 32516 5272 32556 5312
rect 32598 5272 32638 5312
rect 32680 5272 32720 5312
rect 36352 5272 36392 5312
rect 36434 5272 36474 5312
rect 36516 5272 36556 5312
rect 36598 5272 36638 5312
rect 36680 5272 36720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 44352 5272 44392 5312
rect 44434 5272 44474 5312
rect 44516 5272 44556 5312
rect 44598 5272 44638 5312
rect 44680 5272 44720 5312
rect 48352 5272 48392 5312
rect 48434 5272 48474 5312
rect 48516 5272 48556 5312
rect 48598 5272 48638 5312
rect 48680 5272 48720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 56352 5272 56392 5312
rect 56434 5272 56474 5312
rect 56516 5272 56556 5312
rect 56598 5272 56638 5312
rect 56680 5272 56720 5312
rect 60352 5272 60392 5312
rect 60434 5272 60474 5312
rect 60516 5272 60556 5312
rect 60598 5272 60638 5312
rect 60680 5272 60720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 68352 5272 68392 5312
rect 68434 5272 68474 5312
rect 68516 5272 68556 5312
rect 68598 5272 68638 5312
rect 68680 5272 68720 5312
rect 72352 5272 72392 5312
rect 72434 5272 72474 5312
rect 72516 5272 72556 5312
rect 72598 5272 72638 5312
rect 72680 5272 72720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 80352 5272 80392 5312
rect 80434 5272 80474 5312
rect 80516 5272 80556 5312
rect 80598 5272 80638 5312
rect 80680 5272 80720 5312
rect 84352 5272 84392 5312
rect 84434 5272 84474 5312
rect 84516 5272 84556 5312
rect 84598 5272 84638 5312
rect 84680 5272 84720 5312
rect 88352 5272 88392 5312
rect 88434 5272 88474 5312
rect 88516 5272 88556 5312
rect 88598 5272 88638 5312
rect 88680 5272 88720 5312
rect 92352 5272 92392 5312
rect 92434 5272 92474 5312
rect 92516 5272 92556 5312
rect 92598 5272 92638 5312
rect 92680 5272 92720 5312
rect 96352 5272 96392 5312
rect 96434 5272 96474 5312
rect 96516 5272 96556 5312
rect 96598 5272 96638 5312
rect 96680 5272 96720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 7112 4516 7152 4556
rect 7194 4516 7234 4556
rect 7276 4516 7316 4556
rect 7358 4516 7398 4556
rect 7440 4516 7480 4556
rect 11112 4516 11152 4556
rect 11194 4516 11234 4556
rect 11276 4516 11316 4556
rect 11358 4516 11398 4556
rect 11440 4516 11480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 19112 4516 19152 4556
rect 19194 4516 19234 4556
rect 19276 4516 19316 4556
rect 19358 4516 19398 4556
rect 19440 4516 19480 4556
rect 23112 4516 23152 4556
rect 23194 4516 23234 4556
rect 23276 4516 23316 4556
rect 23358 4516 23398 4556
rect 23440 4516 23480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 31112 4516 31152 4556
rect 31194 4516 31234 4556
rect 31276 4516 31316 4556
rect 31358 4516 31398 4556
rect 31440 4516 31480 4556
rect 35112 4516 35152 4556
rect 35194 4516 35234 4556
rect 35276 4516 35316 4556
rect 35358 4516 35398 4556
rect 35440 4516 35480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 43112 4516 43152 4556
rect 43194 4516 43234 4556
rect 43276 4516 43316 4556
rect 43358 4516 43398 4556
rect 43440 4516 43480 4556
rect 47112 4516 47152 4556
rect 47194 4516 47234 4556
rect 47276 4516 47316 4556
rect 47358 4516 47398 4556
rect 47440 4516 47480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 55112 4516 55152 4556
rect 55194 4516 55234 4556
rect 55276 4516 55316 4556
rect 55358 4516 55398 4556
rect 55440 4516 55480 4556
rect 59112 4516 59152 4556
rect 59194 4516 59234 4556
rect 59276 4516 59316 4556
rect 59358 4516 59398 4556
rect 59440 4516 59480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 67112 4516 67152 4556
rect 67194 4516 67234 4556
rect 67276 4516 67316 4556
rect 67358 4516 67398 4556
rect 67440 4516 67480 4556
rect 71112 4516 71152 4556
rect 71194 4516 71234 4556
rect 71276 4516 71316 4556
rect 71358 4516 71398 4556
rect 71440 4516 71480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 79112 4516 79152 4556
rect 79194 4516 79234 4556
rect 79276 4516 79316 4556
rect 79358 4516 79398 4556
rect 79440 4516 79480 4556
rect 83112 4516 83152 4556
rect 83194 4516 83234 4556
rect 83276 4516 83316 4556
rect 83358 4516 83398 4556
rect 83440 4516 83480 4556
rect 87112 4516 87152 4556
rect 87194 4516 87234 4556
rect 87276 4516 87316 4556
rect 87358 4516 87398 4556
rect 87440 4516 87480 4556
rect 91112 4516 91152 4556
rect 91194 4516 91234 4556
rect 91276 4516 91316 4556
rect 91358 4516 91398 4556
rect 91440 4516 91480 4556
rect 95112 4516 95152 4556
rect 95194 4516 95234 4556
rect 95276 4516 95316 4556
rect 95358 4516 95398 4556
rect 95440 4516 95480 4556
rect 99112 4516 99152 4556
rect 99194 4516 99234 4556
rect 99276 4516 99316 4556
rect 99358 4516 99398 4556
rect 99440 4516 99480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 8352 3760 8392 3800
rect 8434 3760 8474 3800
rect 8516 3760 8556 3800
rect 8598 3760 8638 3800
rect 8680 3760 8720 3800
rect 12352 3760 12392 3800
rect 12434 3760 12474 3800
rect 12516 3760 12556 3800
rect 12598 3760 12638 3800
rect 12680 3760 12720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 20352 3760 20392 3800
rect 20434 3760 20474 3800
rect 20516 3760 20556 3800
rect 20598 3760 20638 3800
rect 20680 3760 20720 3800
rect 24352 3760 24392 3800
rect 24434 3760 24474 3800
rect 24516 3760 24556 3800
rect 24598 3760 24638 3800
rect 24680 3760 24720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 32352 3760 32392 3800
rect 32434 3760 32474 3800
rect 32516 3760 32556 3800
rect 32598 3760 32638 3800
rect 32680 3760 32720 3800
rect 36352 3760 36392 3800
rect 36434 3760 36474 3800
rect 36516 3760 36556 3800
rect 36598 3760 36638 3800
rect 36680 3760 36720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 44352 3760 44392 3800
rect 44434 3760 44474 3800
rect 44516 3760 44556 3800
rect 44598 3760 44638 3800
rect 44680 3760 44720 3800
rect 48352 3760 48392 3800
rect 48434 3760 48474 3800
rect 48516 3760 48556 3800
rect 48598 3760 48638 3800
rect 48680 3760 48720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 56352 3760 56392 3800
rect 56434 3760 56474 3800
rect 56516 3760 56556 3800
rect 56598 3760 56638 3800
rect 56680 3760 56720 3800
rect 60352 3760 60392 3800
rect 60434 3760 60474 3800
rect 60516 3760 60556 3800
rect 60598 3760 60638 3800
rect 60680 3760 60720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 68352 3760 68392 3800
rect 68434 3760 68474 3800
rect 68516 3760 68556 3800
rect 68598 3760 68638 3800
rect 68680 3760 68720 3800
rect 72352 3760 72392 3800
rect 72434 3760 72474 3800
rect 72516 3760 72556 3800
rect 72598 3760 72638 3800
rect 72680 3760 72720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 80352 3760 80392 3800
rect 80434 3760 80474 3800
rect 80516 3760 80556 3800
rect 80598 3760 80638 3800
rect 80680 3760 80720 3800
rect 84352 3760 84392 3800
rect 84434 3760 84474 3800
rect 84516 3760 84556 3800
rect 84598 3760 84638 3800
rect 84680 3760 84720 3800
rect 88352 3760 88392 3800
rect 88434 3760 88474 3800
rect 88516 3760 88556 3800
rect 88598 3760 88638 3800
rect 88680 3760 88720 3800
rect 92352 3760 92392 3800
rect 92434 3760 92474 3800
rect 92516 3760 92556 3800
rect 92598 3760 92638 3800
rect 92680 3760 92720 3800
rect 96352 3760 96392 3800
rect 96434 3760 96474 3800
rect 96516 3760 96556 3800
rect 96598 3760 96638 3800
rect 96680 3760 96720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 7112 3004 7152 3044
rect 7194 3004 7234 3044
rect 7276 3004 7316 3044
rect 7358 3004 7398 3044
rect 7440 3004 7480 3044
rect 11112 3004 11152 3044
rect 11194 3004 11234 3044
rect 11276 3004 11316 3044
rect 11358 3004 11398 3044
rect 11440 3004 11480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 19112 3004 19152 3044
rect 19194 3004 19234 3044
rect 19276 3004 19316 3044
rect 19358 3004 19398 3044
rect 19440 3004 19480 3044
rect 23112 3004 23152 3044
rect 23194 3004 23234 3044
rect 23276 3004 23316 3044
rect 23358 3004 23398 3044
rect 23440 3004 23480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 31112 3004 31152 3044
rect 31194 3004 31234 3044
rect 31276 3004 31316 3044
rect 31358 3004 31398 3044
rect 31440 3004 31480 3044
rect 35112 3004 35152 3044
rect 35194 3004 35234 3044
rect 35276 3004 35316 3044
rect 35358 3004 35398 3044
rect 35440 3004 35480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 43112 3004 43152 3044
rect 43194 3004 43234 3044
rect 43276 3004 43316 3044
rect 43358 3004 43398 3044
rect 43440 3004 43480 3044
rect 47112 3004 47152 3044
rect 47194 3004 47234 3044
rect 47276 3004 47316 3044
rect 47358 3004 47398 3044
rect 47440 3004 47480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 55112 3004 55152 3044
rect 55194 3004 55234 3044
rect 55276 3004 55316 3044
rect 55358 3004 55398 3044
rect 55440 3004 55480 3044
rect 59112 3004 59152 3044
rect 59194 3004 59234 3044
rect 59276 3004 59316 3044
rect 59358 3004 59398 3044
rect 59440 3004 59480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 67112 3004 67152 3044
rect 67194 3004 67234 3044
rect 67276 3004 67316 3044
rect 67358 3004 67398 3044
rect 67440 3004 67480 3044
rect 71112 3004 71152 3044
rect 71194 3004 71234 3044
rect 71276 3004 71316 3044
rect 71358 3004 71398 3044
rect 71440 3004 71480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 79112 3004 79152 3044
rect 79194 3004 79234 3044
rect 79276 3004 79316 3044
rect 79358 3004 79398 3044
rect 79440 3004 79480 3044
rect 83112 3004 83152 3044
rect 83194 3004 83234 3044
rect 83276 3004 83316 3044
rect 83358 3004 83398 3044
rect 83440 3004 83480 3044
rect 87112 3004 87152 3044
rect 87194 3004 87234 3044
rect 87276 3004 87316 3044
rect 87358 3004 87398 3044
rect 87440 3004 87480 3044
rect 91112 3004 91152 3044
rect 91194 3004 91234 3044
rect 91276 3004 91316 3044
rect 91358 3004 91398 3044
rect 91440 3004 91480 3044
rect 95112 3004 95152 3044
rect 95194 3004 95234 3044
rect 95276 3004 95316 3044
rect 95358 3004 95398 3044
rect 95440 3004 95480 3044
rect 99112 3004 99152 3044
rect 99194 3004 99234 3044
rect 99276 3004 99316 3044
rect 99358 3004 99398 3044
rect 99440 3004 99480 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 8352 2248 8392 2288
rect 8434 2248 8474 2288
rect 8516 2248 8556 2288
rect 8598 2248 8638 2288
rect 8680 2248 8720 2288
rect 12352 2248 12392 2288
rect 12434 2248 12474 2288
rect 12516 2248 12556 2288
rect 12598 2248 12638 2288
rect 12680 2248 12720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 20352 2248 20392 2288
rect 20434 2248 20474 2288
rect 20516 2248 20556 2288
rect 20598 2248 20638 2288
rect 20680 2248 20720 2288
rect 24352 2248 24392 2288
rect 24434 2248 24474 2288
rect 24516 2248 24556 2288
rect 24598 2248 24638 2288
rect 24680 2248 24720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 32352 2248 32392 2288
rect 32434 2248 32474 2288
rect 32516 2248 32556 2288
rect 32598 2248 32638 2288
rect 32680 2248 32720 2288
rect 36352 2248 36392 2288
rect 36434 2248 36474 2288
rect 36516 2248 36556 2288
rect 36598 2248 36638 2288
rect 36680 2248 36720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 44352 2248 44392 2288
rect 44434 2248 44474 2288
rect 44516 2248 44556 2288
rect 44598 2248 44638 2288
rect 44680 2248 44720 2288
rect 48352 2248 48392 2288
rect 48434 2248 48474 2288
rect 48516 2248 48556 2288
rect 48598 2248 48638 2288
rect 48680 2248 48720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 56352 2248 56392 2288
rect 56434 2248 56474 2288
rect 56516 2248 56556 2288
rect 56598 2248 56638 2288
rect 56680 2248 56720 2288
rect 60352 2248 60392 2288
rect 60434 2248 60474 2288
rect 60516 2248 60556 2288
rect 60598 2248 60638 2288
rect 60680 2248 60720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 68352 2248 68392 2288
rect 68434 2248 68474 2288
rect 68516 2248 68556 2288
rect 68598 2248 68638 2288
rect 68680 2248 68720 2288
rect 72352 2248 72392 2288
rect 72434 2248 72474 2288
rect 72516 2248 72556 2288
rect 72598 2248 72638 2288
rect 72680 2248 72720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 80352 2248 80392 2288
rect 80434 2248 80474 2288
rect 80516 2248 80556 2288
rect 80598 2248 80638 2288
rect 80680 2248 80720 2288
rect 84352 2248 84392 2288
rect 84434 2248 84474 2288
rect 84516 2248 84556 2288
rect 84598 2248 84638 2288
rect 84680 2248 84720 2288
rect 88352 2248 88392 2288
rect 88434 2248 88474 2288
rect 88516 2248 88556 2288
rect 88598 2248 88638 2288
rect 88680 2248 88720 2288
rect 92352 2248 92392 2288
rect 92434 2248 92474 2288
rect 92516 2248 92556 2288
rect 92598 2248 92638 2288
rect 92680 2248 92720 2288
rect 96352 2248 96392 2288
rect 96434 2248 96474 2288
rect 96516 2248 96556 2288
rect 96598 2248 96638 2288
rect 96680 2248 96720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 7112 1492 7152 1532
rect 7194 1492 7234 1532
rect 7276 1492 7316 1532
rect 7358 1492 7398 1532
rect 7440 1492 7480 1532
rect 11112 1492 11152 1532
rect 11194 1492 11234 1532
rect 11276 1492 11316 1532
rect 11358 1492 11398 1532
rect 11440 1492 11480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 19112 1492 19152 1532
rect 19194 1492 19234 1532
rect 19276 1492 19316 1532
rect 19358 1492 19398 1532
rect 19440 1492 19480 1532
rect 23112 1492 23152 1532
rect 23194 1492 23234 1532
rect 23276 1492 23316 1532
rect 23358 1492 23398 1532
rect 23440 1492 23480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 31112 1492 31152 1532
rect 31194 1492 31234 1532
rect 31276 1492 31316 1532
rect 31358 1492 31398 1532
rect 31440 1492 31480 1532
rect 35112 1492 35152 1532
rect 35194 1492 35234 1532
rect 35276 1492 35316 1532
rect 35358 1492 35398 1532
rect 35440 1492 35480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 43112 1492 43152 1532
rect 43194 1492 43234 1532
rect 43276 1492 43316 1532
rect 43358 1492 43398 1532
rect 43440 1492 43480 1532
rect 47112 1492 47152 1532
rect 47194 1492 47234 1532
rect 47276 1492 47316 1532
rect 47358 1492 47398 1532
rect 47440 1492 47480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 55112 1492 55152 1532
rect 55194 1492 55234 1532
rect 55276 1492 55316 1532
rect 55358 1492 55398 1532
rect 55440 1492 55480 1532
rect 59112 1492 59152 1532
rect 59194 1492 59234 1532
rect 59276 1492 59316 1532
rect 59358 1492 59398 1532
rect 59440 1492 59480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 67112 1492 67152 1532
rect 67194 1492 67234 1532
rect 67276 1492 67316 1532
rect 67358 1492 67398 1532
rect 67440 1492 67480 1532
rect 71112 1492 71152 1532
rect 71194 1492 71234 1532
rect 71276 1492 71316 1532
rect 71358 1492 71398 1532
rect 71440 1492 71480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 79112 1492 79152 1532
rect 79194 1492 79234 1532
rect 79276 1492 79316 1532
rect 79358 1492 79398 1532
rect 79440 1492 79480 1532
rect 83112 1492 83152 1532
rect 83194 1492 83234 1532
rect 83276 1492 83316 1532
rect 83358 1492 83398 1532
rect 83440 1492 83480 1532
rect 87112 1492 87152 1532
rect 87194 1492 87234 1532
rect 87276 1492 87316 1532
rect 87358 1492 87398 1532
rect 87440 1492 87480 1532
rect 91112 1492 91152 1532
rect 91194 1492 91234 1532
rect 91276 1492 91316 1532
rect 91358 1492 91398 1532
rect 91440 1492 91480 1532
rect 95112 1492 95152 1532
rect 95194 1492 95234 1532
rect 95276 1492 95316 1532
rect 95358 1492 95398 1532
rect 95440 1492 95480 1532
rect 99112 1492 99152 1532
rect 99194 1492 99234 1532
rect 99276 1492 99316 1532
rect 99358 1492 99398 1532
rect 99440 1492 99480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 8352 736 8392 776
rect 8434 736 8474 776
rect 8516 736 8556 776
rect 8598 736 8638 776
rect 8680 736 8720 776
rect 12352 736 12392 776
rect 12434 736 12474 776
rect 12516 736 12556 776
rect 12598 736 12638 776
rect 12680 736 12720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 20352 736 20392 776
rect 20434 736 20474 776
rect 20516 736 20556 776
rect 20598 736 20638 776
rect 20680 736 20720 776
rect 24352 736 24392 776
rect 24434 736 24474 776
rect 24516 736 24556 776
rect 24598 736 24638 776
rect 24680 736 24720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 32352 736 32392 776
rect 32434 736 32474 776
rect 32516 736 32556 776
rect 32598 736 32638 776
rect 32680 736 32720 776
rect 36352 736 36392 776
rect 36434 736 36474 776
rect 36516 736 36556 776
rect 36598 736 36638 776
rect 36680 736 36720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 44352 736 44392 776
rect 44434 736 44474 776
rect 44516 736 44556 776
rect 44598 736 44638 776
rect 44680 736 44720 776
rect 48352 736 48392 776
rect 48434 736 48474 776
rect 48516 736 48556 776
rect 48598 736 48638 776
rect 48680 736 48720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 56352 736 56392 776
rect 56434 736 56474 776
rect 56516 736 56556 776
rect 56598 736 56638 776
rect 56680 736 56720 776
rect 60352 736 60392 776
rect 60434 736 60474 776
rect 60516 736 60556 776
rect 60598 736 60638 776
rect 60680 736 60720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 68352 736 68392 776
rect 68434 736 68474 776
rect 68516 736 68556 776
rect 68598 736 68638 776
rect 68680 736 68720 776
rect 72352 736 72392 776
rect 72434 736 72474 776
rect 72516 736 72556 776
rect 72598 736 72638 776
rect 72680 736 72720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
rect 80352 736 80392 776
rect 80434 736 80474 776
rect 80516 736 80556 776
rect 80598 736 80638 776
rect 80680 736 80720 776
rect 84352 736 84392 776
rect 84434 736 84474 776
rect 84516 736 84556 776
rect 84598 736 84638 776
rect 84680 736 84720 776
rect 88352 736 88392 776
rect 88434 736 88474 776
rect 88516 736 88556 776
rect 88598 736 88638 776
rect 88680 736 88720 776
rect 92352 736 92392 776
rect 92434 736 92474 776
rect 92516 736 92556 776
rect 92598 736 92638 776
rect 92680 736 92720 776
rect 96352 736 96392 776
rect 96434 736 96474 776
rect 96516 736 96556 776
rect 96598 736 96638 776
rect 96680 736 96720 776
<< metal4 >>
rect 4352 38576 4720 38585
rect 4392 38536 4434 38576
rect 4474 38536 4516 38576
rect 4556 38536 4598 38576
rect 4638 38536 4680 38576
rect 4352 38527 4720 38536
rect 8352 38576 8720 38585
rect 8392 38536 8434 38576
rect 8474 38536 8516 38576
rect 8556 38536 8598 38576
rect 8638 38536 8680 38576
rect 8352 38527 8720 38536
rect 12352 38576 12720 38585
rect 12392 38536 12434 38576
rect 12474 38536 12516 38576
rect 12556 38536 12598 38576
rect 12638 38536 12680 38576
rect 12352 38527 12720 38536
rect 16352 38576 16720 38585
rect 16392 38536 16434 38576
rect 16474 38536 16516 38576
rect 16556 38536 16598 38576
rect 16638 38536 16680 38576
rect 16352 38527 16720 38536
rect 20352 38576 20720 38585
rect 20392 38536 20434 38576
rect 20474 38536 20516 38576
rect 20556 38536 20598 38576
rect 20638 38536 20680 38576
rect 20352 38527 20720 38536
rect 24352 38576 24720 38585
rect 24392 38536 24434 38576
rect 24474 38536 24516 38576
rect 24556 38536 24598 38576
rect 24638 38536 24680 38576
rect 24352 38527 24720 38536
rect 28352 38576 28720 38585
rect 28392 38536 28434 38576
rect 28474 38536 28516 38576
rect 28556 38536 28598 38576
rect 28638 38536 28680 38576
rect 28352 38527 28720 38536
rect 32352 38576 32720 38585
rect 32392 38536 32434 38576
rect 32474 38536 32516 38576
rect 32556 38536 32598 38576
rect 32638 38536 32680 38576
rect 32352 38527 32720 38536
rect 36352 38576 36720 38585
rect 36392 38536 36434 38576
rect 36474 38536 36516 38576
rect 36556 38536 36598 38576
rect 36638 38536 36680 38576
rect 36352 38527 36720 38536
rect 40352 38576 40720 38585
rect 40392 38536 40434 38576
rect 40474 38536 40516 38576
rect 40556 38536 40598 38576
rect 40638 38536 40680 38576
rect 40352 38527 40720 38536
rect 44352 38576 44720 38585
rect 44392 38536 44434 38576
rect 44474 38536 44516 38576
rect 44556 38536 44598 38576
rect 44638 38536 44680 38576
rect 44352 38527 44720 38536
rect 48352 38576 48720 38585
rect 48392 38536 48434 38576
rect 48474 38536 48516 38576
rect 48556 38536 48598 38576
rect 48638 38536 48680 38576
rect 48352 38527 48720 38536
rect 52352 38576 52720 38585
rect 52392 38536 52434 38576
rect 52474 38536 52516 38576
rect 52556 38536 52598 38576
rect 52638 38536 52680 38576
rect 52352 38527 52720 38536
rect 56352 38576 56720 38585
rect 56392 38536 56434 38576
rect 56474 38536 56516 38576
rect 56556 38536 56598 38576
rect 56638 38536 56680 38576
rect 56352 38527 56720 38536
rect 60352 38576 60720 38585
rect 60392 38536 60434 38576
rect 60474 38536 60516 38576
rect 60556 38536 60598 38576
rect 60638 38536 60680 38576
rect 60352 38527 60720 38536
rect 64352 38576 64720 38585
rect 64392 38536 64434 38576
rect 64474 38536 64516 38576
rect 64556 38536 64598 38576
rect 64638 38536 64680 38576
rect 64352 38527 64720 38536
rect 68352 38576 68720 38585
rect 68392 38536 68434 38576
rect 68474 38536 68516 38576
rect 68556 38536 68598 38576
rect 68638 38536 68680 38576
rect 68352 38527 68720 38536
rect 72352 38576 72720 38585
rect 72392 38536 72434 38576
rect 72474 38536 72516 38576
rect 72556 38536 72598 38576
rect 72638 38536 72680 38576
rect 72352 38527 72720 38536
rect 76352 38576 76720 38585
rect 76392 38536 76434 38576
rect 76474 38536 76516 38576
rect 76556 38536 76598 38576
rect 76638 38536 76680 38576
rect 76352 38527 76720 38536
rect 80352 38576 80720 38585
rect 80392 38536 80434 38576
rect 80474 38536 80516 38576
rect 80556 38536 80598 38576
rect 80638 38536 80680 38576
rect 80352 38527 80720 38536
rect 84352 38576 84720 38585
rect 84392 38536 84434 38576
rect 84474 38536 84516 38576
rect 84556 38536 84598 38576
rect 84638 38536 84680 38576
rect 84352 38527 84720 38536
rect 88352 38576 88720 38585
rect 88392 38536 88434 38576
rect 88474 38536 88516 38576
rect 88556 38536 88598 38576
rect 88638 38536 88680 38576
rect 88352 38527 88720 38536
rect 92352 38576 92720 38585
rect 92392 38536 92434 38576
rect 92474 38536 92516 38576
rect 92556 38536 92598 38576
rect 92638 38536 92680 38576
rect 92352 38527 92720 38536
rect 96352 38576 96720 38585
rect 96392 38536 96434 38576
rect 96474 38536 96516 38576
rect 96556 38536 96598 38576
rect 96638 38536 96680 38576
rect 96352 38527 96720 38536
rect 3112 37820 3480 37829
rect 3152 37780 3194 37820
rect 3234 37780 3276 37820
rect 3316 37780 3358 37820
rect 3398 37780 3440 37820
rect 3112 37771 3480 37780
rect 7112 37820 7480 37829
rect 7152 37780 7194 37820
rect 7234 37780 7276 37820
rect 7316 37780 7358 37820
rect 7398 37780 7440 37820
rect 7112 37771 7480 37780
rect 11112 37820 11480 37829
rect 11152 37780 11194 37820
rect 11234 37780 11276 37820
rect 11316 37780 11358 37820
rect 11398 37780 11440 37820
rect 11112 37771 11480 37780
rect 15112 37820 15480 37829
rect 15152 37780 15194 37820
rect 15234 37780 15276 37820
rect 15316 37780 15358 37820
rect 15398 37780 15440 37820
rect 15112 37771 15480 37780
rect 19112 37820 19480 37829
rect 19152 37780 19194 37820
rect 19234 37780 19276 37820
rect 19316 37780 19358 37820
rect 19398 37780 19440 37820
rect 19112 37771 19480 37780
rect 23112 37820 23480 37829
rect 23152 37780 23194 37820
rect 23234 37780 23276 37820
rect 23316 37780 23358 37820
rect 23398 37780 23440 37820
rect 23112 37771 23480 37780
rect 27112 37820 27480 37829
rect 27152 37780 27194 37820
rect 27234 37780 27276 37820
rect 27316 37780 27358 37820
rect 27398 37780 27440 37820
rect 27112 37771 27480 37780
rect 31112 37820 31480 37829
rect 31152 37780 31194 37820
rect 31234 37780 31276 37820
rect 31316 37780 31358 37820
rect 31398 37780 31440 37820
rect 31112 37771 31480 37780
rect 35112 37820 35480 37829
rect 35152 37780 35194 37820
rect 35234 37780 35276 37820
rect 35316 37780 35358 37820
rect 35398 37780 35440 37820
rect 35112 37771 35480 37780
rect 39112 37820 39480 37829
rect 39152 37780 39194 37820
rect 39234 37780 39276 37820
rect 39316 37780 39358 37820
rect 39398 37780 39440 37820
rect 39112 37771 39480 37780
rect 43112 37820 43480 37829
rect 43152 37780 43194 37820
rect 43234 37780 43276 37820
rect 43316 37780 43358 37820
rect 43398 37780 43440 37820
rect 43112 37771 43480 37780
rect 47112 37820 47480 37829
rect 47152 37780 47194 37820
rect 47234 37780 47276 37820
rect 47316 37780 47358 37820
rect 47398 37780 47440 37820
rect 47112 37771 47480 37780
rect 51112 37820 51480 37829
rect 51152 37780 51194 37820
rect 51234 37780 51276 37820
rect 51316 37780 51358 37820
rect 51398 37780 51440 37820
rect 51112 37771 51480 37780
rect 55112 37820 55480 37829
rect 55152 37780 55194 37820
rect 55234 37780 55276 37820
rect 55316 37780 55358 37820
rect 55398 37780 55440 37820
rect 55112 37771 55480 37780
rect 59112 37820 59480 37829
rect 59152 37780 59194 37820
rect 59234 37780 59276 37820
rect 59316 37780 59358 37820
rect 59398 37780 59440 37820
rect 59112 37771 59480 37780
rect 63112 37820 63480 37829
rect 63152 37780 63194 37820
rect 63234 37780 63276 37820
rect 63316 37780 63358 37820
rect 63398 37780 63440 37820
rect 63112 37771 63480 37780
rect 67112 37820 67480 37829
rect 67152 37780 67194 37820
rect 67234 37780 67276 37820
rect 67316 37780 67358 37820
rect 67398 37780 67440 37820
rect 67112 37771 67480 37780
rect 71112 37820 71480 37829
rect 71152 37780 71194 37820
rect 71234 37780 71276 37820
rect 71316 37780 71358 37820
rect 71398 37780 71440 37820
rect 71112 37771 71480 37780
rect 75112 37820 75480 37829
rect 75152 37780 75194 37820
rect 75234 37780 75276 37820
rect 75316 37780 75358 37820
rect 75398 37780 75440 37820
rect 75112 37771 75480 37780
rect 79112 37820 79480 37829
rect 79152 37780 79194 37820
rect 79234 37780 79276 37820
rect 79316 37780 79358 37820
rect 79398 37780 79440 37820
rect 79112 37771 79480 37780
rect 83112 37820 83480 37829
rect 83152 37780 83194 37820
rect 83234 37780 83276 37820
rect 83316 37780 83358 37820
rect 83398 37780 83440 37820
rect 83112 37771 83480 37780
rect 87112 37820 87480 37829
rect 87152 37780 87194 37820
rect 87234 37780 87276 37820
rect 87316 37780 87358 37820
rect 87398 37780 87440 37820
rect 87112 37771 87480 37780
rect 91112 37820 91480 37829
rect 91152 37780 91194 37820
rect 91234 37780 91276 37820
rect 91316 37780 91358 37820
rect 91398 37780 91440 37820
rect 91112 37771 91480 37780
rect 95112 37820 95480 37829
rect 95152 37780 95194 37820
rect 95234 37780 95276 37820
rect 95316 37780 95358 37820
rect 95398 37780 95440 37820
rect 95112 37771 95480 37780
rect 99112 37820 99480 37829
rect 99152 37780 99194 37820
rect 99234 37780 99276 37820
rect 99316 37780 99358 37820
rect 99398 37780 99440 37820
rect 99112 37771 99480 37780
rect 4352 37064 4720 37073
rect 4392 37024 4434 37064
rect 4474 37024 4516 37064
rect 4556 37024 4598 37064
rect 4638 37024 4680 37064
rect 4352 37015 4720 37024
rect 8352 37064 8720 37073
rect 8392 37024 8434 37064
rect 8474 37024 8516 37064
rect 8556 37024 8598 37064
rect 8638 37024 8680 37064
rect 8352 37015 8720 37024
rect 12352 37064 12720 37073
rect 12392 37024 12434 37064
rect 12474 37024 12516 37064
rect 12556 37024 12598 37064
rect 12638 37024 12680 37064
rect 12352 37015 12720 37024
rect 16352 37064 16720 37073
rect 16392 37024 16434 37064
rect 16474 37024 16516 37064
rect 16556 37024 16598 37064
rect 16638 37024 16680 37064
rect 16352 37015 16720 37024
rect 20352 37064 20720 37073
rect 20392 37024 20434 37064
rect 20474 37024 20516 37064
rect 20556 37024 20598 37064
rect 20638 37024 20680 37064
rect 20352 37015 20720 37024
rect 24352 37064 24720 37073
rect 24392 37024 24434 37064
rect 24474 37024 24516 37064
rect 24556 37024 24598 37064
rect 24638 37024 24680 37064
rect 24352 37015 24720 37024
rect 28352 37064 28720 37073
rect 28392 37024 28434 37064
rect 28474 37024 28516 37064
rect 28556 37024 28598 37064
rect 28638 37024 28680 37064
rect 28352 37015 28720 37024
rect 32352 37064 32720 37073
rect 32392 37024 32434 37064
rect 32474 37024 32516 37064
rect 32556 37024 32598 37064
rect 32638 37024 32680 37064
rect 32352 37015 32720 37024
rect 36352 37064 36720 37073
rect 36392 37024 36434 37064
rect 36474 37024 36516 37064
rect 36556 37024 36598 37064
rect 36638 37024 36680 37064
rect 36352 37015 36720 37024
rect 40352 37064 40720 37073
rect 40392 37024 40434 37064
rect 40474 37024 40516 37064
rect 40556 37024 40598 37064
rect 40638 37024 40680 37064
rect 40352 37015 40720 37024
rect 44352 37064 44720 37073
rect 44392 37024 44434 37064
rect 44474 37024 44516 37064
rect 44556 37024 44598 37064
rect 44638 37024 44680 37064
rect 44352 37015 44720 37024
rect 48352 37064 48720 37073
rect 48392 37024 48434 37064
rect 48474 37024 48516 37064
rect 48556 37024 48598 37064
rect 48638 37024 48680 37064
rect 48352 37015 48720 37024
rect 52352 37064 52720 37073
rect 52392 37024 52434 37064
rect 52474 37024 52516 37064
rect 52556 37024 52598 37064
rect 52638 37024 52680 37064
rect 52352 37015 52720 37024
rect 56352 37064 56720 37073
rect 56392 37024 56434 37064
rect 56474 37024 56516 37064
rect 56556 37024 56598 37064
rect 56638 37024 56680 37064
rect 56352 37015 56720 37024
rect 60352 37064 60720 37073
rect 60392 37024 60434 37064
rect 60474 37024 60516 37064
rect 60556 37024 60598 37064
rect 60638 37024 60680 37064
rect 60352 37015 60720 37024
rect 64352 37064 64720 37073
rect 64392 37024 64434 37064
rect 64474 37024 64516 37064
rect 64556 37024 64598 37064
rect 64638 37024 64680 37064
rect 64352 37015 64720 37024
rect 68352 37064 68720 37073
rect 68392 37024 68434 37064
rect 68474 37024 68516 37064
rect 68556 37024 68598 37064
rect 68638 37024 68680 37064
rect 68352 37015 68720 37024
rect 72352 37064 72720 37073
rect 72392 37024 72434 37064
rect 72474 37024 72516 37064
rect 72556 37024 72598 37064
rect 72638 37024 72680 37064
rect 72352 37015 72720 37024
rect 76352 37064 76720 37073
rect 76392 37024 76434 37064
rect 76474 37024 76516 37064
rect 76556 37024 76598 37064
rect 76638 37024 76680 37064
rect 76352 37015 76720 37024
rect 80352 37064 80720 37073
rect 80392 37024 80434 37064
rect 80474 37024 80516 37064
rect 80556 37024 80598 37064
rect 80638 37024 80680 37064
rect 80352 37015 80720 37024
rect 84352 37064 84720 37073
rect 84392 37024 84434 37064
rect 84474 37024 84516 37064
rect 84556 37024 84598 37064
rect 84638 37024 84680 37064
rect 84352 37015 84720 37024
rect 88352 37064 88720 37073
rect 88392 37024 88434 37064
rect 88474 37024 88516 37064
rect 88556 37024 88598 37064
rect 88638 37024 88680 37064
rect 88352 37015 88720 37024
rect 92352 37064 92720 37073
rect 92392 37024 92434 37064
rect 92474 37024 92516 37064
rect 92556 37024 92598 37064
rect 92638 37024 92680 37064
rect 92352 37015 92720 37024
rect 96352 37064 96720 37073
rect 96392 37024 96434 37064
rect 96474 37024 96516 37064
rect 96556 37024 96598 37064
rect 96638 37024 96680 37064
rect 96352 37015 96720 37024
rect 3112 36308 3480 36317
rect 3152 36268 3194 36308
rect 3234 36268 3276 36308
rect 3316 36268 3358 36308
rect 3398 36268 3440 36308
rect 3112 36259 3480 36268
rect 7112 36308 7480 36317
rect 7152 36268 7194 36308
rect 7234 36268 7276 36308
rect 7316 36268 7358 36308
rect 7398 36268 7440 36308
rect 7112 36259 7480 36268
rect 11112 36308 11480 36317
rect 11152 36268 11194 36308
rect 11234 36268 11276 36308
rect 11316 36268 11358 36308
rect 11398 36268 11440 36308
rect 11112 36259 11480 36268
rect 15112 36308 15480 36317
rect 15152 36268 15194 36308
rect 15234 36268 15276 36308
rect 15316 36268 15358 36308
rect 15398 36268 15440 36308
rect 15112 36259 15480 36268
rect 19112 36308 19480 36317
rect 19152 36268 19194 36308
rect 19234 36268 19276 36308
rect 19316 36268 19358 36308
rect 19398 36268 19440 36308
rect 19112 36259 19480 36268
rect 23112 36308 23480 36317
rect 23152 36268 23194 36308
rect 23234 36268 23276 36308
rect 23316 36268 23358 36308
rect 23398 36268 23440 36308
rect 23112 36259 23480 36268
rect 27112 36308 27480 36317
rect 27152 36268 27194 36308
rect 27234 36268 27276 36308
rect 27316 36268 27358 36308
rect 27398 36268 27440 36308
rect 27112 36259 27480 36268
rect 31112 36308 31480 36317
rect 31152 36268 31194 36308
rect 31234 36268 31276 36308
rect 31316 36268 31358 36308
rect 31398 36268 31440 36308
rect 31112 36259 31480 36268
rect 35112 36308 35480 36317
rect 35152 36268 35194 36308
rect 35234 36268 35276 36308
rect 35316 36268 35358 36308
rect 35398 36268 35440 36308
rect 35112 36259 35480 36268
rect 39112 36308 39480 36317
rect 39152 36268 39194 36308
rect 39234 36268 39276 36308
rect 39316 36268 39358 36308
rect 39398 36268 39440 36308
rect 39112 36259 39480 36268
rect 43112 36308 43480 36317
rect 43152 36268 43194 36308
rect 43234 36268 43276 36308
rect 43316 36268 43358 36308
rect 43398 36268 43440 36308
rect 43112 36259 43480 36268
rect 47112 36308 47480 36317
rect 47152 36268 47194 36308
rect 47234 36268 47276 36308
rect 47316 36268 47358 36308
rect 47398 36268 47440 36308
rect 47112 36259 47480 36268
rect 51112 36308 51480 36317
rect 51152 36268 51194 36308
rect 51234 36268 51276 36308
rect 51316 36268 51358 36308
rect 51398 36268 51440 36308
rect 51112 36259 51480 36268
rect 55112 36308 55480 36317
rect 55152 36268 55194 36308
rect 55234 36268 55276 36308
rect 55316 36268 55358 36308
rect 55398 36268 55440 36308
rect 55112 36259 55480 36268
rect 59112 36308 59480 36317
rect 59152 36268 59194 36308
rect 59234 36268 59276 36308
rect 59316 36268 59358 36308
rect 59398 36268 59440 36308
rect 59112 36259 59480 36268
rect 63112 36308 63480 36317
rect 63152 36268 63194 36308
rect 63234 36268 63276 36308
rect 63316 36268 63358 36308
rect 63398 36268 63440 36308
rect 63112 36259 63480 36268
rect 67112 36308 67480 36317
rect 67152 36268 67194 36308
rect 67234 36268 67276 36308
rect 67316 36268 67358 36308
rect 67398 36268 67440 36308
rect 67112 36259 67480 36268
rect 71112 36308 71480 36317
rect 71152 36268 71194 36308
rect 71234 36268 71276 36308
rect 71316 36268 71358 36308
rect 71398 36268 71440 36308
rect 71112 36259 71480 36268
rect 75112 36308 75480 36317
rect 75152 36268 75194 36308
rect 75234 36268 75276 36308
rect 75316 36268 75358 36308
rect 75398 36268 75440 36308
rect 75112 36259 75480 36268
rect 79112 36308 79480 36317
rect 79152 36268 79194 36308
rect 79234 36268 79276 36308
rect 79316 36268 79358 36308
rect 79398 36268 79440 36308
rect 79112 36259 79480 36268
rect 83112 36308 83480 36317
rect 83152 36268 83194 36308
rect 83234 36268 83276 36308
rect 83316 36268 83358 36308
rect 83398 36268 83440 36308
rect 83112 36259 83480 36268
rect 87112 36308 87480 36317
rect 87152 36268 87194 36308
rect 87234 36268 87276 36308
rect 87316 36268 87358 36308
rect 87398 36268 87440 36308
rect 87112 36259 87480 36268
rect 91112 36308 91480 36317
rect 91152 36268 91194 36308
rect 91234 36268 91276 36308
rect 91316 36268 91358 36308
rect 91398 36268 91440 36308
rect 91112 36259 91480 36268
rect 95112 36308 95480 36317
rect 95152 36268 95194 36308
rect 95234 36268 95276 36308
rect 95316 36268 95358 36308
rect 95398 36268 95440 36308
rect 95112 36259 95480 36268
rect 99112 36308 99480 36317
rect 99152 36268 99194 36308
rect 99234 36268 99276 36308
rect 99316 36268 99358 36308
rect 99398 36268 99440 36308
rect 99112 36259 99480 36268
rect 4352 35552 4720 35561
rect 4392 35512 4434 35552
rect 4474 35512 4516 35552
rect 4556 35512 4598 35552
rect 4638 35512 4680 35552
rect 4352 35503 4720 35512
rect 8352 35552 8720 35561
rect 8392 35512 8434 35552
rect 8474 35512 8516 35552
rect 8556 35512 8598 35552
rect 8638 35512 8680 35552
rect 8352 35503 8720 35512
rect 12352 35552 12720 35561
rect 12392 35512 12434 35552
rect 12474 35512 12516 35552
rect 12556 35512 12598 35552
rect 12638 35512 12680 35552
rect 12352 35503 12720 35512
rect 16352 35552 16720 35561
rect 16392 35512 16434 35552
rect 16474 35512 16516 35552
rect 16556 35512 16598 35552
rect 16638 35512 16680 35552
rect 16352 35503 16720 35512
rect 20352 35552 20720 35561
rect 20392 35512 20434 35552
rect 20474 35512 20516 35552
rect 20556 35512 20598 35552
rect 20638 35512 20680 35552
rect 20352 35503 20720 35512
rect 24352 35552 24720 35561
rect 24392 35512 24434 35552
rect 24474 35512 24516 35552
rect 24556 35512 24598 35552
rect 24638 35512 24680 35552
rect 24352 35503 24720 35512
rect 28352 35552 28720 35561
rect 28392 35512 28434 35552
rect 28474 35512 28516 35552
rect 28556 35512 28598 35552
rect 28638 35512 28680 35552
rect 28352 35503 28720 35512
rect 32352 35552 32720 35561
rect 32392 35512 32434 35552
rect 32474 35512 32516 35552
rect 32556 35512 32598 35552
rect 32638 35512 32680 35552
rect 32352 35503 32720 35512
rect 36352 35552 36720 35561
rect 36392 35512 36434 35552
rect 36474 35512 36516 35552
rect 36556 35512 36598 35552
rect 36638 35512 36680 35552
rect 36352 35503 36720 35512
rect 40352 35552 40720 35561
rect 40392 35512 40434 35552
rect 40474 35512 40516 35552
rect 40556 35512 40598 35552
rect 40638 35512 40680 35552
rect 40352 35503 40720 35512
rect 44352 35552 44720 35561
rect 44392 35512 44434 35552
rect 44474 35512 44516 35552
rect 44556 35512 44598 35552
rect 44638 35512 44680 35552
rect 44352 35503 44720 35512
rect 48352 35552 48720 35561
rect 48392 35512 48434 35552
rect 48474 35512 48516 35552
rect 48556 35512 48598 35552
rect 48638 35512 48680 35552
rect 48352 35503 48720 35512
rect 52352 35552 52720 35561
rect 52392 35512 52434 35552
rect 52474 35512 52516 35552
rect 52556 35512 52598 35552
rect 52638 35512 52680 35552
rect 52352 35503 52720 35512
rect 56352 35552 56720 35561
rect 56392 35512 56434 35552
rect 56474 35512 56516 35552
rect 56556 35512 56598 35552
rect 56638 35512 56680 35552
rect 56352 35503 56720 35512
rect 60352 35552 60720 35561
rect 60392 35512 60434 35552
rect 60474 35512 60516 35552
rect 60556 35512 60598 35552
rect 60638 35512 60680 35552
rect 60352 35503 60720 35512
rect 64352 35552 64720 35561
rect 64392 35512 64434 35552
rect 64474 35512 64516 35552
rect 64556 35512 64598 35552
rect 64638 35512 64680 35552
rect 64352 35503 64720 35512
rect 68352 35552 68720 35561
rect 68392 35512 68434 35552
rect 68474 35512 68516 35552
rect 68556 35512 68598 35552
rect 68638 35512 68680 35552
rect 68352 35503 68720 35512
rect 72352 35552 72720 35561
rect 72392 35512 72434 35552
rect 72474 35512 72516 35552
rect 72556 35512 72598 35552
rect 72638 35512 72680 35552
rect 72352 35503 72720 35512
rect 76352 35552 76720 35561
rect 76392 35512 76434 35552
rect 76474 35512 76516 35552
rect 76556 35512 76598 35552
rect 76638 35512 76680 35552
rect 76352 35503 76720 35512
rect 80352 35552 80720 35561
rect 80392 35512 80434 35552
rect 80474 35512 80516 35552
rect 80556 35512 80598 35552
rect 80638 35512 80680 35552
rect 80352 35503 80720 35512
rect 84352 35552 84720 35561
rect 84392 35512 84434 35552
rect 84474 35512 84516 35552
rect 84556 35512 84598 35552
rect 84638 35512 84680 35552
rect 84352 35503 84720 35512
rect 88352 35552 88720 35561
rect 88392 35512 88434 35552
rect 88474 35512 88516 35552
rect 88556 35512 88598 35552
rect 88638 35512 88680 35552
rect 88352 35503 88720 35512
rect 92352 35552 92720 35561
rect 92392 35512 92434 35552
rect 92474 35512 92516 35552
rect 92556 35512 92598 35552
rect 92638 35512 92680 35552
rect 92352 35503 92720 35512
rect 96352 35552 96720 35561
rect 96392 35512 96434 35552
rect 96474 35512 96516 35552
rect 96556 35512 96598 35552
rect 96638 35512 96680 35552
rect 96352 35503 96720 35512
rect 3112 34796 3480 34805
rect 3152 34756 3194 34796
rect 3234 34756 3276 34796
rect 3316 34756 3358 34796
rect 3398 34756 3440 34796
rect 3112 34747 3480 34756
rect 7112 34796 7480 34805
rect 7152 34756 7194 34796
rect 7234 34756 7276 34796
rect 7316 34756 7358 34796
rect 7398 34756 7440 34796
rect 7112 34747 7480 34756
rect 11112 34796 11480 34805
rect 11152 34756 11194 34796
rect 11234 34756 11276 34796
rect 11316 34756 11358 34796
rect 11398 34756 11440 34796
rect 11112 34747 11480 34756
rect 15112 34796 15480 34805
rect 15152 34756 15194 34796
rect 15234 34756 15276 34796
rect 15316 34756 15358 34796
rect 15398 34756 15440 34796
rect 15112 34747 15480 34756
rect 19112 34796 19480 34805
rect 19152 34756 19194 34796
rect 19234 34756 19276 34796
rect 19316 34756 19358 34796
rect 19398 34756 19440 34796
rect 19112 34747 19480 34756
rect 23112 34796 23480 34805
rect 23152 34756 23194 34796
rect 23234 34756 23276 34796
rect 23316 34756 23358 34796
rect 23398 34756 23440 34796
rect 23112 34747 23480 34756
rect 27112 34796 27480 34805
rect 27152 34756 27194 34796
rect 27234 34756 27276 34796
rect 27316 34756 27358 34796
rect 27398 34756 27440 34796
rect 27112 34747 27480 34756
rect 31112 34796 31480 34805
rect 31152 34756 31194 34796
rect 31234 34756 31276 34796
rect 31316 34756 31358 34796
rect 31398 34756 31440 34796
rect 31112 34747 31480 34756
rect 35112 34796 35480 34805
rect 35152 34756 35194 34796
rect 35234 34756 35276 34796
rect 35316 34756 35358 34796
rect 35398 34756 35440 34796
rect 35112 34747 35480 34756
rect 39112 34796 39480 34805
rect 39152 34756 39194 34796
rect 39234 34756 39276 34796
rect 39316 34756 39358 34796
rect 39398 34756 39440 34796
rect 39112 34747 39480 34756
rect 43112 34796 43480 34805
rect 43152 34756 43194 34796
rect 43234 34756 43276 34796
rect 43316 34756 43358 34796
rect 43398 34756 43440 34796
rect 43112 34747 43480 34756
rect 47112 34796 47480 34805
rect 47152 34756 47194 34796
rect 47234 34756 47276 34796
rect 47316 34756 47358 34796
rect 47398 34756 47440 34796
rect 47112 34747 47480 34756
rect 51112 34796 51480 34805
rect 51152 34756 51194 34796
rect 51234 34756 51276 34796
rect 51316 34756 51358 34796
rect 51398 34756 51440 34796
rect 51112 34747 51480 34756
rect 55112 34796 55480 34805
rect 55152 34756 55194 34796
rect 55234 34756 55276 34796
rect 55316 34756 55358 34796
rect 55398 34756 55440 34796
rect 55112 34747 55480 34756
rect 59112 34796 59480 34805
rect 59152 34756 59194 34796
rect 59234 34756 59276 34796
rect 59316 34756 59358 34796
rect 59398 34756 59440 34796
rect 59112 34747 59480 34756
rect 63112 34796 63480 34805
rect 63152 34756 63194 34796
rect 63234 34756 63276 34796
rect 63316 34756 63358 34796
rect 63398 34756 63440 34796
rect 63112 34747 63480 34756
rect 67112 34796 67480 34805
rect 67152 34756 67194 34796
rect 67234 34756 67276 34796
rect 67316 34756 67358 34796
rect 67398 34756 67440 34796
rect 67112 34747 67480 34756
rect 71112 34796 71480 34805
rect 71152 34756 71194 34796
rect 71234 34756 71276 34796
rect 71316 34756 71358 34796
rect 71398 34756 71440 34796
rect 71112 34747 71480 34756
rect 75112 34796 75480 34805
rect 75152 34756 75194 34796
rect 75234 34756 75276 34796
rect 75316 34756 75358 34796
rect 75398 34756 75440 34796
rect 75112 34747 75480 34756
rect 79112 34796 79480 34805
rect 79152 34756 79194 34796
rect 79234 34756 79276 34796
rect 79316 34756 79358 34796
rect 79398 34756 79440 34796
rect 79112 34747 79480 34756
rect 83112 34796 83480 34805
rect 83152 34756 83194 34796
rect 83234 34756 83276 34796
rect 83316 34756 83358 34796
rect 83398 34756 83440 34796
rect 83112 34747 83480 34756
rect 87112 34796 87480 34805
rect 87152 34756 87194 34796
rect 87234 34756 87276 34796
rect 87316 34756 87358 34796
rect 87398 34756 87440 34796
rect 87112 34747 87480 34756
rect 91112 34796 91480 34805
rect 91152 34756 91194 34796
rect 91234 34756 91276 34796
rect 91316 34756 91358 34796
rect 91398 34756 91440 34796
rect 91112 34747 91480 34756
rect 95112 34796 95480 34805
rect 95152 34756 95194 34796
rect 95234 34756 95276 34796
rect 95316 34756 95358 34796
rect 95398 34756 95440 34796
rect 95112 34747 95480 34756
rect 99112 34796 99480 34805
rect 99152 34756 99194 34796
rect 99234 34756 99276 34796
rect 99316 34756 99358 34796
rect 99398 34756 99440 34796
rect 99112 34747 99480 34756
rect 4352 34040 4720 34049
rect 4392 34000 4434 34040
rect 4474 34000 4516 34040
rect 4556 34000 4598 34040
rect 4638 34000 4680 34040
rect 4352 33991 4720 34000
rect 8352 34040 8720 34049
rect 8392 34000 8434 34040
rect 8474 34000 8516 34040
rect 8556 34000 8598 34040
rect 8638 34000 8680 34040
rect 8352 33991 8720 34000
rect 12352 34040 12720 34049
rect 12392 34000 12434 34040
rect 12474 34000 12516 34040
rect 12556 34000 12598 34040
rect 12638 34000 12680 34040
rect 12352 33991 12720 34000
rect 16352 34040 16720 34049
rect 16392 34000 16434 34040
rect 16474 34000 16516 34040
rect 16556 34000 16598 34040
rect 16638 34000 16680 34040
rect 16352 33991 16720 34000
rect 20352 34040 20720 34049
rect 20392 34000 20434 34040
rect 20474 34000 20516 34040
rect 20556 34000 20598 34040
rect 20638 34000 20680 34040
rect 20352 33991 20720 34000
rect 24352 34040 24720 34049
rect 24392 34000 24434 34040
rect 24474 34000 24516 34040
rect 24556 34000 24598 34040
rect 24638 34000 24680 34040
rect 24352 33991 24720 34000
rect 28352 34040 28720 34049
rect 28392 34000 28434 34040
rect 28474 34000 28516 34040
rect 28556 34000 28598 34040
rect 28638 34000 28680 34040
rect 28352 33991 28720 34000
rect 32352 34040 32720 34049
rect 32392 34000 32434 34040
rect 32474 34000 32516 34040
rect 32556 34000 32598 34040
rect 32638 34000 32680 34040
rect 32352 33991 32720 34000
rect 36352 34040 36720 34049
rect 36392 34000 36434 34040
rect 36474 34000 36516 34040
rect 36556 34000 36598 34040
rect 36638 34000 36680 34040
rect 36352 33991 36720 34000
rect 40352 34040 40720 34049
rect 40392 34000 40434 34040
rect 40474 34000 40516 34040
rect 40556 34000 40598 34040
rect 40638 34000 40680 34040
rect 40352 33991 40720 34000
rect 44352 34040 44720 34049
rect 44392 34000 44434 34040
rect 44474 34000 44516 34040
rect 44556 34000 44598 34040
rect 44638 34000 44680 34040
rect 44352 33991 44720 34000
rect 48352 34040 48720 34049
rect 48392 34000 48434 34040
rect 48474 34000 48516 34040
rect 48556 34000 48598 34040
rect 48638 34000 48680 34040
rect 48352 33991 48720 34000
rect 52352 34040 52720 34049
rect 52392 34000 52434 34040
rect 52474 34000 52516 34040
rect 52556 34000 52598 34040
rect 52638 34000 52680 34040
rect 52352 33991 52720 34000
rect 56352 34040 56720 34049
rect 56392 34000 56434 34040
rect 56474 34000 56516 34040
rect 56556 34000 56598 34040
rect 56638 34000 56680 34040
rect 56352 33991 56720 34000
rect 60352 34040 60720 34049
rect 60392 34000 60434 34040
rect 60474 34000 60516 34040
rect 60556 34000 60598 34040
rect 60638 34000 60680 34040
rect 60352 33991 60720 34000
rect 64352 34040 64720 34049
rect 64392 34000 64434 34040
rect 64474 34000 64516 34040
rect 64556 34000 64598 34040
rect 64638 34000 64680 34040
rect 64352 33991 64720 34000
rect 68352 34040 68720 34049
rect 68392 34000 68434 34040
rect 68474 34000 68516 34040
rect 68556 34000 68598 34040
rect 68638 34000 68680 34040
rect 68352 33991 68720 34000
rect 87051 33452 87093 33461
rect 87051 33412 87052 33452
rect 87092 33412 87093 33452
rect 87051 33403 87093 33412
rect 87052 33318 87092 33403
rect 3112 33284 3480 33293
rect 3152 33244 3194 33284
rect 3234 33244 3276 33284
rect 3316 33244 3358 33284
rect 3398 33244 3440 33284
rect 3112 33235 3480 33244
rect 7112 33284 7480 33293
rect 7152 33244 7194 33284
rect 7234 33244 7276 33284
rect 7316 33244 7358 33284
rect 7398 33244 7440 33284
rect 7112 33235 7480 33244
rect 11112 33284 11480 33293
rect 11152 33244 11194 33284
rect 11234 33244 11276 33284
rect 11316 33244 11358 33284
rect 11398 33244 11440 33284
rect 11112 33235 11480 33244
rect 15112 33284 15480 33293
rect 15152 33244 15194 33284
rect 15234 33244 15276 33284
rect 15316 33244 15358 33284
rect 15398 33244 15440 33284
rect 15112 33235 15480 33244
rect 19112 33284 19480 33293
rect 19152 33244 19194 33284
rect 19234 33244 19276 33284
rect 19316 33244 19358 33284
rect 19398 33244 19440 33284
rect 19112 33235 19480 33244
rect 23112 33284 23480 33293
rect 23152 33244 23194 33284
rect 23234 33244 23276 33284
rect 23316 33244 23358 33284
rect 23398 33244 23440 33284
rect 23112 33235 23480 33244
rect 27112 33284 27480 33293
rect 27152 33244 27194 33284
rect 27234 33244 27276 33284
rect 27316 33244 27358 33284
rect 27398 33244 27440 33284
rect 27112 33235 27480 33244
rect 31112 33284 31480 33293
rect 31152 33244 31194 33284
rect 31234 33244 31276 33284
rect 31316 33244 31358 33284
rect 31398 33244 31440 33284
rect 31112 33235 31480 33244
rect 35112 33284 35480 33293
rect 35152 33244 35194 33284
rect 35234 33244 35276 33284
rect 35316 33244 35358 33284
rect 35398 33244 35440 33284
rect 35112 33235 35480 33244
rect 39112 33284 39480 33293
rect 39152 33244 39194 33284
rect 39234 33244 39276 33284
rect 39316 33244 39358 33284
rect 39398 33244 39440 33284
rect 39112 33235 39480 33244
rect 43112 33284 43480 33293
rect 43152 33244 43194 33284
rect 43234 33244 43276 33284
rect 43316 33244 43358 33284
rect 43398 33244 43440 33284
rect 43112 33235 43480 33244
rect 47112 33284 47480 33293
rect 47152 33244 47194 33284
rect 47234 33244 47276 33284
rect 47316 33244 47358 33284
rect 47398 33244 47440 33284
rect 47112 33235 47480 33244
rect 51112 33284 51480 33293
rect 51152 33244 51194 33284
rect 51234 33244 51276 33284
rect 51316 33244 51358 33284
rect 51398 33244 51440 33284
rect 51112 33235 51480 33244
rect 55112 33284 55480 33293
rect 55152 33244 55194 33284
rect 55234 33244 55276 33284
rect 55316 33244 55358 33284
rect 55398 33244 55440 33284
rect 55112 33235 55480 33244
rect 59112 33284 59480 33293
rect 59152 33244 59194 33284
rect 59234 33244 59276 33284
rect 59316 33244 59358 33284
rect 59398 33244 59440 33284
rect 59112 33235 59480 33244
rect 63112 33284 63480 33293
rect 63152 33244 63194 33284
rect 63234 33244 63276 33284
rect 63316 33244 63358 33284
rect 63398 33244 63440 33284
rect 63112 33235 63480 33244
rect 67112 33284 67480 33293
rect 67152 33244 67194 33284
rect 67234 33244 67276 33284
rect 67316 33244 67358 33284
rect 67398 33244 67440 33284
rect 67112 33235 67480 33244
rect 73612 32873 73652 32958
rect 73611 32864 73653 32873
rect 73611 32824 73612 32864
rect 73652 32824 73653 32864
rect 73611 32815 73653 32824
rect 4352 32528 4720 32537
rect 4392 32488 4434 32528
rect 4474 32488 4516 32528
rect 4556 32488 4598 32528
rect 4638 32488 4680 32528
rect 4352 32479 4720 32488
rect 8352 32528 8720 32537
rect 8392 32488 8434 32528
rect 8474 32488 8516 32528
rect 8556 32488 8598 32528
rect 8638 32488 8680 32528
rect 8352 32479 8720 32488
rect 12352 32528 12720 32537
rect 12392 32488 12434 32528
rect 12474 32488 12516 32528
rect 12556 32488 12598 32528
rect 12638 32488 12680 32528
rect 12352 32479 12720 32488
rect 16352 32528 16720 32537
rect 16392 32488 16434 32528
rect 16474 32488 16516 32528
rect 16556 32488 16598 32528
rect 16638 32488 16680 32528
rect 16352 32479 16720 32488
rect 20352 32528 20720 32537
rect 20392 32488 20434 32528
rect 20474 32488 20516 32528
rect 20556 32488 20598 32528
rect 20638 32488 20680 32528
rect 20352 32479 20720 32488
rect 24352 32528 24720 32537
rect 24392 32488 24434 32528
rect 24474 32488 24516 32528
rect 24556 32488 24598 32528
rect 24638 32488 24680 32528
rect 24352 32479 24720 32488
rect 28352 32528 28720 32537
rect 28392 32488 28434 32528
rect 28474 32488 28516 32528
rect 28556 32488 28598 32528
rect 28638 32488 28680 32528
rect 28352 32479 28720 32488
rect 32352 32528 32720 32537
rect 32392 32488 32434 32528
rect 32474 32488 32516 32528
rect 32556 32488 32598 32528
rect 32638 32488 32680 32528
rect 32352 32479 32720 32488
rect 36352 32528 36720 32537
rect 36392 32488 36434 32528
rect 36474 32488 36516 32528
rect 36556 32488 36598 32528
rect 36638 32488 36680 32528
rect 36352 32479 36720 32488
rect 40352 32528 40720 32537
rect 40392 32488 40434 32528
rect 40474 32488 40516 32528
rect 40556 32488 40598 32528
rect 40638 32488 40680 32528
rect 40352 32479 40720 32488
rect 44352 32528 44720 32537
rect 44392 32488 44434 32528
rect 44474 32488 44516 32528
rect 44556 32488 44598 32528
rect 44638 32488 44680 32528
rect 44352 32479 44720 32488
rect 48352 32528 48720 32537
rect 48392 32488 48434 32528
rect 48474 32488 48516 32528
rect 48556 32488 48598 32528
rect 48638 32488 48680 32528
rect 48352 32479 48720 32488
rect 52352 32528 52720 32537
rect 52392 32488 52434 32528
rect 52474 32488 52516 32528
rect 52556 32488 52598 32528
rect 52638 32488 52680 32528
rect 52352 32479 52720 32488
rect 56352 32528 56720 32537
rect 56392 32488 56434 32528
rect 56474 32488 56516 32528
rect 56556 32488 56598 32528
rect 56638 32488 56680 32528
rect 56352 32479 56720 32488
rect 60352 32528 60720 32537
rect 60392 32488 60434 32528
rect 60474 32488 60516 32528
rect 60556 32488 60598 32528
rect 60638 32488 60680 32528
rect 60352 32479 60720 32488
rect 64352 32528 64720 32537
rect 64392 32488 64434 32528
rect 64474 32488 64516 32528
rect 64556 32488 64598 32528
rect 64638 32488 64680 32528
rect 64352 32479 64720 32488
rect 68352 32528 68720 32537
rect 68392 32488 68434 32528
rect 68474 32488 68516 32528
rect 68556 32488 68598 32528
rect 68638 32488 68680 32528
rect 68352 32479 68720 32488
rect 3112 31772 3480 31781
rect 3152 31732 3194 31772
rect 3234 31732 3276 31772
rect 3316 31732 3358 31772
rect 3398 31732 3440 31772
rect 3112 31723 3480 31732
rect 7112 31772 7480 31781
rect 7152 31732 7194 31772
rect 7234 31732 7276 31772
rect 7316 31732 7358 31772
rect 7398 31732 7440 31772
rect 7112 31723 7480 31732
rect 11112 31772 11480 31781
rect 11152 31732 11194 31772
rect 11234 31732 11276 31772
rect 11316 31732 11358 31772
rect 11398 31732 11440 31772
rect 11112 31723 11480 31732
rect 15112 31772 15480 31781
rect 15152 31732 15194 31772
rect 15234 31732 15276 31772
rect 15316 31732 15358 31772
rect 15398 31732 15440 31772
rect 15112 31723 15480 31732
rect 19112 31772 19480 31781
rect 19152 31732 19194 31772
rect 19234 31732 19276 31772
rect 19316 31732 19358 31772
rect 19398 31732 19440 31772
rect 19112 31723 19480 31732
rect 23112 31772 23480 31781
rect 23152 31732 23194 31772
rect 23234 31732 23276 31772
rect 23316 31732 23358 31772
rect 23398 31732 23440 31772
rect 23112 31723 23480 31732
rect 27112 31772 27480 31781
rect 27152 31732 27194 31772
rect 27234 31732 27276 31772
rect 27316 31732 27358 31772
rect 27398 31732 27440 31772
rect 27112 31723 27480 31732
rect 31112 31772 31480 31781
rect 31152 31732 31194 31772
rect 31234 31732 31276 31772
rect 31316 31732 31358 31772
rect 31398 31732 31440 31772
rect 31112 31723 31480 31732
rect 35112 31772 35480 31781
rect 35152 31732 35194 31772
rect 35234 31732 35276 31772
rect 35316 31732 35358 31772
rect 35398 31732 35440 31772
rect 35112 31723 35480 31732
rect 39112 31772 39480 31781
rect 39152 31732 39194 31772
rect 39234 31732 39276 31772
rect 39316 31732 39358 31772
rect 39398 31732 39440 31772
rect 39112 31723 39480 31732
rect 43112 31772 43480 31781
rect 43152 31732 43194 31772
rect 43234 31732 43276 31772
rect 43316 31732 43358 31772
rect 43398 31732 43440 31772
rect 43112 31723 43480 31732
rect 47112 31772 47480 31781
rect 47152 31732 47194 31772
rect 47234 31732 47276 31772
rect 47316 31732 47358 31772
rect 47398 31732 47440 31772
rect 47112 31723 47480 31732
rect 51112 31772 51480 31781
rect 51152 31732 51194 31772
rect 51234 31732 51276 31772
rect 51316 31732 51358 31772
rect 51398 31732 51440 31772
rect 51112 31723 51480 31732
rect 55112 31772 55480 31781
rect 55152 31732 55194 31772
rect 55234 31732 55276 31772
rect 55316 31732 55358 31772
rect 55398 31732 55440 31772
rect 55112 31723 55480 31732
rect 59112 31772 59480 31781
rect 59152 31732 59194 31772
rect 59234 31732 59276 31772
rect 59316 31732 59358 31772
rect 59398 31732 59440 31772
rect 59112 31723 59480 31732
rect 63112 31772 63480 31781
rect 63152 31732 63194 31772
rect 63234 31732 63276 31772
rect 63316 31732 63358 31772
rect 63398 31732 63440 31772
rect 63112 31723 63480 31732
rect 67112 31772 67480 31781
rect 67152 31732 67194 31772
rect 67234 31732 67276 31772
rect 67316 31732 67358 31772
rect 67398 31732 67440 31772
rect 67112 31723 67480 31732
rect 4352 31016 4720 31025
rect 4392 30976 4434 31016
rect 4474 30976 4516 31016
rect 4556 30976 4598 31016
rect 4638 30976 4680 31016
rect 4352 30967 4720 30976
rect 8352 31016 8720 31025
rect 8392 30976 8434 31016
rect 8474 30976 8516 31016
rect 8556 30976 8598 31016
rect 8638 30976 8680 31016
rect 8352 30967 8720 30976
rect 12352 31016 12720 31025
rect 12392 30976 12434 31016
rect 12474 30976 12516 31016
rect 12556 30976 12598 31016
rect 12638 30976 12680 31016
rect 12352 30967 12720 30976
rect 16352 31016 16720 31025
rect 16392 30976 16434 31016
rect 16474 30976 16516 31016
rect 16556 30976 16598 31016
rect 16638 30976 16680 31016
rect 16352 30967 16720 30976
rect 20352 31016 20720 31025
rect 20392 30976 20434 31016
rect 20474 30976 20516 31016
rect 20556 30976 20598 31016
rect 20638 30976 20680 31016
rect 20352 30967 20720 30976
rect 24352 31016 24720 31025
rect 24392 30976 24434 31016
rect 24474 30976 24516 31016
rect 24556 30976 24598 31016
rect 24638 30976 24680 31016
rect 24352 30967 24720 30976
rect 28352 31016 28720 31025
rect 28392 30976 28434 31016
rect 28474 30976 28516 31016
rect 28556 30976 28598 31016
rect 28638 30976 28680 31016
rect 28352 30967 28720 30976
rect 32352 31016 32720 31025
rect 32392 30976 32434 31016
rect 32474 30976 32516 31016
rect 32556 30976 32598 31016
rect 32638 30976 32680 31016
rect 32352 30967 32720 30976
rect 36352 31016 36720 31025
rect 36392 30976 36434 31016
rect 36474 30976 36516 31016
rect 36556 30976 36598 31016
rect 36638 30976 36680 31016
rect 36352 30967 36720 30976
rect 40352 31016 40720 31025
rect 40392 30976 40434 31016
rect 40474 30976 40516 31016
rect 40556 30976 40598 31016
rect 40638 30976 40680 31016
rect 40352 30967 40720 30976
rect 44352 31016 44720 31025
rect 44392 30976 44434 31016
rect 44474 30976 44516 31016
rect 44556 30976 44598 31016
rect 44638 30976 44680 31016
rect 44352 30967 44720 30976
rect 48352 31016 48720 31025
rect 48392 30976 48434 31016
rect 48474 30976 48516 31016
rect 48556 30976 48598 31016
rect 48638 30976 48680 31016
rect 48352 30967 48720 30976
rect 52352 31016 52720 31025
rect 52392 30976 52434 31016
rect 52474 30976 52516 31016
rect 52556 30976 52598 31016
rect 52638 30976 52680 31016
rect 52352 30967 52720 30976
rect 56352 31016 56720 31025
rect 56392 30976 56434 31016
rect 56474 30976 56516 31016
rect 56556 30976 56598 31016
rect 56638 30976 56680 31016
rect 56352 30967 56720 30976
rect 60352 31016 60720 31025
rect 60392 30976 60434 31016
rect 60474 30976 60516 31016
rect 60556 30976 60598 31016
rect 60638 30976 60680 31016
rect 60352 30967 60720 30976
rect 64352 31016 64720 31025
rect 64392 30976 64434 31016
rect 64474 30976 64516 31016
rect 64556 30976 64598 31016
rect 64638 30976 64680 31016
rect 64352 30967 64720 30976
rect 68352 31016 68720 31025
rect 68392 30976 68434 31016
rect 68474 30976 68516 31016
rect 68556 30976 68598 31016
rect 68638 30976 68680 31016
rect 68352 30967 68720 30976
rect 3112 30260 3480 30269
rect 3152 30220 3194 30260
rect 3234 30220 3276 30260
rect 3316 30220 3358 30260
rect 3398 30220 3440 30260
rect 3112 30211 3480 30220
rect 7112 30260 7480 30269
rect 7152 30220 7194 30260
rect 7234 30220 7276 30260
rect 7316 30220 7358 30260
rect 7398 30220 7440 30260
rect 7112 30211 7480 30220
rect 11112 30260 11480 30269
rect 11152 30220 11194 30260
rect 11234 30220 11276 30260
rect 11316 30220 11358 30260
rect 11398 30220 11440 30260
rect 11112 30211 11480 30220
rect 15112 30260 15480 30269
rect 15152 30220 15194 30260
rect 15234 30220 15276 30260
rect 15316 30220 15358 30260
rect 15398 30220 15440 30260
rect 15112 30211 15480 30220
rect 19112 30260 19480 30269
rect 19152 30220 19194 30260
rect 19234 30220 19276 30260
rect 19316 30220 19358 30260
rect 19398 30220 19440 30260
rect 19112 30211 19480 30220
rect 23112 30260 23480 30269
rect 23152 30220 23194 30260
rect 23234 30220 23276 30260
rect 23316 30220 23358 30260
rect 23398 30220 23440 30260
rect 23112 30211 23480 30220
rect 27112 30260 27480 30269
rect 27152 30220 27194 30260
rect 27234 30220 27276 30260
rect 27316 30220 27358 30260
rect 27398 30220 27440 30260
rect 27112 30211 27480 30220
rect 31112 30260 31480 30269
rect 31152 30220 31194 30260
rect 31234 30220 31276 30260
rect 31316 30220 31358 30260
rect 31398 30220 31440 30260
rect 31112 30211 31480 30220
rect 35112 30260 35480 30269
rect 35152 30220 35194 30260
rect 35234 30220 35276 30260
rect 35316 30220 35358 30260
rect 35398 30220 35440 30260
rect 35112 30211 35480 30220
rect 39112 30260 39480 30269
rect 39152 30220 39194 30260
rect 39234 30220 39276 30260
rect 39316 30220 39358 30260
rect 39398 30220 39440 30260
rect 39112 30211 39480 30220
rect 43112 30260 43480 30269
rect 43152 30220 43194 30260
rect 43234 30220 43276 30260
rect 43316 30220 43358 30260
rect 43398 30220 43440 30260
rect 43112 30211 43480 30220
rect 47112 30260 47480 30269
rect 47152 30220 47194 30260
rect 47234 30220 47276 30260
rect 47316 30220 47358 30260
rect 47398 30220 47440 30260
rect 47112 30211 47480 30220
rect 51112 30260 51480 30269
rect 51152 30220 51194 30260
rect 51234 30220 51276 30260
rect 51316 30220 51358 30260
rect 51398 30220 51440 30260
rect 51112 30211 51480 30220
rect 55112 30260 55480 30269
rect 55152 30220 55194 30260
rect 55234 30220 55276 30260
rect 55316 30220 55358 30260
rect 55398 30220 55440 30260
rect 55112 30211 55480 30220
rect 59112 30260 59480 30269
rect 59152 30220 59194 30260
rect 59234 30220 59276 30260
rect 59316 30220 59358 30260
rect 59398 30220 59440 30260
rect 59112 30211 59480 30220
rect 63112 30260 63480 30269
rect 63152 30220 63194 30260
rect 63234 30220 63276 30260
rect 63316 30220 63358 30260
rect 63398 30220 63440 30260
rect 63112 30211 63480 30220
rect 67112 30260 67480 30269
rect 67152 30220 67194 30260
rect 67234 30220 67276 30260
rect 67316 30220 67358 30260
rect 67398 30220 67440 30260
rect 67112 30211 67480 30220
rect 4352 29504 4720 29513
rect 4392 29464 4434 29504
rect 4474 29464 4516 29504
rect 4556 29464 4598 29504
rect 4638 29464 4680 29504
rect 4352 29455 4720 29464
rect 8352 29504 8720 29513
rect 8392 29464 8434 29504
rect 8474 29464 8516 29504
rect 8556 29464 8598 29504
rect 8638 29464 8680 29504
rect 8352 29455 8720 29464
rect 12352 29504 12720 29513
rect 12392 29464 12434 29504
rect 12474 29464 12516 29504
rect 12556 29464 12598 29504
rect 12638 29464 12680 29504
rect 12352 29455 12720 29464
rect 16352 29504 16720 29513
rect 16392 29464 16434 29504
rect 16474 29464 16516 29504
rect 16556 29464 16598 29504
rect 16638 29464 16680 29504
rect 16352 29455 16720 29464
rect 20352 29504 20720 29513
rect 20392 29464 20434 29504
rect 20474 29464 20516 29504
rect 20556 29464 20598 29504
rect 20638 29464 20680 29504
rect 20352 29455 20720 29464
rect 24352 29504 24720 29513
rect 24392 29464 24434 29504
rect 24474 29464 24516 29504
rect 24556 29464 24598 29504
rect 24638 29464 24680 29504
rect 24352 29455 24720 29464
rect 28352 29504 28720 29513
rect 28392 29464 28434 29504
rect 28474 29464 28516 29504
rect 28556 29464 28598 29504
rect 28638 29464 28680 29504
rect 28352 29455 28720 29464
rect 32352 29504 32720 29513
rect 32392 29464 32434 29504
rect 32474 29464 32516 29504
rect 32556 29464 32598 29504
rect 32638 29464 32680 29504
rect 32352 29455 32720 29464
rect 36352 29504 36720 29513
rect 36392 29464 36434 29504
rect 36474 29464 36516 29504
rect 36556 29464 36598 29504
rect 36638 29464 36680 29504
rect 36352 29455 36720 29464
rect 40352 29504 40720 29513
rect 40392 29464 40434 29504
rect 40474 29464 40516 29504
rect 40556 29464 40598 29504
rect 40638 29464 40680 29504
rect 40352 29455 40720 29464
rect 44352 29504 44720 29513
rect 44392 29464 44434 29504
rect 44474 29464 44516 29504
rect 44556 29464 44598 29504
rect 44638 29464 44680 29504
rect 44352 29455 44720 29464
rect 48352 29504 48720 29513
rect 48392 29464 48434 29504
rect 48474 29464 48516 29504
rect 48556 29464 48598 29504
rect 48638 29464 48680 29504
rect 48352 29455 48720 29464
rect 52352 29504 52720 29513
rect 52392 29464 52434 29504
rect 52474 29464 52516 29504
rect 52556 29464 52598 29504
rect 52638 29464 52680 29504
rect 52352 29455 52720 29464
rect 56352 29504 56720 29513
rect 56392 29464 56434 29504
rect 56474 29464 56516 29504
rect 56556 29464 56598 29504
rect 56638 29464 56680 29504
rect 56352 29455 56720 29464
rect 60352 29504 60720 29513
rect 60392 29464 60434 29504
rect 60474 29464 60516 29504
rect 60556 29464 60598 29504
rect 60638 29464 60680 29504
rect 60352 29455 60720 29464
rect 64352 29504 64720 29513
rect 64392 29464 64434 29504
rect 64474 29464 64516 29504
rect 64556 29464 64598 29504
rect 64638 29464 64680 29504
rect 64352 29455 64720 29464
rect 68352 29504 68720 29513
rect 68392 29464 68434 29504
rect 68474 29464 68516 29504
rect 68556 29464 68598 29504
rect 68638 29464 68680 29504
rect 68352 29455 68720 29464
rect 3112 28748 3480 28757
rect 3152 28708 3194 28748
rect 3234 28708 3276 28748
rect 3316 28708 3358 28748
rect 3398 28708 3440 28748
rect 3112 28699 3480 28708
rect 7112 28748 7480 28757
rect 7152 28708 7194 28748
rect 7234 28708 7276 28748
rect 7316 28708 7358 28748
rect 7398 28708 7440 28748
rect 7112 28699 7480 28708
rect 11112 28748 11480 28757
rect 11152 28708 11194 28748
rect 11234 28708 11276 28748
rect 11316 28708 11358 28748
rect 11398 28708 11440 28748
rect 11112 28699 11480 28708
rect 15112 28748 15480 28757
rect 15152 28708 15194 28748
rect 15234 28708 15276 28748
rect 15316 28708 15358 28748
rect 15398 28708 15440 28748
rect 15112 28699 15480 28708
rect 19112 28748 19480 28757
rect 19152 28708 19194 28748
rect 19234 28708 19276 28748
rect 19316 28708 19358 28748
rect 19398 28708 19440 28748
rect 19112 28699 19480 28708
rect 23112 28748 23480 28757
rect 23152 28708 23194 28748
rect 23234 28708 23276 28748
rect 23316 28708 23358 28748
rect 23398 28708 23440 28748
rect 23112 28699 23480 28708
rect 27112 28748 27480 28757
rect 27152 28708 27194 28748
rect 27234 28708 27276 28748
rect 27316 28708 27358 28748
rect 27398 28708 27440 28748
rect 27112 28699 27480 28708
rect 31112 28748 31480 28757
rect 31152 28708 31194 28748
rect 31234 28708 31276 28748
rect 31316 28708 31358 28748
rect 31398 28708 31440 28748
rect 31112 28699 31480 28708
rect 35112 28748 35480 28757
rect 35152 28708 35194 28748
rect 35234 28708 35276 28748
rect 35316 28708 35358 28748
rect 35398 28708 35440 28748
rect 35112 28699 35480 28708
rect 39112 28748 39480 28757
rect 39152 28708 39194 28748
rect 39234 28708 39276 28748
rect 39316 28708 39358 28748
rect 39398 28708 39440 28748
rect 39112 28699 39480 28708
rect 43112 28748 43480 28757
rect 43152 28708 43194 28748
rect 43234 28708 43276 28748
rect 43316 28708 43358 28748
rect 43398 28708 43440 28748
rect 43112 28699 43480 28708
rect 47112 28748 47480 28757
rect 47152 28708 47194 28748
rect 47234 28708 47276 28748
rect 47316 28708 47358 28748
rect 47398 28708 47440 28748
rect 47112 28699 47480 28708
rect 51112 28748 51480 28757
rect 51152 28708 51194 28748
rect 51234 28708 51276 28748
rect 51316 28708 51358 28748
rect 51398 28708 51440 28748
rect 51112 28699 51480 28708
rect 55112 28748 55480 28757
rect 55152 28708 55194 28748
rect 55234 28708 55276 28748
rect 55316 28708 55358 28748
rect 55398 28708 55440 28748
rect 55112 28699 55480 28708
rect 59112 28748 59480 28757
rect 59152 28708 59194 28748
rect 59234 28708 59276 28748
rect 59316 28708 59358 28748
rect 59398 28708 59440 28748
rect 59112 28699 59480 28708
rect 63112 28748 63480 28757
rect 63152 28708 63194 28748
rect 63234 28708 63276 28748
rect 63316 28708 63358 28748
rect 63398 28708 63440 28748
rect 63112 28699 63480 28708
rect 67112 28748 67480 28757
rect 67152 28708 67194 28748
rect 67234 28708 67276 28748
rect 67316 28708 67358 28748
rect 67398 28708 67440 28748
rect 67112 28699 67480 28708
rect 4352 27992 4720 28001
rect 4392 27952 4434 27992
rect 4474 27952 4516 27992
rect 4556 27952 4598 27992
rect 4638 27952 4680 27992
rect 4352 27943 4720 27952
rect 8352 27992 8720 28001
rect 8392 27952 8434 27992
rect 8474 27952 8516 27992
rect 8556 27952 8598 27992
rect 8638 27952 8680 27992
rect 8352 27943 8720 27952
rect 12352 27992 12720 28001
rect 12392 27952 12434 27992
rect 12474 27952 12516 27992
rect 12556 27952 12598 27992
rect 12638 27952 12680 27992
rect 12352 27943 12720 27952
rect 16352 27992 16720 28001
rect 16392 27952 16434 27992
rect 16474 27952 16516 27992
rect 16556 27952 16598 27992
rect 16638 27952 16680 27992
rect 16352 27943 16720 27952
rect 20352 27992 20720 28001
rect 20392 27952 20434 27992
rect 20474 27952 20516 27992
rect 20556 27952 20598 27992
rect 20638 27952 20680 27992
rect 20352 27943 20720 27952
rect 24352 27992 24720 28001
rect 24392 27952 24434 27992
rect 24474 27952 24516 27992
rect 24556 27952 24598 27992
rect 24638 27952 24680 27992
rect 24352 27943 24720 27952
rect 28352 27992 28720 28001
rect 28392 27952 28434 27992
rect 28474 27952 28516 27992
rect 28556 27952 28598 27992
rect 28638 27952 28680 27992
rect 28352 27943 28720 27952
rect 32352 27992 32720 28001
rect 32392 27952 32434 27992
rect 32474 27952 32516 27992
rect 32556 27952 32598 27992
rect 32638 27952 32680 27992
rect 32352 27943 32720 27952
rect 36352 27992 36720 28001
rect 36392 27952 36434 27992
rect 36474 27952 36516 27992
rect 36556 27952 36598 27992
rect 36638 27952 36680 27992
rect 36352 27943 36720 27952
rect 40352 27992 40720 28001
rect 40392 27952 40434 27992
rect 40474 27952 40516 27992
rect 40556 27952 40598 27992
rect 40638 27952 40680 27992
rect 40352 27943 40720 27952
rect 44352 27992 44720 28001
rect 44392 27952 44434 27992
rect 44474 27952 44516 27992
rect 44556 27952 44598 27992
rect 44638 27952 44680 27992
rect 44352 27943 44720 27952
rect 48352 27992 48720 28001
rect 48392 27952 48434 27992
rect 48474 27952 48516 27992
rect 48556 27952 48598 27992
rect 48638 27952 48680 27992
rect 48352 27943 48720 27952
rect 52352 27992 52720 28001
rect 52392 27952 52434 27992
rect 52474 27952 52516 27992
rect 52556 27952 52598 27992
rect 52638 27952 52680 27992
rect 52352 27943 52720 27952
rect 56352 27992 56720 28001
rect 56392 27952 56434 27992
rect 56474 27952 56516 27992
rect 56556 27952 56598 27992
rect 56638 27952 56680 27992
rect 56352 27943 56720 27952
rect 60352 27992 60720 28001
rect 60392 27952 60434 27992
rect 60474 27952 60516 27992
rect 60556 27952 60598 27992
rect 60638 27952 60680 27992
rect 60352 27943 60720 27952
rect 64352 27992 64720 28001
rect 64392 27952 64434 27992
rect 64474 27952 64516 27992
rect 64556 27952 64598 27992
rect 64638 27952 64680 27992
rect 64352 27943 64720 27952
rect 68352 27992 68720 28001
rect 68392 27952 68434 27992
rect 68474 27952 68516 27992
rect 68556 27952 68598 27992
rect 68638 27952 68680 27992
rect 68352 27943 68720 27952
rect 3112 27236 3480 27245
rect 3152 27196 3194 27236
rect 3234 27196 3276 27236
rect 3316 27196 3358 27236
rect 3398 27196 3440 27236
rect 3112 27187 3480 27196
rect 7112 27236 7480 27245
rect 7152 27196 7194 27236
rect 7234 27196 7276 27236
rect 7316 27196 7358 27236
rect 7398 27196 7440 27236
rect 7112 27187 7480 27196
rect 11112 27236 11480 27245
rect 11152 27196 11194 27236
rect 11234 27196 11276 27236
rect 11316 27196 11358 27236
rect 11398 27196 11440 27236
rect 11112 27187 11480 27196
rect 15112 27236 15480 27245
rect 15152 27196 15194 27236
rect 15234 27196 15276 27236
rect 15316 27196 15358 27236
rect 15398 27196 15440 27236
rect 15112 27187 15480 27196
rect 19112 27236 19480 27245
rect 19152 27196 19194 27236
rect 19234 27196 19276 27236
rect 19316 27196 19358 27236
rect 19398 27196 19440 27236
rect 19112 27187 19480 27196
rect 23112 27236 23480 27245
rect 23152 27196 23194 27236
rect 23234 27196 23276 27236
rect 23316 27196 23358 27236
rect 23398 27196 23440 27236
rect 23112 27187 23480 27196
rect 27112 27236 27480 27245
rect 27152 27196 27194 27236
rect 27234 27196 27276 27236
rect 27316 27196 27358 27236
rect 27398 27196 27440 27236
rect 27112 27187 27480 27196
rect 31112 27236 31480 27245
rect 31152 27196 31194 27236
rect 31234 27196 31276 27236
rect 31316 27196 31358 27236
rect 31398 27196 31440 27236
rect 31112 27187 31480 27196
rect 35112 27236 35480 27245
rect 35152 27196 35194 27236
rect 35234 27196 35276 27236
rect 35316 27196 35358 27236
rect 35398 27196 35440 27236
rect 35112 27187 35480 27196
rect 39112 27236 39480 27245
rect 39152 27196 39194 27236
rect 39234 27196 39276 27236
rect 39316 27196 39358 27236
rect 39398 27196 39440 27236
rect 39112 27187 39480 27196
rect 43112 27236 43480 27245
rect 43152 27196 43194 27236
rect 43234 27196 43276 27236
rect 43316 27196 43358 27236
rect 43398 27196 43440 27236
rect 43112 27187 43480 27196
rect 47112 27236 47480 27245
rect 47152 27196 47194 27236
rect 47234 27196 47276 27236
rect 47316 27196 47358 27236
rect 47398 27196 47440 27236
rect 47112 27187 47480 27196
rect 51112 27236 51480 27245
rect 51152 27196 51194 27236
rect 51234 27196 51276 27236
rect 51316 27196 51358 27236
rect 51398 27196 51440 27236
rect 51112 27187 51480 27196
rect 55112 27236 55480 27245
rect 55152 27196 55194 27236
rect 55234 27196 55276 27236
rect 55316 27196 55358 27236
rect 55398 27196 55440 27236
rect 55112 27187 55480 27196
rect 59112 27236 59480 27245
rect 59152 27196 59194 27236
rect 59234 27196 59276 27236
rect 59316 27196 59358 27236
rect 59398 27196 59440 27236
rect 59112 27187 59480 27196
rect 63112 27236 63480 27245
rect 63152 27196 63194 27236
rect 63234 27196 63276 27236
rect 63316 27196 63358 27236
rect 63398 27196 63440 27236
rect 63112 27187 63480 27196
rect 67112 27236 67480 27245
rect 67152 27196 67194 27236
rect 67234 27196 67276 27236
rect 67316 27196 67358 27236
rect 67398 27196 67440 27236
rect 67112 27187 67480 27196
rect 71884 26816 71924 26825
rect 71884 26573 71924 26776
rect 71883 26564 71925 26573
rect 71883 26524 71884 26564
rect 71924 26524 71925 26564
rect 71883 26515 71925 26524
rect 73227 26564 73269 26573
rect 73227 26524 73228 26564
rect 73268 26524 73269 26564
rect 73227 26515 73269 26524
rect 4352 26480 4720 26489
rect 4392 26440 4434 26480
rect 4474 26440 4516 26480
rect 4556 26440 4598 26480
rect 4638 26440 4680 26480
rect 4352 26431 4720 26440
rect 8352 26480 8720 26489
rect 8392 26440 8434 26480
rect 8474 26440 8516 26480
rect 8556 26440 8598 26480
rect 8638 26440 8680 26480
rect 8352 26431 8720 26440
rect 12352 26480 12720 26489
rect 12392 26440 12434 26480
rect 12474 26440 12516 26480
rect 12556 26440 12598 26480
rect 12638 26440 12680 26480
rect 12352 26431 12720 26440
rect 16352 26480 16720 26489
rect 16392 26440 16434 26480
rect 16474 26440 16516 26480
rect 16556 26440 16598 26480
rect 16638 26440 16680 26480
rect 16352 26431 16720 26440
rect 20352 26480 20720 26489
rect 20392 26440 20434 26480
rect 20474 26440 20516 26480
rect 20556 26440 20598 26480
rect 20638 26440 20680 26480
rect 20352 26431 20720 26440
rect 24352 26480 24720 26489
rect 24392 26440 24434 26480
rect 24474 26440 24516 26480
rect 24556 26440 24598 26480
rect 24638 26440 24680 26480
rect 24352 26431 24720 26440
rect 28352 26480 28720 26489
rect 28392 26440 28434 26480
rect 28474 26440 28516 26480
rect 28556 26440 28598 26480
rect 28638 26440 28680 26480
rect 28352 26431 28720 26440
rect 32352 26480 32720 26489
rect 32392 26440 32434 26480
rect 32474 26440 32516 26480
rect 32556 26440 32598 26480
rect 32638 26440 32680 26480
rect 32352 26431 32720 26440
rect 36352 26480 36720 26489
rect 36392 26440 36434 26480
rect 36474 26440 36516 26480
rect 36556 26440 36598 26480
rect 36638 26440 36680 26480
rect 36352 26431 36720 26440
rect 40352 26480 40720 26489
rect 40392 26440 40434 26480
rect 40474 26440 40516 26480
rect 40556 26440 40598 26480
rect 40638 26440 40680 26480
rect 40352 26431 40720 26440
rect 44352 26480 44720 26489
rect 44392 26440 44434 26480
rect 44474 26440 44516 26480
rect 44556 26440 44598 26480
rect 44638 26440 44680 26480
rect 44352 26431 44720 26440
rect 48352 26480 48720 26489
rect 48392 26440 48434 26480
rect 48474 26440 48516 26480
rect 48556 26440 48598 26480
rect 48638 26440 48680 26480
rect 48352 26431 48720 26440
rect 52352 26480 52720 26489
rect 52392 26440 52434 26480
rect 52474 26440 52516 26480
rect 52556 26440 52598 26480
rect 52638 26440 52680 26480
rect 52352 26431 52720 26440
rect 56352 26480 56720 26489
rect 56392 26440 56434 26480
rect 56474 26440 56516 26480
rect 56556 26440 56598 26480
rect 56638 26440 56680 26480
rect 56352 26431 56720 26440
rect 60352 26480 60720 26489
rect 60392 26440 60434 26480
rect 60474 26440 60516 26480
rect 60556 26440 60598 26480
rect 60638 26440 60680 26480
rect 60352 26431 60720 26440
rect 64352 26480 64720 26489
rect 64392 26440 64434 26480
rect 64474 26440 64516 26480
rect 64556 26440 64598 26480
rect 64638 26440 64680 26480
rect 64352 26431 64720 26440
rect 68352 26480 68720 26489
rect 68392 26440 68434 26480
rect 68474 26440 68516 26480
rect 68556 26440 68598 26480
rect 68638 26440 68680 26480
rect 68352 26431 68720 26440
rect 3112 25724 3480 25733
rect 3152 25684 3194 25724
rect 3234 25684 3276 25724
rect 3316 25684 3358 25724
rect 3398 25684 3440 25724
rect 3112 25675 3480 25684
rect 7112 25724 7480 25733
rect 7152 25684 7194 25724
rect 7234 25684 7276 25724
rect 7316 25684 7358 25724
rect 7398 25684 7440 25724
rect 7112 25675 7480 25684
rect 11112 25724 11480 25733
rect 11152 25684 11194 25724
rect 11234 25684 11276 25724
rect 11316 25684 11358 25724
rect 11398 25684 11440 25724
rect 11112 25675 11480 25684
rect 15112 25724 15480 25733
rect 15152 25684 15194 25724
rect 15234 25684 15276 25724
rect 15316 25684 15358 25724
rect 15398 25684 15440 25724
rect 15112 25675 15480 25684
rect 19112 25724 19480 25733
rect 19152 25684 19194 25724
rect 19234 25684 19276 25724
rect 19316 25684 19358 25724
rect 19398 25684 19440 25724
rect 19112 25675 19480 25684
rect 23112 25724 23480 25733
rect 23152 25684 23194 25724
rect 23234 25684 23276 25724
rect 23316 25684 23358 25724
rect 23398 25684 23440 25724
rect 23112 25675 23480 25684
rect 27112 25724 27480 25733
rect 27152 25684 27194 25724
rect 27234 25684 27276 25724
rect 27316 25684 27358 25724
rect 27398 25684 27440 25724
rect 27112 25675 27480 25684
rect 31112 25724 31480 25733
rect 31152 25684 31194 25724
rect 31234 25684 31276 25724
rect 31316 25684 31358 25724
rect 31398 25684 31440 25724
rect 31112 25675 31480 25684
rect 35112 25724 35480 25733
rect 35152 25684 35194 25724
rect 35234 25684 35276 25724
rect 35316 25684 35358 25724
rect 35398 25684 35440 25724
rect 35112 25675 35480 25684
rect 39112 25724 39480 25733
rect 39152 25684 39194 25724
rect 39234 25684 39276 25724
rect 39316 25684 39358 25724
rect 39398 25684 39440 25724
rect 39112 25675 39480 25684
rect 43112 25724 43480 25733
rect 43152 25684 43194 25724
rect 43234 25684 43276 25724
rect 43316 25684 43358 25724
rect 43398 25684 43440 25724
rect 43112 25675 43480 25684
rect 47112 25724 47480 25733
rect 47152 25684 47194 25724
rect 47234 25684 47276 25724
rect 47316 25684 47358 25724
rect 47398 25684 47440 25724
rect 47112 25675 47480 25684
rect 51112 25724 51480 25733
rect 51152 25684 51194 25724
rect 51234 25684 51276 25724
rect 51316 25684 51358 25724
rect 51398 25684 51440 25724
rect 51112 25675 51480 25684
rect 55112 25724 55480 25733
rect 55152 25684 55194 25724
rect 55234 25684 55276 25724
rect 55316 25684 55358 25724
rect 55398 25684 55440 25724
rect 55112 25675 55480 25684
rect 59112 25724 59480 25733
rect 59152 25684 59194 25724
rect 59234 25684 59276 25724
rect 59316 25684 59358 25724
rect 59398 25684 59440 25724
rect 59112 25675 59480 25684
rect 63112 25724 63480 25733
rect 63152 25684 63194 25724
rect 63234 25684 63276 25724
rect 63316 25684 63358 25724
rect 63398 25684 63440 25724
rect 63112 25675 63480 25684
rect 67112 25724 67480 25733
rect 67152 25684 67194 25724
rect 67234 25684 67276 25724
rect 67316 25684 67358 25724
rect 67398 25684 67440 25724
rect 67112 25675 67480 25684
rect 4352 24968 4720 24977
rect 4392 24928 4434 24968
rect 4474 24928 4516 24968
rect 4556 24928 4598 24968
rect 4638 24928 4680 24968
rect 4352 24919 4720 24928
rect 8352 24968 8720 24977
rect 8392 24928 8434 24968
rect 8474 24928 8516 24968
rect 8556 24928 8598 24968
rect 8638 24928 8680 24968
rect 8352 24919 8720 24928
rect 12352 24968 12720 24977
rect 12392 24928 12434 24968
rect 12474 24928 12516 24968
rect 12556 24928 12598 24968
rect 12638 24928 12680 24968
rect 12352 24919 12720 24928
rect 16352 24968 16720 24977
rect 16392 24928 16434 24968
rect 16474 24928 16516 24968
rect 16556 24928 16598 24968
rect 16638 24928 16680 24968
rect 16352 24919 16720 24928
rect 20352 24968 20720 24977
rect 20392 24928 20434 24968
rect 20474 24928 20516 24968
rect 20556 24928 20598 24968
rect 20638 24928 20680 24968
rect 20352 24919 20720 24928
rect 24352 24968 24720 24977
rect 24392 24928 24434 24968
rect 24474 24928 24516 24968
rect 24556 24928 24598 24968
rect 24638 24928 24680 24968
rect 24352 24919 24720 24928
rect 28352 24968 28720 24977
rect 28392 24928 28434 24968
rect 28474 24928 28516 24968
rect 28556 24928 28598 24968
rect 28638 24928 28680 24968
rect 28352 24919 28720 24928
rect 32352 24968 32720 24977
rect 32392 24928 32434 24968
rect 32474 24928 32516 24968
rect 32556 24928 32598 24968
rect 32638 24928 32680 24968
rect 32352 24919 32720 24928
rect 36352 24968 36720 24977
rect 36392 24928 36434 24968
rect 36474 24928 36516 24968
rect 36556 24928 36598 24968
rect 36638 24928 36680 24968
rect 36352 24919 36720 24928
rect 40352 24968 40720 24977
rect 40392 24928 40434 24968
rect 40474 24928 40516 24968
rect 40556 24928 40598 24968
rect 40638 24928 40680 24968
rect 40352 24919 40720 24928
rect 44352 24968 44720 24977
rect 44392 24928 44434 24968
rect 44474 24928 44516 24968
rect 44556 24928 44598 24968
rect 44638 24928 44680 24968
rect 44352 24919 44720 24928
rect 48352 24968 48720 24977
rect 48392 24928 48434 24968
rect 48474 24928 48516 24968
rect 48556 24928 48598 24968
rect 48638 24928 48680 24968
rect 48352 24919 48720 24928
rect 52352 24968 52720 24977
rect 52392 24928 52434 24968
rect 52474 24928 52516 24968
rect 52556 24928 52598 24968
rect 52638 24928 52680 24968
rect 52352 24919 52720 24928
rect 56352 24968 56720 24977
rect 56392 24928 56434 24968
rect 56474 24928 56516 24968
rect 56556 24928 56598 24968
rect 56638 24928 56680 24968
rect 56352 24919 56720 24928
rect 60352 24968 60720 24977
rect 60392 24928 60434 24968
rect 60474 24928 60516 24968
rect 60556 24928 60598 24968
rect 60638 24928 60680 24968
rect 60352 24919 60720 24928
rect 64352 24968 64720 24977
rect 64392 24928 64434 24968
rect 64474 24928 64516 24968
rect 64556 24928 64598 24968
rect 64638 24928 64680 24968
rect 64352 24919 64720 24928
rect 68352 24968 68720 24977
rect 68392 24928 68434 24968
rect 68474 24928 68516 24968
rect 68556 24928 68598 24968
rect 68638 24928 68680 24968
rect 68352 24919 68720 24928
rect 73228 24632 73268 26515
rect 85708 25724 85748 25733
rect 85708 25397 85748 25684
rect 85707 25388 85749 25397
rect 85707 25348 85708 25388
rect 85748 25348 85749 25388
rect 85707 25339 85749 25348
rect 86859 25388 86901 25397
rect 86859 25348 86860 25388
rect 86900 25348 86901 25388
rect 86859 25339 86901 25348
rect 86860 25254 86900 25339
rect 73228 24583 73268 24592
rect 3112 24212 3480 24221
rect 3152 24172 3194 24212
rect 3234 24172 3276 24212
rect 3316 24172 3358 24212
rect 3398 24172 3440 24212
rect 3112 24163 3480 24172
rect 7112 24212 7480 24221
rect 7152 24172 7194 24212
rect 7234 24172 7276 24212
rect 7316 24172 7358 24212
rect 7398 24172 7440 24212
rect 7112 24163 7480 24172
rect 11112 24212 11480 24221
rect 11152 24172 11194 24212
rect 11234 24172 11276 24212
rect 11316 24172 11358 24212
rect 11398 24172 11440 24212
rect 11112 24163 11480 24172
rect 15112 24212 15480 24221
rect 15152 24172 15194 24212
rect 15234 24172 15276 24212
rect 15316 24172 15358 24212
rect 15398 24172 15440 24212
rect 15112 24163 15480 24172
rect 19112 24212 19480 24221
rect 19152 24172 19194 24212
rect 19234 24172 19276 24212
rect 19316 24172 19358 24212
rect 19398 24172 19440 24212
rect 19112 24163 19480 24172
rect 23112 24212 23480 24221
rect 23152 24172 23194 24212
rect 23234 24172 23276 24212
rect 23316 24172 23358 24212
rect 23398 24172 23440 24212
rect 23112 24163 23480 24172
rect 27112 24212 27480 24221
rect 27152 24172 27194 24212
rect 27234 24172 27276 24212
rect 27316 24172 27358 24212
rect 27398 24172 27440 24212
rect 27112 24163 27480 24172
rect 31112 24212 31480 24221
rect 31152 24172 31194 24212
rect 31234 24172 31276 24212
rect 31316 24172 31358 24212
rect 31398 24172 31440 24212
rect 31112 24163 31480 24172
rect 35112 24212 35480 24221
rect 35152 24172 35194 24212
rect 35234 24172 35276 24212
rect 35316 24172 35358 24212
rect 35398 24172 35440 24212
rect 35112 24163 35480 24172
rect 39112 24212 39480 24221
rect 39152 24172 39194 24212
rect 39234 24172 39276 24212
rect 39316 24172 39358 24212
rect 39398 24172 39440 24212
rect 39112 24163 39480 24172
rect 43112 24212 43480 24221
rect 43152 24172 43194 24212
rect 43234 24172 43276 24212
rect 43316 24172 43358 24212
rect 43398 24172 43440 24212
rect 43112 24163 43480 24172
rect 47112 24212 47480 24221
rect 47152 24172 47194 24212
rect 47234 24172 47276 24212
rect 47316 24172 47358 24212
rect 47398 24172 47440 24212
rect 47112 24163 47480 24172
rect 51112 24212 51480 24221
rect 51152 24172 51194 24212
rect 51234 24172 51276 24212
rect 51316 24172 51358 24212
rect 51398 24172 51440 24212
rect 51112 24163 51480 24172
rect 55112 24212 55480 24221
rect 55152 24172 55194 24212
rect 55234 24172 55276 24212
rect 55316 24172 55358 24212
rect 55398 24172 55440 24212
rect 55112 24163 55480 24172
rect 59112 24212 59480 24221
rect 59152 24172 59194 24212
rect 59234 24172 59276 24212
rect 59316 24172 59358 24212
rect 59398 24172 59440 24212
rect 59112 24163 59480 24172
rect 63112 24212 63480 24221
rect 63152 24172 63194 24212
rect 63234 24172 63276 24212
rect 63316 24172 63358 24212
rect 63398 24172 63440 24212
rect 63112 24163 63480 24172
rect 67112 24212 67480 24221
rect 67152 24172 67194 24212
rect 67234 24172 67276 24212
rect 67316 24172 67358 24212
rect 67398 24172 67440 24212
rect 67112 24163 67480 24172
rect 71112 24212 71480 24221
rect 71152 24172 71194 24212
rect 71234 24172 71276 24212
rect 71316 24172 71358 24212
rect 71398 24172 71440 24212
rect 71112 24163 71480 24172
rect 75112 24212 75480 24221
rect 75152 24172 75194 24212
rect 75234 24172 75276 24212
rect 75316 24172 75358 24212
rect 75398 24172 75440 24212
rect 75112 24163 75480 24172
rect 79112 24212 79480 24221
rect 79152 24172 79194 24212
rect 79234 24172 79276 24212
rect 79316 24172 79358 24212
rect 79398 24172 79440 24212
rect 79112 24163 79480 24172
rect 83112 24212 83480 24221
rect 83152 24172 83194 24212
rect 83234 24172 83276 24212
rect 83316 24172 83358 24212
rect 83398 24172 83440 24212
rect 83112 24163 83480 24172
rect 87112 24212 87480 24221
rect 87152 24172 87194 24212
rect 87234 24172 87276 24212
rect 87316 24172 87358 24212
rect 87398 24172 87440 24212
rect 87112 24163 87480 24172
rect 91112 24212 91480 24221
rect 91152 24172 91194 24212
rect 91234 24172 91276 24212
rect 91316 24172 91358 24212
rect 91398 24172 91440 24212
rect 91112 24163 91480 24172
rect 95112 24212 95480 24221
rect 95152 24172 95194 24212
rect 95234 24172 95276 24212
rect 95316 24172 95358 24212
rect 95398 24172 95440 24212
rect 95112 24163 95480 24172
rect 99112 24212 99480 24221
rect 99152 24172 99194 24212
rect 99234 24172 99276 24212
rect 99316 24172 99358 24212
rect 99398 24172 99440 24212
rect 99112 24163 99480 24172
rect 4352 23456 4720 23465
rect 4392 23416 4434 23456
rect 4474 23416 4516 23456
rect 4556 23416 4598 23456
rect 4638 23416 4680 23456
rect 4352 23407 4720 23416
rect 8352 23456 8720 23465
rect 8392 23416 8434 23456
rect 8474 23416 8516 23456
rect 8556 23416 8598 23456
rect 8638 23416 8680 23456
rect 8352 23407 8720 23416
rect 12352 23456 12720 23465
rect 12392 23416 12434 23456
rect 12474 23416 12516 23456
rect 12556 23416 12598 23456
rect 12638 23416 12680 23456
rect 12352 23407 12720 23416
rect 16352 23456 16720 23465
rect 16392 23416 16434 23456
rect 16474 23416 16516 23456
rect 16556 23416 16598 23456
rect 16638 23416 16680 23456
rect 16352 23407 16720 23416
rect 20352 23456 20720 23465
rect 20392 23416 20434 23456
rect 20474 23416 20516 23456
rect 20556 23416 20598 23456
rect 20638 23416 20680 23456
rect 20352 23407 20720 23416
rect 24352 23456 24720 23465
rect 24392 23416 24434 23456
rect 24474 23416 24516 23456
rect 24556 23416 24598 23456
rect 24638 23416 24680 23456
rect 24352 23407 24720 23416
rect 28352 23456 28720 23465
rect 28392 23416 28434 23456
rect 28474 23416 28516 23456
rect 28556 23416 28598 23456
rect 28638 23416 28680 23456
rect 28352 23407 28720 23416
rect 32352 23456 32720 23465
rect 32392 23416 32434 23456
rect 32474 23416 32516 23456
rect 32556 23416 32598 23456
rect 32638 23416 32680 23456
rect 32352 23407 32720 23416
rect 36352 23456 36720 23465
rect 36392 23416 36434 23456
rect 36474 23416 36516 23456
rect 36556 23416 36598 23456
rect 36638 23416 36680 23456
rect 36352 23407 36720 23416
rect 40352 23456 40720 23465
rect 40392 23416 40434 23456
rect 40474 23416 40516 23456
rect 40556 23416 40598 23456
rect 40638 23416 40680 23456
rect 40352 23407 40720 23416
rect 44352 23456 44720 23465
rect 44392 23416 44434 23456
rect 44474 23416 44516 23456
rect 44556 23416 44598 23456
rect 44638 23416 44680 23456
rect 44352 23407 44720 23416
rect 48352 23456 48720 23465
rect 48392 23416 48434 23456
rect 48474 23416 48516 23456
rect 48556 23416 48598 23456
rect 48638 23416 48680 23456
rect 48352 23407 48720 23416
rect 52352 23456 52720 23465
rect 52392 23416 52434 23456
rect 52474 23416 52516 23456
rect 52556 23416 52598 23456
rect 52638 23416 52680 23456
rect 52352 23407 52720 23416
rect 56352 23456 56720 23465
rect 56392 23416 56434 23456
rect 56474 23416 56516 23456
rect 56556 23416 56598 23456
rect 56638 23416 56680 23456
rect 56352 23407 56720 23416
rect 60352 23456 60720 23465
rect 60392 23416 60434 23456
rect 60474 23416 60516 23456
rect 60556 23416 60598 23456
rect 60638 23416 60680 23456
rect 60352 23407 60720 23416
rect 64352 23456 64720 23465
rect 64392 23416 64434 23456
rect 64474 23416 64516 23456
rect 64556 23416 64598 23456
rect 64638 23416 64680 23456
rect 64352 23407 64720 23416
rect 68352 23456 68720 23465
rect 68392 23416 68434 23456
rect 68474 23416 68516 23456
rect 68556 23416 68598 23456
rect 68638 23416 68680 23456
rect 68352 23407 68720 23416
rect 72352 23456 72720 23465
rect 72392 23416 72434 23456
rect 72474 23416 72516 23456
rect 72556 23416 72598 23456
rect 72638 23416 72680 23456
rect 72352 23407 72720 23416
rect 76352 23456 76720 23465
rect 76392 23416 76434 23456
rect 76474 23416 76516 23456
rect 76556 23416 76598 23456
rect 76638 23416 76680 23456
rect 76352 23407 76720 23416
rect 80352 23456 80720 23465
rect 80392 23416 80434 23456
rect 80474 23416 80516 23456
rect 80556 23416 80598 23456
rect 80638 23416 80680 23456
rect 80352 23407 80720 23416
rect 84352 23456 84720 23465
rect 84392 23416 84434 23456
rect 84474 23416 84516 23456
rect 84556 23416 84598 23456
rect 84638 23416 84680 23456
rect 84352 23407 84720 23416
rect 88352 23456 88720 23465
rect 88392 23416 88434 23456
rect 88474 23416 88516 23456
rect 88556 23416 88598 23456
rect 88638 23416 88680 23456
rect 88352 23407 88720 23416
rect 92352 23456 92720 23465
rect 92392 23416 92434 23456
rect 92474 23416 92516 23456
rect 92556 23416 92598 23456
rect 92638 23416 92680 23456
rect 92352 23407 92720 23416
rect 96352 23456 96720 23465
rect 96392 23416 96434 23456
rect 96474 23416 96516 23456
rect 96556 23416 96598 23456
rect 96638 23416 96680 23456
rect 96352 23407 96720 23416
rect 3112 22700 3480 22709
rect 3152 22660 3194 22700
rect 3234 22660 3276 22700
rect 3316 22660 3358 22700
rect 3398 22660 3440 22700
rect 3112 22651 3480 22660
rect 7112 22700 7480 22709
rect 7152 22660 7194 22700
rect 7234 22660 7276 22700
rect 7316 22660 7358 22700
rect 7398 22660 7440 22700
rect 7112 22651 7480 22660
rect 11112 22700 11480 22709
rect 11152 22660 11194 22700
rect 11234 22660 11276 22700
rect 11316 22660 11358 22700
rect 11398 22660 11440 22700
rect 11112 22651 11480 22660
rect 15112 22700 15480 22709
rect 15152 22660 15194 22700
rect 15234 22660 15276 22700
rect 15316 22660 15358 22700
rect 15398 22660 15440 22700
rect 15112 22651 15480 22660
rect 19112 22700 19480 22709
rect 19152 22660 19194 22700
rect 19234 22660 19276 22700
rect 19316 22660 19358 22700
rect 19398 22660 19440 22700
rect 19112 22651 19480 22660
rect 23112 22700 23480 22709
rect 23152 22660 23194 22700
rect 23234 22660 23276 22700
rect 23316 22660 23358 22700
rect 23398 22660 23440 22700
rect 23112 22651 23480 22660
rect 27112 22700 27480 22709
rect 27152 22660 27194 22700
rect 27234 22660 27276 22700
rect 27316 22660 27358 22700
rect 27398 22660 27440 22700
rect 27112 22651 27480 22660
rect 31112 22700 31480 22709
rect 31152 22660 31194 22700
rect 31234 22660 31276 22700
rect 31316 22660 31358 22700
rect 31398 22660 31440 22700
rect 31112 22651 31480 22660
rect 35112 22700 35480 22709
rect 35152 22660 35194 22700
rect 35234 22660 35276 22700
rect 35316 22660 35358 22700
rect 35398 22660 35440 22700
rect 35112 22651 35480 22660
rect 39112 22700 39480 22709
rect 39152 22660 39194 22700
rect 39234 22660 39276 22700
rect 39316 22660 39358 22700
rect 39398 22660 39440 22700
rect 39112 22651 39480 22660
rect 43112 22700 43480 22709
rect 43152 22660 43194 22700
rect 43234 22660 43276 22700
rect 43316 22660 43358 22700
rect 43398 22660 43440 22700
rect 43112 22651 43480 22660
rect 47112 22700 47480 22709
rect 47152 22660 47194 22700
rect 47234 22660 47276 22700
rect 47316 22660 47358 22700
rect 47398 22660 47440 22700
rect 47112 22651 47480 22660
rect 51112 22700 51480 22709
rect 51152 22660 51194 22700
rect 51234 22660 51276 22700
rect 51316 22660 51358 22700
rect 51398 22660 51440 22700
rect 51112 22651 51480 22660
rect 55112 22700 55480 22709
rect 55152 22660 55194 22700
rect 55234 22660 55276 22700
rect 55316 22660 55358 22700
rect 55398 22660 55440 22700
rect 55112 22651 55480 22660
rect 59112 22700 59480 22709
rect 59152 22660 59194 22700
rect 59234 22660 59276 22700
rect 59316 22660 59358 22700
rect 59398 22660 59440 22700
rect 59112 22651 59480 22660
rect 63112 22700 63480 22709
rect 63152 22660 63194 22700
rect 63234 22660 63276 22700
rect 63316 22660 63358 22700
rect 63398 22660 63440 22700
rect 63112 22651 63480 22660
rect 67112 22700 67480 22709
rect 67152 22660 67194 22700
rect 67234 22660 67276 22700
rect 67316 22660 67358 22700
rect 67398 22660 67440 22700
rect 67112 22651 67480 22660
rect 71112 22700 71480 22709
rect 71152 22660 71194 22700
rect 71234 22660 71276 22700
rect 71316 22660 71358 22700
rect 71398 22660 71440 22700
rect 71112 22651 71480 22660
rect 75112 22700 75480 22709
rect 75152 22660 75194 22700
rect 75234 22660 75276 22700
rect 75316 22660 75358 22700
rect 75398 22660 75440 22700
rect 75112 22651 75480 22660
rect 79112 22700 79480 22709
rect 79152 22660 79194 22700
rect 79234 22660 79276 22700
rect 79316 22660 79358 22700
rect 79398 22660 79440 22700
rect 79112 22651 79480 22660
rect 83112 22700 83480 22709
rect 83152 22660 83194 22700
rect 83234 22660 83276 22700
rect 83316 22660 83358 22700
rect 83398 22660 83440 22700
rect 83112 22651 83480 22660
rect 87112 22700 87480 22709
rect 87152 22660 87194 22700
rect 87234 22660 87276 22700
rect 87316 22660 87358 22700
rect 87398 22660 87440 22700
rect 87112 22651 87480 22660
rect 91112 22700 91480 22709
rect 91152 22660 91194 22700
rect 91234 22660 91276 22700
rect 91316 22660 91358 22700
rect 91398 22660 91440 22700
rect 91112 22651 91480 22660
rect 95112 22700 95480 22709
rect 95152 22660 95194 22700
rect 95234 22660 95276 22700
rect 95316 22660 95358 22700
rect 95398 22660 95440 22700
rect 95112 22651 95480 22660
rect 99112 22700 99480 22709
rect 99152 22660 99194 22700
rect 99234 22660 99276 22700
rect 99316 22660 99358 22700
rect 99398 22660 99440 22700
rect 99112 22651 99480 22660
rect 4352 21944 4720 21953
rect 4392 21904 4434 21944
rect 4474 21904 4516 21944
rect 4556 21904 4598 21944
rect 4638 21904 4680 21944
rect 4352 21895 4720 21904
rect 8352 21944 8720 21953
rect 8392 21904 8434 21944
rect 8474 21904 8516 21944
rect 8556 21904 8598 21944
rect 8638 21904 8680 21944
rect 8352 21895 8720 21904
rect 12352 21944 12720 21953
rect 12392 21904 12434 21944
rect 12474 21904 12516 21944
rect 12556 21904 12598 21944
rect 12638 21904 12680 21944
rect 12352 21895 12720 21904
rect 16352 21944 16720 21953
rect 16392 21904 16434 21944
rect 16474 21904 16516 21944
rect 16556 21904 16598 21944
rect 16638 21904 16680 21944
rect 16352 21895 16720 21904
rect 20352 21944 20720 21953
rect 20392 21904 20434 21944
rect 20474 21904 20516 21944
rect 20556 21904 20598 21944
rect 20638 21904 20680 21944
rect 20352 21895 20720 21904
rect 24352 21944 24720 21953
rect 24392 21904 24434 21944
rect 24474 21904 24516 21944
rect 24556 21904 24598 21944
rect 24638 21904 24680 21944
rect 24352 21895 24720 21904
rect 28352 21944 28720 21953
rect 28392 21904 28434 21944
rect 28474 21904 28516 21944
rect 28556 21904 28598 21944
rect 28638 21904 28680 21944
rect 28352 21895 28720 21904
rect 32352 21944 32720 21953
rect 32392 21904 32434 21944
rect 32474 21904 32516 21944
rect 32556 21904 32598 21944
rect 32638 21904 32680 21944
rect 32352 21895 32720 21904
rect 36352 21944 36720 21953
rect 36392 21904 36434 21944
rect 36474 21904 36516 21944
rect 36556 21904 36598 21944
rect 36638 21904 36680 21944
rect 36352 21895 36720 21904
rect 40352 21944 40720 21953
rect 40392 21904 40434 21944
rect 40474 21904 40516 21944
rect 40556 21904 40598 21944
rect 40638 21904 40680 21944
rect 40352 21895 40720 21904
rect 44352 21944 44720 21953
rect 44392 21904 44434 21944
rect 44474 21904 44516 21944
rect 44556 21904 44598 21944
rect 44638 21904 44680 21944
rect 44352 21895 44720 21904
rect 48352 21944 48720 21953
rect 48392 21904 48434 21944
rect 48474 21904 48516 21944
rect 48556 21904 48598 21944
rect 48638 21904 48680 21944
rect 48352 21895 48720 21904
rect 52352 21944 52720 21953
rect 52392 21904 52434 21944
rect 52474 21904 52516 21944
rect 52556 21904 52598 21944
rect 52638 21904 52680 21944
rect 52352 21895 52720 21904
rect 56352 21944 56720 21953
rect 56392 21904 56434 21944
rect 56474 21904 56516 21944
rect 56556 21904 56598 21944
rect 56638 21904 56680 21944
rect 56352 21895 56720 21904
rect 60352 21944 60720 21953
rect 60392 21904 60434 21944
rect 60474 21904 60516 21944
rect 60556 21904 60598 21944
rect 60638 21904 60680 21944
rect 60352 21895 60720 21904
rect 64352 21944 64720 21953
rect 64392 21904 64434 21944
rect 64474 21904 64516 21944
rect 64556 21904 64598 21944
rect 64638 21904 64680 21944
rect 64352 21895 64720 21904
rect 68352 21944 68720 21953
rect 68392 21904 68434 21944
rect 68474 21904 68516 21944
rect 68556 21904 68598 21944
rect 68638 21904 68680 21944
rect 68352 21895 68720 21904
rect 72352 21944 72720 21953
rect 72392 21904 72434 21944
rect 72474 21904 72516 21944
rect 72556 21904 72598 21944
rect 72638 21904 72680 21944
rect 72352 21895 72720 21904
rect 76352 21944 76720 21953
rect 76392 21904 76434 21944
rect 76474 21904 76516 21944
rect 76556 21904 76598 21944
rect 76638 21904 76680 21944
rect 76352 21895 76720 21904
rect 80352 21944 80720 21953
rect 80392 21904 80434 21944
rect 80474 21904 80516 21944
rect 80556 21904 80598 21944
rect 80638 21904 80680 21944
rect 80352 21895 80720 21904
rect 84352 21944 84720 21953
rect 84392 21904 84434 21944
rect 84474 21904 84516 21944
rect 84556 21904 84598 21944
rect 84638 21904 84680 21944
rect 84352 21895 84720 21904
rect 88352 21944 88720 21953
rect 88392 21904 88434 21944
rect 88474 21904 88516 21944
rect 88556 21904 88598 21944
rect 88638 21904 88680 21944
rect 88352 21895 88720 21904
rect 92352 21944 92720 21953
rect 92392 21904 92434 21944
rect 92474 21904 92516 21944
rect 92556 21904 92598 21944
rect 92638 21904 92680 21944
rect 92352 21895 92720 21904
rect 96352 21944 96720 21953
rect 96392 21904 96434 21944
rect 96474 21904 96516 21944
rect 96556 21904 96598 21944
rect 96638 21904 96680 21944
rect 96352 21895 96720 21904
rect 3112 21188 3480 21197
rect 3152 21148 3194 21188
rect 3234 21148 3276 21188
rect 3316 21148 3358 21188
rect 3398 21148 3440 21188
rect 3112 21139 3480 21148
rect 7112 21188 7480 21197
rect 7152 21148 7194 21188
rect 7234 21148 7276 21188
rect 7316 21148 7358 21188
rect 7398 21148 7440 21188
rect 7112 21139 7480 21148
rect 11112 21188 11480 21197
rect 11152 21148 11194 21188
rect 11234 21148 11276 21188
rect 11316 21148 11358 21188
rect 11398 21148 11440 21188
rect 11112 21139 11480 21148
rect 15112 21188 15480 21197
rect 15152 21148 15194 21188
rect 15234 21148 15276 21188
rect 15316 21148 15358 21188
rect 15398 21148 15440 21188
rect 15112 21139 15480 21148
rect 19112 21188 19480 21197
rect 19152 21148 19194 21188
rect 19234 21148 19276 21188
rect 19316 21148 19358 21188
rect 19398 21148 19440 21188
rect 19112 21139 19480 21148
rect 23112 21188 23480 21197
rect 23152 21148 23194 21188
rect 23234 21148 23276 21188
rect 23316 21148 23358 21188
rect 23398 21148 23440 21188
rect 23112 21139 23480 21148
rect 27112 21188 27480 21197
rect 27152 21148 27194 21188
rect 27234 21148 27276 21188
rect 27316 21148 27358 21188
rect 27398 21148 27440 21188
rect 27112 21139 27480 21148
rect 31112 21188 31480 21197
rect 31152 21148 31194 21188
rect 31234 21148 31276 21188
rect 31316 21148 31358 21188
rect 31398 21148 31440 21188
rect 31112 21139 31480 21148
rect 35112 21188 35480 21197
rect 35152 21148 35194 21188
rect 35234 21148 35276 21188
rect 35316 21148 35358 21188
rect 35398 21148 35440 21188
rect 35112 21139 35480 21148
rect 39112 21188 39480 21197
rect 39152 21148 39194 21188
rect 39234 21148 39276 21188
rect 39316 21148 39358 21188
rect 39398 21148 39440 21188
rect 39112 21139 39480 21148
rect 43112 21188 43480 21197
rect 43152 21148 43194 21188
rect 43234 21148 43276 21188
rect 43316 21148 43358 21188
rect 43398 21148 43440 21188
rect 43112 21139 43480 21148
rect 47112 21188 47480 21197
rect 47152 21148 47194 21188
rect 47234 21148 47276 21188
rect 47316 21148 47358 21188
rect 47398 21148 47440 21188
rect 47112 21139 47480 21148
rect 51112 21188 51480 21197
rect 51152 21148 51194 21188
rect 51234 21148 51276 21188
rect 51316 21148 51358 21188
rect 51398 21148 51440 21188
rect 51112 21139 51480 21148
rect 55112 21188 55480 21197
rect 55152 21148 55194 21188
rect 55234 21148 55276 21188
rect 55316 21148 55358 21188
rect 55398 21148 55440 21188
rect 55112 21139 55480 21148
rect 59112 21188 59480 21197
rect 59152 21148 59194 21188
rect 59234 21148 59276 21188
rect 59316 21148 59358 21188
rect 59398 21148 59440 21188
rect 59112 21139 59480 21148
rect 63112 21188 63480 21197
rect 63152 21148 63194 21188
rect 63234 21148 63276 21188
rect 63316 21148 63358 21188
rect 63398 21148 63440 21188
rect 63112 21139 63480 21148
rect 67112 21188 67480 21197
rect 67152 21148 67194 21188
rect 67234 21148 67276 21188
rect 67316 21148 67358 21188
rect 67398 21148 67440 21188
rect 67112 21139 67480 21148
rect 71112 21188 71480 21197
rect 71152 21148 71194 21188
rect 71234 21148 71276 21188
rect 71316 21148 71358 21188
rect 71398 21148 71440 21188
rect 71112 21139 71480 21148
rect 75112 21188 75480 21197
rect 75152 21148 75194 21188
rect 75234 21148 75276 21188
rect 75316 21148 75358 21188
rect 75398 21148 75440 21188
rect 75112 21139 75480 21148
rect 79112 21188 79480 21197
rect 79152 21148 79194 21188
rect 79234 21148 79276 21188
rect 79316 21148 79358 21188
rect 79398 21148 79440 21188
rect 79112 21139 79480 21148
rect 83112 21188 83480 21197
rect 83152 21148 83194 21188
rect 83234 21148 83276 21188
rect 83316 21148 83358 21188
rect 83398 21148 83440 21188
rect 83112 21139 83480 21148
rect 87112 21188 87480 21197
rect 87152 21148 87194 21188
rect 87234 21148 87276 21188
rect 87316 21148 87358 21188
rect 87398 21148 87440 21188
rect 87112 21139 87480 21148
rect 91112 21188 91480 21197
rect 91152 21148 91194 21188
rect 91234 21148 91276 21188
rect 91316 21148 91358 21188
rect 91398 21148 91440 21188
rect 91112 21139 91480 21148
rect 95112 21188 95480 21197
rect 95152 21148 95194 21188
rect 95234 21148 95276 21188
rect 95316 21148 95358 21188
rect 95398 21148 95440 21188
rect 95112 21139 95480 21148
rect 99112 21188 99480 21197
rect 99152 21148 99194 21188
rect 99234 21148 99276 21188
rect 99316 21148 99358 21188
rect 99398 21148 99440 21188
rect 99112 21139 99480 21148
rect 4352 20432 4720 20441
rect 4392 20392 4434 20432
rect 4474 20392 4516 20432
rect 4556 20392 4598 20432
rect 4638 20392 4680 20432
rect 4352 20383 4720 20392
rect 8352 20432 8720 20441
rect 8392 20392 8434 20432
rect 8474 20392 8516 20432
rect 8556 20392 8598 20432
rect 8638 20392 8680 20432
rect 8352 20383 8720 20392
rect 12352 20432 12720 20441
rect 12392 20392 12434 20432
rect 12474 20392 12516 20432
rect 12556 20392 12598 20432
rect 12638 20392 12680 20432
rect 12352 20383 12720 20392
rect 16352 20432 16720 20441
rect 16392 20392 16434 20432
rect 16474 20392 16516 20432
rect 16556 20392 16598 20432
rect 16638 20392 16680 20432
rect 16352 20383 16720 20392
rect 20352 20432 20720 20441
rect 20392 20392 20434 20432
rect 20474 20392 20516 20432
rect 20556 20392 20598 20432
rect 20638 20392 20680 20432
rect 20352 20383 20720 20392
rect 24352 20432 24720 20441
rect 24392 20392 24434 20432
rect 24474 20392 24516 20432
rect 24556 20392 24598 20432
rect 24638 20392 24680 20432
rect 24352 20383 24720 20392
rect 28352 20432 28720 20441
rect 28392 20392 28434 20432
rect 28474 20392 28516 20432
rect 28556 20392 28598 20432
rect 28638 20392 28680 20432
rect 28352 20383 28720 20392
rect 32352 20432 32720 20441
rect 32392 20392 32434 20432
rect 32474 20392 32516 20432
rect 32556 20392 32598 20432
rect 32638 20392 32680 20432
rect 32352 20383 32720 20392
rect 36352 20432 36720 20441
rect 36392 20392 36434 20432
rect 36474 20392 36516 20432
rect 36556 20392 36598 20432
rect 36638 20392 36680 20432
rect 36352 20383 36720 20392
rect 40352 20432 40720 20441
rect 40392 20392 40434 20432
rect 40474 20392 40516 20432
rect 40556 20392 40598 20432
rect 40638 20392 40680 20432
rect 40352 20383 40720 20392
rect 44352 20432 44720 20441
rect 44392 20392 44434 20432
rect 44474 20392 44516 20432
rect 44556 20392 44598 20432
rect 44638 20392 44680 20432
rect 44352 20383 44720 20392
rect 48352 20432 48720 20441
rect 48392 20392 48434 20432
rect 48474 20392 48516 20432
rect 48556 20392 48598 20432
rect 48638 20392 48680 20432
rect 48352 20383 48720 20392
rect 52352 20432 52720 20441
rect 52392 20392 52434 20432
rect 52474 20392 52516 20432
rect 52556 20392 52598 20432
rect 52638 20392 52680 20432
rect 52352 20383 52720 20392
rect 56352 20432 56720 20441
rect 56392 20392 56434 20432
rect 56474 20392 56516 20432
rect 56556 20392 56598 20432
rect 56638 20392 56680 20432
rect 56352 20383 56720 20392
rect 60352 20432 60720 20441
rect 60392 20392 60434 20432
rect 60474 20392 60516 20432
rect 60556 20392 60598 20432
rect 60638 20392 60680 20432
rect 60352 20383 60720 20392
rect 64352 20432 64720 20441
rect 64392 20392 64434 20432
rect 64474 20392 64516 20432
rect 64556 20392 64598 20432
rect 64638 20392 64680 20432
rect 64352 20383 64720 20392
rect 68352 20432 68720 20441
rect 68392 20392 68434 20432
rect 68474 20392 68516 20432
rect 68556 20392 68598 20432
rect 68638 20392 68680 20432
rect 68352 20383 68720 20392
rect 72352 20432 72720 20441
rect 72392 20392 72434 20432
rect 72474 20392 72516 20432
rect 72556 20392 72598 20432
rect 72638 20392 72680 20432
rect 72352 20383 72720 20392
rect 76352 20432 76720 20441
rect 76392 20392 76434 20432
rect 76474 20392 76516 20432
rect 76556 20392 76598 20432
rect 76638 20392 76680 20432
rect 76352 20383 76720 20392
rect 80352 20432 80720 20441
rect 80392 20392 80434 20432
rect 80474 20392 80516 20432
rect 80556 20392 80598 20432
rect 80638 20392 80680 20432
rect 80352 20383 80720 20392
rect 84352 20432 84720 20441
rect 84392 20392 84434 20432
rect 84474 20392 84516 20432
rect 84556 20392 84598 20432
rect 84638 20392 84680 20432
rect 84352 20383 84720 20392
rect 88352 20432 88720 20441
rect 88392 20392 88434 20432
rect 88474 20392 88516 20432
rect 88556 20392 88598 20432
rect 88638 20392 88680 20432
rect 88352 20383 88720 20392
rect 92352 20432 92720 20441
rect 92392 20392 92434 20432
rect 92474 20392 92516 20432
rect 92556 20392 92598 20432
rect 92638 20392 92680 20432
rect 92352 20383 92720 20392
rect 96352 20432 96720 20441
rect 96392 20392 96434 20432
rect 96474 20392 96516 20432
rect 96556 20392 96598 20432
rect 96638 20392 96680 20432
rect 96352 20383 96720 20392
rect 3112 19676 3480 19685
rect 3152 19636 3194 19676
rect 3234 19636 3276 19676
rect 3316 19636 3358 19676
rect 3398 19636 3440 19676
rect 3112 19627 3480 19636
rect 7112 19676 7480 19685
rect 7152 19636 7194 19676
rect 7234 19636 7276 19676
rect 7316 19636 7358 19676
rect 7398 19636 7440 19676
rect 7112 19627 7480 19636
rect 11112 19676 11480 19685
rect 11152 19636 11194 19676
rect 11234 19636 11276 19676
rect 11316 19636 11358 19676
rect 11398 19636 11440 19676
rect 11112 19627 11480 19636
rect 15112 19676 15480 19685
rect 15152 19636 15194 19676
rect 15234 19636 15276 19676
rect 15316 19636 15358 19676
rect 15398 19636 15440 19676
rect 15112 19627 15480 19636
rect 19112 19676 19480 19685
rect 19152 19636 19194 19676
rect 19234 19636 19276 19676
rect 19316 19636 19358 19676
rect 19398 19636 19440 19676
rect 19112 19627 19480 19636
rect 23112 19676 23480 19685
rect 23152 19636 23194 19676
rect 23234 19636 23276 19676
rect 23316 19636 23358 19676
rect 23398 19636 23440 19676
rect 23112 19627 23480 19636
rect 27112 19676 27480 19685
rect 27152 19636 27194 19676
rect 27234 19636 27276 19676
rect 27316 19636 27358 19676
rect 27398 19636 27440 19676
rect 27112 19627 27480 19636
rect 31112 19676 31480 19685
rect 31152 19636 31194 19676
rect 31234 19636 31276 19676
rect 31316 19636 31358 19676
rect 31398 19636 31440 19676
rect 31112 19627 31480 19636
rect 35112 19676 35480 19685
rect 35152 19636 35194 19676
rect 35234 19636 35276 19676
rect 35316 19636 35358 19676
rect 35398 19636 35440 19676
rect 35112 19627 35480 19636
rect 39112 19676 39480 19685
rect 39152 19636 39194 19676
rect 39234 19636 39276 19676
rect 39316 19636 39358 19676
rect 39398 19636 39440 19676
rect 39112 19627 39480 19636
rect 43112 19676 43480 19685
rect 43152 19636 43194 19676
rect 43234 19636 43276 19676
rect 43316 19636 43358 19676
rect 43398 19636 43440 19676
rect 43112 19627 43480 19636
rect 47112 19676 47480 19685
rect 47152 19636 47194 19676
rect 47234 19636 47276 19676
rect 47316 19636 47358 19676
rect 47398 19636 47440 19676
rect 47112 19627 47480 19636
rect 51112 19676 51480 19685
rect 51152 19636 51194 19676
rect 51234 19636 51276 19676
rect 51316 19636 51358 19676
rect 51398 19636 51440 19676
rect 51112 19627 51480 19636
rect 55112 19676 55480 19685
rect 55152 19636 55194 19676
rect 55234 19636 55276 19676
rect 55316 19636 55358 19676
rect 55398 19636 55440 19676
rect 55112 19627 55480 19636
rect 59112 19676 59480 19685
rect 59152 19636 59194 19676
rect 59234 19636 59276 19676
rect 59316 19636 59358 19676
rect 59398 19636 59440 19676
rect 59112 19627 59480 19636
rect 63112 19676 63480 19685
rect 63152 19636 63194 19676
rect 63234 19636 63276 19676
rect 63316 19636 63358 19676
rect 63398 19636 63440 19676
rect 63112 19627 63480 19636
rect 67112 19676 67480 19685
rect 67152 19636 67194 19676
rect 67234 19636 67276 19676
rect 67316 19636 67358 19676
rect 67398 19636 67440 19676
rect 67112 19627 67480 19636
rect 71112 19676 71480 19685
rect 71152 19636 71194 19676
rect 71234 19636 71276 19676
rect 71316 19636 71358 19676
rect 71398 19636 71440 19676
rect 71112 19627 71480 19636
rect 75112 19676 75480 19685
rect 75152 19636 75194 19676
rect 75234 19636 75276 19676
rect 75316 19636 75358 19676
rect 75398 19636 75440 19676
rect 75112 19627 75480 19636
rect 79112 19676 79480 19685
rect 79152 19636 79194 19676
rect 79234 19636 79276 19676
rect 79316 19636 79358 19676
rect 79398 19636 79440 19676
rect 79112 19627 79480 19636
rect 83112 19676 83480 19685
rect 83152 19636 83194 19676
rect 83234 19636 83276 19676
rect 83316 19636 83358 19676
rect 83398 19636 83440 19676
rect 83112 19627 83480 19636
rect 87112 19676 87480 19685
rect 87152 19636 87194 19676
rect 87234 19636 87276 19676
rect 87316 19636 87358 19676
rect 87398 19636 87440 19676
rect 87112 19627 87480 19636
rect 91112 19676 91480 19685
rect 91152 19636 91194 19676
rect 91234 19636 91276 19676
rect 91316 19636 91358 19676
rect 91398 19636 91440 19676
rect 91112 19627 91480 19636
rect 95112 19676 95480 19685
rect 95152 19636 95194 19676
rect 95234 19636 95276 19676
rect 95316 19636 95358 19676
rect 95398 19636 95440 19676
rect 95112 19627 95480 19636
rect 99112 19676 99480 19685
rect 99152 19636 99194 19676
rect 99234 19636 99276 19676
rect 99316 19636 99358 19676
rect 99398 19636 99440 19676
rect 99112 19627 99480 19636
rect 4352 18920 4720 18929
rect 4392 18880 4434 18920
rect 4474 18880 4516 18920
rect 4556 18880 4598 18920
rect 4638 18880 4680 18920
rect 4352 18871 4720 18880
rect 8352 18920 8720 18929
rect 8392 18880 8434 18920
rect 8474 18880 8516 18920
rect 8556 18880 8598 18920
rect 8638 18880 8680 18920
rect 8352 18871 8720 18880
rect 12352 18920 12720 18929
rect 12392 18880 12434 18920
rect 12474 18880 12516 18920
rect 12556 18880 12598 18920
rect 12638 18880 12680 18920
rect 12352 18871 12720 18880
rect 16352 18920 16720 18929
rect 16392 18880 16434 18920
rect 16474 18880 16516 18920
rect 16556 18880 16598 18920
rect 16638 18880 16680 18920
rect 16352 18871 16720 18880
rect 20352 18920 20720 18929
rect 20392 18880 20434 18920
rect 20474 18880 20516 18920
rect 20556 18880 20598 18920
rect 20638 18880 20680 18920
rect 20352 18871 20720 18880
rect 24352 18920 24720 18929
rect 24392 18880 24434 18920
rect 24474 18880 24516 18920
rect 24556 18880 24598 18920
rect 24638 18880 24680 18920
rect 24352 18871 24720 18880
rect 28352 18920 28720 18929
rect 28392 18880 28434 18920
rect 28474 18880 28516 18920
rect 28556 18880 28598 18920
rect 28638 18880 28680 18920
rect 28352 18871 28720 18880
rect 32352 18920 32720 18929
rect 32392 18880 32434 18920
rect 32474 18880 32516 18920
rect 32556 18880 32598 18920
rect 32638 18880 32680 18920
rect 32352 18871 32720 18880
rect 36352 18920 36720 18929
rect 36392 18880 36434 18920
rect 36474 18880 36516 18920
rect 36556 18880 36598 18920
rect 36638 18880 36680 18920
rect 36352 18871 36720 18880
rect 40352 18920 40720 18929
rect 40392 18880 40434 18920
rect 40474 18880 40516 18920
rect 40556 18880 40598 18920
rect 40638 18880 40680 18920
rect 40352 18871 40720 18880
rect 44352 18920 44720 18929
rect 44392 18880 44434 18920
rect 44474 18880 44516 18920
rect 44556 18880 44598 18920
rect 44638 18880 44680 18920
rect 44352 18871 44720 18880
rect 48352 18920 48720 18929
rect 48392 18880 48434 18920
rect 48474 18880 48516 18920
rect 48556 18880 48598 18920
rect 48638 18880 48680 18920
rect 48352 18871 48720 18880
rect 52352 18920 52720 18929
rect 52392 18880 52434 18920
rect 52474 18880 52516 18920
rect 52556 18880 52598 18920
rect 52638 18880 52680 18920
rect 52352 18871 52720 18880
rect 56352 18920 56720 18929
rect 56392 18880 56434 18920
rect 56474 18880 56516 18920
rect 56556 18880 56598 18920
rect 56638 18880 56680 18920
rect 56352 18871 56720 18880
rect 60352 18920 60720 18929
rect 60392 18880 60434 18920
rect 60474 18880 60516 18920
rect 60556 18880 60598 18920
rect 60638 18880 60680 18920
rect 60352 18871 60720 18880
rect 64352 18920 64720 18929
rect 64392 18880 64434 18920
rect 64474 18880 64516 18920
rect 64556 18880 64598 18920
rect 64638 18880 64680 18920
rect 64352 18871 64720 18880
rect 68352 18920 68720 18929
rect 68392 18880 68434 18920
rect 68474 18880 68516 18920
rect 68556 18880 68598 18920
rect 68638 18880 68680 18920
rect 68352 18871 68720 18880
rect 72352 18920 72720 18929
rect 72392 18880 72434 18920
rect 72474 18880 72516 18920
rect 72556 18880 72598 18920
rect 72638 18880 72680 18920
rect 72352 18871 72720 18880
rect 76352 18920 76720 18929
rect 76392 18880 76434 18920
rect 76474 18880 76516 18920
rect 76556 18880 76598 18920
rect 76638 18880 76680 18920
rect 76352 18871 76720 18880
rect 80352 18920 80720 18929
rect 80392 18880 80434 18920
rect 80474 18880 80516 18920
rect 80556 18880 80598 18920
rect 80638 18880 80680 18920
rect 80352 18871 80720 18880
rect 84352 18920 84720 18929
rect 84392 18880 84434 18920
rect 84474 18880 84516 18920
rect 84556 18880 84598 18920
rect 84638 18880 84680 18920
rect 84352 18871 84720 18880
rect 88352 18920 88720 18929
rect 88392 18880 88434 18920
rect 88474 18880 88516 18920
rect 88556 18880 88598 18920
rect 88638 18880 88680 18920
rect 88352 18871 88720 18880
rect 92352 18920 92720 18929
rect 92392 18880 92434 18920
rect 92474 18880 92516 18920
rect 92556 18880 92598 18920
rect 92638 18880 92680 18920
rect 92352 18871 92720 18880
rect 96352 18920 96720 18929
rect 96392 18880 96434 18920
rect 96474 18880 96516 18920
rect 96556 18880 96598 18920
rect 96638 18880 96680 18920
rect 96352 18871 96720 18880
rect 3112 18164 3480 18173
rect 3152 18124 3194 18164
rect 3234 18124 3276 18164
rect 3316 18124 3358 18164
rect 3398 18124 3440 18164
rect 3112 18115 3480 18124
rect 7112 18164 7480 18173
rect 7152 18124 7194 18164
rect 7234 18124 7276 18164
rect 7316 18124 7358 18164
rect 7398 18124 7440 18164
rect 7112 18115 7480 18124
rect 11112 18164 11480 18173
rect 11152 18124 11194 18164
rect 11234 18124 11276 18164
rect 11316 18124 11358 18164
rect 11398 18124 11440 18164
rect 11112 18115 11480 18124
rect 15112 18164 15480 18173
rect 15152 18124 15194 18164
rect 15234 18124 15276 18164
rect 15316 18124 15358 18164
rect 15398 18124 15440 18164
rect 15112 18115 15480 18124
rect 19112 18164 19480 18173
rect 19152 18124 19194 18164
rect 19234 18124 19276 18164
rect 19316 18124 19358 18164
rect 19398 18124 19440 18164
rect 19112 18115 19480 18124
rect 23112 18164 23480 18173
rect 23152 18124 23194 18164
rect 23234 18124 23276 18164
rect 23316 18124 23358 18164
rect 23398 18124 23440 18164
rect 23112 18115 23480 18124
rect 27112 18164 27480 18173
rect 27152 18124 27194 18164
rect 27234 18124 27276 18164
rect 27316 18124 27358 18164
rect 27398 18124 27440 18164
rect 27112 18115 27480 18124
rect 31112 18164 31480 18173
rect 31152 18124 31194 18164
rect 31234 18124 31276 18164
rect 31316 18124 31358 18164
rect 31398 18124 31440 18164
rect 31112 18115 31480 18124
rect 35112 18164 35480 18173
rect 35152 18124 35194 18164
rect 35234 18124 35276 18164
rect 35316 18124 35358 18164
rect 35398 18124 35440 18164
rect 35112 18115 35480 18124
rect 39112 18164 39480 18173
rect 39152 18124 39194 18164
rect 39234 18124 39276 18164
rect 39316 18124 39358 18164
rect 39398 18124 39440 18164
rect 39112 18115 39480 18124
rect 43112 18164 43480 18173
rect 43152 18124 43194 18164
rect 43234 18124 43276 18164
rect 43316 18124 43358 18164
rect 43398 18124 43440 18164
rect 43112 18115 43480 18124
rect 47112 18164 47480 18173
rect 47152 18124 47194 18164
rect 47234 18124 47276 18164
rect 47316 18124 47358 18164
rect 47398 18124 47440 18164
rect 47112 18115 47480 18124
rect 51112 18164 51480 18173
rect 51152 18124 51194 18164
rect 51234 18124 51276 18164
rect 51316 18124 51358 18164
rect 51398 18124 51440 18164
rect 51112 18115 51480 18124
rect 55112 18164 55480 18173
rect 55152 18124 55194 18164
rect 55234 18124 55276 18164
rect 55316 18124 55358 18164
rect 55398 18124 55440 18164
rect 55112 18115 55480 18124
rect 59112 18164 59480 18173
rect 59152 18124 59194 18164
rect 59234 18124 59276 18164
rect 59316 18124 59358 18164
rect 59398 18124 59440 18164
rect 59112 18115 59480 18124
rect 63112 18164 63480 18173
rect 63152 18124 63194 18164
rect 63234 18124 63276 18164
rect 63316 18124 63358 18164
rect 63398 18124 63440 18164
rect 63112 18115 63480 18124
rect 67112 18164 67480 18173
rect 67152 18124 67194 18164
rect 67234 18124 67276 18164
rect 67316 18124 67358 18164
rect 67398 18124 67440 18164
rect 67112 18115 67480 18124
rect 71112 18164 71480 18173
rect 71152 18124 71194 18164
rect 71234 18124 71276 18164
rect 71316 18124 71358 18164
rect 71398 18124 71440 18164
rect 71112 18115 71480 18124
rect 75112 18164 75480 18173
rect 75152 18124 75194 18164
rect 75234 18124 75276 18164
rect 75316 18124 75358 18164
rect 75398 18124 75440 18164
rect 75112 18115 75480 18124
rect 79112 18164 79480 18173
rect 79152 18124 79194 18164
rect 79234 18124 79276 18164
rect 79316 18124 79358 18164
rect 79398 18124 79440 18164
rect 79112 18115 79480 18124
rect 83112 18164 83480 18173
rect 83152 18124 83194 18164
rect 83234 18124 83276 18164
rect 83316 18124 83358 18164
rect 83398 18124 83440 18164
rect 83112 18115 83480 18124
rect 87112 18164 87480 18173
rect 87152 18124 87194 18164
rect 87234 18124 87276 18164
rect 87316 18124 87358 18164
rect 87398 18124 87440 18164
rect 87112 18115 87480 18124
rect 91112 18164 91480 18173
rect 91152 18124 91194 18164
rect 91234 18124 91276 18164
rect 91316 18124 91358 18164
rect 91398 18124 91440 18164
rect 91112 18115 91480 18124
rect 95112 18164 95480 18173
rect 95152 18124 95194 18164
rect 95234 18124 95276 18164
rect 95316 18124 95358 18164
rect 95398 18124 95440 18164
rect 95112 18115 95480 18124
rect 99112 18164 99480 18173
rect 99152 18124 99194 18164
rect 99234 18124 99276 18164
rect 99316 18124 99358 18164
rect 99398 18124 99440 18164
rect 99112 18115 99480 18124
rect 4352 17408 4720 17417
rect 4392 17368 4434 17408
rect 4474 17368 4516 17408
rect 4556 17368 4598 17408
rect 4638 17368 4680 17408
rect 4352 17359 4720 17368
rect 8352 17408 8720 17417
rect 8392 17368 8434 17408
rect 8474 17368 8516 17408
rect 8556 17368 8598 17408
rect 8638 17368 8680 17408
rect 8352 17359 8720 17368
rect 12352 17408 12720 17417
rect 12392 17368 12434 17408
rect 12474 17368 12516 17408
rect 12556 17368 12598 17408
rect 12638 17368 12680 17408
rect 12352 17359 12720 17368
rect 16352 17408 16720 17417
rect 16392 17368 16434 17408
rect 16474 17368 16516 17408
rect 16556 17368 16598 17408
rect 16638 17368 16680 17408
rect 16352 17359 16720 17368
rect 20352 17408 20720 17417
rect 20392 17368 20434 17408
rect 20474 17368 20516 17408
rect 20556 17368 20598 17408
rect 20638 17368 20680 17408
rect 20352 17359 20720 17368
rect 24352 17408 24720 17417
rect 24392 17368 24434 17408
rect 24474 17368 24516 17408
rect 24556 17368 24598 17408
rect 24638 17368 24680 17408
rect 24352 17359 24720 17368
rect 28352 17408 28720 17417
rect 28392 17368 28434 17408
rect 28474 17368 28516 17408
rect 28556 17368 28598 17408
rect 28638 17368 28680 17408
rect 28352 17359 28720 17368
rect 32352 17408 32720 17417
rect 32392 17368 32434 17408
rect 32474 17368 32516 17408
rect 32556 17368 32598 17408
rect 32638 17368 32680 17408
rect 32352 17359 32720 17368
rect 36352 17408 36720 17417
rect 36392 17368 36434 17408
rect 36474 17368 36516 17408
rect 36556 17368 36598 17408
rect 36638 17368 36680 17408
rect 36352 17359 36720 17368
rect 40352 17408 40720 17417
rect 40392 17368 40434 17408
rect 40474 17368 40516 17408
rect 40556 17368 40598 17408
rect 40638 17368 40680 17408
rect 40352 17359 40720 17368
rect 44352 17408 44720 17417
rect 44392 17368 44434 17408
rect 44474 17368 44516 17408
rect 44556 17368 44598 17408
rect 44638 17368 44680 17408
rect 44352 17359 44720 17368
rect 48352 17408 48720 17417
rect 48392 17368 48434 17408
rect 48474 17368 48516 17408
rect 48556 17368 48598 17408
rect 48638 17368 48680 17408
rect 48352 17359 48720 17368
rect 52352 17408 52720 17417
rect 52392 17368 52434 17408
rect 52474 17368 52516 17408
rect 52556 17368 52598 17408
rect 52638 17368 52680 17408
rect 52352 17359 52720 17368
rect 56352 17408 56720 17417
rect 56392 17368 56434 17408
rect 56474 17368 56516 17408
rect 56556 17368 56598 17408
rect 56638 17368 56680 17408
rect 56352 17359 56720 17368
rect 60352 17408 60720 17417
rect 60392 17368 60434 17408
rect 60474 17368 60516 17408
rect 60556 17368 60598 17408
rect 60638 17368 60680 17408
rect 60352 17359 60720 17368
rect 64352 17408 64720 17417
rect 64392 17368 64434 17408
rect 64474 17368 64516 17408
rect 64556 17368 64598 17408
rect 64638 17368 64680 17408
rect 64352 17359 64720 17368
rect 68352 17408 68720 17417
rect 68392 17368 68434 17408
rect 68474 17368 68516 17408
rect 68556 17368 68598 17408
rect 68638 17368 68680 17408
rect 68352 17359 68720 17368
rect 72352 17408 72720 17417
rect 72392 17368 72434 17408
rect 72474 17368 72516 17408
rect 72556 17368 72598 17408
rect 72638 17368 72680 17408
rect 72352 17359 72720 17368
rect 76352 17408 76720 17417
rect 76392 17368 76434 17408
rect 76474 17368 76516 17408
rect 76556 17368 76598 17408
rect 76638 17368 76680 17408
rect 76352 17359 76720 17368
rect 80352 17408 80720 17417
rect 80392 17368 80434 17408
rect 80474 17368 80516 17408
rect 80556 17368 80598 17408
rect 80638 17368 80680 17408
rect 80352 17359 80720 17368
rect 84352 17408 84720 17417
rect 84392 17368 84434 17408
rect 84474 17368 84516 17408
rect 84556 17368 84598 17408
rect 84638 17368 84680 17408
rect 84352 17359 84720 17368
rect 88352 17408 88720 17417
rect 88392 17368 88434 17408
rect 88474 17368 88516 17408
rect 88556 17368 88598 17408
rect 88638 17368 88680 17408
rect 88352 17359 88720 17368
rect 92352 17408 92720 17417
rect 92392 17368 92434 17408
rect 92474 17368 92516 17408
rect 92556 17368 92598 17408
rect 92638 17368 92680 17408
rect 92352 17359 92720 17368
rect 96352 17408 96720 17417
rect 96392 17368 96434 17408
rect 96474 17368 96516 17408
rect 96556 17368 96598 17408
rect 96638 17368 96680 17408
rect 96352 17359 96720 17368
rect 3112 16652 3480 16661
rect 3152 16612 3194 16652
rect 3234 16612 3276 16652
rect 3316 16612 3358 16652
rect 3398 16612 3440 16652
rect 3112 16603 3480 16612
rect 7112 16652 7480 16661
rect 7152 16612 7194 16652
rect 7234 16612 7276 16652
rect 7316 16612 7358 16652
rect 7398 16612 7440 16652
rect 7112 16603 7480 16612
rect 11112 16652 11480 16661
rect 11152 16612 11194 16652
rect 11234 16612 11276 16652
rect 11316 16612 11358 16652
rect 11398 16612 11440 16652
rect 11112 16603 11480 16612
rect 15112 16652 15480 16661
rect 15152 16612 15194 16652
rect 15234 16612 15276 16652
rect 15316 16612 15358 16652
rect 15398 16612 15440 16652
rect 15112 16603 15480 16612
rect 19112 16652 19480 16661
rect 19152 16612 19194 16652
rect 19234 16612 19276 16652
rect 19316 16612 19358 16652
rect 19398 16612 19440 16652
rect 19112 16603 19480 16612
rect 23112 16652 23480 16661
rect 23152 16612 23194 16652
rect 23234 16612 23276 16652
rect 23316 16612 23358 16652
rect 23398 16612 23440 16652
rect 23112 16603 23480 16612
rect 27112 16652 27480 16661
rect 27152 16612 27194 16652
rect 27234 16612 27276 16652
rect 27316 16612 27358 16652
rect 27398 16612 27440 16652
rect 27112 16603 27480 16612
rect 31112 16652 31480 16661
rect 31152 16612 31194 16652
rect 31234 16612 31276 16652
rect 31316 16612 31358 16652
rect 31398 16612 31440 16652
rect 31112 16603 31480 16612
rect 35112 16652 35480 16661
rect 35152 16612 35194 16652
rect 35234 16612 35276 16652
rect 35316 16612 35358 16652
rect 35398 16612 35440 16652
rect 35112 16603 35480 16612
rect 39112 16652 39480 16661
rect 39152 16612 39194 16652
rect 39234 16612 39276 16652
rect 39316 16612 39358 16652
rect 39398 16612 39440 16652
rect 39112 16603 39480 16612
rect 43112 16652 43480 16661
rect 43152 16612 43194 16652
rect 43234 16612 43276 16652
rect 43316 16612 43358 16652
rect 43398 16612 43440 16652
rect 43112 16603 43480 16612
rect 47112 16652 47480 16661
rect 47152 16612 47194 16652
rect 47234 16612 47276 16652
rect 47316 16612 47358 16652
rect 47398 16612 47440 16652
rect 47112 16603 47480 16612
rect 51112 16652 51480 16661
rect 51152 16612 51194 16652
rect 51234 16612 51276 16652
rect 51316 16612 51358 16652
rect 51398 16612 51440 16652
rect 51112 16603 51480 16612
rect 55112 16652 55480 16661
rect 55152 16612 55194 16652
rect 55234 16612 55276 16652
rect 55316 16612 55358 16652
rect 55398 16612 55440 16652
rect 55112 16603 55480 16612
rect 59112 16652 59480 16661
rect 59152 16612 59194 16652
rect 59234 16612 59276 16652
rect 59316 16612 59358 16652
rect 59398 16612 59440 16652
rect 59112 16603 59480 16612
rect 63112 16652 63480 16661
rect 63152 16612 63194 16652
rect 63234 16612 63276 16652
rect 63316 16612 63358 16652
rect 63398 16612 63440 16652
rect 63112 16603 63480 16612
rect 67112 16652 67480 16661
rect 67152 16612 67194 16652
rect 67234 16612 67276 16652
rect 67316 16612 67358 16652
rect 67398 16612 67440 16652
rect 67112 16603 67480 16612
rect 71112 16652 71480 16661
rect 71152 16612 71194 16652
rect 71234 16612 71276 16652
rect 71316 16612 71358 16652
rect 71398 16612 71440 16652
rect 71112 16603 71480 16612
rect 75112 16652 75480 16661
rect 75152 16612 75194 16652
rect 75234 16612 75276 16652
rect 75316 16612 75358 16652
rect 75398 16612 75440 16652
rect 75112 16603 75480 16612
rect 79112 16652 79480 16661
rect 79152 16612 79194 16652
rect 79234 16612 79276 16652
rect 79316 16612 79358 16652
rect 79398 16612 79440 16652
rect 79112 16603 79480 16612
rect 83112 16652 83480 16661
rect 83152 16612 83194 16652
rect 83234 16612 83276 16652
rect 83316 16612 83358 16652
rect 83398 16612 83440 16652
rect 83112 16603 83480 16612
rect 87112 16652 87480 16661
rect 87152 16612 87194 16652
rect 87234 16612 87276 16652
rect 87316 16612 87358 16652
rect 87398 16612 87440 16652
rect 87112 16603 87480 16612
rect 91112 16652 91480 16661
rect 91152 16612 91194 16652
rect 91234 16612 91276 16652
rect 91316 16612 91358 16652
rect 91398 16612 91440 16652
rect 91112 16603 91480 16612
rect 95112 16652 95480 16661
rect 95152 16612 95194 16652
rect 95234 16612 95276 16652
rect 95316 16612 95358 16652
rect 95398 16612 95440 16652
rect 95112 16603 95480 16612
rect 99112 16652 99480 16661
rect 99152 16612 99194 16652
rect 99234 16612 99276 16652
rect 99316 16612 99358 16652
rect 99398 16612 99440 16652
rect 99112 16603 99480 16612
rect 86187 16400 86229 16409
rect 86187 16360 86188 16400
rect 86228 16360 86229 16400
rect 86187 16351 86229 16360
rect 86188 16266 86228 16351
rect 4352 15896 4720 15905
rect 4392 15856 4434 15896
rect 4474 15856 4516 15896
rect 4556 15856 4598 15896
rect 4638 15856 4680 15896
rect 4352 15847 4720 15856
rect 8352 15896 8720 15905
rect 8392 15856 8434 15896
rect 8474 15856 8516 15896
rect 8556 15856 8598 15896
rect 8638 15856 8680 15896
rect 8352 15847 8720 15856
rect 12352 15896 12720 15905
rect 12392 15856 12434 15896
rect 12474 15856 12516 15896
rect 12556 15856 12598 15896
rect 12638 15856 12680 15896
rect 12352 15847 12720 15856
rect 16352 15896 16720 15905
rect 16392 15856 16434 15896
rect 16474 15856 16516 15896
rect 16556 15856 16598 15896
rect 16638 15856 16680 15896
rect 16352 15847 16720 15856
rect 20352 15896 20720 15905
rect 20392 15856 20434 15896
rect 20474 15856 20516 15896
rect 20556 15856 20598 15896
rect 20638 15856 20680 15896
rect 20352 15847 20720 15856
rect 24352 15896 24720 15905
rect 24392 15856 24434 15896
rect 24474 15856 24516 15896
rect 24556 15856 24598 15896
rect 24638 15856 24680 15896
rect 24352 15847 24720 15856
rect 28352 15896 28720 15905
rect 28392 15856 28434 15896
rect 28474 15856 28516 15896
rect 28556 15856 28598 15896
rect 28638 15856 28680 15896
rect 28352 15847 28720 15856
rect 32352 15896 32720 15905
rect 32392 15856 32434 15896
rect 32474 15856 32516 15896
rect 32556 15856 32598 15896
rect 32638 15856 32680 15896
rect 32352 15847 32720 15856
rect 36352 15896 36720 15905
rect 36392 15856 36434 15896
rect 36474 15856 36516 15896
rect 36556 15856 36598 15896
rect 36638 15856 36680 15896
rect 36352 15847 36720 15856
rect 40352 15896 40720 15905
rect 40392 15856 40434 15896
rect 40474 15856 40516 15896
rect 40556 15856 40598 15896
rect 40638 15856 40680 15896
rect 40352 15847 40720 15856
rect 44352 15896 44720 15905
rect 44392 15856 44434 15896
rect 44474 15856 44516 15896
rect 44556 15856 44598 15896
rect 44638 15856 44680 15896
rect 44352 15847 44720 15856
rect 48352 15896 48720 15905
rect 48392 15856 48434 15896
rect 48474 15856 48516 15896
rect 48556 15856 48598 15896
rect 48638 15856 48680 15896
rect 48352 15847 48720 15856
rect 52352 15896 52720 15905
rect 52392 15856 52434 15896
rect 52474 15856 52516 15896
rect 52556 15856 52598 15896
rect 52638 15856 52680 15896
rect 52352 15847 52720 15856
rect 56352 15896 56720 15905
rect 56392 15856 56434 15896
rect 56474 15856 56516 15896
rect 56556 15856 56598 15896
rect 56638 15856 56680 15896
rect 56352 15847 56720 15856
rect 60352 15896 60720 15905
rect 60392 15856 60434 15896
rect 60474 15856 60516 15896
rect 60556 15856 60598 15896
rect 60638 15856 60680 15896
rect 60352 15847 60720 15856
rect 64352 15896 64720 15905
rect 64392 15856 64434 15896
rect 64474 15856 64516 15896
rect 64556 15856 64598 15896
rect 64638 15856 64680 15896
rect 64352 15847 64720 15856
rect 68352 15896 68720 15905
rect 68392 15856 68434 15896
rect 68474 15856 68516 15896
rect 68556 15856 68598 15896
rect 68638 15856 68680 15896
rect 68352 15847 68720 15856
rect 72352 15896 72720 15905
rect 72392 15856 72434 15896
rect 72474 15856 72516 15896
rect 72556 15856 72598 15896
rect 72638 15856 72680 15896
rect 72352 15847 72720 15856
rect 76352 15896 76720 15905
rect 76392 15856 76434 15896
rect 76474 15856 76516 15896
rect 76556 15856 76598 15896
rect 76638 15856 76680 15896
rect 76352 15847 76720 15856
rect 80352 15896 80720 15905
rect 80392 15856 80434 15896
rect 80474 15856 80516 15896
rect 80556 15856 80598 15896
rect 80638 15856 80680 15896
rect 80352 15847 80720 15856
rect 84352 15896 84720 15905
rect 84392 15856 84434 15896
rect 84474 15856 84516 15896
rect 84556 15856 84598 15896
rect 84638 15856 84680 15896
rect 84352 15847 84720 15856
rect 88352 15896 88720 15905
rect 88392 15856 88434 15896
rect 88474 15856 88516 15896
rect 88556 15856 88598 15896
rect 88638 15856 88680 15896
rect 88352 15847 88720 15856
rect 92352 15896 92720 15905
rect 92392 15856 92434 15896
rect 92474 15856 92516 15896
rect 92556 15856 92598 15896
rect 92638 15856 92680 15896
rect 92352 15847 92720 15856
rect 96352 15896 96720 15905
rect 96392 15856 96434 15896
rect 96474 15856 96516 15896
rect 96556 15856 96598 15896
rect 96638 15856 96680 15896
rect 96352 15847 96720 15856
rect 90892 15308 90932 15317
rect 3112 15140 3480 15149
rect 3152 15100 3194 15140
rect 3234 15100 3276 15140
rect 3316 15100 3358 15140
rect 3398 15100 3440 15140
rect 3112 15091 3480 15100
rect 7112 15140 7480 15149
rect 7152 15100 7194 15140
rect 7234 15100 7276 15140
rect 7316 15100 7358 15140
rect 7398 15100 7440 15140
rect 7112 15091 7480 15100
rect 11112 15140 11480 15149
rect 11152 15100 11194 15140
rect 11234 15100 11276 15140
rect 11316 15100 11358 15140
rect 11398 15100 11440 15140
rect 11112 15091 11480 15100
rect 15112 15140 15480 15149
rect 15152 15100 15194 15140
rect 15234 15100 15276 15140
rect 15316 15100 15358 15140
rect 15398 15100 15440 15140
rect 15112 15091 15480 15100
rect 19112 15140 19480 15149
rect 19152 15100 19194 15140
rect 19234 15100 19276 15140
rect 19316 15100 19358 15140
rect 19398 15100 19440 15140
rect 19112 15091 19480 15100
rect 23112 15140 23480 15149
rect 23152 15100 23194 15140
rect 23234 15100 23276 15140
rect 23316 15100 23358 15140
rect 23398 15100 23440 15140
rect 23112 15091 23480 15100
rect 27112 15140 27480 15149
rect 27152 15100 27194 15140
rect 27234 15100 27276 15140
rect 27316 15100 27358 15140
rect 27398 15100 27440 15140
rect 27112 15091 27480 15100
rect 31112 15140 31480 15149
rect 31152 15100 31194 15140
rect 31234 15100 31276 15140
rect 31316 15100 31358 15140
rect 31398 15100 31440 15140
rect 31112 15091 31480 15100
rect 35112 15140 35480 15149
rect 35152 15100 35194 15140
rect 35234 15100 35276 15140
rect 35316 15100 35358 15140
rect 35398 15100 35440 15140
rect 35112 15091 35480 15100
rect 39112 15140 39480 15149
rect 39152 15100 39194 15140
rect 39234 15100 39276 15140
rect 39316 15100 39358 15140
rect 39398 15100 39440 15140
rect 39112 15091 39480 15100
rect 43112 15140 43480 15149
rect 43152 15100 43194 15140
rect 43234 15100 43276 15140
rect 43316 15100 43358 15140
rect 43398 15100 43440 15140
rect 43112 15091 43480 15100
rect 47112 15140 47480 15149
rect 47152 15100 47194 15140
rect 47234 15100 47276 15140
rect 47316 15100 47358 15140
rect 47398 15100 47440 15140
rect 47112 15091 47480 15100
rect 51112 15140 51480 15149
rect 51152 15100 51194 15140
rect 51234 15100 51276 15140
rect 51316 15100 51358 15140
rect 51398 15100 51440 15140
rect 51112 15091 51480 15100
rect 55112 15140 55480 15149
rect 55152 15100 55194 15140
rect 55234 15100 55276 15140
rect 55316 15100 55358 15140
rect 55398 15100 55440 15140
rect 55112 15091 55480 15100
rect 59112 15140 59480 15149
rect 59152 15100 59194 15140
rect 59234 15100 59276 15140
rect 59316 15100 59358 15140
rect 59398 15100 59440 15140
rect 59112 15091 59480 15100
rect 63112 15140 63480 15149
rect 63152 15100 63194 15140
rect 63234 15100 63276 15140
rect 63316 15100 63358 15140
rect 63398 15100 63440 15140
rect 63112 15091 63480 15100
rect 67112 15140 67480 15149
rect 67152 15100 67194 15140
rect 67234 15100 67276 15140
rect 67316 15100 67358 15140
rect 67398 15100 67440 15140
rect 67112 15091 67480 15100
rect 4352 14384 4720 14393
rect 4392 14344 4434 14384
rect 4474 14344 4516 14384
rect 4556 14344 4598 14384
rect 4638 14344 4680 14384
rect 4352 14335 4720 14344
rect 8352 14384 8720 14393
rect 8392 14344 8434 14384
rect 8474 14344 8516 14384
rect 8556 14344 8598 14384
rect 8638 14344 8680 14384
rect 8352 14335 8720 14344
rect 12352 14384 12720 14393
rect 12392 14344 12434 14384
rect 12474 14344 12516 14384
rect 12556 14344 12598 14384
rect 12638 14344 12680 14384
rect 12352 14335 12720 14344
rect 16352 14384 16720 14393
rect 16392 14344 16434 14384
rect 16474 14344 16516 14384
rect 16556 14344 16598 14384
rect 16638 14344 16680 14384
rect 16352 14335 16720 14344
rect 20352 14384 20720 14393
rect 20392 14344 20434 14384
rect 20474 14344 20516 14384
rect 20556 14344 20598 14384
rect 20638 14344 20680 14384
rect 20352 14335 20720 14344
rect 24352 14384 24720 14393
rect 24392 14344 24434 14384
rect 24474 14344 24516 14384
rect 24556 14344 24598 14384
rect 24638 14344 24680 14384
rect 24352 14335 24720 14344
rect 28352 14384 28720 14393
rect 28392 14344 28434 14384
rect 28474 14344 28516 14384
rect 28556 14344 28598 14384
rect 28638 14344 28680 14384
rect 28352 14335 28720 14344
rect 32352 14384 32720 14393
rect 32392 14344 32434 14384
rect 32474 14344 32516 14384
rect 32556 14344 32598 14384
rect 32638 14344 32680 14384
rect 32352 14335 32720 14344
rect 36352 14384 36720 14393
rect 36392 14344 36434 14384
rect 36474 14344 36516 14384
rect 36556 14344 36598 14384
rect 36638 14344 36680 14384
rect 36352 14335 36720 14344
rect 40352 14384 40720 14393
rect 40392 14344 40434 14384
rect 40474 14344 40516 14384
rect 40556 14344 40598 14384
rect 40638 14344 40680 14384
rect 40352 14335 40720 14344
rect 44352 14384 44720 14393
rect 44392 14344 44434 14384
rect 44474 14344 44516 14384
rect 44556 14344 44598 14384
rect 44638 14344 44680 14384
rect 44352 14335 44720 14344
rect 48352 14384 48720 14393
rect 48392 14344 48434 14384
rect 48474 14344 48516 14384
rect 48556 14344 48598 14384
rect 48638 14344 48680 14384
rect 48352 14335 48720 14344
rect 52352 14384 52720 14393
rect 52392 14344 52434 14384
rect 52474 14344 52516 14384
rect 52556 14344 52598 14384
rect 52638 14344 52680 14384
rect 52352 14335 52720 14344
rect 56352 14384 56720 14393
rect 56392 14344 56434 14384
rect 56474 14344 56516 14384
rect 56556 14344 56598 14384
rect 56638 14344 56680 14384
rect 56352 14335 56720 14344
rect 60352 14384 60720 14393
rect 60392 14344 60434 14384
rect 60474 14344 60516 14384
rect 60556 14344 60598 14384
rect 60638 14344 60680 14384
rect 60352 14335 60720 14344
rect 64352 14384 64720 14393
rect 64392 14344 64434 14384
rect 64474 14344 64516 14384
rect 64556 14344 64598 14384
rect 64638 14344 64680 14384
rect 64352 14335 64720 14344
rect 68352 14384 68720 14393
rect 68392 14344 68434 14384
rect 68474 14344 68516 14384
rect 68556 14344 68598 14384
rect 68638 14344 68680 14384
rect 68352 14335 68720 14344
rect 3112 13628 3480 13637
rect 3152 13588 3194 13628
rect 3234 13588 3276 13628
rect 3316 13588 3358 13628
rect 3398 13588 3440 13628
rect 3112 13579 3480 13588
rect 7112 13628 7480 13637
rect 7152 13588 7194 13628
rect 7234 13588 7276 13628
rect 7316 13588 7358 13628
rect 7398 13588 7440 13628
rect 7112 13579 7480 13588
rect 11112 13628 11480 13637
rect 11152 13588 11194 13628
rect 11234 13588 11276 13628
rect 11316 13588 11358 13628
rect 11398 13588 11440 13628
rect 11112 13579 11480 13588
rect 15112 13628 15480 13637
rect 15152 13588 15194 13628
rect 15234 13588 15276 13628
rect 15316 13588 15358 13628
rect 15398 13588 15440 13628
rect 15112 13579 15480 13588
rect 19112 13628 19480 13637
rect 19152 13588 19194 13628
rect 19234 13588 19276 13628
rect 19316 13588 19358 13628
rect 19398 13588 19440 13628
rect 19112 13579 19480 13588
rect 23112 13628 23480 13637
rect 23152 13588 23194 13628
rect 23234 13588 23276 13628
rect 23316 13588 23358 13628
rect 23398 13588 23440 13628
rect 23112 13579 23480 13588
rect 27112 13628 27480 13637
rect 27152 13588 27194 13628
rect 27234 13588 27276 13628
rect 27316 13588 27358 13628
rect 27398 13588 27440 13628
rect 27112 13579 27480 13588
rect 31112 13628 31480 13637
rect 31152 13588 31194 13628
rect 31234 13588 31276 13628
rect 31316 13588 31358 13628
rect 31398 13588 31440 13628
rect 31112 13579 31480 13588
rect 35112 13628 35480 13637
rect 35152 13588 35194 13628
rect 35234 13588 35276 13628
rect 35316 13588 35358 13628
rect 35398 13588 35440 13628
rect 35112 13579 35480 13588
rect 39112 13628 39480 13637
rect 39152 13588 39194 13628
rect 39234 13588 39276 13628
rect 39316 13588 39358 13628
rect 39398 13588 39440 13628
rect 39112 13579 39480 13588
rect 43112 13628 43480 13637
rect 43152 13588 43194 13628
rect 43234 13588 43276 13628
rect 43316 13588 43358 13628
rect 43398 13588 43440 13628
rect 43112 13579 43480 13588
rect 47112 13628 47480 13637
rect 47152 13588 47194 13628
rect 47234 13588 47276 13628
rect 47316 13588 47358 13628
rect 47398 13588 47440 13628
rect 47112 13579 47480 13588
rect 51112 13628 51480 13637
rect 51152 13588 51194 13628
rect 51234 13588 51276 13628
rect 51316 13588 51358 13628
rect 51398 13588 51440 13628
rect 51112 13579 51480 13588
rect 55112 13628 55480 13637
rect 55152 13588 55194 13628
rect 55234 13588 55276 13628
rect 55316 13588 55358 13628
rect 55398 13588 55440 13628
rect 55112 13579 55480 13588
rect 59112 13628 59480 13637
rect 59152 13588 59194 13628
rect 59234 13588 59276 13628
rect 59316 13588 59358 13628
rect 59398 13588 59440 13628
rect 59112 13579 59480 13588
rect 63112 13628 63480 13637
rect 63152 13588 63194 13628
rect 63234 13588 63276 13628
rect 63316 13588 63358 13628
rect 63398 13588 63440 13628
rect 63112 13579 63480 13588
rect 67112 13628 67480 13637
rect 67152 13588 67194 13628
rect 67234 13588 67276 13628
rect 67316 13588 67358 13628
rect 67398 13588 67440 13628
rect 67112 13579 67480 13588
rect 90892 13460 90932 15268
rect 90892 13411 90932 13420
rect 72460 13376 72500 13385
rect 71884 13336 72460 13376
rect 71884 13292 71924 13336
rect 72460 13327 72500 13336
rect 71884 13243 71924 13252
rect 4352 12872 4720 12881
rect 4392 12832 4434 12872
rect 4474 12832 4516 12872
rect 4556 12832 4598 12872
rect 4638 12832 4680 12872
rect 4352 12823 4720 12832
rect 8352 12872 8720 12881
rect 8392 12832 8434 12872
rect 8474 12832 8516 12872
rect 8556 12832 8598 12872
rect 8638 12832 8680 12872
rect 8352 12823 8720 12832
rect 12352 12872 12720 12881
rect 12392 12832 12434 12872
rect 12474 12832 12516 12872
rect 12556 12832 12598 12872
rect 12638 12832 12680 12872
rect 12352 12823 12720 12832
rect 16352 12872 16720 12881
rect 16392 12832 16434 12872
rect 16474 12832 16516 12872
rect 16556 12832 16598 12872
rect 16638 12832 16680 12872
rect 16352 12823 16720 12832
rect 20352 12872 20720 12881
rect 20392 12832 20434 12872
rect 20474 12832 20516 12872
rect 20556 12832 20598 12872
rect 20638 12832 20680 12872
rect 20352 12823 20720 12832
rect 24352 12872 24720 12881
rect 24392 12832 24434 12872
rect 24474 12832 24516 12872
rect 24556 12832 24598 12872
rect 24638 12832 24680 12872
rect 24352 12823 24720 12832
rect 28352 12872 28720 12881
rect 28392 12832 28434 12872
rect 28474 12832 28516 12872
rect 28556 12832 28598 12872
rect 28638 12832 28680 12872
rect 28352 12823 28720 12832
rect 32352 12872 32720 12881
rect 32392 12832 32434 12872
rect 32474 12832 32516 12872
rect 32556 12832 32598 12872
rect 32638 12832 32680 12872
rect 32352 12823 32720 12832
rect 36352 12872 36720 12881
rect 36392 12832 36434 12872
rect 36474 12832 36516 12872
rect 36556 12832 36598 12872
rect 36638 12832 36680 12872
rect 36352 12823 36720 12832
rect 40352 12872 40720 12881
rect 40392 12832 40434 12872
rect 40474 12832 40516 12872
rect 40556 12832 40598 12872
rect 40638 12832 40680 12872
rect 40352 12823 40720 12832
rect 44352 12872 44720 12881
rect 44392 12832 44434 12872
rect 44474 12832 44516 12872
rect 44556 12832 44598 12872
rect 44638 12832 44680 12872
rect 44352 12823 44720 12832
rect 48352 12872 48720 12881
rect 48392 12832 48434 12872
rect 48474 12832 48516 12872
rect 48556 12832 48598 12872
rect 48638 12832 48680 12872
rect 48352 12823 48720 12832
rect 52352 12872 52720 12881
rect 52392 12832 52434 12872
rect 52474 12832 52516 12872
rect 52556 12832 52598 12872
rect 52638 12832 52680 12872
rect 52352 12823 52720 12832
rect 56352 12872 56720 12881
rect 56392 12832 56434 12872
rect 56474 12832 56516 12872
rect 56556 12832 56598 12872
rect 56638 12832 56680 12872
rect 56352 12823 56720 12832
rect 60352 12872 60720 12881
rect 60392 12832 60434 12872
rect 60474 12832 60516 12872
rect 60556 12832 60598 12872
rect 60638 12832 60680 12872
rect 60352 12823 60720 12832
rect 64352 12872 64720 12881
rect 64392 12832 64434 12872
rect 64474 12832 64516 12872
rect 64556 12832 64598 12872
rect 64638 12832 64680 12872
rect 64352 12823 64720 12832
rect 68352 12872 68720 12881
rect 68392 12832 68434 12872
rect 68474 12832 68516 12872
rect 68556 12832 68598 12872
rect 68638 12832 68680 12872
rect 68352 12823 68720 12832
rect 3112 12116 3480 12125
rect 3152 12076 3194 12116
rect 3234 12076 3276 12116
rect 3316 12076 3358 12116
rect 3398 12076 3440 12116
rect 3112 12067 3480 12076
rect 7112 12116 7480 12125
rect 7152 12076 7194 12116
rect 7234 12076 7276 12116
rect 7316 12076 7358 12116
rect 7398 12076 7440 12116
rect 7112 12067 7480 12076
rect 11112 12116 11480 12125
rect 11152 12076 11194 12116
rect 11234 12076 11276 12116
rect 11316 12076 11358 12116
rect 11398 12076 11440 12116
rect 11112 12067 11480 12076
rect 15112 12116 15480 12125
rect 15152 12076 15194 12116
rect 15234 12076 15276 12116
rect 15316 12076 15358 12116
rect 15398 12076 15440 12116
rect 15112 12067 15480 12076
rect 19112 12116 19480 12125
rect 19152 12076 19194 12116
rect 19234 12076 19276 12116
rect 19316 12076 19358 12116
rect 19398 12076 19440 12116
rect 19112 12067 19480 12076
rect 23112 12116 23480 12125
rect 23152 12076 23194 12116
rect 23234 12076 23276 12116
rect 23316 12076 23358 12116
rect 23398 12076 23440 12116
rect 23112 12067 23480 12076
rect 27112 12116 27480 12125
rect 27152 12076 27194 12116
rect 27234 12076 27276 12116
rect 27316 12076 27358 12116
rect 27398 12076 27440 12116
rect 27112 12067 27480 12076
rect 31112 12116 31480 12125
rect 31152 12076 31194 12116
rect 31234 12076 31276 12116
rect 31316 12076 31358 12116
rect 31398 12076 31440 12116
rect 31112 12067 31480 12076
rect 35112 12116 35480 12125
rect 35152 12076 35194 12116
rect 35234 12076 35276 12116
rect 35316 12076 35358 12116
rect 35398 12076 35440 12116
rect 35112 12067 35480 12076
rect 39112 12116 39480 12125
rect 39152 12076 39194 12116
rect 39234 12076 39276 12116
rect 39316 12076 39358 12116
rect 39398 12076 39440 12116
rect 39112 12067 39480 12076
rect 43112 12116 43480 12125
rect 43152 12076 43194 12116
rect 43234 12076 43276 12116
rect 43316 12076 43358 12116
rect 43398 12076 43440 12116
rect 43112 12067 43480 12076
rect 47112 12116 47480 12125
rect 47152 12076 47194 12116
rect 47234 12076 47276 12116
rect 47316 12076 47358 12116
rect 47398 12076 47440 12116
rect 47112 12067 47480 12076
rect 51112 12116 51480 12125
rect 51152 12076 51194 12116
rect 51234 12076 51276 12116
rect 51316 12076 51358 12116
rect 51398 12076 51440 12116
rect 51112 12067 51480 12076
rect 55112 12116 55480 12125
rect 55152 12076 55194 12116
rect 55234 12076 55276 12116
rect 55316 12076 55358 12116
rect 55398 12076 55440 12116
rect 55112 12067 55480 12076
rect 59112 12116 59480 12125
rect 59152 12076 59194 12116
rect 59234 12076 59276 12116
rect 59316 12076 59358 12116
rect 59398 12076 59440 12116
rect 59112 12067 59480 12076
rect 63112 12116 63480 12125
rect 63152 12076 63194 12116
rect 63234 12076 63276 12116
rect 63316 12076 63358 12116
rect 63398 12076 63440 12116
rect 63112 12067 63480 12076
rect 67112 12116 67480 12125
rect 67152 12076 67194 12116
rect 67234 12076 67276 12116
rect 67316 12076 67358 12116
rect 67398 12076 67440 12116
rect 67112 12067 67480 12076
rect 4352 11360 4720 11369
rect 4392 11320 4434 11360
rect 4474 11320 4516 11360
rect 4556 11320 4598 11360
rect 4638 11320 4680 11360
rect 4352 11311 4720 11320
rect 8352 11360 8720 11369
rect 8392 11320 8434 11360
rect 8474 11320 8516 11360
rect 8556 11320 8598 11360
rect 8638 11320 8680 11360
rect 8352 11311 8720 11320
rect 12352 11360 12720 11369
rect 12392 11320 12434 11360
rect 12474 11320 12516 11360
rect 12556 11320 12598 11360
rect 12638 11320 12680 11360
rect 12352 11311 12720 11320
rect 16352 11360 16720 11369
rect 16392 11320 16434 11360
rect 16474 11320 16516 11360
rect 16556 11320 16598 11360
rect 16638 11320 16680 11360
rect 16352 11311 16720 11320
rect 20352 11360 20720 11369
rect 20392 11320 20434 11360
rect 20474 11320 20516 11360
rect 20556 11320 20598 11360
rect 20638 11320 20680 11360
rect 20352 11311 20720 11320
rect 24352 11360 24720 11369
rect 24392 11320 24434 11360
rect 24474 11320 24516 11360
rect 24556 11320 24598 11360
rect 24638 11320 24680 11360
rect 24352 11311 24720 11320
rect 28352 11360 28720 11369
rect 28392 11320 28434 11360
rect 28474 11320 28516 11360
rect 28556 11320 28598 11360
rect 28638 11320 28680 11360
rect 28352 11311 28720 11320
rect 32352 11360 32720 11369
rect 32392 11320 32434 11360
rect 32474 11320 32516 11360
rect 32556 11320 32598 11360
rect 32638 11320 32680 11360
rect 32352 11311 32720 11320
rect 36352 11360 36720 11369
rect 36392 11320 36434 11360
rect 36474 11320 36516 11360
rect 36556 11320 36598 11360
rect 36638 11320 36680 11360
rect 36352 11311 36720 11320
rect 40352 11360 40720 11369
rect 40392 11320 40434 11360
rect 40474 11320 40516 11360
rect 40556 11320 40598 11360
rect 40638 11320 40680 11360
rect 40352 11311 40720 11320
rect 44352 11360 44720 11369
rect 44392 11320 44434 11360
rect 44474 11320 44516 11360
rect 44556 11320 44598 11360
rect 44638 11320 44680 11360
rect 44352 11311 44720 11320
rect 48352 11360 48720 11369
rect 48392 11320 48434 11360
rect 48474 11320 48516 11360
rect 48556 11320 48598 11360
rect 48638 11320 48680 11360
rect 48352 11311 48720 11320
rect 52352 11360 52720 11369
rect 52392 11320 52434 11360
rect 52474 11320 52516 11360
rect 52556 11320 52598 11360
rect 52638 11320 52680 11360
rect 52352 11311 52720 11320
rect 56352 11360 56720 11369
rect 56392 11320 56434 11360
rect 56474 11320 56516 11360
rect 56556 11320 56598 11360
rect 56638 11320 56680 11360
rect 56352 11311 56720 11320
rect 60352 11360 60720 11369
rect 60392 11320 60434 11360
rect 60474 11320 60516 11360
rect 60556 11320 60598 11360
rect 60638 11320 60680 11360
rect 60352 11311 60720 11320
rect 64352 11360 64720 11369
rect 64392 11320 64434 11360
rect 64474 11320 64516 11360
rect 64556 11320 64598 11360
rect 64638 11320 64680 11360
rect 64352 11311 64720 11320
rect 68352 11360 68720 11369
rect 68392 11320 68434 11360
rect 68474 11320 68516 11360
rect 68556 11320 68598 11360
rect 68638 11320 68680 11360
rect 68352 11311 68720 11320
rect 3112 10604 3480 10613
rect 3152 10564 3194 10604
rect 3234 10564 3276 10604
rect 3316 10564 3358 10604
rect 3398 10564 3440 10604
rect 3112 10555 3480 10564
rect 7112 10604 7480 10613
rect 7152 10564 7194 10604
rect 7234 10564 7276 10604
rect 7316 10564 7358 10604
rect 7398 10564 7440 10604
rect 7112 10555 7480 10564
rect 11112 10604 11480 10613
rect 11152 10564 11194 10604
rect 11234 10564 11276 10604
rect 11316 10564 11358 10604
rect 11398 10564 11440 10604
rect 11112 10555 11480 10564
rect 15112 10604 15480 10613
rect 15152 10564 15194 10604
rect 15234 10564 15276 10604
rect 15316 10564 15358 10604
rect 15398 10564 15440 10604
rect 15112 10555 15480 10564
rect 19112 10604 19480 10613
rect 19152 10564 19194 10604
rect 19234 10564 19276 10604
rect 19316 10564 19358 10604
rect 19398 10564 19440 10604
rect 19112 10555 19480 10564
rect 23112 10604 23480 10613
rect 23152 10564 23194 10604
rect 23234 10564 23276 10604
rect 23316 10564 23358 10604
rect 23398 10564 23440 10604
rect 23112 10555 23480 10564
rect 27112 10604 27480 10613
rect 27152 10564 27194 10604
rect 27234 10564 27276 10604
rect 27316 10564 27358 10604
rect 27398 10564 27440 10604
rect 27112 10555 27480 10564
rect 31112 10604 31480 10613
rect 31152 10564 31194 10604
rect 31234 10564 31276 10604
rect 31316 10564 31358 10604
rect 31398 10564 31440 10604
rect 31112 10555 31480 10564
rect 35112 10604 35480 10613
rect 35152 10564 35194 10604
rect 35234 10564 35276 10604
rect 35316 10564 35358 10604
rect 35398 10564 35440 10604
rect 35112 10555 35480 10564
rect 39112 10604 39480 10613
rect 39152 10564 39194 10604
rect 39234 10564 39276 10604
rect 39316 10564 39358 10604
rect 39398 10564 39440 10604
rect 39112 10555 39480 10564
rect 43112 10604 43480 10613
rect 43152 10564 43194 10604
rect 43234 10564 43276 10604
rect 43316 10564 43358 10604
rect 43398 10564 43440 10604
rect 43112 10555 43480 10564
rect 47112 10604 47480 10613
rect 47152 10564 47194 10604
rect 47234 10564 47276 10604
rect 47316 10564 47358 10604
rect 47398 10564 47440 10604
rect 47112 10555 47480 10564
rect 51112 10604 51480 10613
rect 51152 10564 51194 10604
rect 51234 10564 51276 10604
rect 51316 10564 51358 10604
rect 51398 10564 51440 10604
rect 51112 10555 51480 10564
rect 55112 10604 55480 10613
rect 55152 10564 55194 10604
rect 55234 10564 55276 10604
rect 55316 10564 55358 10604
rect 55398 10564 55440 10604
rect 55112 10555 55480 10564
rect 59112 10604 59480 10613
rect 59152 10564 59194 10604
rect 59234 10564 59276 10604
rect 59316 10564 59358 10604
rect 59398 10564 59440 10604
rect 59112 10555 59480 10564
rect 63112 10604 63480 10613
rect 63152 10564 63194 10604
rect 63234 10564 63276 10604
rect 63316 10564 63358 10604
rect 63398 10564 63440 10604
rect 63112 10555 63480 10564
rect 67112 10604 67480 10613
rect 67152 10564 67194 10604
rect 67234 10564 67276 10604
rect 67316 10564 67358 10604
rect 67398 10564 67440 10604
rect 67112 10555 67480 10564
rect 4352 9848 4720 9857
rect 4392 9808 4434 9848
rect 4474 9808 4516 9848
rect 4556 9808 4598 9848
rect 4638 9808 4680 9848
rect 4352 9799 4720 9808
rect 8352 9848 8720 9857
rect 8392 9808 8434 9848
rect 8474 9808 8516 9848
rect 8556 9808 8598 9848
rect 8638 9808 8680 9848
rect 8352 9799 8720 9808
rect 12352 9848 12720 9857
rect 12392 9808 12434 9848
rect 12474 9808 12516 9848
rect 12556 9808 12598 9848
rect 12638 9808 12680 9848
rect 12352 9799 12720 9808
rect 16352 9848 16720 9857
rect 16392 9808 16434 9848
rect 16474 9808 16516 9848
rect 16556 9808 16598 9848
rect 16638 9808 16680 9848
rect 16352 9799 16720 9808
rect 20352 9848 20720 9857
rect 20392 9808 20434 9848
rect 20474 9808 20516 9848
rect 20556 9808 20598 9848
rect 20638 9808 20680 9848
rect 20352 9799 20720 9808
rect 24352 9848 24720 9857
rect 24392 9808 24434 9848
rect 24474 9808 24516 9848
rect 24556 9808 24598 9848
rect 24638 9808 24680 9848
rect 24352 9799 24720 9808
rect 28352 9848 28720 9857
rect 28392 9808 28434 9848
rect 28474 9808 28516 9848
rect 28556 9808 28598 9848
rect 28638 9808 28680 9848
rect 28352 9799 28720 9808
rect 32352 9848 32720 9857
rect 32392 9808 32434 9848
rect 32474 9808 32516 9848
rect 32556 9808 32598 9848
rect 32638 9808 32680 9848
rect 32352 9799 32720 9808
rect 36352 9848 36720 9857
rect 36392 9808 36434 9848
rect 36474 9808 36516 9848
rect 36556 9808 36598 9848
rect 36638 9808 36680 9848
rect 36352 9799 36720 9808
rect 40352 9848 40720 9857
rect 40392 9808 40434 9848
rect 40474 9808 40516 9848
rect 40556 9808 40598 9848
rect 40638 9808 40680 9848
rect 40352 9799 40720 9808
rect 44352 9848 44720 9857
rect 44392 9808 44434 9848
rect 44474 9808 44516 9848
rect 44556 9808 44598 9848
rect 44638 9808 44680 9848
rect 44352 9799 44720 9808
rect 48352 9848 48720 9857
rect 48392 9808 48434 9848
rect 48474 9808 48516 9848
rect 48556 9808 48598 9848
rect 48638 9808 48680 9848
rect 48352 9799 48720 9808
rect 52352 9848 52720 9857
rect 52392 9808 52434 9848
rect 52474 9808 52516 9848
rect 52556 9808 52598 9848
rect 52638 9808 52680 9848
rect 52352 9799 52720 9808
rect 56352 9848 56720 9857
rect 56392 9808 56434 9848
rect 56474 9808 56516 9848
rect 56556 9808 56598 9848
rect 56638 9808 56680 9848
rect 56352 9799 56720 9808
rect 60352 9848 60720 9857
rect 60392 9808 60434 9848
rect 60474 9808 60516 9848
rect 60556 9808 60598 9848
rect 60638 9808 60680 9848
rect 60352 9799 60720 9808
rect 64352 9848 64720 9857
rect 64392 9808 64434 9848
rect 64474 9808 64516 9848
rect 64556 9808 64598 9848
rect 64638 9808 64680 9848
rect 64352 9799 64720 9808
rect 68352 9848 68720 9857
rect 68392 9808 68434 9848
rect 68474 9808 68516 9848
rect 68556 9808 68598 9848
rect 68638 9808 68680 9848
rect 68352 9799 68720 9808
rect 3112 9092 3480 9101
rect 3152 9052 3194 9092
rect 3234 9052 3276 9092
rect 3316 9052 3358 9092
rect 3398 9052 3440 9092
rect 3112 9043 3480 9052
rect 7112 9092 7480 9101
rect 7152 9052 7194 9092
rect 7234 9052 7276 9092
rect 7316 9052 7358 9092
rect 7398 9052 7440 9092
rect 7112 9043 7480 9052
rect 11112 9092 11480 9101
rect 11152 9052 11194 9092
rect 11234 9052 11276 9092
rect 11316 9052 11358 9092
rect 11398 9052 11440 9092
rect 11112 9043 11480 9052
rect 15112 9092 15480 9101
rect 15152 9052 15194 9092
rect 15234 9052 15276 9092
rect 15316 9052 15358 9092
rect 15398 9052 15440 9092
rect 15112 9043 15480 9052
rect 19112 9092 19480 9101
rect 19152 9052 19194 9092
rect 19234 9052 19276 9092
rect 19316 9052 19358 9092
rect 19398 9052 19440 9092
rect 19112 9043 19480 9052
rect 23112 9092 23480 9101
rect 23152 9052 23194 9092
rect 23234 9052 23276 9092
rect 23316 9052 23358 9092
rect 23398 9052 23440 9092
rect 23112 9043 23480 9052
rect 27112 9092 27480 9101
rect 27152 9052 27194 9092
rect 27234 9052 27276 9092
rect 27316 9052 27358 9092
rect 27398 9052 27440 9092
rect 27112 9043 27480 9052
rect 31112 9092 31480 9101
rect 31152 9052 31194 9092
rect 31234 9052 31276 9092
rect 31316 9052 31358 9092
rect 31398 9052 31440 9092
rect 31112 9043 31480 9052
rect 35112 9092 35480 9101
rect 35152 9052 35194 9092
rect 35234 9052 35276 9092
rect 35316 9052 35358 9092
rect 35398 9052 35440 9092
rect 35112 9043 35480 9052
rect 39112 9092 39480 9101
rect 39152 9052 39194 9092
rect 39234 9052 39276 9092
rect 39316 9052 39358 9092
rect 39398 9052 39440 9092
rect 39112 9043 39480 9052
rect 43112 9092 43480 9101
rect 43152 9052 43194 9092
rect 43234 9052 43276 9092
rect 43316 9052 43358 9092
rect 43398 9052 43440 9092
rect 43112 9043 43480 9052
rect 47112 9092 47480 9101
rect 47152 9052 47194 9092
rect 47234 9052 47276 9092
rect 47316 9052 47358 9092
rect 47398 9052 47440 9092
rect 47112 9043 47480 9052
rect 51112 9092 51480 9101
rect 51152 9052 51194 9092
rect 51234 9052 51276 9092
rect 51316 9052 51358 9092
rect 51398 9052 51440 9092
rect 51112 9043 51480 9052
rect 55112 9092 55480 9101
rect 55152 9052 55194 9092
rect 55234 9052 55276 9092
rect 55316 9052 55358 9092
rect 55398 9052 55440 9092
rect 55112 9043 55480 9052
rect 59112 9092 59480 9101
rect 59152 9052 59194 9092
rect 59234 9052 59276 9092
rect 59316 9052 59358 9092
rect 59398 9052 59440 9092
rect 59112 9043 59480 9052
rect 63112 9092 63480 9101
rect 63152 9052 63194 9092
rect 63234 9052 63276 9092
rect 63316 9052 63358 9092
rect 63398 9052 63440 9092
rect 63112 9043 63480 9052
rect 67112 9092 67480 9101
rect 67152 9052 67194 9092
rect 67234 9052 67276 9092
rect 67316 9052 67358 9092
rect 67398 9052 67440 9092
rect 67112 9043 67480 9052
rect 4352 8336 4720 8345
rect 4392 8296 4434 8336
rect 4474 8296 4516 8336
rect 4556 8296 4598 8336
rect 4638 8296 4680 8336
rect 4352 8287 4720 8296
rect 8352 8336 8720 8345
rect 8392 8296 8434 8336
rect 8474 8296 8516 8336
rect 8556 8296 8598 8336
rect 8638 8296 8680 8336
rect 8352 8287 8720 8296
rect 12352 8336 12720 8345
rect 12392 8296 12434 8336
rect 12474 8296 12516 8336
rect 12556 8296 12598 8336
rect 12638 8296 12680 8336
rect 12352 8287 12720 8296
rect 16352 8336 16720 8345
rect 16392 8296 16434 8336
rect 16474 8296 16516 8336
rect 16556 8296 16598 8336
rect 16638 8296 16680 8336
rect 16352 8287 16720 8296
rect 20352 8336 20720 8345
rect 20392 8296 20434 8336
rect 20474 8296 20516 8336
rect 20556 8296 20598 8336
rect 20638 8296 20680 8336
rect 20352 8287 20720 8296
rect 24352 8336 24720 8345
rect 24392 8296 24434 8336
rect 24474 8296 24516 8336
rect 24556 8296 24598 8336
rect 24638 8296 24680 8336
rect 24352 8287 24720 8296
rect 28352 8336 28720 8345
rect 28392 8296 28434 8336
rect 28474 8296 28516 8336
rect 28556 8296 28598 8336
rect 28638 8296 28680 8336
rect 28352 8287 28720 8296
rect 32352 8336 32720 8345
rect 32392 8296 32434 8336
rect 32474 8296 32516 8336
rect 32556 8296 32598 8336
rect 32638 8296 32680 8336
rect 32352 8287 32720 8296
rect 36352 8336 36720 8345
rect 36392 8296 36434 8336
rect 36474 8296 36516 8336
rect 36556 8296 36598 8336
rect 36638 8296 36680 8336
rect 36352 8287 36720 8296
rect 40352 8336 40720 8345
rect 40392 8296 40434 8336
rect 40474 8296 40516 8336
rect 40556 8296 40598 8336
rect 40638 8296 40680 8336
rect 40352 8287 40720 8296
rect 44352 8336 44720 8345
rect 44392 8296 44434 8336
rect 44474 8296 44516 8336
rect 44556 8296 44598 8336
rect 44638 8296 44680 8336
rect 44352 8287 44720 8296
rect 48352 8336 48720 8345
rect 48392 8296 48434 8336
rect 48474 8296 48516 8336
rect 48556 8296 48598 8336
rect 48638 8296 48680 8336
rect 48352 8287 48720 8296
rect 52352 8336 52720 8345
rect 52392 8296 52434 8336
rect 52474 8296 52516 8336
rect 52556 8296 52598 8336
rect 52638 8296 52680 8336
rect 52352 8287 52720 8296
rect 56352 8336 56720 8345
rect 56392 8296 56434 8336
rect 56474 8296 56516 8336
rect 56556 8296 56598 8336
rect 56638 8296 56680 8336
rect 56352 8287 56720 8296
rect 60352 8336 60720 8345
rect 60392 8296 60434 8336
rect 60474 8296 60516 8336
rect 60556 8296 60598 8336
rect 60638 8296 60680 8336
rect 60352 8287 60720 8296
rect 64352 8336 64720 8345
rect 64392 8296 64434 8336
rect 64474 8296 64516 8336
rect 64556 8296 64598 8336
rect 64638 8296 64680 8336
rect 64352 8287 64720 8296
rect 68352 8336 68720 8345
rect 68392 8296 68434 8336
rect 68474 8296 68516 8336
rect 68556 8296 68598 8336
rect 68638 8296 68680 8336
rect 68352 8287 68720 8296
rect 93772 7832 93812 7841
rect 3112 7580 3480 7589
rect 3152 7540 3194 7580
rect 3234 7540 3276 7580
rect 3316 7540 3358 7580
rect 3398 7540 3440 7580
rect 3112 7531 3480 7540
rect 7112 7580 7480 7589
rect 7152 7540 7194 7580
rect 7234 7540 7276 7580
rect 7316 7540 7358 7580
rect 7398 7540 7440 7580
rect 7112 7531 7480 7540
rect 11112 7580 11480 7589
rect 11152 7540 11194 7580
rect 11234 7540 11276 7580
rect 11316 7540 11358 7580
rect 11398 7540 11440 7580
rect 11112 7531 11480 7540
rect 15112 7580 15480 7589
rect 15152 7540 15194 7580
rect 15234 7540 15276 7580
rect 15316 7540 15358 7580
rect 15398 7540 15440 7580
rect 15112 7531 15480 7540
rect 19112 7580 19480 7589
rect 19152 7540 19194 7580
rect 19234 7540 19276 7580
rect 19316 7540 19358 7580
rect 19398 7540 19440 7580
rect 19112 7531 19480 7540
rect 23112 7580 23480 7589
rect 23152 7540 23194 7580
rect 23234 7540 23276 7580
rect 23316 7540 23358 7580
rect 23398 7540 23440 7580
rect 23112 7531 23480 7540
rect 27112 7580 27480 7589
rect 27152 7540 27194 7580
rect 27234 7540 27276 7580
rect 27316 7540 27358 7580
rect 27398 7540 27440 7580
rect 27112 7531 27480 7540
rect 31112 7580 31480 7589
rect 31152 7540 31194 7580
rect 31234 7540 31276 7580
rect 31316 7540 31358 7580
rect 31398 7540 31440 7580
rect 31112 7531 31480 7540
rect 35112 7580 35480 7589
rect 35152 7540 35194 7580
rect 35234 7540 35276 7580
rect 35316 7540 35358 7580
rect 35398 7540 35440 7580
rect 35112 7531 35480 7540
rect 39112 7580 39480 7589
rect 39152 7540 39194 7580
rect 39234 7540 39276 7580
rect 39316 7540 39358 7580
rect 39398 7540 39440 7580
rect 39112 7531 39480 7540
rect 43112 7580 43480 7589
rect 43152 7540 43194 7580
rect 43234 7540 43276 7580
rect 43316 7540 43358 7580
rect 43398 7540 43440 7580
rect 43112 7531 43480 7540
rect 47112 7580 47480 7589
rect 47152 7540 47194 7580
rect 47234 7540 47276 7580
rect 47316 7540 47358 7580
rect 47398 7540 47440 7580
rect 47112 7531 47480 7540
rect 51112 7580 51480 7589
rect 51152 7540 51194 7580
rect 51234 7540 51276 7580
rect 51316 7540 51358 7580
rect 51398 7540 51440 7580
rect 51112 7531 51480 7540
rect 55112 7580 55480 7589
rect 55152 7540 55194 7580
rect 55234 7540 55276 7580
rect 55316 7540 55358 7580
rect 55398 7540 55440 7580
rect 55112 7531 55480 7540
rect 59112 7580 59480 7589
rect 59152 7540 59194 7580
rect 59234 7540 59276 7580
rect 59316 7540 59358 7580
rect 59398 7540 59440 7580
rect 59112 7531 59480 7540
rect 63112 7580 63480 7589
rect 63152 7540 63194 7580
rect 63234 7540 63276 7580
rect 63316 7540 63358 7580
rect 63398 7540 63440 7580
rect 63112 7531 63480 7540
rect 67112 7580 67480 7589
rect 67152 7540 67194 7580
rect 67234 7540 67276 7580
rect 67316 7540 67358 7580
rect 67398 7540 67440 7580
rect 67112 7531 67480 7540
rect 86667 7496 86709 7505
rect 86667 7456 86668 7496
rect 86708 7456 86709 7496
rect 86667 7447 86709 7456
rect 86668 7362 86708 7447
rect 4352 6824 4720 6833
rect 4392 6784 4434 6824
rect 4474 6784 4516 6824
rect 4556 6784 4598 6824
rect 4638 6784 4680 6824
rect 4352 6775 4720 6784
rect 8352 6824 8720 6833
rect 8392 6784 8434 6824
rect 8474 6784 8516 6824
rect 8556 6784 8598 6824
rect 8638 6784 8680 6824
rect 8352 6775 8720 6784
rect 12352 6824 12720 6833
rect 12392 6784 12434 6824
rect 12474 6784 12516 6824
rect 12556 6784 12598 6824
rect 12638 6784 12680 6824
rect 12352 6775 12720 6784
rect 16352 6824 16720 6833
rect 16392 6784 16434 6824
rect 16474 6784 16516 6824
rect 16556 6784 16598 6824
rect 16638 6784 16680 6824
rect 16352 6775 16720 6784
rect 20352 6824 20720 6833
rect 20392 6784 20434 6824
rect 20474 6784 20516 6824
rect 20556 6784 20598 6824
rect 20638 6784 20680 6824
rect 20352 6775 20720 6784
rect 24352 6824 24720 6833
rect 24392 6784 24434 6824
rect 24474 6784 24516 6824
rect 24556 6784 24598 6824
rect 24638 6784 24680 6824
rect 24352 6775 24720 6784
rect 28352 6824 28720 6833
rect 28392 6784 28434 6824
rect 28474 6784 28516 6824
rect 28556 6784 28598 6824
rect 28638 6784 28680 6824
rect 28352 6775 28720 6784
rect 32352 6824 32720 6833
rect 32392 6784 32434 6824
rect 32474 6784 32516 6824
rect 32556 6784 32598 6824
rect 32638 6784 32680 6824
rect 32352 6775 32720 6784
rect 36352 6824 36720 6833
rect 36392 6784 36434 6824
rect 36474 6784 36516 6824
rect 36556 6784 36598 6824
rect 36638 6784 36680 6824
rect 36352 6775 36720 6784
rect 40352 6824 40720 6833
rect 40392 6784 40434 6824
rect 40474 6784 40516 6824
rect 40556 6784 40598 6824
rect 40638 6784 40680 6824
rect 40352 6775 40720 6784
rect 44352 6824 44720 6833
rect 44392 6784 44434 6824
rect 44474 6784 44516 6824
rect 44556 6784 44598 6824
rect 44638 6784 44680 6824
rect 44352 6775 44720 6784
rect 48352 6824 48720 6833
rect 48392 6784 48434 6824
rect 48474 6784 48516 6824
rect 48556 6784 48598 6824
rect 48638 6784 48680 6824
rect 48352 6775 48720 6784
rect 52352 6824 52720 6833
rect 52392 6784 52434 6824
rect 52474 6784 52516 6824
rect 52556 6784 52598 6824
rect 52638 6784 52680 6824
rect 52352 6775 52720 6784
rect 56352 6824 56720 6833
rect 56392 6784 56434 6824
rect 56474 6784 56516 6824
rect 56556 6784 56598 6824
rect 56638 6784 56680 6824
rect 56352 6775 56720 6784
rect 60352 6824 60720 6833
rect 60392 6784 60434 6824
rect 60474 6784 60516 6824
rect 60556 6784 60598 6824
rect 60638 6784 60680 6824
rect 60352 6775 60720 6784
rect 64352 6824 64720 6833
rect 64392 6784 64434 6824
rect 64474 6784 64516 6824
rect 64556 6784 64598 6824
rect 64638 6784 64680 6824
rect 64352 6775 64720 6784
rect 68352 6824 68720 6833
rect 68392 6784 68434 6824
rect 68474 6784 68516 6824
rect 68556 6784 68598 6824
rect 68638 6784 68680 6824
rect 68352 6775 68720 6784
rect 93772 6656 93812 7792
rect 93772 6607 93812 6616
rect 3112 6068 3480 6077
rect 3152 6028 3194 6068
rect 3234 6028 3276 6068
rect 3316 6028 3358 6068
rect 3398 6028 3440 6068
rect 3112 6019 3480 6028
rect 7112 6068 7480 6077
rect 7152 6028 7194 6068
rect 7234 6028 7276 6068
rect 7316 6028 7358 6068
rect 7398 6028 7440 6068
rect 7112 6019 7480 6028
rect 11112 6068 11480 6077
rect 11152 6028 11194 6068
rect 11234 6028 11276 6068
rect 11316 6028 11358 6068
rect 11398 6028 11440 6068
rect 11112 6019 11480 6028
rect 15112 6068 15480 6077
rect 15152 6028 15194 6068
rect 15234 6028 15276 6068
rect 15316 6028 15358 6068
rect 15398 6028 15440 6068
rect 15112 6019 15480 6028
rect 19112 6068 19480 6077
rect 19152 6028 19194 6068
rect 19234 6028 19276 6068
rect 19316 6028 19358 6068
rect 19398 6028 19440 6068
rect 19112 6019 19480 6028
rect 23112 6068 23480 6077
rect 23152 6028 23194 6068
rect 23234 6028 23276 6068
rect 23316 6028 23358 6068
rect 23398 6028 23440 6068
rect 23112 6019 23480 6028
rect 27112 6068 27480 6077
rect 27152 6028 27194 6068
rect 27234 6028 27276 6068
rect 27316 6028 27358 6068
rect 27398 6028 27440 6068
rect 27112 6019 27480 6028
rect 31112 6068 31480 6077
rect 31152 6028 31194 6068
rect 31234 6028 31276 6068
rect 31316 6028 31358 6068
rect 31398 6028 31440 6068
rect 31112 6019 31480 6028
rect 35112 6068 35480 6077
rect 35152 6028 35194 6068
rect 35234 6028 35276 6068
rect 35316 6028 35358 6068
rect 35398 6028 35440 6068
rect 35112 6019 35480 6028
rect 39112 6068 39480 6077
rect 39152 6028 39194 6068
rect 39234 6028 39276 6068
rect 39316 6028 39358 6068
rect 39398 6028 39440 6068
rect 39112 6019 39480 6028
rect 43112 6068 43480 6077
rect 43152 6028 43194 6068
rect 43234 6028 43276 6068
rect 43316 6028 43358 6068
rect 43398 6028 43440 6068
rect 43112 6019 43480 6028
rect 47112 6068 47480 6077
rect 47152 6028 47194 6068
rect 47234 6028 47276 6068
rect 47316 6028 47358 6068
rect 47398 6028 47440 6068
rect 47112 6019 47480 6028
rect 51112 6068 51480 6077
rect 51152 6028 51194 6068
rect 51234 6028 51276 6068
rect 51316 6028 51358 6068
rect 51398 6028 51440 6068
rect 51112 6019 51480 6028
rect 55112 6068 55480 6077
rect 55152 6028 55194 6068
rect 55234 6028 55276 6068
rect 55316 6028 55358 6068
rect 55398 6028 55440 6068
rect 55112 6019 55480 6028
rect 59112 6068 59480 6077
rect 59152 6028 59194 6068
rect 59234 6028 59276 6068
rect 59316 6028 59358 6068
rect 59398 6028 59440 6068
rect 59112 6019 59480 6028
rect 63112 6068 63480 6077
rect 63152 6028 63194 6068
rect 63234 6028 63276 6068
rect 63316 6028 63358 6068
rect 63398 6028 63440 6068
rect 63112 6019 63480 6028
rect 67112 6068 67480 6077
rect 67152 6028 67194 6068
rect 67234 6028 67276 6068
rect 67316 6028 67358 6068
rect 67398 6028 67440 6068
rect 67112 6019 67480 6028
rect 4352 5312 4720 5321
rect 4392 5272 4434 5312
rect 4474 5272 4516 5312
rect 4556 5272 4598 5312
rect 4638 5272 4680 5312
rect 4352 5263 4720 5272
rect 8352 5312 8720 5321
rect 8392 5272 8434 5312
rect 8474 5272 8516 5312
rect 8556 5272 8598 5312
rect 8638 5272 8680 5312
rect 8352 5263 8720 5272
rect 12352 5312 12720 5321
rect 12392 5272 12434 5312
rect 12474 5272 12516 5312
rect 12556 5272 12598 5312
rect 12638 5272 12680 5312
rect 12352 5263 12720 5272
rect 16352 5312 16720 5321
rect 16392 5272 16434 5312
rect 16474 5272 16516 5312
rect 16556 5272 16598 5312
rect 16638 5272 16680 5312
rect 16352 5263 16720 5272
rect 20352 5312 20720 5321
rect 20392 5272 20434 5312
rect 20474 5272 20516 5312
rect 20556 5272 20598 5312
rect 20638 5272 20680 5312
rect 20352 5263 20720 5272
rect 24352 5312 24720 5321
rect 24392 5272 24434 5312
rect 24474 5272 24516 5312
rect 24556 5272 24598 5312
rect 24638 5272 24680 5312
rect 24352 5263 24720 5272
rect 28352 5312 28720 5321
rect 28392 5272 28434 5312
rect 28474 5272 28516 5312
rect 28556 5272 28598 5312
rect 28638 5272 28680 5312
rect 28352 5263 28720 5272
rect 32352 5312 32720 5321
rect 32392 5272 32434 5312
rect 32474 5272 32516 5312
rect 32556 5272 32598 5312
rect 32638 5272 32680 5312
rect 32352 5263 32720 5272
rect 36352 5312 36720 5321
rect 36392 5272 36434 5312
rect 36474 5272 36516 5312
rect 36556 5272 36598 5312
rect 36638 5272 36680 5312
rect 36352 5263 36720 5272
rect 40352 5312 40720 5321
rect 40392 5272 40434 5312
rect 40474 5272 40516 5312
rect 40556 5272 40598 5312
rect 40638 5272 40680 5312
rect 40352 5263 40720 5272
rect 44352 5312 44720 5321
rect 44392 5272 44434 5312
rect 44474 5272 44516 5312
rect 44556 5272 44598 5312
rect 44638 5272 44680 5312
rect 44352 5263 44720 5272
rect 48352 5312 48720 5321
rect 48392 5272 48434 5312
rect 48474 5272 48516 5312
rect 48556 5272 48598 5312
rect 48638 5272 48680 5312
rect 48352 5263 48720 5272
rect 52352 5312 52720 5321
rect 52392 5272 52434 5312
rect 52474 5272 52516 5312
rect 52556 5272 52598 5312
rect 52638 5272 52680 5312
rect 52352 5263 52720 5272
rect 56352 5312 56720 5321
rect 56392 5272 56434 5312
rect 56474 5272 56516 5312
rect 56556 5272 56598 5312
rect 56638 5272 56680 5312
rect 56352 5263 56720 5272
rect 60352 5312 60720 5321
rect 60392 5272 60434 5312
rect 60474 5272 60516 5312
rect 60556 5272 60598 5312
rect 60638 5272 60680 5312
rect 60352 5263 60720 5272
rect 64352 5312 64720 5321
rect 64392 5272 64434 5312
rect 64474 5272 64516 5312
rect 64556 5272 64598 5312
rect 64638 5272 64680 5312
rect 64352 5263 64720 5272
rect 68352 5312 68720 5321
rect 68392 5272 68434 5312
rect 68474 5272 68516 5312
rect 68556 5272 68598 5312
rect 68638 5272 68680 5312
rect 68352 5263 68720 5272
rect 72352 5312 72720 5321
rect 72392 5272 72434 5312
rect 72474 5272 72516 5312
rect 72556 5272 72598 5312
rect 72638 5272 72680 5312
rect 72352 5263 72720 5272
rect 76352 5312 76720 5321
rect 76392 5272 76434 5312
rect 76474 5272 76516 5312
rect 76556 5272 76598 5312
rect 76638 5272 76680 5312
rect 76352 5263 76720 5272
rect 80352 5312 80720 5321
rect 80392 5272 80434 5312
rect 80474 5272 80516 5312
rect 80556 5272 80598 5312
rect 80638 5272 80680 5312
rect 80352 5263 80720 5272
rect 84352 5312 84720 5321
rect 84392 5272 84434 5312
rect 84474 5272 84516 5312
rect 84556 5272 84598 5312
rect 84638 5272 84680 5312
rect 84352 5263 84720 5272
rect 88352 5312 88720 5321
rect 88392 5272 88434 5312
rect 88474 5272 88516 5312
rect 88556 5272 88598 5312
rect 88638 5272 88680 5312
rect 88352 5263 88720 5272
rect 92352 5312 92720 5321
rect 92392 5272 92434 5312
rect 92474 5272 92516 5312
rect 92556 5272 92598 5312
rect 92638 5272 92680 5312
rect 92352 5263 92720 5272
rect 96352 5312 96720 5321
rect 96392 5272 96434 5312
rect 96474 5272 96516 5312
rect 96556 5272 96598 5312
rect 96638 5272 96680 5312
rect 96352 5263 96720 5272
rect 3112 4556 3480 4565
rect 3152 4516 3194 4556
rect 3234 4516 3276 4556
rect 3316 4516 3358 4556
rect 3398 4516 3440 4556
rect 3112 4507 3480 4516
rect 7112 4556 7480 4565
rect 7152 4516 7194 4556
rect 7234 4516 7276 4556
rect 7316 4516 7358 4556
rect 7398 4516 7440 4556
rect 7112 4507 7480 4516
rect 11112 4556 11480 4565
rect 11152 4516 11194 4556
rect 11234 4516 11276 4556
rect 11316 4516 11358 4556
rect 11398 4516 11440 4556
rect 11112 4507 11480 4516
rect 15112 4556 15480 4565
rect 15152 4516 15194 4556
rect 15234 4516 15276 4556
rect 15316 4516 15358 4556
rect 15398 4516 15440 4556
rect 15112 4507 15480 4516
rect 19112 4556 19480 4565
rect 19152 4516 19194 4556
rect 19234 4516 19276 4556
rect 19316 4516 19358 4556
rect 19398 4516 19440 4556
rect 19112 4507 19480 4516
rect 23112 4556 23480 4565
rect 23152 4516 23194 4556
rect 23234 4516 23276 4556
rect 23316 4516 23358 4556
rect 23398 4516 23440 4556
rect 23112 4507 23480 4516
rect 27112 4556 27480 4565
rect 27152 4516 27194 4556
rect 27234 4516 27276 4556
rect 27316 4516 27358 4556
rect 27398 4516 27440 4556
rect 27112 4507 27480 4516
rect 31112 4556 31480 4565
rect 31152 4516 31194 4556
rect 31234 4516 31276 4556
rect 31316 4516 31358 4556
rect 31398 4516 31440 4556
rect 31112 4507 31480 4516
rect 35112 4556 35480 4565
rect 35152 4516 35194 4556
rect 35234 4516 35276 4556
rect 35316 4516 35358 4556
rect 35398 4516 35440 4556
rect 35112 4507 35480 4516
rect 39112 4556 39480 4565
rect 39152 4516 39194 4556
rect 39234 4516 39276 4556
rect 39316 4516 39358 4556
rect 39398 4516 39440 4556
rect 39112 4507 39480 4516
rect 43112 4556 43480 4565
rect 43152 4516 43194 4556
rect 43234 4516 43276 4556
rect 43316 4516 43358 4556
rect 43398 4516 43440 4556
rect 43112 4507 43480 4516
rect 47112 4556 47480 4565
rect 47152 4516 47194 4556
rect 47234 4516 47276 4556
rect 47316 4516 47358 4556
rect 47398 4516 47440 4556
rect 47112 4507 47480 4516
rect 51112 4556 51480 4565
rect 51152 4516 51194 4556
rect 51234 4516 51276 4556
rect 51316 4516 51358 4556
rect 51398 4516 51440 4556
rect 51112 4507 51480 4516
rect 55112 4556 55480 4565
rect 55152 4516 55194 4556
rect 55234 4516 55276 4556
rect 55316 4516 55358 4556
rect 55398 4516 55440 4556
rect 55112 4507 55480 4516
rect 59112 4556 59480 4565
rect 59152 4516 59194 4556
rect 59234 4516 59276 4556
rect 59316 4516 59358 4556
rect 59398 4516 59440 4556
rect 59112 4507 59480 4516
rect 63112 4556 63480 4565
rect 63152 4516 63194 4556
rect 63234 4516 63276 4556
rect 63316 4516 63358 4556
rect 63398 4516 63440 4556
rect 63112 4507 63480 4516
rect 67112 4556 67480 4565
rect 67152 4516 67194 4556
rect 67234 4516 67276 4556
rect 67316 4516 67358 4556
rect 67398 4516 67440 4556
rect 67112 4507 67480 4516
rect 71112 4556 71480 4565
rect 71152 4516 71194 4556
rect 71234 4516 71276 4556
rect 71316 4516 71358 4556
rect 71398 4516 71440 4556
rect 71112 4507 71480 4516
rect 75112 4556 75480 4565
rect 75152 4516 75194 4556
rect 75234 4516 75276 4556
rect 75316 4516 75358 4556
rect 75398 4516 75440 4556
rect 75112 4507 75480 4516
rect 79112 4556 79480 4565
rect 79152 4516 79194 4556
rect 79234 4516 79276 4556
rect 79316 4516 79358 4556
rect 79398 4516 79440 4556
rect 79112 4507 79480 4516
rect 83112 4556 83480 4565
rect 83152 4516 83194 4556
rect 83234 4516 83276 4556
rect 83316 4516 83358 4556
rect 83398 4516 83440 4556
rect 83112 4507 83480 4516
rect 87112 4556 87480 4565
rect 87152 4516 87194 4556
rect 87234 4516 87276 4556
rect 87316 4516 87358 4556
rect 87398 4516 87440 4556
rect 87112 4507 87480 4516
rect 91112 4556 91480 4565
rect 91152 4516 91194 4556
rect 91234 4516 91276 4556
rect 91316 4516 91358 4556
rect 91398 4516 91440 4556
rect 91112 4507 91480 4516
rect 95112 4556 95480 4565
rect 95152 4516 95194 4556
rect 95234 4516 95276 4556
rect 95316 4516 95358 4556
rect 95398 4516 95440 4556
rect 95112 4507 95480 4516
rect 99112 4556 99480 4565
rect 99152 4516 99194 4556
rect 99234 4516 99276 4556
rect 99316 4516 99358 4556
rect 99398 4516 99440 4556
rect 99112 4507 99480 4516
rect 4352 3800 4720 3809
rect 4392 3760 4434 3800
rect 4474 3760 4516 3800
rect 4556 3760 4598 3800
rect 4638 3760 4680 3800
rect 4352 3751 4720 3760
rect 8352 3800 8720 3809
rect 8392 3760 8434 3800
rect 8474 3760 8516 3800
rect 8556 3760 8598 3800
rect 8638 3760 8680 3800
rect 8352 3751 8720 3760
rect 12352 3800 12720 3809
rect 12392 3760 12434 3800
rect 12474 3760 12516 3800
rect 12556 3760 12598 3800
rect 12638 3760 12680 3800
rect 12352 3751 12720 3760
rect 16352 3800 16720 3809
rect 16392 3760 16434 3800
rect 16474 3760 16516 3800
rect 16556 3760 16598 3800
rect 16638 3760 16680 3800
rect 16352 3751 16720 3760
rect 20352 3800 20720 3809
rect 20392 3760 20434 3800
rect 20474 3760 20516 3800
rect 20556 3760 20598 3800
rect 20638 3760 20680 3800
rect 20352 3751 20720 3760
rect 24352 3800 24720 3809
rect 24392 3760 24434 3800
rect 24474 3760 24516 3800
rect 24556 3760 24598 3800
rect 24638 3760 24680 3800
rect 24352 3751 24720 3760
rect 28352 3800 28720 3809
rect 28392 3760 28434 3800
rect 28474 3760 28516 3800
rect 28556 3760 28598 3800
rect 28638 3760 28680 3800
rect 28352 3751 28720 3760
rect 32352 3800 32720 3809
rect 32392 3760 32434 3800
rect 32474 3760 32516 3800
rect 32556 3760 32598 3800
rect 32638 3760 32680 3800
rect 32352 3751 32720 3760
rect 36352 3800 36720 3809
rect 36392 3760 36434 3800
rect 36474 3760 36516 3800
rect 36556 3760 36598 3800
rect 36638 3760 36680 3800
rect 36352 3751 36720 3760
rect 40352 3800 40720 3809
rect 40392 3760 40434 3800
rect 40474 3760 40516 3800
rect 40556 3760 40598 3800
rect 40638 3760 40680 3800
rect 40352 3751 40720 3760
rect 44352 3800 44720 3809
rect 44392 3760 44434 3800
rect 44474 3760 44516 3800
rect 44556 3760 44598 3800
rect 44638 3760 44680 3800
rect 44352 3751 44720 3760
rect 48352 3800 48720 3809
rect 48392 3760 48434 3800
rect 48474 3760 48516 3800
rect 48556 3760 48598 3800
rect 48638 3760 48680 3800
rect 48352 3751 48720 3760
rect 52352 3800 52720 3809
rect 52392 3760 52434 3800
rect 52474 3760 52516 3800
rect 52556 3760 52598 3800
rect 52638 3760 52680 3800
rect 52352 3751 52720 3760
rect 56352 3800 56720 3809
rect 56392 3760 56434 3800
rect 56474 3760 56516 3800
rect 56556 3760 56598 3800
rect 56638 3760 56680 3800
rect 56352 3751 56720 3760
rect 60352 3800 60720 3809
rect 60392 3760 60434 3800
rect 60474 3760 60516 3800
rect 60556 3760 60598 3800
rect 60638 3760 60680 3800
rect 60352 3751 60720 3760
rect 64352 3800 64720 3809
rect 64392 3760 64434 3800
rect 64474 3760 64516 3800
rect 64556 3760 64598 3800
rect 64638 3760 64680 3800
rect 64352 3751 64720 3760
rect 68352 3800 68720 3809
rect 68392 3760 68434 3800
rect 68474 3760 68516 3800
rect 68556 3760 68598 3800
rect 68638 3760 68680 3800
rect 68352 3751 68720 3760
rect 72352 3800 72720 3809
rect 72392 3760 72434 3800
rect 72474 3760 72516 3800
rect 72556 3760 72598 3800
rect 72638 3760 72680 3800
rect 72352 3751 72720 3760
rect 76352 3800 76720 3809
rect 76392 3760 76434 3800
rect 76474 3760 76516 3800
rect 76556 3760 76598 3800
rect 76638 3760 76680 3800
rect 76352 3751 76720 3760
rect 80352 3800 80720 3809
rect 80392 3760 80434 3800
rect 80474 3760 80516 3800
rect 80556 3760 80598 3800
rect 80638 3760 80680 3800
rect 80352 3751 80720 3760
rect 84352 3800 84720 3809
rect 84392 3760 84434 3800
rect 84474 3760 84516 3800
rect 84556 3760 84598 3800
rect 84638 3760 84680 3800
rect 84352 3751 84720 3760
rect 88352 3800 88720 3809
rect 88392 3760 88434 3800
rect 88474 3760 88516 3800
rect 88556 3760 88598 3800
rect 88638 3760 88680 3800
rect 88352 3751 88720 3760
rect 92352 3800 92720 3809
rect 92392 3760 92434 3800
rect 92474 3760 92516 3800
rect 92556 3760 92598 3800
rect 92638 3760 92680 3800
rect 92352 3751 92720 3760
rect 96352 3800 96720 3809
rect 96392 3760 96434 3800
rect 96474 3760 96516 3800
rect 96556 3760 96598 3800
rect 96638 3760 96680 3800
rect 96352 3751 96720 3760
rect 3112 3044 3480 3053
rect 3152 3004 3194 3044
rect 3234 3004 3276 3044
rect 3316 3004 3358 3044
rect 3398 3004 3440 3044
rect 3112 2995 3480 3004
rect 7112 3044 7480 3053
rect 7152 3004 7194 3044
rect 7234 3004 7276 3044
rect 7316 3004 7358 3044
rect 7398 3004 7440 3044
rect 7112 2995 7480 3004
rect 11112 3044 11480 3053
rect 11152 3004 11194 3044
rect 11234 3004 11276 3044
rect 11316 3004 11358 3044
rect 11398 3004 11440 3044
rect 11112 2995 11480 3004
rect 15112 3044 15480 3053
rect 15152 3004 15194 3044
rect 15234 3004 15276 3044
rect 15316 3004 15358 3044
rect 15398 3004 15440 3044
rect 15112 2995 15480 3004
rect 19112 3044 19480 3053
rect 19152 3004 19194 3044
rect 19234 3004 19276 3044
rect 19316 3004 19358 3044
rect 19398 3004 19440 3044
rect 19112 2995 19480 3004
rect 23112 3044 23480 3053
rect 23152 3004 23194 3044
rect 23234 3004 23276 3044
rect 23316 3004 23358 3044
rect 23398 3004 23440 3044
rect 23112 2995 23480 3004
rect 27112 3044 27480 3053
rect 27152 3004 27194 3044
rect 27234 3004 27276 3044
rect 27316 3004 27358 3044
rect 27398 3004 27440 3044
rect 27112 2995 27480 3004
rect 31112 3044 31480 3053
rect 31152 3004 31194 3044
rect 31234 3004 31276 3044
rect 31316 3004 31358 3044
rect 31398 3004 31440 3044
rect 31112 2995 31480 3004
rect 35112 3044 35480 3053
rect 35152 3004 35194 3044
rect 35234 3004 35276 3044
rect 35316 3004 35358 3044
rect 35398 3004 35440 3044
rect 35112 2995 35480 3004
rect 39112 3044 39480 3053
rect 39152 3004 39194 3044
rect 39234 3004 39276 3044
rect 39316 3004 39358 3044
rect 39398 3004 39440 3044
rect 39112 2995 39480 3004
rect 43112 3044 43480 3053
rect 43152 3004 43194 3044
rect 43234 3004 43276 3044
rect 43316 3004 43358 3044
rect 43398 3004 43440 3044
rect 43112 2995 43480 3004
rect 47112 3044 47480 3053
rect 47152 3004 47194 3044
rect 47234 3004 47276 3044
rect 47316 3004 47358 3044
rect 47398 3004 47440 3044
rect 47112 2995 47480 3004
rect 51112 3044 51480 3053
rect 51152 3004 51194 3044
rect 51234 3004 51276 3044
rect 51316 3004 51358 3044
rect 51398 3004 51440 3044
rect 51112 2995 51480 3004
rect 55112 3044 55480 3053
rect 55152 3004 55194 3044
rect 55234 3004 55276 3044
rect 55316 3004 55358 3044
rect 55398 3004 55440 3044
rect 55112 2995 55480 3004
rect 59112 3044 59480 3053
rect 59152 3004 59194 3044
rect 59234 3004 59276 3044
rect 59316 3004 59358 3044
rect 59398 3004 59440 3044
rect 59112 2995 59480 3004
rect 63112 3044 63480 3053
rect 63152 3004 63194 3044
rect 63234 3004 63276 3044
rect 63316 3004 63358 3044
rect 63398 3004 63440 3044
rect 63112 2995 63480 3004
rect 67112 3044 67480 3053
rect 67152 3004 67194 3044
rect 67234 3004 67276 3044
rect 67316 3004 67358 3044
rect 67398 3004 67440 3044
rect 67112 2995 67480 3004
rect 71112 3044 71480 3053
rect 71152 3004 71194 3044
rect 71234 3004 71276 3044
rect 71316 3004 71358 3044
rect 71398 3004 71440 3044
rect 71112 2995 71480 3004
rect 75112 3044 75480 3053
rect 75152 3004 75194 3044
rect 75234 3004 75276 3044
rect 75316 3004 75358 3044
rect 75398 3004 75440 3044
rect 75112 2995 75480 3004
rect 79112 3044 79480 3053
rect 79152 3004 79194 3044
rect 79234 3004 79276 3044
rect 79316 3004 79358 3044
rect 79398 3004 79440 3044
rect 79112 2995 79480 3004
rect 83112 3044 83480 3053
rect 83152 3004 83194 3044
rect 83234 3004 83276 3044
rect 83316 3004 83358 3044
rect 83398 3004 83440 3044
rect 83112 2995 83480 3004
rect 87112 3044 87480 3053
rect 87152 3004 87194 3044
rect 87234 3004 87276 3044
rect 87316 3004 87358 3044
rect 87398 3004 87440 3044
rect 87112 2995 87480 3004
rect 91112 3044 91480 3053
rect 91152 3004 91194 3044
rect 91234 3004 91276 3044
rect 91316 3004 91358 3044
rect 91398 3004 91440 3044
rect 91112 2995 91480 3004
rect 95112 3044 95480 3053
rect 95152 3004 95194 3044
rect 95234 3004 95276 3044
rect 95316 3004 95358 3044
rect 95398 3004 95440 3044
rect 95112 2995 95480 3004
rect 99112 3044 99480 3053
rect 99152 3004 99194 3044
rect 99234 3004 99276 3044
rect 99316 3004 99358 3044
rect 99398 3004 99440 3044
rect 99112 2995 99480 3004
rect 4352 2288 4720 2297
rect 4392 2248 4434 2288
rect 4474 2248 4516 2288
rect 4556 2248 4598 2288
rect 4638 2248 4680 2288
rect 4352 2239 4720 2248
rect 8352 2288 8720 2297
rect 8392 2248 8434 2288
rect 8474 2248 8516 2288
rect 8556 2248 8598 2288
rect 8638 2248 8680 2288
rect 8352 2239 8720 2248
rect 12352 2288 12720 2297
rect 12392 2248 12434 2288
rect 12474 2248 12516 2288
rect 12556 2248 12598 2288
rect 12638 2248 12680 2288
rect 12352 2239 12720 2248
rect 16352 2288 16720 2297
rect 16392 2248 16434 2288
rect 16474 2248 16516 2288
rect 16556 2248 16598 2288
rect 16638 2248 16680 2288
rect 16352 2239 16720 2248
rect 20352 2288 20720 2297
rect 20392 2248 20434 2288
rect 20474 2248 20516 2288
rect 20556 2248 20598 2288
rect 20638 2248 20680 2288
rect 20352 2239 20720 2248
rect 24352 2288 24720 2297
rect 24392 2248 24434 2288
rect 24474 2248 24516 2288
rect 24556 2248 24598 2288
rect 24638 2248 24680 2288
rect 24352 2239 24720 2248
rect 28352 2288 28720 2297
rect 28392 2248 28434 2288
rect 28474 2248 28516 2288
rect 28556 2248 28598 2288
rect 28638 2248 28680 2288
rect 28352 2239 28720 2248
rect 32352 2288 32720 2297
rect 32392 2248 32434 2288
rect 32474 2248 32516 2288
rect 32556 2248 32598 2288
rect 32638 2248 32680 2288
rect 32352 2239 32720 2248
rect 36352 2288 36720 2297
rect 36392 2248 36434 2288
rect 36474 2248 36516 2288
rect 36556 2248 36598 2288
rect 36638 2248 36680 2288
rect 36352 2239 36720 2248
rect 40352 2288 40720 2297
rect 40392 2248 40434 2288
rect 40474 2248 40516 2288
rect 40556 2248 40598 2288
rect 40638 2248 40680 2288
rect 40352 2239 40720 2248
rect 44352 2288 44720 2297
rect 44392 2248 44434 2288
rect 44474 2248 44516 2288
rect 44556 2248 44598 2288
rect 44638 2248 44680 2288
rect 44352 2239 44720 2248
rect 48352 2288 48720 2297
rect 48392 2248 48434 2288
rect 48474 2248 48516 2288
rect 48556 2248 48598 2288
rect 48638 2248 48680 2288
rect 48352 2239 48720 2248
rect 52352 2288 52720 2297
rect 52392 2248 52434 2288
rect 52474 2248 52516 2288
rect 52556 2248 52598 2288
rect 52638 2248 52680 2288
rect 52352 2239 52720 2248
rect 56352 2288 56720 2297
rect 56392 2248 56434 2288
rect 56474 2248 56516 2288
rect 56556 2248 56598 2288
rect 56638 2248 56680 2288
rect 56352 2239 56720 2248
rect 60352 2288 60720 2297
rect 60392 2248 60434 2288
rect 60474 2248 60516 2288
rect 60556 2248 60598 2288
rect 60638 2248 60680 2288
rect 60352 2239 60720 2248
rect 64352 2288 64720 2297
rect 64392 2248 64434 2288
rect 64474 2248 64516 2288
rect 64556 2248 64598 2288
rect 64638 2248 64680 2288
rect 64352 2239 64720 2248
rect 68352 2288 68720 2297
rect 68392 2248 68434 2288
rect 68474 2248 68516 2288
rect 68556 2248 68598 2288
rect 68638 2248 68680 2288
rect 68352 2239 68720 2248
rect 72352 2288 72720 2297
rect 72392 2248 72434 2288
rect 72474 2248 72516 2288
rect 72556 2248 72598 2288
rect 72638 2248 72680 2288
rect 72352 2239 72720 2248
rect 76352 2288 76720 2297
rect 76392 2248 76434 2288
rect 76474 2248 76516 2288
rect 76556 2248 76598 2288
rect 76638 2248 76680 2288
rect 76352 2239 76720 2248
rect 80352 2288 80720 2297
rect 80392 2248 80434 2288
rect 80474 2248 80516 2288
rect 80556 2248 80598 2288
rect 80638 2248 80680 2288
rect 80352 2239 80720 2248
rect 84352 2288 84720 2297
rect 84392 2248 84434 2288
rect 84474 2248 84516 2288
rect 84556 2248 84598 2288
rect 84638 2248 84680 2288
rect 84352 2239 84720 2248
rect 88352 2288 88720 2297
rect 88392 2248 88434 2288
rect 88474 2248 88516 2288
rect 88556 2248 88598 2288
rect 88638 2248 88680 2288
rect 88352 2239 88720 2248
rect 92352 2288 92720 2297
rect 92392 2248 92434 2288
rect 92474 2248 92516 2288
rect 92556 2248 92598 2288
rect 92638 2248 92680 2288
rect 92352 2239 92720 2248
rect 96352 2288 96720 2297
rect 96392 2248 96434 2288
rect 96474 2248 96516 2288
rect 96556 2248 96598 2288
rect 96638 2248 96680 2288
rect 96352 2239 96720 2248
rect 3112 1532 3480 1541
rect 3152 1492 3194 1532
rect 3234 1492 3276 1532
rect 3316 1492 3358 1532
rect 3398 1492 3440 1532
rect 3112 1483 3480 1492
rect 7112 1532 7480 1541
rect 7152 1492 7194 1532
rect 7234 1492 7276 1532
rect 7316 1492 7358 1532
rect 7398 1492 7440 1532
rect 7112 1483 7480 1492
rect 11112 1532 11480 1541
rect 11152 1492 11194 1532
rect 11234 1492 11276 1532
rect 11316 1492 11358 1532
rect 11398 1492 11440 1532
rect 11112 1483 11480 1492
rect 15112 1532 15480 1541
rect 15152 1492 15194 1532
rect 15234 1492 15276 1532
rect 15316 1492 15358 1532
rect 15398 1492 15440 1532
rect 15112 1483 15480 1492
rect 19112 1532 19480 1541
rect 19152 1492 19194 1532
rect 19234 1492 19276 1532
rect 19316 1492 19358 1532
rect 19398 1492 19440 1532
rect 19112 1483 19480 1492
rect 23112 1532 23480 1541
rect 23152 1492 23194 1532
rect 23234 1492 23276 1532
rect 23316 1492 23358 1532
rect 23398 1492 23440 1532
rect 23112 1483 23480 1492
rect 27112 1532 27480 1541
rect 27152 1492 27194 1532
rect 27234 1492 27276 1532
rect 27316 1492 27358 1532
rect 27398 1492 27440 1532
rect 27112 1483 27480 1492
rect 31112 1532 31480 1541
rect 31152 1492 31194 1532
rect 31234 1492 31276 1532
rect 31316 1492 31358 1532
rect 31398 1492 31440 1532
rect 31112 1483 31480 1492
rect 35112 1532 35480 1541
rect 35152 1492 35194 1532
rect 35234 1492 35276 1532
rect 35316 1492 35358 1532
rect 35398 1492 35440 1532
rect 35112 1483 35480 1492
rect 39112 1532 39480 1541
rect 39152 1492 39194 1532
rect 39234 1492 39276 1532
rect 39316 1492 39358 1532
rect 39398 1492 39440 1532
rect 39112 1483 39480 1492
rect 43112 1532 43480 1541
rect 43152 1492 43194 1532
rect 43234 1492 43276 1532
rect 43316 1492 43358 1532
rect 43398 1492 43440 1532
rect 43112 1483 43480 1492
rect 47112 1532 47480 1541
rect 47152 1492 47194 1532
rect 47234 1492 47276 1532
rect 47316 1492 47358 1532
rect 47398 1492 47440 1532
rect 47112 1483 47480 1492
rect 51112 1532 51480 1541
rect 51152 1492 51194 1532
rect 51234 1492 51276 1532
rect 51316 1492 51358 1532
rect 51398 1492 51440 1532
rect 51112 1483 51480 1492
rect 55112 1532 55480 1541
rect 55152 1492 55194 1532
rect 55234 1492 55276 1532
rect 55316 1492 55358 1532
rect 55398 1492 55440 1532
rect 55112 1483 55480 1492
rect 59112 1532 59480 1541
rect 59152 1492 59194 1532
rect 59234 1492 59276 1532
rect 59316 1492 59358 1532
rect 59398 1492 59440 1532
rect 59112 1483 59480 1492
rect 63112 1532 63480 1541
rect 63152 1492 63194 1532
rect 63234 1492 63276 1532
rect 63316 1492 63358 1532
rect 63398 1492 63440 1532
rect 63112 1483 63480 1492
rect 67112 1532 67480 1541
rect 67152 1492 67194 1532
rect 67234 1492 67276 1532
rect 67316 1492 67358 1532
rect 67398 1492 67440 1532
rect 67112 1483 67480 1492
rect 71112 1532 71480 1541
rect 71152 1492 71194 1532
rect 71234 1492 71276 1532
rect 71316 1492 71358 1532
rect 71398 1492 71440 1532
rect 71112 1483 71480 1492
rect 75112 1532 75480 1541
rect 75152 1492 75194 1532
rect 75234 1492 75276 1532
rect 75316 1492 75358 1532
rect 75398 1492 75440 1532
rect 75112 1483 75480 1492
rect 79112 1532 79480 1541
rect 79152 1492 79194 1532
rect 79234 1492 79276 1532
rect 79316 1492 79358 1532
rect 79398 1492 79440 1532
rect 79112 1483 79480 1492
rect 83112 1532 83480 1541
rect 83152 1492 83194 1532
rect 83234 1492 83276 1532
rect 83316 1492 83358 1532
rect 83398 1492 83440 1532
rect 83112 1483 83480 1492
rect 87112 1532 87480 1541
rect 87152 1492 87194 1532
rect 87234 1492 87276 1532
rect 87316 1492 87358 1532
rect 87398 1492 87440 1532
rect 87112 1483 87480 1492
rect 91112 1532 91480 1541
rect 91152 1492 91194 1532
rect 91234 1492 91276 1532
rect 91316 1492 91358 1532
rect 91398 1492 91440 1532
rect 91112 1483 91480 1492
rect 95112 1532 95480 1541
rect 95152 1492 95194 1532
rect 95234 1492 95276 1532
rect 95316 1492 95358 1532
rect 95398 1492 95440 1532
rect 95112 1483 95480 1492
rect 99112 1532 99480 1541
rect 99152 1492 99194 1532
rect 99234 1492 99276 1532
rect 99316 1492 99358 1532
rect 99398 1492 99440 1532
rect 99112 1483 99480 1492
rect 4352 776 4720 785
rect 4392 736 4434 776
rect 4474 736 4516 776
rect 4556 736 4598 776
rect 4638 736 4680 776
rect 4352 727 4720 736
rect 8352 776 8720 785
rect 8392 736 8434 776
rect 8474 736 8516 776
rect 8556 736 8598 776
rect 8638 736 8680 776
rect 8352 727 8720 736
rect 12352 776 12720 785
rect 12392 736 12434 776
rect 12474 736 12516 776
rect 12556 736 12598 776
rect 12638 736 12680 776
rect 12352 727 12720 736
rect 16352 776 16720 785
rect 16392 736 16434 776
rect 16474 736 16516 776
rect 16556 736 16598 776
rect 16638 736 16680 776
rect 16352 727 16720 736
rect 20352 776 20720 785
rect 20392 736 20434 776
rect 20474 736 20516 776
rect 20556 736 20598 776
rect 20638 736 20680 776
rect 20352 727 20720 736
rect 24352 776 24720 785
rect 24392 736 24434 776
rect 24474 736 24516 776
rect 24556 736 24598 776
rect 24638 736 24680 776
rect 24352 727 24720 736
rect 28352 776 28720 785
rect 28392 736 28434 776
rect 28474 736 28516 776
rect 28556 736 28598 776
rect 28638 736 28680 776
rect 28352 727 28720 736
rect 32352 776 32720 785
rect 32392 736 32434 776
rect 32474 736 32516 776
rect 32556 736 32598 776
rect 32638 736 32680 776
rect 32352 727 32720 736
rect 36352 776 36720 785
rect 36392 736 36434 776
rect 36474 736 36516 776
rect 36556 736 36598 776
rect 36638 736 36680 776
rect 36352 727 36720 736
rect 40352 776 40720 785
rect 40392 736 40434 776
rect 40474 736 40516 776
rect 40556 736 40598 776
rect 40638 736 40680 776
rect 40352 727 40720 736
rect 44352 776 44720 785
rect 44392 736 44434 776
rect 44474 736 44516 776
rect 44556 736 44598 776
rect 44638 736 44680 776
rect 44352 727 44720 736
rect 48352 776 48720 785
rect 48392 736 48434 776
rect 48474 736 48516 776
rect 48556 736 48598 776
rect 48638 736 48680 776
rect 48352 727 48720 736
rect 52352 776 52720 785
rect 52392 736 52434 776
rect 52474 736 52516 776
rect 52556 736 52598 776
rect 52638 736 52680 776
rect 52352 727 52720 736
rect 56352 776 56720 785
rect 56392 736 56434 776
rect 56474 736 56516 776
rect 56556 736 56598 776
rect 56638 736 56680 776
rect 56352 727 56720 736
rect 60352 776 60720 785
rect 60392 736 60434 776
rect 60474 736 60516 776
rect 60556 736 60598 776
rect 60638 736 60680 776
rect 60352 727 60720 736
rect 64352 776 64720 785
rect 64392 736 64434 776
rect 64474 736 64516 776
rect 64556 736 64598 776
rect 64638 736 64680 776
rect 64352 727 64720 736
rect 68352 776 68720 785
rect 68392 736 68434 776
rect 68474 736 68516 776
rect 68556 736 68598 776
rect 68638 736 68680 776
rect 68352 727 68720 736
rect 72352 776 72720 785
rect 72392 736 72434 776
rect 72474 736 72516 776
rect 72556 736 72598 776
rect 72638 736 72680 776
rect 72352 727 72720 736
rect 76352 776 76720 785
rect 76392 736 76434 776
rect 76474 736 76516 776
rect 76556 736 76598 776
rect 76638 736 76680 776
rect 76352 727 76720 736
rect 80352 776 80720 785
rect 80392 736 80434 776
rect 80474 736 80516 776
rect 80556 736 80598 776
rect 80638 736 80680 776
rect 80352 727 80720 736
rect 84352 776 84720 785
rect 84392 736 84434 776
rect 84474 736 84516 776
rect 84556 736 84598 776
rect 84638 736 84680 776
rect 84352 727 84720 736
rect 88352 776 88720 785
rect 88392 736 88434 776
rect 88474 736 88516 776
rect 88556 736 88598 776
rect 88638 736 88680 776
rect 88352 727 88720 736
rect 92352 776 92720 785
rect 92392 736 92434 776
rect 92474 736 92516 776
rect 92556 736 92598 776
rect 92638 736 92680 776
rect 92352 727 92720 736
rect 96352 776 96720 785
rect 96392 736 96434 776
rect 96474 736 96516 776
rect 96556 736 96598 776
rect 96638 736 96680 776
rect 96352 727 96720 736
<< via4 >>
rect 4352 38536 4392 38576
rect 4434 38536 4474 38576
rect 4516 38536 4556 38576
rect 4598 38536 4638 38576
rect 4680 38536 4720 38576
rect 8352 38536 8392 38576
rect 8434 38536 8474 38576
rect 8516 38536 8556 38576
rect 8598 38536 8638 38576
rect 8680 38536 8720 38576
rect 12352 38536 12392 38576
rect 12434 38536 12474 38576
rect 12516 38536 12556 38576
rect 12598 38536 12638 38576
rect 12680 38536 12720 38576
rect 16352 38536 16392 38576
rect 16434 38536 16474 38576
rect 16516 38536 16556 38576
rect 16598 38536 16638 38576
rect 16680 38536 16720 38576
rect 20352 38536 20392 38576
rect 20434 38536 20474 38576
rect 20516 38536 20556 38576
rect 20598 38536 20638 38576
rect 20680 38536 20720 38576
rect 24352 38536 24392 38576
rect 24434 38536 24474 38576
rect 24516 38536 24556 38576
rect 24598 38536 24638 38576
rect 24680 38536 24720 38576
rect 28352 38536 28392 38576
rect 28434 38536 28474 38576
rect 28516 38536 28556 38576
rect 28598 38536 28638 38576
rect 28680 38536 28720 38576
rect 32352 38536 32392 38576
rect 32434 38536 32474 38576
rect 32516 38536 32556 38576
rect 32598 38536 32638 38576
rect 32680 38536 32720 38576
rect 36352 38536 36392 38576
rect 36434 38536 36474 38576
rect 36516 38536 36556 38576
rect 36598 38536 36638 38576
rect 36680 38536 36720 38576
rect 40352 38536 40392 38576
rect 40434 38536 40474 38576
rect 40516 38536 40556 38576
rect 40598 38536 40638 38576
rect 40680 38536 40720 38576
rect 44352 38536 44392 38576
rect 44434 38536 44474 38576
rect 44516 38536 44556 38576
rect 44598 38536 44638 38576
rect 44680 38536 44720 38576
rect 48352 38536 48392 38576
rect 48434 38536 48474 38576
rect 48516 38536 48556 38576
rect 48598 38536 48638 38576
rect 48680 38536 48720 38576
rect 52352 38536 52392 38576
rect 52434 38536 52474 38576
rect 52516 38536 52556 38576
rect 52598 38536 52638 38576
rect 52680 38536 52720 38576
rect 56352 38536 56392 38576
rect 56434 38536 56474 38576
rect 56516 38536 56556 38576
rect 56598 38536 56638 38576
rect 56680 38536 56720 38576
rect 60352 38536 60392 38576
rect 60434 38536 60474 38576
rect 60516 38536 60556 38576
rect 60598 38536 60638 38576
rect 60680 38536 60720 38576
rect 64352 38536 64392 38576
rect 64434 38536 64474 38576
rect 64516 38536 64556 38576
rect 64598 38536 64638 38576
rect 64680 38536 64720 38576
rect 68352 38536 68392 38576
rect 68434 38536 68474 38576
rect 68516 38536 68556 38576
rect 68598 38536 68638 38576
rect 68680 38536 68720 38576
rect 72352 38536 72392 38576
rect 72434 38536 72474 38576
rect 72516 38536 72556 38576
rect 72598 38536 72638 38576
rect 72680 38536 72720 38576
rect 76352 38536 76392 38576
rect 76434 38536 76474 38576
rect 76516 38536 76556 38576
rect 76598 38536 76638 38576
rect 76680 38536 76720 38576
rect 80352 38536 80392 38576
rect 80434 38536 80474 38576
rect 80516 38536 80556 38576
rect 80598 38536 80638 38576
rect 80680 38536 80720 38576
rect 84352 38536 84392 38576
rect 84434 38536 84474 38576
rect 84516 38536 84556 38576
rect 84598 38536 84638 38576
rect 84680 38536 84720 38576
rect 88352 38536 88392 38576
rect 88434 38536 88474 38576
rect 88516 38536 88556 38576
rect 88598 38536 88638 38576
rect 88680 38536 88720 38576
rect 92352 38536 92392 38576
rect 92434 38536 92474 38576
rect 92516 38536 92556 38576
rect 92598 38536 92638 38576
rect 92680 38536 92720 38576
rect 96352 38536 96392 38576
rect 96434 38536 96474 38576
rect 96516 38536 96556 38576
rect 96598 38536 96638 38576
rect 96680 38536 96720 38576
rect 3112 37780 3152 37820
rect 3194 37780 3234 37820
rect 3276 37780 3316 37820
rect 3358 37780 3398 37820
rect 3440 37780 3480 37820
rect 7112 37780 7152 37820
rect 7194 37780 7234 37820
rect 7276 37780 7316 37820
rect 7358 37780 7398 37820
rect 7440 37780 7480 37820
rect 11112 37780 11152 37820
rect 11194 37780 11234 37820
rect 11276 37780 11316 37820
rect 11358 37780 11398 37820
rect 11440 37780 11480 37820
rect 15112 37780 15152 37820
rect 15194 37780 15234 37820
rect 15276 37780 15316 37820
rect 15358 37780 15398 37820
rect 15440 37780 15480 37820
rect 19112 37780 19152 37820
rect 19194 37780 19234 37820
rect 19276 37780 19316 37820
rect 19358 37780 19398 37820
rect 19440 37780 19480 37820
rect 23112 37780 23152 37820
rect 23194 37780 23234 37820
rect 23276 37780 23316 37820
rect 23358 37780 23398 37820
rect 23440 37780 23480 37820
rect 27112 37780 27152 37820
rect 27194 37780 27234 37820
rect 27276 37780 27316 37820
rect 27358 37780 27398 37820
rect 27440 37780 27480 37820
rect 31112 37780 31152 37820
rect 31194 37780 31234 37820
rect 31276 37780 31316 37820
rect 31358 37780 31398 37820
rect 31440 37780 31480 37820
rect 35112 37780 35152 37820
rect 35194 37780 35234 37820
rect 35276 37780 35316 37820
rect 35358 37780 35398 37820
rect 35440 37780 35480 37820
rect 39112 37780 39152 37820
rect 39194 37780 39234 37820
rect 39276 37780 39316 37820
rect 39358 37780 39398 37820
rect 39440 37780 39480 37820
rect 43112 37780 43152 37820
rect 43194 37780 43234 37820
rect 43276 37780 43316 37820
rect 43358 37780 43398 37820
rect 43440 37780 43480 37820
rect 47112 37780 47152 37820
rect 47194 37780 47234 37820
rect 47276 37780 47316 37820
rect 47358 37780 47398 37820
rect 47440 37780 47480 37820
rect 51112 37780 51152 37820
rect 51194 37780 51234 37820
rect 51276 37780 51316 37820
rect 51358 37780 51398 37820
rect 51440 37780 51480 37820
rect 55112 37780 55152 37820
rect 55194 37780 55234 37820
rect 55276 37780 55316 37820
rect 55358 37780 55398 37820
rect 55440 37780 55480 37820
rect 59112 37780 59152 37820
rect 59194 37780 59234 37820
rect 59276 37780 59316 37820
rect 59358 37780 59398 37820
rect 59440 37780 59480 37820
rect 63112 37780 63152 37820
rect 63194 37780 63234 37820
rect 63276 37780 63316 37820
rect 63358 37780 63398 37820
rect 63440 37780 63480 37820
rect 67112 37780 67152 37820
rect 67194 37780 67234 37820
rect 67276 37780 67316 37820
rect 67358 37780 67398 37820
rect 67440 37780 67480 37820
rect 71112 37780 71152 37820
rect 71194 37780 71234 37820
rect 71276 37780 71316 37820
rect 71358 37780 71398 37820
rect 71440 37780 71480 37820
rect 75112 37780 75152 37820
rect 75194 37780 75234 37820
rect 75276 37780 75316 37820
rect 75358 37780 75398 37820
rect 75440 37780 75480 37820
rect 79112 37780 79152 37820
rect 79194 37780 79234 37820
rect 79276 37780 79316 37820
rect 79358 37780 79398 37820
rect 79440 37780 79480 37820
rect 83112 37780 83152 37820
rect 83194 37780 83234 37820
rect 83276 37780 83316 37820
rect 83358 37780 83398 37820
rect 83440 37780 83480 37820
rect 87112 37780 87152 37820
rect 87194 37780 87234 37820
rect 87276 37780 87316 37820
rect 87358 37780 87398 37820
rect 87440 37780 87480 37820
rect 91112 37780 91152 37820
rect 91194 37780 91234 37820
rect 91276 37780 91316 37820
rect 91358 37780 91398 37820
rect 91440 37780 91480 37820
rect 95112 37780 95152 37820
rect 95194 37780 95234 37820
rect 95276 37780 95316 37820
rect 95358 37780 95398 37820
rect 95440 37780 95480 37820
rect 99112 37780 99152 37820
rect 99194 37780 99234 37820
rect 99276 37780 99316 37820
rect 99358 37780 99398 37820
rect 99440 37780 99480 37820
rect 4352 37024 4392 37064
rect 4434 37024 4474 37064
rect 4516 37024 4556 37064
rect 4598 37024 4638 37064
rect 4680 37024 4720 37064
rect 8352 37024 8392 37064
rect 8434 37024 8474 37064
rect 8516 37024 8556 37064
rect 8598 37024 8638 37064
rect 8680 37024 8720 37064
rect 12352 37024 12392 37064
rect 12434 37024 12474 37064
rect 12516 37024 12556 37064
rect 12598 37024 12638 37064
rect 12680 37024 12720 37064
rect 16352 37024 16392 37064
rect 16434 37024 16474 37064
rect 16516 37024 16556 37064
rect 16598 37024 16638 37064
rect 16680 37024 16720 37064
rect 20352 37024 20392 37064
rect 20434 37024 20474 37064
rect 20516 37024 20556 37064
rect 20598 37024 20638 37064
rect 20680 37024 20720 37064
rect 24352 37024 24392 37064
rect 24434 37024 24474 37064
rect 24516 37024 24556 37064
rect 24598 37024 24638 37064
rect 24680 37024 24720 37064
rect 28352 37024 28392 37064
rect 28434 37024 28474 37064
rect 28516 37024 28556 37064
rect 28598 37024 28638 37064
rect 28680 37024 28720 37064
rect 32352 37024 32392 37064
rect 32434 37024 32474 37064
rect 32516 37024 32556 37064
rect 32598 37024 32638 37064
rect 32680 37024 32720 37064
rect 36352 37024 36392 37064
rect 36434 37024 36474 37064
rect 36516 37024 36556 37064
rect 36598 37024 36638 37064
rect 36680 37024 36720 37064
rect 40352 37024 40392 37064
rect 40434 37024 40474 37064
rect 40516 37024 40556 37064
rect 40598 37024 40638 37064
rect 40680 37024 40720 37064
rect 44352 37024 44392 37064
rect 44434 37024 44474 37064
rect 44516 37024 44556 37064
rect 44598 37024 44638 37064
rect 44680 37024 44720 37064
rect 48352 37024 48392 37064
rect 48434 37024 48474 37064
rect 48516 37024 48556 37064
rect 48598 37024 48638 37064
rect 48680 37024 48720 37064
rect 52352 37024 52392 37064
rect 52434 37024 52474 37064
rect 52516 37024 52556 37064
rect 52598 37024 52638 37064
rect 52680 37024 52720 37064
rect 56352 37024 56392 37064
rect 56434 37024 56474 37064
rect 56516 37024 56556 37064
rect 56598 37024 56638 37064
rect 56680 37024 56720 37064
rect 60352 37024 60392 37064
rect 60434 37024 60474 37064
rect 60516 37024 60556 37064
rect 60598 37024 60638 37064
rect 60680 37024 60720 37064
rect 64352 37024 64392 37064
rect 64434 37024 64474 37064
rect 64516 37024 64556 37064
rect 64598 37024 64638 37064
rect 64680 37024 64720 37064
rect 68352 37024 68392 37064
rect 68434 37024 68474 37064
rect 68516 37024 68556 37064
rect 68598 37024 68638 37064
rect 68680 37024 68720 37064
rect 72352 37024 72392 37064
rect 72434 37024 72474 37064
rect 72516 37024 72556 37064
rect 72598 37024 72638 37064
rect 72680 37024 72720 37064
rect 76352 37024 76392 37064
rect 76434 37024 76474 37064
rect 76516 37024 76556 37064
rect 76598 37024 76638 37064
rect 76680 37024 76720 37064
rect 80352 37024 80392 37064
rect 80434 37024 80474 37064
rect 80516 37024 80556 37064
rect 80598 37024 80638 37064
rect 80680 37024 80720 37064
rect 84352 37024 84392 37064
rect 84434 37024 84474 37064
rect 84516 37024 84556 37064
rect 84598 37024 84638 37064
rect 84680 37024 84720 37064
rect 88352 37024 88392 37064
rect 88434 37024 88474 37064
rect 88516 37024 88556 37064
rect 88598 37024 88638 37064
rect 88680 37024 88720 37064
rect 92352 37024 92392 37064
rect 92434 37024 92474 37064
rect 92516 37024 92556 37064
rect 92598 37024 92638 37064
rect 92680 37024 92720 37064
rect 96352 37024 96392 37064
rect 96434 37024 96474 37064
rect 96516 37024 96556 37064
rect 96598 37024 96638 37064
rect 96680 37024 96720 37064
rect 3112 36268 3152 36308
rect 3194 36268 3234 36308
rect 3276 36268 3316 36308
rect 3358 36268 3398 36308
rect 3440 36268 3480 36308
rect 7112 36268 7152 36308
rect 7194 36268 7234 36308
rect 7276 36268 7316 36308
rect 7358 36268 7398 36308
rect 7440 36268 7480 36308
rect 11112 36268 11152 36308
rect 11194 36268 11234 36308
rect 11276 36268 11316 36308
rect 11358 36268 11398 36308
rect 11440 36268 11480 36308
rect 15112 36268 15152 36308
rect 15194 36268 15234 36308
rect 15276 36268 15316 36308
rect 15358 36268 15398 36308
rect 15440 36268 15480 36308
rect 19112 36268 19152 36308
rect 19194 36268 19234 36308
rect 19276 36268 19316 36308
rect 19358 36268 19398 36308
rect 19440 36268 19480 36308
rect 23112 36268 23152 36308
rect 23194 36268 23234 36308
rect 23276 36268 23316 36308
rect 23358 36268 23398 36308
rect 23440 36268 23480 36308
rect 27112 36268 27152 36308
rect 27194 36268 27234 36308
rect 27276 36268 27316 36308
rect 27358 36268 27398 36308
rect 27440 36268 27480 36308
rect 31112 36268 31152 36308
rect 31194 36268 31234 36308
rect 31276 36268 31316 36308
rect 31358 36268 31398 36308
rect 31440 36268 31480 36308
rect 35112 36268 35152 36308
rect 35194 36268 35234 36308
rect 35276 36268 35316 36308
rect 35358 36268 35398 36308
rect 35440 36268 35480 36308
rect 39112 36268 39152 36308
rect 39194 36268 39234 36308
rect 39276 36268 39316 36308
rect 39358 36268 39398 36308
rect 39440 36268 39480 36308
rect 43112 36268 43152 36308
rect 43194 36268 43234 36308
rect 43276 36268 43316 36308
rect 43358 36268 43398 36308
rect 43440 36268 43480 36308
rect 47112 36268 47152 36308
rect 47194 36268 47234 36308
rect 47276 36268 47316 36308
rect 47358 36268 47398 36308
rect 47440 36268 47480 36308
rect 51112 36268 51152 36308
rect 51194 36268 51234 36308
rect 51276 36268 51316 36308
rect 51358 36268 51398 36308
rect 51440 36268 51480 36308
rect 55112 36268 55152 36308
rect 55194 36268 55234 36308
rect 55276 36268 55316 36308
rect 55358 36268 55398 36308
rect 55440 36268 55480 36308
rect 59112 36268 59152 36308
rect 59194 36268 59234 36308
rect 59276 36268 59316 36308
rect 59358 36268 59398 36308
rect 59440 36268 59480 36308
rect 63112 36268 63152 36308
rect 63194 36268 63234 36308
rect 63276 36268 63316 36308
rect 63358 36268 63398 36308
rect 63440 36268 63480 36308
rect 67112 36268 67152 36308
rect 67194 36268 67234 36308
rect 67276 36268 67316 36308
rect 67358 36268 67398 36308
rect 67440 36268 67480 36308
rect 71112 36268 71152 36308
rect 71194 36268 71234 36308
rect 71276 36268 71316 36308
rect 71358 36268 71398 36308
rect 71440 36268 71480 36308
rect 75112 36268 75152 36308
rect 75194 36268 75234 36308
rect 75276 36268 75316 36308
rect 75358 36268 75398 36308
rect 75440 36268 75480 36308
rect 79112 36268 79152 36308
rect 79194 36268 79234 36308
rect 79276 36268 79316 36308
rect 79358 36268 79398 36308
rect 79440 36268 79480 36308
rect 83112 36268 83152 36308
rect 83194 36268 83234 36308
rect 83276 36268 83316 36308
rect 83358 36268 83398 36308
rect 83440 36268 83480 36308
rect 87112 36268 87152 36308
rect 87194 36268 87234 36308
rect 87276 36268 87316 36308
rect 87358 36268 87398 36308
rect 87440 36268 87480 36308
rect 91112 36268 91152 36308
rect 91194 36268 91234 36308
rect 91276 36268 91316 36308
rect 91358 36268 91398 36308
rect 91440 36268 91480 36308
rect 95112 36268 95152 36308
rect 95194 36268 95234 36308
rect 95276 36268 95316 36308
rect 95358 36268 95398 36308
rect 95440 36268 95480 36308
rect 99112 36268 99152 36308
rect 99194 36268 99234 36308
rect 99276 36268 99316 36308
rect 99358 36268 99398 36308
rect 99440 36268 99480 36308
rect 4352 35512 4392 35552
rect 4434 35512 4474 35552
rect 4516 35512 4556 35552
rect 4598 35512 4638 35552
rect 4680 35512 4720 35552
rect 8352 35512 8392 35552
rect 8434 35512 8474 35552
rect 8516 35512 8556 35552
rect 8598 35512 8638 35552
rect 8680 35512 8720 35552
rect 12352 35512 12392 35552
rect 12434 35512 12474 35552
rect 12516 35512 12556 35552
rect 12598 35512 12638 35552
rect 12680 35512 12720 35552
rect 16352 35512 16392 35552
rect 16434 35512 16474 35552
rect 16516 35512 16556 35552
rect 16598 35512 16638 35552
rect 16680 35512 16720 35552
rect 20352 35512 20392 35552
rect 20434 35512 20474 35552
rect 20516 35512 20556 35552
rect 20598 35512 20638 35552
rect 20680 35512 20720 35552
rect 24352 35512 24392 35552
rect 24434 35512 24474 35552
rect 24516 35512 24556 35552
rect 24598 35512 24638 35552
rect 24680 35512 24720 35552
rect 28352 35512 28392 35552
rect 28434 35512 28474 35552
rect 28516 35512 28556 35552
rect 28598 35512 28638 35552
rect 28680 35512 28720 35552
rect 32352 35512 32392 35552
rect 32434 35512 32474 35552
rect 32516 35512 32556 35552
rect 32598 35512 32638 35552
rect 32680 35512 32720 35552
rect 36352 35512 36392 35552
rect 36434 35512 36474 35552
rect 36516 35512 36556 35552
rect 36598 35512 36638 35552
rect 36680 35512 36720 35552
rect 40352 35512 40392 35552
rect 40434 35512 40474 35552
rect 40516 35512 40556 35552
rect 40598 35512 40638 35552
rect 40680 35512 40720 35552
rect 44352 35512 44392 35552
rect 44434 35512 44474 35552
rect 44516 35512 44556 35552
rect 44598 35512 44638 35552
rect 44680 35512 44720 35552
rect 48352 35512 48392 35552
rect 48434 35512 48474 35552
rect 48516 35512 48556 35552
rect 48598 35512 48638 35552
rect 48680 35512 48720 35552
rect 52352 35512 52392 35552
rect 52434 35512 52474 35552
rect 52516 35512 52556 35552
rect 52598 35512 52638 35552
rect 52680 35512 52720 35552
rect 56352 35512 56392 35552
rect 56434 35512 56474 35552
rect 56516 35512 56556 35552
rect 56598 35512 56638 35552
rect 56680 35512 56720 35552
rect 60352 35512 60392 35552
rect 60434 35512 60474 35552
rect 60516 35512 60556 35552
rect 60598 35512 60638 35552
rect 60680 35512 60720 35552
rect 64352 35512 64392 35552
rect 64434 35512 64474 35552
rect 64516 35512 64556 35552
rect 64598 35512 64638 35552
rect 64680 35512 64720 35552
rect 68352 35512 68392 35552
rect 68434 35512 68474 35552
rect 68516 35512 68556 35552
rect 68598 35512 68638 35552
rect 68680 35512 68720 35552
rect 72352 35512 72392 35552
rect 72434 35512 72474 35552
rect 72516 35512 72556 35552
rect 72598 35512 72638 35552
rect 72680 35512 72720 35552
rect 76352 35512 76392 35552
rect 76434 35512 76474 35552
rect 76516 35512 76556 35552
rect 76598 35512 76638 35552
rect 76680 35512 76720 35552
rect 80352 35512 80392 35552
rect 80434 35512 80474 35552
rect 80516 35512 80556 35552
rect 80598 35512 80638 35552
rect 80680 35512 80720 35552
rect 84352 35512 84392 35552
rect 84434 35512 84474 35552
rect 84516 35512 84556 35552
rect 84598 35512 84638 35552
rect 84680 35512 84720 35552
rect 88352 35512 88392 35552
rect 88434 35512 88474 35552
rect 88516 35512 88556 35552
rect 88598 35512 88638 35552
rect 88680 35512 88720 35552
rect 92352 35512 92392 35552
rect 92434 35512 92474 35552
rect 92516 35512 92556 35552
rect 92598 35512 92638 35552
rect 92680 35512 92720 35552
rect 96352 35512 96392 35552
rect 96434 35512 96474 35552
rect 96516 35512 96556 35552
rect 96598 35512 96638 35552
rect 96680 35512 96720 35552
rect 3112 34756 3152 34796
rect 3194 34756 3234 34796
rect 3276 34756 3316 34796
rect 3358 34756 3398 34796
rect 3440 34756 3480 34796
rect 7112 34756 7152 34796
rect 7194 34756 7234 34796
rect 7276 34756 7316 34796
rect 7358 34756 7398 34796
rect 7440 34756 7480 34796
rect 11112 34756 11152 34796
rect 11194 34756 11234 34796
rect 11276 34756 11316 34796
rect 11358 34756 11398 34796
rect 11440 34756 11480 34796
rect 15112 34756 15152 34796
rect 15194 34756 15234 34796
rect 15276 34756 15316 34796
rect 15358 34756 15398 34796
rect 15440 34756 15480 34796
rect 19112 34756 19152 34796
rect 19194 34756 19234 34796
rect 19276 34756 19316 34796
rect 19358 34756 19398 34796
rect 19440 34756 19480 34796
rect 23112 34756 23152 34796
rect 23194 34756 23234 34796
rect 23276 34756 23316 34796
rect 23358 34756 23398 34796
rect 23440 34756 23480 34796
rect 27112 34756 27152 34796
rect 27194 34756 27234 34796
rect 27276 34756 27316 34796
rect 27358 34756 27398 34796
rect 27440 34756 27480 34796
rect 31112 34756 31152 34796
rect 31194 34756 31234 34796
rect 31276 34756 31316 34796
rect 31358 34756 31398 34796
rect 31440 34756 31480 34796
rect 35112 34756 35152 34796
rect 35194 34756 35234 34796
rect 35276 34756 35316 34796
rect 35358 34756 35398 34796
rect 35440 34756 35480 34796
rect 39112 34756 39152 34796
rect 39194 34756 39234 34796
rect 39276 34756 39316 34796
rect 39358 34756 39398 34796
rect 39440 34756 39480 34796
rect 43112 34756 43152 34796
rect 43194 34756 43234 34796
rect 43276 34756 43316 34796
rect 43358 34756 43398 34796
rect 43440 34756 43480 34796
rect 47112 34756 47152 34796
rect 47194 34756 47234 34796
rect 47276 34756 47316 34796
rect 47358 34756 47398 34796
rect 47440 34756 47480 34796
rect 51112 34756 51152 34796
rect 51194 34756 51234 34796
rect 51276 34756 51316 34796
rect 51358 34756 51398 34796
rect 51440 34756 51480 34796
rect 55112 34756 55152 34796
rect 55194 34756 55234 34796
rect 55276 34756 55316 34796
rect 55358 34756 55398 34796
rect 55440 34756 55480 34796
rect 59112 34756 59152 34796
rect 59194 34756 59234 34796
rect 59276 34756 59316 34796
rect 59358 34756 59398 34796
rect 59440 34756 59480 34796
rect 63112 34756 63152 34796
rect 63194 34756 63234 34796
rect 63276 34756 63316 34796
rect 63358 34756 63398 34796
rect 63440 34756 63480 34796
rect 67112 34756 67152 34796
rect 67194 34756 67234 34796
rect 67276 34756 67316 34796
rect 67358 34756 67398 34796
rect 67440 34756 67480 34796
rect 71112 34756 71152 34796
rect 71194 34756 71234 34796
rect 71276 34756 71316 34796
rect 71358 34756 71398 34796
rect 71440 34756 71480 34796
rect 75112 34756 75152 34796
rect 75194 34756 75234 34796
rect 75276 34756 75316 34796
rect 75358 34756 75398 34796
rect 75440 34756 75480 34796
rect 79112 34756 79152 34796
rect 79194 34756 79234 34796
rect 79276 34756 79316 34796
rect 79358 34756 79398 34796
rect 79440 34756 79480 34796
rect 83112 34756 83152 34796
rect 83194 34756 83234 34796
rect 83276 34756 83316 34796
rect 83358 34756 83398 34796
rect 83440 34756 83480 34796
rect 87112 34756 87152 34796
rect 87194 34756 87234 34796
rect 87276 34756 87316 34796
rect 87358 34756 87398 34796
rect 87440 34756 87480 34796
rect 91112 34756 91152 34796
rect 91194 34756 91234 34796
rect 91276 34756 91316 34796
rect 91358 34756 91398 34796
rect 91440 34756 91480 34796
rect 95112 34756 95152 34796
rect 95194 34756 95234 34796
rect 95276 34756 95316 34796
rect 95358 34756 95398 34796
rect 95440 34756 95480 34796
rect 99112 34756 99152 34796
rect 99194 34756 99234 34796
rect 99276 34756 99316 34796
rect 99358 34756 99398 34796
rect 99440 34756 99480 34796
rect 4352 34000 4392 34040
rect 4434 34000 4474 34040
rect 4516 34000 4556 34040
rect 4598 34000 4638 34040
rect 4680 34000 4720 34040
rect 8352 34000 8392 34040
rect 8434 34000 8474 34040
rect 8516 34000 8556 34040
rect 8598 34000 8638 34040
rect 8680 34000 8720 34040
rect 12352 34000 12392 34040
rect 12434 34000 12474 34040
rect 12516 34000 12556 34040
rect 12598 34000 12638 34040
rect 12680 34000 12720 34040
rect 16352 34000 16392 34040
rect 16434 34000 16474 34040
rect 16516 34000 16556 34040
rect 16598 34000 16638 34040
rect 16680 34000 16720 34040
rect 20352 34000 20392 34040
rect 20434 34000 20474 34040
rect 20516 34000 20556 34040
rect 20598 34000 20638 34040
rect 20680 34000 20720 34040
rect 24352 34000 24392 34040
rect 24434 34000 24474 34040
rect 24516 34000 24556 34040
rect 24598 34000 24638 34040
rect 24680 34000 24720 34040
rect 28352 34000 28392 34040
rect 28434 34000 28474 34040
rect 28516 34000 28556 34040
rect 28598 34000 28638 34040
rect 28680 34000 28720 34040
rect 32352 34000 32392 34040
rect 32434 34000 32474 34040
rect 32516 34000 32556 34040
rect 32598 34000 32638 34040
rect 32680 34000 32720 34040
rect 36352 34000 36392 34040
rect 36434 34000 36474 34040
rect 36516 34000 36556 34040
rect 36598 34000 36638 34040
rect 36680 34000 36720 34040
rect 40352 34000 40392 34040
rect 40434 34000 40474 34040
rect 40516 34000 40556 34040
rect 40598 34000 40638 34040
rect 40680 34000 40720 34040
rect 44352 34000 44392 34040
rect 44434 34000 44474 34040
rect 44516 34000 44556 34040
rect 44598 34000 44638 34040
rect 44680 34000 44720 34040
rect 48352 34000 48392 34040
rect 48434 34000 48474 34040
rect 48516 34000 48556 34040
rect 48598 34000 48638 34040
rect 48680 34000 48720 34040
rect 52352 34000 52392 34040
rect 52434 34000 52474 34040
rect 52516 34000 52556 34040
rect 52598 34000 52638 34040
rect 52680 34000 52720 34040
rect 56352 34000 56392 34040
rect 56434 34000 56474 34040
rect 56516 34000 56556 34040
rect 56598 34000 56638 34040
rect 56680 34000 56720 34040
rect 60352 34000 60392 34040
rect 60434 34000 60474 34040
rect 60516 34000 60556 34040
rect 60598 34000 60638 34040
rect 60680 34000 60720 34040
rect 64352 34000 64392 34040
rect 64434 34000 64474 34040
rect 64516 34000 64556 34040
rect 64598 34000 64638 34040
rect 64680 34000 64720 34040
rect 68352 34000 68392 34040
rect 68434 34000 68474 34040
rect 68516 34000 68556 34040
rect 68598 34000 68638 34040
rect 68680 34000 68720 34040
rect 87052 33412 87092 33452
rect 3112 33244 3152 33284
rect 3194 33244 3234 33284
rect 3276 33244 3316 33284
rect 3358 33244 3398 33284
rect 3440 33244 3480 33284
rect 7112 33244 7152 33284
rect 7194 33244 7234 33284
rect 7276 33244 7316 33284
rect 7358 33244 7398 33284
rect 7440 33244 7480 33284
rect 11112 33244 11152 33284
rect 11194 33244 11234 33284
rect 11276 33244 11316 33284
rect 11358 33244 11398 33284
rect 11440 33244 11480 33284
rect 15112 33244 15152 33284
rect 15194 33244 15234 33284
rect 15276 33244 15316 33284
rect 15358 33244 15398 33284
rect 15440 33244 15480 33284
rect 19112 33244 19152 33284
rect 19194 33244 19234 33284
rect 19276 33244 19316 33284
rect 19358 33244 19398 33284
rect 19440 33244 19480 33284
rect 23112 33244 23152 33284
rect 23194 33244 23234 33284
rect 23276 33244 23316 33284
rect 23358 33244 23398 33284
rect 23440 33244 23480 33284
rect 27112 33244 27152 33284
rect 27194 33244 27234 33284
rect 27276 33244 27316 33284
rect 27358 33244 27398 33284
rect 27440 33244 27480 33284
rect 31112 33244 31152 33284
rect 31194 33244 31234 33284
rect 31276 33244 31316 33284
rect 31358 33244 31398 33284
rect 31440 33244 31480 33284
rect 35112 33244 35152 33284
rect 35194 33244 35234 33284
rect 35276 33244 35316 33284
rect 35358 33244 35398 33284
rect 35440 33244 35480 33284
rect 39112 33244 39152 33284
rect 39194 33244 39234 33284
rect 39276 33244 39316 33284
rect 39358 33244 39398 33284
rect 39440 33244 39480 33284
rect 43112 33244 43152 33284
rect 43194 33244 43234 33284
rect 43276 33244 43316 33284
rect 43358 33244 43398 33284
rect 43440 33244 43480 33284
rect 47112 33244 47152 33284
rect 47194 33244 47234 33284
rect 47276 33244 47316 33284
rect 47358 33244 47398 33284
rect 47440 33244 47480 33284
rect 51112 33244 51152 33284
rect 51194 33244 51234 33284
rect 51276 33244 51316 33284
rect 51358 33244 51398 33284
rect 51440 33244 51480 33284
rect 55112 33244 55152 33284
rect 55194 33244 55234 33284
rect 55276 33244 55316 33284
rect 55358 33244 55398 33284
rect 55440 33244 55480 33284
rect 59112 33244 59152 33284
rect 59194 33244 59234 33284
rect 59276 33244 59316 33284
rect 59358 33244 59398 33284
rect 59440 33244 59480 33284
rect 63112 33244 63152 33284
rect 63194 33244 63234 33284
rect 63276 33244 63316 33284
rect 63358 33244 63398 33284
rect 63440 33244 63480 33284
rect 67112 33244 67152 33284
rect 67194 33244 67234 33284
rect 67276 33244 67316 33284
rect 67358 33244 67398 33284
rect 67440 33244 67480 33284
rect 73612 32824 73652 32864
rect 4352 32488 4392 32528
rect 4434 32488 4474 32528
rect 4516 32488 4556 32528
rect 4598 32488 4638 32528
rect 4680 32488 4720 32528
rect 8352 32488 8392 32528
rect 8434 32488 8474 32528
rect 8516 32488 8556 32528
rect 8598 32488 8638 32528
rect 8680 32488 8720 32528
rect 12352 32488 12392 32528
rect 12434 32488 12474 32528
rect 12516 32488 12556 32528
rect 12598 32488 12638 32528
rect 12680 32488 12720 32528
rect 16352 32488 16392 32528
rect 16434 32488 16474 32528
rect 16516 32488 16556 32528
rect 16598 32488 16638 32528
rect 16680 32488 16720 32528
rect 20352 32488 20392 32528
rect 20434 32488 20474 32528
rect 20516 32488 20556 32528
rect 20598 32488 20638 32528
rect 20680 32488 20720 32528
rect 24352 32488 24392 32528
rect 24434 32488 24474 32528
rect 24516 32488 24556 32528
rect 24598 32488 24638 32528
rect 24680 32488 24720 32528
rect 28352 32488 28392 32528
rect 28434 32488 28474 32528
rect 28516 32488 28556 32528
rect 28598 32488 28638 32528
rect 28680 32488 28720 32528
rect 32352 32488 32392 32528
rect 32434 32488 32474 32528
rect 32516 32488 32556 32528
rect 32598 32488 32638 32528
rect 32680 32488 32720 32528
rect 36352 32488 36392 32528
rect 36434 32488 36474 32528
rect 36516 32488 36556 32528
rect 36598 32488 36638 32528
rect 36680 32488 36720 32528
rect 40352 32488 40392 32528
rect 40434 32488 40474 32528
rect 40516 32488 40556 32528
rect 40598 32488 40638 32528
rect 40680 32488 40720 32528
rect 44352 32488 44392 32528
rect 44434 32488 44474 32528
rect 44516 32488 44556 32528
rect 44598 32488 44638 32528
rect 44680 32488 44720 32528
rect 48352 32488 48392 32528
rect 48434 32488 48474 32528
rect 48516 32488 48556 32528
rect 48598 32488 48638 32528
rect 48680 32488 48720 32528
rect 52352 32488 52392 32528
rect 52434 32488 52474 32528
rect 52516 32488 52556 32528
rect 52598 32488 52638 32528
rect 52680 32488 52720 32528
rect 56352 32488 56392 32528
rect 56434 32488 56474 32528
rect 56516 32488 56556 32528
rect 56598 32488 56638 32528
rect 56680 32488 56720 32528
rect 60352 32488 60392 32528
rect 60434 32488 60474 32528
rect 60516 32488 60556 32528
rect 60598 32488 60638 32528
rect 60680 32488 60720 32528
rect 64352 32488 64392 32528
rect 64434 32488 64474 32528
rect 64516 32488 64556 32528
rect 64598 32488 64638 32528
rect 64680 32488 64720 32528
rect 68352 32488 68392 32528
rect 68434 32488 68474 32528
rect 68516 32488 68556 32528
rect 68598 32488 68638 32528
rect 68680 32488 68720 32528
rect 3112 31732 3152 31772
rect 3194 31732 3234 31772
rect 3276 31732 3316 31772
rect 3358 31732 3398 31772
rect 3440 31732 3480 31772
rect 7112 31732 7152 31772
rect 7194 31732 7234 31772
rect 7276 31732 7316 31772
rect 7358 31732 7398 31772
rect 7440 31732 7480 31772
rect 11112 31732 11152 31772
rect 11194 31732 11234 31772
rect 11276 31732 11316 31772
rect 11358 31732 11398 31772
rect 11440 31732 11480 31772
rect 15112 31732 15152 31772
rect 15194 31732 15234 31772
rect 15276 31732 15316 31772
rect 15358 31732 15398 31772
rect 15440 31732 15480 31772
rect 19112 31732 19152 31772
rect 19194 31732 19234 31772
rect 19276 31732 19316 31772
rect 19358 31732 19398 31772
rect 19440 31732 19480 31772
rect 23112 31732 23152 31772
rect 23194 31732 23234 31772
rect 23276 31732 23316 31772
rect 23358 31732 23398 31772
rect 23440 31732 23480 31772
rect 27112 31732 27152 31772
rect 27194 31732 27234 31772
rect 27276 31732 27316 31772
rect 27358 31732 27398 31772
rect 27440 31732 27480 31772
rect 31112 31732 31152 31772
rect 31194 31732 31234 31772
rect 31276 31732 31316 31772
rect 31358 31732 31398 31772
rect 31440 31732 31480 31772
rect 35112 31732 35152 31772
rect 35194 31732 35234 31772
rect 35276 31732 35316 31772
rect 35358 31732 35398 31772
rect 35440 31732 35480 31772
rect 39112 31732 39152 31772
rect 39194 31732 39234 31772
rect 39276 31732 39316 31772
rect 39358 31732 39398 31772
rect 39440 31732 39480 31772
rect 43112 31732 43152 31772
rect 43194 31732 43234 31772
rect 43276 31732 43316 31772
rect 43358 31732 43398 31772
rect 43440 31732 43480 31772
rect 47112 31732 47152 31772
rect 47194 31732 47234 31772
rect 47276 31732 47316 31772
rect 47358 31732 47398 31772
rect 47440 31732 47480 31772
rect 51112 31732 51152 31772
rect 51194 31732 51234 31772
rect 51276 31732 51316 31772
rect 51358 31732 51398 31772
rect 51440 31732 51480 31772
rect 55112 31732 55152 31772
rect 55194 31732 55234 31772
rect 55276 31732 55316 31772
rect 55358 31732 55398 31772
rect 55440 31732 55480 31772
rect 59112 31732 59152 31772
rect 59194 31732 59234 31772
rect 59276 31732 59316 31772
rect 59358 31732 59398 31772
rect 59440 31732 59480 31772
rect 63112 31732 63152 31772
rect 63194 31732 63234 31772
rect 63276 31732 63316 31772
rect 63358 31732 63398 31772
rect 63440 31732 63480 31772
rect 67112 31732 67152 31772
rect 67194 31732 67234 31772
rect 67276 31732 67316 31772
rect 67358 31732 67398 31772
rect 67440 31732 67480 31772
rect 4352 30976 4392 31016
rect 4434 30976 4474 31016
rect 4516 30976 4556 31016
rect 4598 30976 4638 31016
rect 4680 30976 4720 31016
rect 8352 30976 8392 31016
rect 8434 30976 8474 31016
rect 8516 30976 8556 31016
rect 8598 30976 8638 31016
rect 8680 30976 8720 31016
rect 12352 30976 12392 31016
rect 12434 30976 12474 31016
rect 12516 30976 12556 31016
rect 12598 30976 12638 31016
rect 12680 30976 12720 31016
rect 16352 30976 16392 31016
rect 16434 30976 16474 31016
rect 16516 30976 16556 31016
rect 16598 30976 16638 31016
rect 16680 30976 16720 31016
rect 20352 30976 20392 31016
rect 20434 30976 20474 31016
rect 20516 30976 20556 31016
rect 20598 30976 20638 31016
rect 20680 30976 20720 31016
rect 24352 30976 24392 31016
rect 24434 30976 24474 31016
rect 24516 30976 24556 31016
rect 24598 30976 24638 31016
rect 24680 30976 24720 31016
rect 28352 30976 28392 31016
rect 28434 30976 28474 31016
rect 28516 30976 28556 31016
rect 28598 30976 28638 31016
rect 28680 30976 28720 31016
rect 32352 30976 32392 31016
rect 32434 30976 32474 31016
rect 32516 30976 32556 31016
rect 32598 30976 32638 31016
rect 32680 30976 32720 31016
rect 36352 30976 36392 31016
rect 36434 30976 36474 31016
rect 36516 30976 36556 31016
rect 36598 30976 36638 31016
rect 36680 30976 36720 31016
rect 40352 30976 40392 31016
rect 40434 30976 40474 31016
rect 40516 30976 40556 31016
rect 40598 30976 40638 31016
rect 40680 30976 40720 31016
rect 44352 30976 44392 31016
rect 44434 30976 44474 31016
rect 44516 30976 44556 31016
rect 44598 30976 44638 31016
rect 44680 30976 44720 31016
rect 48352 30976 48392 31016
rect 48434 30976 48474 31016
rect 48516 30976 48556 31016
rect 48598 30976 48638 31016
rect 48680 30976 48720 31016
rect 52352 30976 52392 31016
rect 52434 30976 52474 31016
rect 52516 30976 52556 31016
rect 52598 30976 52638 31016
rect 52680 30976 52720 31016
rect 56352 30976 56392 31016
rect 56434 30976 56474 31016
rect 56516 30976 56556 31016
rect 56598 30976 56638 31016
rect 56680 30976 56720 31016
rect 60352 30976 60392 31016
rect 60434 30976 60474 31016
rect 60516 30976 60556 31016
rect 60598 30976 60638 31016
rect 60680 30976 60720 31016
rect 64352 30976 64392 31016
rect 64434 30976 64474 31016
rect 64516 30976 64556 31016
rect 64598 30976 64638 31016
rect 64680 30976 64720 31016
rect 68352 30976 68392 31016
rect 68434 30976 68474 31016
rect 68516 30976 68556 31016
rect 68598 30976 68638 31016
rect 68680 30976 68720 31016
rect 3112 30220 3152 30260
rect 3194 30220 3234 30260
rect 3276 30220 3316 30260
rect 3358 30220 3398 30260
rect 3440 30220 3480 30260
rect 7112 30220 7152 30260
rect 7194 30220 7234 30260
rect 7276 30220 7316 30260
rect 7358 30220 7398 30260
rect 7440 30220 7480 30260
rect 11112 30220 11152 30260
rect 11194 30220 11234 30260
rect 11276 30220 11316 30260
rect 11358 30220 11398 30260
rect 11440 30220 11480 30260
rect 15112 30220 15152 30260
rect 15194 30220 15234 30260
rect 15276 30220 15316 30260
rect 15358 30220 15398 30260
rect 15440 30220 15480 30260
rect 19112 30220 19152 30260
rect 19194 30220 19234 30260
rect 19276 30220 19316 30260
rect 19358 30220 19398 30260
rect 19440 30220 19480 30260
rect 23112 30220 23152 30260
rect 23194 30220 23234 30260
rect 23276 30220 23316 30260
rect 23358 30220 23398 30260
rect 23440 30220 23480 30260
rect 27112 30220 27152 30260
rect 27194 30220 27234 30260
rect 27276 30220 27316 30260
rect 27358 30220 27398 30260
rect 27440 30220 27480 30260
rect 31112 30220 31152 30260
rect 31194 30220 31234 30260
rect 31276 30220 31316 30260
rect 31358 30220 31398 30260
rect 31440 30220 31480 30260
rect 35112 30220 35152 30260
rect 35194 30220 35234 30260
rect 35276 30220 35316 30260
rect 35358 30220 35398 30260
rect 35440 30220 35480 30260
rect 39112 30220 39152 30260
rect 39194 30220 39234 30260
rect 39276 30220 39316 30260
rect 39358 30220 39398 30260
rect 39440 30220 39480 30260
rect 43112 30220 43152 30260
rect 43194 30220 43234 30260
rect 43276 30220 43316 30260
rect 43358 30220 43398 30260
rect 43440 30220 43480 30260
rect 47112 30220 47152 30260
rect 47194 30220 47234 30260
rect 47276 30220 47316 30260
rect 47358 30220 47398 30260
rect 47440 30220 47480 30260
rect 51112 30220 51152 30260
rect 51194 30220 51234 30260
rect 51276 30220 51316 30260
rect 51358 30220 51398 30260
rect 51440 30220 51480 30260
rect 55112 30220 55152 30260
rect 55194 30220 55234 30260
rect 55276 30220 55316 30260
rect 55358 30220 55398 30260
rect 55440 30220 55480 30260
rect 59112 30220 59152 30260
rect 59194 30220 59234 30260
rect 59276 30220 59316 30260
rect 59358 30220 59398 30260
rect 59440 30220 59480 30260
rect 63112 30220 63152 30260
rect 63194 30220 63234 30260
rect 63276 30220 63316 30260
rect 63358 30220 63398 30260
rect 63440 30220 63480 30260
rect 67112 30220 67152 30260
rect 67194 30220 67234 30260
rect 67276 30220 67316 30260
rect 67358 30220 67398 30260
rect 67440 30220 67480 30260
rect 4352 29464 4392 29504
rect 4434 29464 4474 29504
rect 4516 29464 4556 29504
rect 4598 29464 4638 29504
rect 4680 29464 4720 29504
rect 8352 29464 8392 29504
rect 8434 29464 8474 29504
rect 8516 29464 8556 29504
rect 8598 29464 8638 29504
rect 8680 29464 8720 29504
rect 12352 29464 12392 29504
rect 12434 29464 12474 29504
rect 12516 29464 12556 29504
rect 12598 29464 12638 29504
rect 12680 29464 12720 29504
rect 16352 29464 16392 29504
rect 16434 29464 16474 29504
rect 16516 29464 16556 29504
rect 16598 29464 16638 29504
rect 16680 29464 16720 29504
rect 20352 29464 20392 29504
rect 20434 29464 20474 29504
rect 20516 29464 20556 29504
rect 20598 29464 20638 29504
rect 20680 29464 20720 29504
rect 24352 29464 24392 29504
rect 24434 29464 24474 29504
rect 24516 29464 24556 29504
rect 24598 29464 24638 29504
rect 24680 29464 24720 29504
rect 28352 29464 28392 29504
rect 28434 29464 28474 29504
rect 28516 29464 28556 29504
rect 28598 29464 28638 29504
rect 28680 29464 28720 29504
rect 32352 29464 32392 29504
rect 32434 29464 32474 29504
rect 32516 29464 32556 29504
rect 32598 29464 32638 29504
rect 32680 29464 32720 29504
rect 36352 29464 36392 29504
rect 36434 29464 36474 29504
rect 36516 29464 36556 29504
rect 36598 29464 36638 29504
rect 36680 29464 36720 29504
rect 40352 29464 40392 29504
rect 40434 29464 40474 29504
rect 40516 29464 40556 29504
rect 40598 29464 40638 29504
rect 40680 29464 40720 29504
rect 44352 29464 44392 29504
rect 44434 29464 44474 29504
rect 44516 29464 44556 29504
rect 44598 29464 44638 29504
rect 44680 29464 44720 29504
rect 48352 29464 48392 29504
rect 48434 29464 48474 29504
rect 48516 29464 48556 29504
rect 48598 29464 48638 29504
rect 48680 29464 48720 29504
rect 52352 29464 52392 29504
rect 52434 29464 52474 29504
rect 52516 29464 52556 29504
rect 52598 29464 52638 29504
rect 52680 29464 52720 29504
rect 56352 29464 56392 29504
rect 56434 29464 56474 29504
rect 56516 29464 56556 29504
rect 56598 29464 56638 29504
rect 56680 29464 56720 29504
rect 60352 29464 60392 29504
rect 60434 29464 60474 29504
rect 60516 29464 60556 29504
rect 60598 29464 60638 29504
rect 60680 29464 60720 29504
rect 64352 29464 64392 29504
rect 64434 29464 64474 29504
rect 64516 29464 64556 29504
rect 64598 29464 64638 29504
rect 64680 29464 64720 29504
rect 68352 29464 68392 29504
rect 68434 29464 68474 29504
rect 68516 29464 68556 29504
rect 68598 29464 68638 29504
rect 68680 29464 68720 29504
rect 3112 28708 3152 28748
rect 3194 28708 3234 28748
rect 3276 28708 3316 28748
rect 3358 28708 3398 28748
rect 3440 28708 3480 28748
rect 7112 28708 7152 28748
rect 7194 28708 7234 28748
rect 7276 28708 7316 28748
rect 7358 28708 7398 28748
rect 7440 28708 7480 28748
rect 11112 28708 11152 28748
rect 11194 28708 11234 28748
rect 11276 28708 11316 28748
rect 11358 28708 11398 28748
rect 11440 28708 11480 28748
rect 15112 28708 15152 28748
rect 15194 28708 15234 28748
rect 15276 28708 15316 28748
rect 15358 28708 15398 28748
rect 15440 28708 15480 28748
rect 19112 28708 19152 28748
rect 19194 28708 19234 28748
rect 19276 28708 19316 28748
rect 19358 28708 19398 28748
rect 19440 28708 19480 28748
rect 23112 28708 23152 28748
rect 23194 28708 23234 28748
rect 23276 28708 23316 28748
rect 23358 28708 23398 28748
rect 23440 28708 23480 28748
rect 27112 28708 27152 28748
rect 27194 28708 27234 28748
rect 27276 28708 27316 28748
rect 27358 28708 27398 28748
rect 27440 28708 27480 28748
rect 31112 28708 31152 28748
rect 31194 28708 31234 28748
rect 31276 28708 31316 28748
rect 31358 28708 31398 28748
rect 31440 28708 31480 28748
rect 35112 28708 35152 28748
rect 35194 28708 35234 28748
rect 35276 28708 35316 28748
rect 35358 28708 35398 28748
rect 35440 28708 35480 28748
rect 39112 28708 39152 28748
rect 39194 28708 39234 28748
rect 39276 28708 39316 28748
rect 39358 28708 39398 28748
rect 39440 28708 39480 28748
rect 43112 28708 43152 28748
rect 43194 28708 43234 28748
rect 43276 28708 43316 28748
rect 43358 28708 43398 28748
rect 43440 28708 43480 28748
rect 47112 28708 47152 28748
rect 47194 28708 47234 28748
rect 47276 28708 47316 28748
rect 47358 28708 47398 28748
rect 47440 28708 47480 28748
rect 51112 28708 51152 28748
rect 51194 28708 51234 28748
rect 51276 28708 51316 28748
rect 51358 28708 51398 28748
rect 51440 28708 51480 28748
rect 55112 28708 55152 28748
rect 55194 28708 55234 28748
rect 55276 28708 55316 28748
rect 55358 28708 55398 28748
rect 55440 28708 55480 28748
rect 59112 28708 59152 28748
rect 59194 28708 59234 28748
rect 59276 28708 59316 28748
rect 59358 28708 59398 28748
rect 59440 28708 59480 28748
rect 63112 28708 63152 28748
rect 63194 28708 63234 28748
rect 63276 28708 63316 28748
rect 63358 28708 63398 28748
rect 63440 28708 63480 28748
rect 67112 28708 67152 28748
rect 67194 28708 67234 28748
rect 67276 28708 67316 28748
rect 67358 28708 67398 28748
rect 67440 28708 67480 28748
rect 4352 27952 4392 27992
rect 4434 27952 4474 27992
rect 4516 27952 4556 27992
rect 4598 27952 4638 27992
rect 4680 27952 4720 27992
rect 8352 27952 8392 27992
rect 8434 27952 8474 27992
rect 8516 27952 8556 27992
rect 8598 27952 8638 27992
rect 8680 27952 8720 27992
rect 12352 27952 12392 27992
rect 12434 27952 12474 27992
rect 12516 27952 12556 27992
rect 12598 27952 12638 27992
rect 12680 27952 12720 27992
rect 16352 27952 16392 27992
rect 16434 27952 16474 27992
rect 16516 27952 16556 27992
rect 16598 27952 16638 27992
rect 16680 27952 16720 27992
rect 20352 27952 20392 27992
rect 20434 27952 20474 27992
rect 20516 27952 20556 27992
rect 20598 27952 20638 27992
rect 20680 27952 20720 27992
rect 24352 27952 24392 27992
rect 24434 27952 24474 27992
rect 24516 27952 24556 27992
rect 24598 27952 24638 27992
rect 24680 27952 24720 27992
rect 28352 27952 28392 27992
rect 28434 27952 28474 27992
rect 28516 27952 28556 27992
rect 28598 27952 28638 27992
rect 28680 27952 28720 27992
rect 32352 27952 32392 27992
rect 32434 27952 32474 27992
rect 32516 27952 32556 27992
rect 32598 27952 32638 27992
rect 32680 27952 32720 27992
rect 36352 27952 36392 27992
rect 36434 27952 36474 27992
rect 36516 27952 36556 27992
rect 36598 27952 36638 27992
rect 36680 27952 36720 27992
rect 40352 27952 40392 27992
rect 40434 27952 40474 27992
rect 40516 27952 40556 27992
rect 40598 27952 40638 27992
rect 40680 27952 40720 27992
rect 44352 27952 44392 27992
rect 44434 27952 44474 27992
rect 44516 27952 44556 27992
rect 44598 27952 44638 27992
rect 44680 27952 44720 27992
rect 48352 27952 48392 27992
rect 48434 27952 48474 27992
rect 48516 27952 48556 27992
rect 48598 27952 48638 27992
rect 48680 27952 48720 27992
rect 52352 27952 52392 27992
rect 52434 27952 52474 27992
rect 52516 27952 52556 27992
rect 52598 27952 52638 27992
rect 52680 27952 52720 27992
rect 56352 27952 56392 27992
rect 56434 27952 56474 27992
rect 56516 27952 56556 27992
rect 56598 27952 56638 27992
rect 56680 27952 56720 27992
rect 60352 27952 60392 27992
rect 60434 27952 60474 27992
rect 60516 27952 60556 27992
rect 60598 27952 60638 27992
rect 60680 27952 60720 27992
rect 64352 27952 64392 27992
rect 64434 27952 64474 27992
rect 64516 27952 64556 27992
rect 64598 27952 64638 27992
rect 64680 27952 64720 27992
rect 68352 27952 68392 27992
rect 68434 27952 68474 27992
rect 68516 27952 68556 27992
rect 68598 27952 68638 27992
rect 68680 27952 68720 27992
rect 3112 27196 3152 27236
rect 3194 27196 3234 27236
rect 3276 27196 3316 27236
rect 3358 27196 3398 27236
rect 3440 27196 3480 27236
rect 7112 27196 7152 27236
rect 7194 27196 7234 27236
rect 7276 27196 7316 27236
rect 7358 27196 7398 27236
rect 7440 27196 7480 27236
rect 11112 27196 11152 27236
rect 11194 27196 11234 27236
rect 11276 27196 11316 27236
rect 11358 27196 11398 27236
rect 11440 27196 11480 27236
rect 15112 27196 15152 27236
rect 15194 27196 15234 27236
rect 15276 27196 15316 27236
rect 15358 27196 15398 27236
rect 15440 27196 15480 27236
rect 19112 27196 19152 27236
rect 19194 27196 19234 27236
rect 19276 27196 19316 27236
rect 19358 27196 19398 27236
rect 19440 27196 19480 27236
rect 23112 27196 23152 27236
rect 23194 27196 23234 27236
rect 23276 27196 23316 27236
rect 23358 27196 23398 27236
rect 23440 27196 23480 27236
rect 27112 27196 27152 27236
rect 27194 27196 27234 27236
rect 27276 27196 27316 27236
rect 27358 27196 27398 27236
rect 27440 27196 27480 27236
rect 31112 27196 31152 27236
rect 31194 27196 31234 27236
rect 31276 27196 31316 27236
rect 31358 27196 31398 27236
rect 31440 27196 31480 27236
rect 35112 27196 35152 27236
rect 35194 27196 35234 27236
rect 35276 27196 35316 27236
rect 35358 27196 35398 27236
rect 35440 27196 35480 27236
rect 39112 27196 39152 27236
rect 39194 27196 39234 27236
rect 39276 27196 39316 27236
rect 39358 27196 39398 27236
rect 39440 27196 39480 27236
rect 43112 27196 43152 27236
rect 43194 27196 43234 27236
rect 43276 27196 43316 27236
rect 43358 27196 43398 27236
rect 43440 27196 43480 27236
rect 47112 27196 47152 27236
rect 47194 27196 47234 27236
rect 47276 27196 47316 27236
rect 47358 27196 47398 27236
rect 47440 27196 47480 27236
rect 51112 27196 51152 27236
rect 51194 27196 51234 27236
rect 51276 27196 51316 27236
rect 51358 27196 51398 27236
rect 51440 27196 51480 27236
rect 55112 27196 55152 27236
rect 55194 27196 55234 27236
rect 55276 27196 55316 27236
rect 55358 27196 55398 27236
rect 55440 27196 55480 27236
rect 59112 27196 59152 27236
rect 59194 27196 59234 27236
rect 59276 27196 59316 27236
rect 59358 27196 59398 27236
rect 59440 27196 59480 27236
rect 63112 27196 63152 27236
rect 63194 27196 63234 27236
rect 63276 27196 63316 27236
rect 63358 27196 63398 27236
rect 63440 27196 63480 27236
rect 67112 27196 67152 27236
rect 67194 27196 67234 27236
rect 67276 27196 67316 27236
rect 67358 27196 67398 27236
rect 67440 27196 67480 27236
rect 71884 26524 71924 26564
rect 73228 26524 73268 26564
rect 4352 26440 4392 26480
rect 4434 26440 4474 26480
rect 4516 26440 4556 26480
rect 4598 26440 4638 26480
rect 4680 26440 4720 26480
rect 8352 26440 8392 26480
rect 8434 26440 8474 26480
rect 8516 26440 8556 26480
rect 8598 26440 8638 26480
rect 8680 26440 8720 26480
rect 12352 26440 12392 26480
rect 12434 26440 12474 26480
rect 12516 26440 12556 26480
rect 12598 26440 12638 26480
rect 12680 26440 12720 26480
rect 16352 26440 16392 26480
rect 16434 26440 16474 26480
rect 16516 26440 16556 26480
rect 16598 26440 16638 26480
rect 16680 26440 16720 26480
rect 20352 26440 20392 26480
rect 20434 26440 20474 26480
rect 20516 26440 20556 26480
rect 20598 26440 20638 26480
rect 20680 26440 20720 26480
rect 24352 26440 24392 26480
rect 24434 26440 24474 26480
rect 24516 26440 24556 26480
rect 24598 26440 24638 26480
rect 24680 26440 24720 26480
rect 28352 26440 28392 26480
rect 28434 26440 28474 26480
rect 28516 26440 28556 26480
rect 28598 26440 28638 26480
rect 28680 26440 28720 26480
rect 32352 26440 32392 26480
rect 32434 26440 32474 26480
rect 32516 26440 32556 26480
rect 32598 26440 32638 26480
rect 32680 26440 32720 26480
rect 36352 26440 36392 26480
rect 36434 26440 36474 26480
rect 36516 26440 36556 26480
rect 36598 26440 36638 26480
rect 36680 26440 36720 26480
rect 40352 26440 40392 26480
rect 40434 26440 40474 26480
rect 40516 26440 40556 26480
rect 40598 26440 40638 26480
rect 40680 26440 40720 26480
rect 44352 26440 44392 26480
rect 44434 26440 44474 26480
rect 44516 26440 44556 26480
rect 44598 26440 44638 26480
rect 44680 26440 44720 26480
rect 48352 26440 48392 26480
rect 48434 26440 48474 26480
rect 48516 26440 48556 26480
rect 48598 26440 48638 26480
rect 48680 26440 48720 26480
rect 52352 26440 52392 26480
rect 52434 26440 52474 26480
rect 52516 26440 52556 26480
rect 52598 26440 52638 26480
rect 52680 26440 52720 26480
rect 56352 26440 56392 26480
rect 56434 26440 56474 26480
rect 56516 26440 56556 26480
rect 56598 26440 56638 26480
rect 56680 26440 56720 26480
rect 60352 26440 60392 26480
rect 60434 26440 60474 26480
rect 60516 26440 60556 26480
rect 60598 26440 60638 26480
rect 60680 26440 60720 26480
rect 64352 26440 64392 26480
rect 64434 26440 64474 26480
rect 64516 26440 64556 26480
rect 64598 26440 64638 26480
rect 64680 26440 64720 26480
rect 68352 26440 68392 26480
rect 68434 26440 68474 26480
rect 68516 26440 68556 26480
rect 68598 26440 68638 26480
rect 68680 26440 68720 26480
rect 3112 25684 3152 25724
rect 3194 25684 3234 25724
rect 3276 25684 3316 25724
rect 3358 25684 3398 25724
rect 3440 25684 3480 25724
rect 7112 25684 7152 25724
rect 7194 25684 7234 25724
rect 7276 25684 7316 25724
rect 7358 25684 7398 25724
rect 7440 25684 7480 25724
rect 11112 25684 11152 25724
rect 11194 25684 11234 25724
rect 11276 25684 11316 25724
rect 11358 25684 11398 25724
rect 11440 25684 11480 25724
rect 15112 25684 15152 25724
rect 15194 25684 15234 25724
rect 15276 25684 15316 25724
rect 15358 25684 15398 25724
rect 15440 25684 15480 25724
rect 19112 25684 19152 25724
rect 19194 25684 19234 25724
rect 19276 25684 19316 25724
rect 19358 25684 19398 25724
rect 19440 25684 19480 25724
rect 23112 25684 23152 25724
rect 23194 25684 23234 25724
rect 23276 25684 23316 25724
rect 23358 25684 23398 25724
rect 23440 25684 23480 25724
rect 27112 25684 27152 25724
rect 27194 25684 27234 25724
rect 27276 25684 27316 25724
rect 27358 25684 27398 25724
rect 27440 25684 27480 25724
rect 31112 25684 31152 25724
rect 31194 25684 31234 25724
rect 31276 25684 31316 25724
rect 31358 25684 31398 25724
rect 31440 25684 31480 25724
rect 35112 25684 35152 25724
rect 35194 25684 35234 25724
rect 35276 25684 35316 25724
rect 35358 25684 35398 25724
rect 35440 25684 35480 25724
rect 39112 25684 39152 25724
rect 39194 25684 39234 25724
rect 39276 25684 39316 25724
rect 39358 25684 39398 25724
rect 39440 25684 39480 25724
rect 43112 25684 43152 25724
rect 43194 25684 43234 25724
rect 43276 25684 43316 25724
rect 43358 25684 43398 25724
rect 43440 25684 43480 25724
rect 47112 25684 47152 25724
rect 47194 25684 47234 25724
rect 47276 25684 47316 25724
rect 47358 25684 47398 25724
rect 47440 25684 47480 25724
rect 51112 25684 51152 25724
rect 51194 25684 51234 25724
rect 51276 25684 51316 25724
rect 51358 25684 51398 25724
rect 51440 25684 51480 25724
rect 55112 25684 55152 25724
rect 55194 25684 55234 25724
rect 55276 25684 55316 25724
rect 55358 25684 55398 25724
rect 55440 25684 55480 25724
rect 59112 25684 59152 25724
rect 59194 25684 59234 25724
rect 59276 25684 59316 25724
rect 59358 25684 59398 25724
rect 59440 25684 59480 25724
rect 63112 25684 63152 25724
rect 63194 25684 63234 25724
rect 63276 25684 63316 25724
rect 63358 25684 63398 25724
rect 63440 25684 63480 25724
rect 67112 25684 67152 25724
rect 67194 25684 67234 25724
rect 67276 25684 67316 25724
rect 67358 25684 67398 25724
rect 67440 25684 67480 25724
rect 4352 24928 4392 24968
rect 4434 24928 4474 24968
rect 4516 24928 4556 24968
rect 4598 24928 4638 24968
rect 4680 24928 4720 24968
rect 8352 24928 8392 24968
rect 8434 24928 8474 24968
rect 8516 24928 8556 24968
rect 8598 24928 8638 24968
rect 8680 24928 8720 24968
rect 12352 24928 12392 24968
rect 12434 24928 12474 24968
rect 12516 24928 12556 24968
rect 12598 24928 12638 24968
rect 12680 24928 12720 24968
rect 16352 24928 16392 24968
rect 16434 24928 16474 24968
rect 16516 24928 16556 24968
rect 16598 24928 16638 24968
rect 16680 24928 16720 24968
rect 20352 24928 20392 24968
rect 20434 24928 20474 24968
rect 20516 24928 20556 24968
rect 20598 24928 20638 24968
rect 20680 24928 20720 24968
rect 24352 24928 24392 24968
rect 24434 24928 24474 24968
rect 24516 24928 24556 24968
rect 24598 24928 24638 24968
rect 24680 24928 24720 24968
rect 28352 24928 28392 24968
rect 28434 24928 28474 24968
rect 28516 24928 28556 24968
rect 28598 24928 28638 24968
rect 28680 24928 28720 24968
rect 32352 24928 32392 24968
rect 32434 24928 32474 24968
rect 32516 24928 32556 24968
rect 32598 24928 32638 24968
rect 32680 24928 32720 24968
rect 36352 24928 36392 24968
rect 36434 24928 36474 24968
rect 36516 24928 36556 24968
rect 36598 24928 36638 24968
rect 36680 24928 36720 24968
rect 40352 24928 40392 24968
rect 40434 24928 40474 24968
rect 40516 24928 40556 24968
rect 40598 24928 40638 24968
rect 40680 24928 40720 24968
rect 44352 24928 44392 24968
rect 44434 24928 44474 24968
rect 44516 24928 44556 24968
rect 44598 24928 44638 24968
rect 44680 24928 44720 24968
rect 48352 24928 48392 24968
rect 48434 24928 48474 24968
rect 48516 24928 48556 24968
rect 48598 24928 48638 24968
rect 48680 24928 48720 24968
rect 52352 24928 52392 24968
rect 52434 24928 52474 24968
rect 52516 24928 52556 24968
rect 52598 24928 52638 24968
rect 52680 24928 52720 24968
rect 56352 24928 56392 24968
rect 56434 24928 56474 24968
rect 56516 24928 56556 24968
rect 56598 24928 56638 24968
rect 56680 24928 56720 24968
rect 60352 24928 60392 24968
rect 60434 24928 60474 24968
rect 60516 24928 60556 24968
rect 60598 24928 60638 24968
rect 60680 24928 60720 24968
rect 64352 24928 64392 24968
rect 64434 24928 64474 24968
rect 64516 24928 64556 24968
rect 64598 24928 64638 24968
rect 64680 24928 64720 24968
rect 68352 24928 68392 24968
rect 68434 24928 68474 24968
rect 68516 24928 68556 24968
rect 68598 24928 68638 24968
rect 68680 24928 68720 24968
rect 85708 25348 85748 25388
rect 86860 25348 86900 25388
rect 3112 24172 3152 24212
rect 3194 24172 3234 24212
rect 3276 24172 3316 24212
rect 3358 24172 3398 24212
rect 3440 24172 3480 24212
rect 7112 24172 7152 24212
rect 7194 24172 7234 24212
rect 7276 24172 7316 24212
rect 7358 24172 7398 24212
rect 7440 24172 7480 24212
rect 11112 24172 11152 24212
rect 11194 24172 11234 24212
rect 11276 24172 11316 24212
rect 11358 24172 11398 24212
rect 11440 24172 11480 24212
rect 15112 24172 15152 24212
rect 15194 24172 15234 24212
rect 15276 24172 15316 24212
rect 15358 24172 15398 24212
rect 15440 24172 15480 24212
rect 19112 24172 19152 24212
rect 19194 24172 19234 24212
rect 19276 24172 19316 24212
rect 19358 24172 19398 24212
rect 19440 24172 19480 24212
rect 23112 24172 23152 24212
rect 23194 24172 23234 24212
rect 23276 24172 23316 24212
rect 23358 24172 23398 24212
rect 23440 24172 23480 24212
rect 27112 24172 27152 24212
rect 27194 24172 27234 24212
rect 27276 24172 27316 24212
rect 27358 24172 27398 24212
rect 27440 24172 27480 24212
rect 31112 24172 31152 24212
rect 31194 24172 31234 24212
rect 31276 24172 31316 24212
rect 31358 24172 31398 24212
rect 31440 24172 31480 24212
rect 35112 24172 35152 24212
rect 35194 24172 35234 24212
rect 35276 24172 35316 24212
rect 35358 24172 35398 24212
rect 35440 24172 35480 24212
rect 39112 24172 39152 24212
rect 39194 24172 39234 24212
rect 39276 24172 39316 24212
rect 39358 24172 39398 24212
rect 39440 24172 39480 24212
rect 43112 24172 43152 24212
rect 43194 24172 43234 24212
rect 43276 24172 43316 24212
rect 43358 24172 43398 24212
rect 43440 24172 43480 24212
rect 47112 24172 47152 24212
rect 47194 24172 47234 24212
rect 47276 24172 47316 24212
rect 47358 24172 47398 24212
rect 47440 24172 47480 24212
rect 51112 24172 51152 24212
rect 51194 24172 51234 24212
rect 51276 24172 51316 24212
rect 51358 24172 51398 24212
rect 51440 24172 51480 24212
rect 55112 24172 55152 24212
rect 55194 24172 55234 24212
rect 55276 24172 55316 24212
rect 55358 24172 55398 24212
rect 55440 24172 55480 24212
rect 59112 24172 59152 24212
rect 59194 24172 59234 24212
rect 59276 24172 59316 24212
rect 59358 24172 59398 24212
rect 59440 24172 59480 24212
rect 63112 24172 63152 24212
rect 63194 24172 63234 24212
rect 63276 24172 63316 24212
rect 63358 24172 63398 24212
rect 63440 24172 63480 24212
rect 67112 24172 67152 24212
rect 67194 24172 67234 24212
rect 67276 24172 67316 24212
rect 67358 24172 67398 24212
rect 67440 24172 67480 24212
rect 71112 24172 71152 24212
rect 71194 24172 71234 24212
rect 71276 24172 71316 24212
rect 71358 24172 71398 24212
rect 71440 24172 71480 24212
rect 75112 24172 75152 24212
rect 75194 24172 75234 24212
rect 75276 24172 75316 24212
rect 75358 24172 75398 24212
rect 75440 24172 75480 24212
rect 79112 24172 79152 24212
rect 79194 24172 79234 24212
rect 79276 24172 79316 24212
rect 79358 24172 79398 24212
rect 79440 24172 79480 24212
rect 83112 24172 83152 24212
rect 83194 24172 83234 24212
rect 83276 24172 83316 24212
rect 83358 24172 83398 24212
rect 83440 24172 83480 24212
rect 87112 24172 87152 24212
rect 87194 24172 87234 24212
rect 87276 24172 87316 24212
rect 87358 24172 87398 24212
rect 87440 24172 87480 24212
rect 91112 24172 91152 24212
rect 91194 24172 91234 24212
rect 91276 24172 91316 24212
rect 91358 24172 91398 24212
rect 91440 24172 91480 24212
rect 95112 24172 95152 24212
rect 95194 24172 95234 24212
rect 95276 24172 95316 24212
rect 95358 24172 95398 24212
rect 95440 24172 95480 24212
rect 99112 24172 99152 24212
rect 99194 24172 99234 24212
rect 99276 24172 99316 24212
rect 99358 24172 99398 24212
rect 99440 24172 99480 24212
rect 4352 23416 4392 23456
rect 4434 23416 4474 23456
rect 4516 23416 4556 23456
rect 4598 23416 4638 23456
rect 4680 23416 4720 23456
rect 8352 23416 8392 23456
rect 8434 23416 8474 23456
rect 8516 23416 8556 23456
rect 8598 23416 8638 23456
rect 8680 23416 8720 23456
rect 12352 23416 12392 23456
rect 12434 23416 12474 23456
rect 12516 23416 12556 23456
rect 12598 23416 12638 23456
rect 12680 23416 12720 23456
rect 16352 23416 16392 23456
rect 16434 23416 16474 23456
rect 16516 23416 16556 23456
rect 16598 23416 16638 23456
rect 16680 23416 16720 23456
rect 20352 23416 20392 23456
rect 20434 23416 20474 23456
rect 20516 23416 20556 23456
rect 20598 23416 20638 23456
rect 20680 23416 20720 23456
rect 24352 23416 24392 23456
rect 24434 23416 24474 23456
rect 24516 23416 24556 23456
rect 24598 23416 24638 23456
rect 24680 23416 24720 23456
rect 28352 23416 28392 23456
rect 28434 23416 28474 23456
rect 28516 23416 28556 23456
rect 28598 23416 28638 23456
rect 28680 23416 28720 23456
rect 32352 23416 32392 23456
rect 32434 23416 32474 23456
rect 32516 23416 32556 23456
rect 32598 23416 32638 23456
rect 32680 23416 32720 23456
rect 36352 23416 36392 23456
rect 36434 23416 36474 23456
rect 36516 23416 36556 23456
rect 36598 23416 36638 23456
rect 36680 23416 36720 23456
rect 40352 23416 40392 23456
rect 40434 23416 40474 23456
rect 40516 23416 40556 23456
rect 40598 23416 40638 23456
rect 40680 23416 40720 23456
rect 44352 23416 44392 23456
rect 44434 23416 44474 23456
rect 44516 23416 44556 23456
rect 44598 23416 44638 23456
rect 44680 23416 44720 23456
rect 48352 23416 48392 23456
rect 48434 23416 48474 23456
rect 48516 23416 48556 23456
rect 48598 23416 48638 23456
rect 48680 23416 48720 23456
rect 52352 23416 52392 23456
rect 52434 23416 52474 23456
rect 52516 23416 52556 23456
rect 52598 23416 52638 23456
rect 52680 23416 52720 23456
rect 56352 23416 56392 23456
rect 56434 23416 56474 23456
rect 56516 23416 56556 23456
rect 56598 23416 56638 23456
rect 56680 23416 56720 23456
rect 60352 23416 60392 23456
rect 60434 23416 60474 23456
rect 60516 23416 60556 23456
rect 60598 23416 60638 23456
rect 60680 23416 60720 23456
rect 64352 23416 64392 23456
rect 64434 23416 64474 23456
rect 64516 23416 64556 23456
rect 64598 23416 64638 23456
rect 64680 23416 64720 23456
rect 68352 23416 68392 23456
rect 68434 23416 68474 23456
rect 68516 23416 68556 23456
rect 68598 23416 68638 23456
rect 68680 23416 68720 23456
rect 72352 23416 72392 23456
rect 72434 23416 72474 23456
rect 72516 23416 72556 23456
rect 72598 23416 72638 23456
rect 72680 23416 72720 23456
rect 76352 23416 76392 23456
rect 76434 23416 76474 23456
rect 76516 23416 76556 23456
rect 76598 23416 76638 23456
rect 76680 23416 76720 23456
rect 80352 23416 80392 23456
rect 80434 23416 80474 23456
rect 80516 23416 80556 23456
rect 80598 23416 80638 23456
rect 80680 23416 80720 23456
rect 84352 23416 84392 23456
rect 84434 23416 84474 23456
rect 84516 23416 84556 23456
rect 84598 23416 84638 23456
rect 84680 23416 84720 23456
rect 88352 23416 88392 23456
rect 88434 23416 88474 23456
rect 88516 23416 88556 23456
rect 88598 23416 88638 23456
rect 88680 23416 88720 23456
rect 92352 23416 92392 23456
rect 92434 23416 92474 23456
rect 92516 23416 92556 23456
rect 92598 23416 92638 23456
rect 92680 23416 92720 23456
rect 96352 23416 96392 23456
rect 96434 23416 96474 23456
rect 96516 23416 96556 23456
rect 96598 23416 96638 23456
rect 96680 23416 96720 23456
rect 3112 22660 3152 22700
rect 3194 22660 3234 22700
rect 3276 22660 3316 22700
rect 3358 22660 3398 22700
rect 3440 22660 3480 22700
rect 7112 22660 7152 22700
rect 7194 22660 7234 22700
rect 7276 22660 7316 22700
rect 7358 22660 7398 22700
rect 7440 22660 7480 22700
rect 11112 22660 11152 22700
rect 11194 22660 11234 22700
rect 11276 22660 11316 22700
rect 11358 22660 11398 22700
rect 11440 22660 11480 22700
rect 15112 22660 15152 22700
rect 15194 22660 15234 22700
rect 15276 22660 15316 22700
rect 15358 22660 15398 22700
rect 15440 22660 15480 22700
rect 19112 22660 19152 22700
rect 19194 22660 19234 22700
rect 19276 22660 19316 22700
rect 19358 22660 19398 22700
rect 19440 22660 19480 22700
rect 23112 22660 23152 22700
rect 23194 22660 23234 22700
rect 23276 22660 23316 22700
rect 23358 22660 23398 22700
rect 23440 22660 23480 22700
rect 27112 22660 27152 22700
rect 27194 22660 27234 22700
rect 27276 22660 27316 22700
rect 27358 22660 27398 22700
rect 27440 22660 27480 22700
rect 31112 22660 31152 22700
rect 31194 22660 31234 22700
rect 31276 22660 31316 22700
rect 31358 22660 31398 22700
rect 31440 22660 31480 22700
rect 35112 22660 35152 22700
rect 35194 22660 35234 22700
rect 35276 22660 35316 22700
rect 35358 22660 35398 22700
rect 35440 22660 35480 22700
rect 39112 22660 39152 22700
rect 39194 22660 39234 22700
rect 39276 22660 39316 22700
rect 39358 22660 39398 22700
rect 39440 22660 39480 22700
rect 43112 22660 43152 22700
rect 43194 22660 43234 22700
rect 43276 22660 43316 22700
rect 43358 22660 43398 22700
rect 43440 22660 43480 22700
rect 47112 22660 47152 22700
rect 47194 22660 47234 22700
rect 47276 22660 47316 22700
rect 47358 22660 47398 22700
rect 47440 22660 47480 22700
rect 51112 22660 51152 22700
rect 51194 22660 51234 22700
rect 51276 22660 51316 22700
rect 51358 22660 51398 22700
rect 51440 22660 51480 22700
rect 55112 22660 55152 22700
rect 55194 22660 55234 22700
rect 55276 22660 55316 22700
rect 55358 22660 55398 22700
rect 55440 22660 55480 22700
rect 59112 22660 59152 22700
rect 59194 22660 59234 22700
rect 59276 22660 59316 22700
rect 59358 22660 59398 22700
rect 59440 22660 59480 22700
rect 63112 22660 63152 22700
rect 63194 22660 63234 22700
rect 63276 22660 63316 22700
rect 63358 22660 63398 22700
rect 63440 22660 63480 22700
rect 67112 22660 67152 22700
rect 67194 22660 67234 22700
rect 67276 22660 67316 22700
rect 67358 22660 67398 22700
rect 67440 22660 67480 22700
rect 71112 22660 71152 22700
rect 71194 22660 71234 22700
rect 71276 22660 71316 22700
rect 71358 22660 71398 22700
rect 71440 22660 71480 22700
rect 75112 22660 75152 22700
rect 75194 22660 75234 22700
rect 75276 22660 75316 22700
rect 75358 22660 75398 22700
rect 75440 22660 75480 22700
rect 79112 22660 79152 22700
rect 79194 22660 79234 22700
rect 79276 22660 79316 22700
rect 79358 22660 79398 22700
rect 79440 22660 79480 22700
rect 83112 22660 83152 22700
rect 83194 22660 83234 22700
rect 83276 22660 83316 22700
rect 83358 22660 83398 22700
rect 83440 22660 83480 22700
rect 87112 22660 87152 22700
rect 87194 22660 87234 22700
rect 87276 22660 87316 22700
rect 87358 22660 87398 22700
rect 87440 22660 87480 22700
rect 91112 22660 91152 22700
rect 91194 22660 91234 22700
rect 91276 22660 91316 22700
rect 91358 22660 91398 22700
rect 91440 22660 91480 22700
rect 95112 22660 95152 22700
rect 95194 22660 95234 22700
rect 95276 22660 95316 22700
rect 95358 22660 95398 22700
rect 95440 22660 95480 22700
rect 99112 22660 99152 22700
rect 99194 22660 99234 22700
rect 99276 22660 99316 22700
rect 99358 22660 99398 22700
rect 99440 22660 99480 22700
rect 4352 21904 4392 21944
rect 4434 21904 4474 21944
rect 4516 21904 4556 21944
rect 4598 21904 4638 21944
rect 4680 21904 4720 21944
rect 8352 21904 8392 21944
rect 8434 21904 8474 21944
rect 8516 21904 8556 21944
rect 8598 21904 8638 21944
rect 8680 21904 8720 21944
rect 12352 21904 12392 21944
rect 12434 21904 12474 21944
rect 12516 21904 12556 21944
rect 12598 21904 12638 21944
rect 12680 21904 12720 21944
rect 16352 21904 16392 21944
rect 16434 21904 16474 21944
rect 16516 21904 16556 21944
rect 16598 21904 16638 21944
rect 16680 21904 16720 21944
rect 20352 21904 20392 21944
rect 20434 21904 20474 21944
rect 20516 21904 20556 21944
rect 20598 21904 20638 21944
rect 20680 21904 20720 21944
rect 24352 21904 24392 21944
rect 24434 21904 24474 21944
rect 24516 21904 24556 21944
rect 24598 21904 24638 21944
rect 24680 21904 24720 21944
rect 28352 21904 28392 21944
rect 28434 21904 28474 21944
rect 28516 21904 28556 21944
rect 28598 21904 28638 21944
rect 28680 21904 28720 21944
rect 32352 21904 32392 21944
rect 32434 21904 32474 21944
rect 32516 21904 32556 21944
rect 32598 21904 32638 21944
rect 32680 21904 32720 21944
rect 36352 21904 36392 21944
rect 36434 21904 36474 21944
rect 36516 21904 36556 21944
rect 36598 21904 36638 21944
rect 36680 21904 36720 21944
rect 40352 21904 40392 21944
rect 40434 21904 40474 21944
rect 40516 21904 40556 21944
rect 40598 21904 40638 21944
rect 40680 21904 40720 21944
rect 44352 21904 44392 21944
rect 44434 21904 44474 21944
rect 44516 21904 44556 21944
rect 44598 21904 44638 21944
rect 44680 21904 44720 21944
rect 48352 21904 48392 21944
rect 48434 21904 48474 21944
rect 48516 21904 48556 21944
rect 48598 21904 48638 21944
rect 48680 21904 48720 21944
rect 52352 21904 52392 21944
rect 52434 21904 52474 21944
rect 52516 21904 52556 21944
rect 52598 21904 52638 21944
rect 52680 21904 52720 21944
rect 56352 21904 56392 21944
rect 56434 21904 56474 21944
rect 56516 21904 56556 21944
rect 56598 21904 56638 21944
rect 56680 21904 56720 21944
rect 60352 21904 60392 21944
rect 60434 21904 60474 21944
rect 60516 21904 60556 21944
rect 60598 21904 60638 21944
rect 60680 21904 60720 21944
rect 64352 21904 64392 21944
rect 64434 21904 64474 21944
rect 64516 21904 64556 21944
rect 64598 21904 64638 21944
rect 64680 21904 64720 21944
rect 68352 21904 68392 21944
rect 68434 21904 68474 21944
rect 68516 21904 68556 21944
rect 68598 21904 68638 21944
rect 68680 21904 68720 21944
rect 72352 21904 72392 21944
rect 72434 21904 72474 21944
rect 72516 21904 72556 21944
rect 72598 21904 72638 21944
rect 72680 21904 72720 21944
rect 76352 21904 76392 21944
rect 76434 21904 76474 21944
rect 76516 21904 76556 21944
rect 76598 21904 76638 21944
rect 76680 21904 76720 21944
rect 80352 21904 80392 21944
rect 80434 21904 80474 21944
rect 80516 21904 80556 21944
rect 80598 21904 80638 21944
rect 80680 21904 80720 21944
rect 84352 21904 84392 21944
rect 84434 21904 84474 21944
rect 84516 21904 84556 21944
rect 84598 21904 84638 21944
rect 84680 21904 84720 21944
rect 88352 21904 88392 21944
rect 88434 21904 88474 21944
rect 88516 21904 88556 21944
rect 88598 21904 88638 21944
rect 88680 21904 88720 21944
rect 92352 21904 92392 21944
rect 92434 21904 92474 21944
rect 92516 21904 92556 21944
rect 92598 21904 92638 21944
rect 92680 21904 92720 21944
rect 96352 21904 96392 21944
rect 96434 21904 96474 21944
rect 96516 21904 96556 21944
rect 96598 21904 96638 21944
rect 96680 21904 96720 21944
rect 3112 21148 3152 21188
rect 3194 21148 3234 21188
rect 3276 21148 3316 21188
rect 3358 21148 3398 21188
rect 3440 21148 3480 21188
rect 7112 21148 7152 21188
rect 7194 21148 7234 21188
rect 7276 21148 7316 21188
rect 7358 21148 7398 21188
rect 7440 21148 7480 21188
rect 11112 21148 11152 21188
rect 11194 21148 11234 21188
rect 11276 21148 11316 21188
rect 11358 21148 11398 21188
rect 11440 21148 11480 21188
rect 15112 21148 15152 21188
rect 15194 21148 15234 21188
rect 15276 21148 15316 21188
rect 15358 21148 15398 21188
rect 15440 21148 15480 21188
rect 19112 21148 19152 21188
rect 19194 21148 19234 21188
rect 19276 21148 19316 21188
rect 19358 21148 19398 21188
rect 19440 21148 19480 21188
rect 23112 21148 23152 21188
rect 23194 21148 23234 21188
rect 23276 21148 23316 21188
rect 23358 21148 23398 21188
rect 23440 21148 23480 21188
rect 27112 21148 27152 21188
rect 27194 21148 27234 21188
rect 27276 21148 27316 21188
rect 27358 21148 27398 21188
rect 27440 21148 27480 21188
rect 31112 21148 31152 21188
rect 31194 21148 31234 21188
rect 31276 21148 31316 21188
rect 31358 21148 31398 21188
rect 31440 21148 31480 21188
rect 35112 21148 35152 21188
rect 35194 21148 35234 21188
rect 35276 21148 35316 21188
rect 35358 21148 35398 21188
rect 35440 21148 35480 21188
rect 39112 21148 39152 21188
rect 39194 21148 39234 21188
rect 39276 21148 39316 21188
rect 39358 21148 39398 21188
rect 39440 21148 39480 21188
rect 43112 21148 43152 21188
rect 43194 21148 43234 21188
rect 43276 21148 43316 21188
rect 43358 21148 43398 21188
rect 43440 21148 43480 21188
rect 47112 21148 47152 21188
rect 47194 21148 47234 21188
rect 47276 21148 47316 21188
rect 47358 21148 47398 21188
rect 47440 21148 47480 21188
rect 51112 21148 51152 21188
rect 51194 21148 51234 21188
rect 51276 21148 51316 21188
rect 51358 21148 51398 21188
rect 51440 21148 51480 21188
rect 55112 21148 55152 21188
rect 55194 21148 55234 21188
rect 55276 21148 55316 21188
rect 55358 21148 55398 21188
rect 55440 21148 55480 21188
rect 59112 21148 59152 21188
rect 59194 21148 59234 21188
rect 59276 21148 59316 21188
rect 59358 21148 59398 21188
rect 59440 21148 59480 21188
rect 63112 21148 63152 21188
rect 63194 21148 63234 21188
rect 63276 21148 63316 21188
rect 63358 21148 63398 21188
rect 63440 21148 63480 21188
rect 67112 21148 67152 21188
rect 67194 21148 67234 21188
rect 67276 21148 67316 21188
rect 67358 21148 67398 21188
rect 67440 21148 67480 21188
rect 71112 21148 71152 21188
rect 71194 21148 71234 21188
rect 71276 21148 71316 21188
rect 71358 21148 71398 21188
rect 71440 21148 71480 21188
rect 75112 21148 75152 21188
rect 75194 21148 75234 21188
rect 75276 21148 75316 21188
rect 75358 21148 75398 21188
rect 75440 21148 75480 21188
rect 79112 21148 79152 21188
rect 79194 21148 79234 21188
rect 79276 21148 79316 21188
rect 79358 21148 79398 21188
rect 79440 21148 79480 21188
rect 83112 21148 83152 21188
rect 83194 21148 83234 21188
rect 83276 21148 83316 21188
rect 83358 21148 83398 21188
rect 83440 21148 83480 21188
rect 87112 21148 87152 21188
rect 87194 21148 87234 21188
rect 87276 21148 87316 21188
rect 87358 21148 87398 21188
rect 87440 21148 87480 21188
rect 91112 21148 91152 21188
rect 91194 21148 91234 21188
rect 91276 21148 91316 21188
rect 91358 21148 91398 21188
rect 91440 21148 91480 21188
rect 95112 21148 95152 21188
rect 95194 21148 95234 21188
rect 95276 21148 95316 21188
rect 95358 21148 95398 21188
rect 95440 21148 95480 21188
rect 99112 21148 99152 21188
rect 99194 21148 99234 21188
rect 99276 21148 99316 21188
rect 99358 21148 99398 21188
rect 99440 21148 99480 21188
rect 4352 20392 4392 20432
rect 4434 20392 4474 20432
rect 4516 20392 4556 20432
rect 4598 20392 4638 20432
rect 4680 20392 4720 20432
rect 8352 20392 8392 20432
rect 8434 20392 8474 20432
rect 8516 20392 8556 20432
rect 8598 20392 8638 20432
rect 8680 20392 8720 20432
rect 12352 20392 12392 20432
rect 12434 20392 12474 20432
rect 12516 20392 12556 20432
rect 12598 20392 12638 20432
rect 12680 20392 12720 20432
rect 16352 20392 16392 20432
rect 16434 20392 16474 20432
rect 16516 20392 16556 20432
rect 16598 20392 16638 20432
rect 16680 20392 16720 20432
rect 20352 20392 20392 20432
rect 20434 20392 20474 20432
rect 20516 20392 20556 20432
rect 20598 20392 20638 20432
rect 20680 20392 20720 20432
rect 24352 20392 24392 20432
rect 24434 20392 24474 20432
rect 24516 20392 24556 20432
rect 24598 20392 24638 20432
rect 24680 20392 24720 20432
rect 28352 20392 28392 20432
rect 28434 20392 28474 20432
rect 28516 20392 28556 20432
rect 28598 20392 28638 20432
rect 28680 20392 28720 20432
rect 32352 20392 32392 20432
rect 32434 20392 32474 20432
rect 32516 20392 32556 20432
rect 32598 20392 32638 20432
rect 32680 20392 32720 20432
rect 36352 20392 36392 20432
rect 36434 20392 36474 20432
rect 36516 20392 36556 20432
rect 36598 20392 36638 20432
rect 36680 20392 36720 20432
rect 40352 20392 40392 20432
rect 40434 20392 40474 20432
rect 40516 20392 40556 20432
rect 40598 20392 40638 20432
rect 40680 20392 40720 20432
rect 44352 20392 44392 20432
rect 44434 20392 44474 20432
rect 44516 20392 44556 20432
rect 44598 20392 44638 20432
rect 44680 20392 44720 20432
rect 48352 20392 48392 20432
rect 48434 20392 48474 20432
rect 48516 20392 48556 20432
rect 48598 20392 48638 20432
rect 48680 20392 48720 20432
rect 52352 20392 52392 20432
rect 52434 20392 52474 20432
rect 52516 20392 52556 20432
rect 52598 20392 52638 20432
rect 52680 20392 52720 20432
rect 56352 20392 56392 20432
rect 56434 20392 56474 20432
rect 56516 20392 56556 20432
rect 56598 20392 56638 20432
rect 56680 20392 56720 20432
rect 60352 20392 60392 20432
rect 60434 20392 60474 20432
rect 60516 20392 60556 20432
rect 60598 20392 60638 20432
rect 60680 20392 60720 20432
rect 64352 20392 64392 20432
rect 64434 20392 64474 20432
rect 64516 20392 64556 20432
rect 64598 20392 64638 20432
rect 64680 20392 64720 20432
rect 68352 20392 68392 20432
rect 68434 20392 68474 20432
rect 68516 20392 68556 20432
rect 68598 20392 68638 20432
rect 68680 20392 68720 20432
rect 72352 20392 72392 20432
rect 72434 20392 72474 20432
rect 72516 20392 72556 20432
rect 72598 20392 72638 20432
rect 72680 20392 72720 20432
rect 76352 20392 76392 20432
rect 76434 20392 76474 20432
rect 76516 20392 76556 20432
rect 76598 20392 76638 20432
rect 76680 20392 76720 20432
rect 80352 20392 80392 20432
rect 80434 20392 80474 20432
rect 80516 20392 80556 20432
rect 80598 20392 80638 20432
rect 80680 20392 80720 20432
rect 84352 20392 84392 20432
rect 84434 20392 84474 20432
rect 84516 20392 84556 20432
rect 84598 20392 84638 20432
rect 84680 20392 84720 20432
rect 88352 20392 88392 20432
rect 88434 20392 88474 20432
rect 88516 20392 88556 20432
rect 88598 20392 88638 20432
rect 88680 20392 88720 20432
rect 92352 20392 92392 20432
rect 92434 20392 92474 20432
rect 92516 20392 92556 20432
rect 92598 20392 92638 20432
rect 92680 20392 92720 20432
rect 96352 20392 96392 20432
rect 96434 20392 96474 20432
rect 96516 20392 96556 20432
rect 96598 20392 96638 20432
rect 96680 20392 96720 20432
rect 3112 19636 3152 19676
rect 3194 19636 3234 19676
rect 3276 19636 3316 19676
rect 3358 19636 3398 19676
rect 3440 19636 3480 19676
rect 7112 19636 7152 19676
rect 7194 19636 7234 19676
rect 7276 19636 7316 19676
rect 7358 19636 7398 19676
rect 7440 19636 7480 19676
rect 11112 19636 11152 19676
rect 11194 19636 11234 19676
rect 11276 19636 11316 19676
rect 11358 19636 11398 19676
rect 11440 19636 11480 19676
rect 15112 19636 15152 19676
rect 15194 19636 15234 19676
rect 15276 19636 15316 19676
rect 15358 19636 15398 19676
rect 15440 19636 15480 19676
rect 19112 19636 19152 19676
rect 19194 19636 19234 19676
rect 19276 19636 19316 19676
rect 19358 19636 19398 19676
rect 19440 19636 19480 19676
rect 23112 19636 23152 19676
rect 23194 19636 23234 19676
rect 23276 19636 23316 19676
rect 23358 19636 23398 19676
rect 23440 19636 23480 19676
rect 27112 19636 27152 19676
rect 27194 19636 27234 19676
rect 27276 19636 27316 19676
rect 27358 19636 27398 19676
rect 27440 19636 27480 19676
rect 31112 19636 31152 19676
rect 31194 19636 31234 19676
rect 31276 19636 31316 19676
rect 31358 19636 31398 19676
rect 31440 19636 31480 19676
rect 35112 19636 35152 19676
rect 35194 19636 35234 19676
rect 35276 19636 35316 19676
rect 35358 19636 35398 19676
rect 35440 19636 35480 19676
rect 39112 19636 39152 19676
rect 39194 19636 39234 19676
rect 39276 19636 39316 19676
rect 39358 19636 39398 19676
rect 39440 19636 39480 19676
rect 43112 19636 43152 19676
rect 43194 19636 43234 19676
rect 43276 19636 43316 19676
rect 43358 19636 43398 19676
rect 43440 19636 43480 19676
rect 47112 19636 47152 19676
rect 47194 19636 47234 19676
rect 47276 19636 47316 19676
rect 47358 19636 47398 19676
rect 47440 19636 47480 19676
rect 51112 19636 51152 19676
rect 51194 19636 51234 19676
rect 51276 19636 51316 19676
rect 51358 19636 51398 19676
rect 51440 19636 51480 19676
rect 55112 19636 55152 19676
rect 55194 19636 55234 19676
rect 55276 19636 55316 19676
rect 55358 19636 55398 19676
rect 55440 19636 55480 19676
rect 59112 19636 59152 19676
rect 59194 19636 59234 19676
rect 59276 19636 59316 19676
rect 59358 19636 59398 19676
rect 59440 19636 59480 19676
rect 63112 19636 63152 19676
rect 63194 19636 63234 19676
rect 63276 19636 63316 19676
rect 63358 19636 63398 19676
rect 63440 19636 63480 19676
rect 67112 19636 67152 19676
rect 67194 19636 67234 19676
rect 67276 19636 67316 19676
rect 67358 19636 67398 19676
rect 67440 19636 67480 19676
rect 71112 19636 71152 19676
rect 71194 19636 71234 19676
rect 71276 19636 71316 19676
rect 71358 19636 71398 19676
rect 71440 19636 71480 19676
rect 75112 19636 75152 19676
rect 75194 19636 75234 19676
rect 75276 19636 75316 19676
rect 75358 19636 75398 19676
rect 75440 19636 75480 19676
rect 79112 19636 79152 19676
rect 79194 19636 79234 19676
rect 79276 19636 79316 19676
rect 79358 19636 79398 19676
rect 79440 19636 79480 19676
rect 83112 19636 83152 19676
rect 83194 19636 83234 19676
rect 83276 19636 83316 19676
rect 83358 19636 83398 19676
rect 83440 19636 83480 19676
rect 87112 19636 87152 19676
rect 87194 19636 87234 19676
rect 87276 19636 87316 19676
rect 87358 19636 87398 19676
rect 87440 19636 87480 19676
rect 91112 19636 91152 19676
rect 91194 19636 91234 19676
rect 91276 19636 91316 19676
rect 91358 19636 91398 19676
rect 91440 19636 91480 19676
rect 95112 19636 95152 19676
rect 95194 19636 95234 19676
rect 95276 19636 95316 19676
rect 95358 19636 95398 19676
rect 95440 19636 95480 19676
rect 99112 19636 99152 19676
rect 99194 19636 99234 19676
rect 99276 19636 99316 19676
rect 99358 19636 99398 19676
rect 99440 19636 99480 19676
rect 4352 18880 4392 18920
rect 4434 18880 4474 18920
rect 4516 18880 4556 18920
rect 4598 18880 4638 18920
rect 4680 18880 4720 18920
rect 8352 18880 8392 18920
rect 8434 18880 8474 18920
rect 8516 18880 8556 18920
rect 8598 18880 8638 18920
rect 8680 18880 8720 18920
rect 12352 18880 12392 18920
rect 12434 18880 12474 18920
rect 12516 18880 12556 18920
rect 12598 18880 12638 18920
rect 12680 18880 12720 18920
rect 16352 18880 16392 18920
rect 16434 18880 16474 18920
rect 16516 18880 16556 18920
rect 16598 18880 16638 18920
rect 16680 18880 16720 18920
rect 20352 18880 20392 18920
rect 20434 18880 20474 18920
rect 20516 18880 20556 18920
rect 20598 18880 20638 18920
rect 20680 18880 20720 18920
rect 24352 18880 24392 18920
rect 24434 18880 24474 18920
rect 24516 18880 24556 18920
rect 24598 18880 24638 18920
rect 24680 18880 24720 18920
rect 28352 18880 28392 18920
rect 28434 18880 28474 18920
rect 28516 18880 28556 18920
rect 28598 18880 28638 18920
rect 28680 18880 28720 18920
rect 32352 18880 32392 18920
rect 32434 18880 32474 18920
rect 32516 18880 32556 18920
rect 32598 18880 32638 18920
rect 32680 18880 32720 18920
rect 36352 18880 36392 18920
rect 36434 18880 36474 18920
rect 36516 18880 36556 18920
rect 36598 18880 36638 18920
rect 36680 18880 36720 18920
rect 40352 18880 40392 18920
rect 40434 18880 40474 18920
rect 40516 18880 40556 18920
rect 40598 18880 40638 18920
rect 40680 18880 40720 18920
rect 44352 18880 44392 18920
rect 44434 18880 44474 18920
rect 44516 18880 44556 18920
rect 44598 18880 44638 18920
rect 44680 18880 44720 18920
rect 48352 18880 48392 18920
rect 48434 18880 48474 18920
rect 48516 18880 48556 18920
rect 48598 18880 48638 18920
rect 48680 18880 48720 18920
rect 52352 18880 52392 18920
rect 52434 18880 52474 18920
rect 52516 18880 52556 18920
rect 52598 18880 52638 18920
rect 52680 18880 52720 18920
rect 56352 18880 56392 18920
rect 56434 18880 56474 18920
rect 56516 18880 56556 18920
rect 56598 18880 56638 18920
rect 56680 18880 56720 18920
rect 60352 18880 60392 18920
rect 60434 18880 60474 18920
rect 60516 18880 60556 18920
rect 60598 18880 60638 18920
rect 60680 18880 60720 18920
rect 64352 18880 64392 18920
rect 64434 18880 64474 18920
rect 64516 18880 64556 18920
rect 64598 18880 64638 18920
rect 64680 18880 64720 18920
rect 68352 18880 68392 18920
rect 68434 18880 68474 18920
rect 68516 18880 68556 18920
rect 68598 18880 68638 18920
rect 68680 18880 68720 18920
rect 72352 18880 72392 18920
rect 72434 18880 72474 18920
rect 72516 18880 72556 18920
rect 72598 18880 72638 18920
rect 72680 18880 72720 18920
rect 76352 18880 76392 18920
rect 76434 18880 76474 18920
rect 76516 18880 76556 18920
rect 76598 18880 76638 18920
rect 76680 18880 76720 18920
rect 80352 18880 80392 18920
rect 80434 18880 80474 18920
rect 80516 18880 80556 18920
rect 80598 18880 80638 18920
rect 80680 18880 80720 18920
rect 84352 18880 84392 18920
rect 84434 18880 84474 18920
rect 84516 18880 84556 18920
rect 84598 18880 84638 18920
rect 84680 18880 84720 18920
rect 88352 18880 88392 18920
rect 88434 18880 88474 18920
rect 88516 18880 88556 18920
rect 88598 18880 88638 18920
rect 88680 18880 88720 18920
rect 92352 18880 92392 18920
rect 92434 18880 92474 18920
rect 92516 18880 92556 18920
rect 92598 18880 92638 18920
rect 92680 18880 92720 18920
rect 96352 18880 96392 18920
rect 96434 18880 96474 18920
rect 96516 18880 96556 18920
rect 96598 18880 96638 18920
rect 96680 18880 96720 18920
rect 3112 18124 3152 18164
rect 3194 18124 3234 18164
rect 3276 18124 3316 18164
rect 3358 18124 3398 18164
rect 3440 18124 3480 18164
rect 7112 18124 7152 18164
rect 7194 18124 7234 18164
rect 7276 18124 7316 18164
rect 7358 18124 7398 18164
rect 7440 18124 7480 18164
rect 11112 18124 11152 18164
rect 11194 18124 11234 18164
rect 11276 18124 11316 18164
rect 11358 18124 11398 18164
rect 11440 18124 11480 18164
rect 15112 18124 15152 18164
rect 15194 18124 15234 18164
rect 15276 18124 15316 18164
rect 15358 18124 15398 18164
rect 15440 18124 15480 18164
rect 19112 18124 19152 18164
rect 19194 18124 19234 18164
rect 19276 18124 19316 18164
rect 19358 18124 19398 18164
rect 19440 18124 19480 18164
rect 23112 18124 23152 18164
rect 23194 18124 23234 18164
rect 23276 18124 23316 18164
rect 23358 18124 23398 18164
rect 23440 18124 23480 18164
rect 27112 18124 27152 18164
rect 27194 18124 27234 18164
rect 27276 18124 27316 18164
rect 27358 18124 27398 18164
rect 27440 18124 27480 18164
rect 31112 18124 31152 18164
rect 31194 18124 31234 18164
rect 31276 18124 31316 18164
rect 31358 18124 31398 18164
rect 31440 18124 31480 18164
rect 35112 18124 35152 18164
rect 35194 18124 35234 18164
rect 35276 18124 35316 18164
rect 35358 18124 35398 18164
rect 35440 18124 35480 18164
rect 39112 18124 39152 18164
rect 39194 18124 39234 18164
rect 39276 18124 39316 18164
rect 39358 18124 39398 18164
rect 39440 18124 39480 18164
rect 43112 18124 43152 18164
rect 43194 18124 43234 18164
rect 43276 18124 43316 18164
rect 43358 18124 43398 18164
rect 43440 18124 43480 18164
rect 47112 18124 47152 18164
rect 47194 18124 47234 18164
rect 47276 18124 47316 18164
rect 47358 18124 47398 18164
rect 47440 18124 47480 18164
rect 51112 18124 51152 18164
rect 51194 18124 51234 18164
rect 51276 18124 51316 18164
rect 51358 18124 51398 18164
rect 51440 18124 51480 18164
rect 55112 18124 55152 18164
rect 55194 18124 55234 18164
rect 55276 18124 55316 18164
rect 55358 18124 55398 18164
rect 55440 18124 55480 18164
rect 59112 18124 59152 18164
rect 59194 18124 59234 18164
rect 59276 18124 59316 18164
rect 59358 18124 59398 18164
rect 59440 18124 59480 18164
rect 63112 18124 63152 18164
rect 63194 18124 63234 18164
rect 63276 18124 63316 18164
rect 63358 18124 63398 18164
rect 63440 18124 63480 18164
rect 67112 18124 67152 18164
rect 67194 18124 67234 18164
rect 67276 18124 67316 18164
rect 67358 18124 67398 18164
rect 67440 18124 67480 18164
rect 71112 18124 71152 18164
rect 71194 18124 71234 18164
rect 71276 18124 71316 18164
rect 71358 18124 71398 18164
rect 71440 18124 71480 18164
rect 75112 18124 75152 18164
rect 75194 18124 75234 18164
rect 75276 18124 75316 18164
rect 75358 18124 75398 18164
rect 75440 18124 75480 18164
rect 79112 18124 79152 18164
rect 79194 18124 79234 18164
rect 79276 18124 79316 18164
rect 79358 18124 79398 18164
rect 79440 18124 79480 18164
rect 83112 18124 83152 18164
rect 83194 18124 83234 18164
rect 83276 18124 83316 18164
rect 83358 18124 83398 18164
rect 83440 18124 83480 18164
rect 87112 18124 87152 18164
rect 87194 18124 87234 18164
rect 87276 18124 87316 18164
rect 87358 18124 87398 18164
rect 87440 18124 87480 18164
rect 91112 18124 91152 18164
rect 91194 18124 91234 18164
rect 91276 18124 91316 18164
rect 91358 18124 91398 18164
rect 91440 18124 91480 18164
rect 95112 18124 95152 18164
rect 95194 18124 95234 18164
rect 95276 18124 95316 18164
rect 95358 18124 95398 18164
rect 95440 18124 95480 18164
rect 99112 18124 99152 18164
rect 99194 18124 99234 18164
rect 99276 18124 99316 18164
rect 99358 18124 99398 18164
rect 99440 18124 99480 18164
rect 4352 17368 4392 17408
rect 4434 17368 4474 17408
rect 4516 17368 4556 17408
rect 4598 17368 4638 17408
rect 4680 17368 4720 17408
rect 8352 17368 8392 17408
rect 8434 17368 8474 17408
rect 8516 17368 8556 17408
rect 8598 17368 8638 17408
rect 8680 17368 8720 17408
rect 12352 17368 12392 17408
rect 12434 17368 12474 17408
rect 12516 17368 12556 17408
rect 12598 17368 12638 17408
rect 12680 17368 12720 17408
rect 16352 17368 16392 17408
rect 16434 17368 16474 17408
rect 16516 17368 16556 17408
rect 16598 17368 16638 17408
rect 16680 17368 16720 17408
rect 20352 17368 20392 17408
rect 20434 17368 20474 17408
rect 20516 17368 20556 17408
rect 20598 17368 20638 17408
rect 20680 17368 20720 17408
rect 24352 17368 24392 17408
rect 24434 17368 24474 17408
rect 24516 17368 24556 17408
rect 24598 17368 24638 17408
rect 24680 17368 24720 17408
rect 28352 17368 28392 17408
rect 28434 17368 28474 17408
rect 28516 17368 28556 17408
rect 28598 17368 28638 17408
rect 28680 17368 28720 17408
rect 32352 17368 32392 17408
rect 32434 17368 32474 17408
rect 32516 17368 32556 17408
rect 32598 17368 32638 17408
rect 32680 17368 32720 17408
rect 36352 17368 36392 17408
rect 36434 17368 36474 17408
rect 36516 17368 36556 17408
rect 36598 17368 36638 17408
rect 36680 17368 36720 17408
rect 40352 17368 40392 17408
rect 40434 17368 40474 17408
rect 40516 17368 40556 17408
rect 40598 17368 40638 17408
rect 40680 17368 40720 17408
rect 44352 17368 44392 17408
rect 44434 17368 44474 17408
rect 44516 17368 44556 17408
rect 44598 17368 44638 17408
rect 44680 17368 44720 17408
rect 48352 17368 48392 17408
rect 48434 17368 48474 17408
rect 48516 17368 48556 17408
rect 48598 17368 48638 17408
rect 48680 17368 48720 17408
rect 52352 17368 52392 17408
rect 52434 17368 52474 17408
rect 52516 17368 52556 17408
rect 52598 17368 52638 17408
rect 52680 17368 52720 17408
rect 56352 17368 56392 17408
rect 56434 17368 56474 17408
rect 56516 17368 56556 17408
rect 56598 17368 56638 17408
rect 56680 17368 56720 17408
rect 60352 17368 60392 17408
rect 60434 17368 60474 17408
rect 60516 17368 60556 17408
rect 60598 17368 60638 17408
rect 60680 17368 60720 17408
rect 64352 17368 64392 17408
rect 64434 17368 64474 17408
rect 64516 17368 64556 17408
rect 64598 17368 64638 17408
rect 64680 17368 64720 17408
rect 68352 17368 68392 17408
rect 68434 17368 68474 17408
rect 68516 17368 68556 17408
rect 68598 17368 68638 17408
rect 68680 17368 68720 17408
rect 72352 17368 72392 17408
rect 72434 17368 72474 17408
rect 72516 17368 72556 17408
rect 72598 17368 72638 17408
rect 72680 17368 72720 17408
rect 76352 17368 76392 17408
rect 76434 17368 76474 17408
rect 76516 17368 76556 17408
rect 76598 17368 76638 17408
rect 76680 17368 76720 17408
rect 80352 17368 80392 17408
rect 80434 17368 80474 17408
rect 80516 17368 80556 17408
rect 80598 17368 80638 17408
rect 80680 17368 80720 17408
rect 84352 17368 84392 17408
rect 84434 17368 84474 17408
rect 84516 17368 84556 17408
rect 84598 17368 84638 17408
rect 84680 17368 84720 17408
rect 88352 17368 88392 17408
rect 88434 17368 88474 17408
rect 88516 17368 88556 17408
rect 88598 17368 88638 17408
rect 88680 17368 88720 17408
rect 92352 17368 92392 17408
rect 92434 17368 92474 17408
rect 92516 17368 92556 17408
rect 92598 17368 92638 17408
rect 92680 17368 92720 17408
rect 96352 17368 96392 17408
rect 96434 17368 96474 17408
rect 96516 17368 96556 17408
rect 96598 17368 96638 17408
rect 96680 17368 96720 17408
rect 3112 16612 3152 16652
rect 3194 16612 3234 16652
rect 3276 16612 3316 16652
rect 3358 16612 3398 16652
rect 3440 16612 3480 16652
rect 7112 16612 7152 16652
rect 7194 16612 7234 16652
rect 7276 16612 7316 16652
rect 7358 16612 7398 16652
rect 7440 16612 7480 16652
rect 11112 16612 11152 16652
rect 11194 16612 11234 16652
rect 11276 16612 11316 16652
rect 11358 16612 11398 16652
rect 11440 16612 11480 16652
rect 15112 16612 15152 16652
rect 15194 16612 15234 16652
rect 15276 16612 15316 16652
rect 15358 16612 15398 16652
rect 15440 16612 15480 16652
rect 19112 16612 19152 16652
rect 19194 16612 19234 16652
rect 19276 16612 19316 16652
rect 19358 16612 19398 16652
rect 19440 16612 19480 16652
rect 23112 16612 23152 16652
rect 23194 16612 23234 16652
rect 23276 16612 23316 16652
rect 23358 16612 23398 16652
rect 23440 16612 23480 16652
rect 27112 16612 27152 16652
rect 27194 16612 27234 16652
rect 27276 16612 27316 16652
rect 27358 16612 27398 16652
rect 27440 16612 27480 16652
rect 31112 16612 31152 16652
rect 31194 16612 31234 16652
rect 31276 16612 31316 16652
rect 31358 16612 31398 16652
rect 31440 16612 31480 16652
rect 35112 16612 35152 16652
rect 35194 16612 35234 16652
rect 35276 16612 35316 16652
rect 35358 16612 35398 16652
rect 35440 16612 35480 16652
rect 39112 16612 39152 16652
rect 39194 16612 39234 16652
rect 39276 16612 39316 16652
rect 39358 16612 39398 16652
rect 39440 16612 39480 16652
rect 43112 16612 43152 16652
rect 43194 16612 43234 16652
rect 43276 16612 43316 16652
rect 43358 16612 43398 16652
rect 43440 16612 43480 16652
rect 47112 16612 47152 16652
rect 47194 16612 47234 16652
rect 47276 16612 47316 16652
rect 47358 16612 47398 16652
rect 47440 16612 47480 16652
rect 51112 16612 51152 16652
rect 51194 16612 51234 16652
rect 51276 16612 51316 16652
rect 51358 16612 51398 16652
rect 51440 16612 51480 16652
rect 55112 16612 55152 16652
rect 55194 16612 55234 16652
rect 55276 16612 55316 16652
rect 55358 16612 55398 16652
rect 55440 16612 55480 16652
rect 59112 16612 59152 16652
rect 59194 16612 59234 16652
rect 59276 16612 59316 16652
rect 59358 16612 59398 16652
rect 59440 16612 59480 16652
rect 63112 16612 63152 16652
rect 63194 16612 63234 16652
rect 63276 16612 63316 16652
rect 63358 16612 63398 16652
rect 63440 16612 63480 16652
rect 67112 16612 67152 16652
rect 67194 16612 67234 16652
rect 67276 16612 67316 16652
rect 67358 16612 67398 16652
rect 67440 16612 67480 16652
rect 71112 16612 71152 16652
rect 71194 16612 71234 16652
rect 71276 16612 71316 16652
rect 71358 16612 71398 16652
rect 71440 16612 71480 16652
rect 75112 16612 75152 16652
rect 75194 16612 75234 16652
rect 75276 16612 75316 16652
rect 75358 16612 75398 16652
rect 75440 16612 75480 16652
rect 79112 16612 79152 16652
rect 79194 16612 79234 16652
rect 79276 16612 79316 16652
rect 79358 16612 79398 16652
rect 79440 16612 79480 16652
rect 83112 16612 83152 16652
rect 83194 16612 83234 16652
rect 83276 16612 83316 16652
rect 83358 16612 83398 16652
rect 83440 16612 83480 16652
rect 87112 16612 87152 16652
rect 87194 16612 87234 16652
rect 87276 16612 87316 16652
rect 87358 16612 87398 16652
rect 87440 16612 87480 16652
rect 91112 16612 91152 16652
rect 91194 16612 91234 16652
rect 91276 16612 91316 16652
rect 91358 16612 91398 16652
rect 91440 16612 91480 16652
rect 95112 16612 95152 16652
rect 95194 16612 95234 16652
rect 95276 16612 95316 16652
rect 95358 16612 95398 16652
rect 95440 16612 95480 16652
rect 99112 16612 99152 16652
rect 99194 16612 99234 16652
rect 99276 16612 99316 16652
rect 99358 16612 99398 16652
rect 99440 16612 99480 16652
rect 86188 16360 86228 16400
rect 4352 15856 4392 15896
rect 4434 15856 4474 15896
rect 4516 15856 4556 15896
rect 4598 15856 4638 15896
rect 4680 15856 4720 15896
rect 8352 15856 8392 15896
rect 8434 15856 8474 15896
rect 8516 15856 8556 15896
rect 8598 15856 8638 15896
rect 8680 15856 8720 15896
rect 12352 15856 12392 15896
rect 12434 15856 12474 15896
rect 12516 15856 12556 15896
rect 12598 15856 12638 15896
rect 12680 15856 12720 15896
rect 16352 15856 16392 15896
rect 16434 15856 16474 15896
rect 16516 15856 16556 15896
rect 16598 15856 16638 15896
rect 16680 15856 16720 15896
rect 20352 15856 20392 15896
rect 20434 15856 20474 15896
rect 20516 15856 20556 15896
rect 20598 15856 20638 15896
rect 20680 15856 20720 15896
rect 24352 15856 24392 15896
rect 24434 15856 24474 15896
rect 24516 15856 24556 15896
rect 24598 15856 24638 15896
rect 24680 15856 24720 15896
rect 28352 15856 28392 15896
rect 28434 15856 28474 15896
rect 28516 15856 28556 15896
rect 28598 15856 28638 15896
rect 28680 15856 28720 15896
rect 32352 15856 32392 15896
rect 32434 15856 32474 15896
rect 32516 15856 32556 15896
rect 32598 15856 32638 15896
rect 32680 15856 32720 15896
rect 36352 15856 36392 15896
rect 36434 15856 36474 15896
rect 36516 15856 36556 15896
rect 36598 15856 36638 15896
rect 36680 15856 36720 15896
rect 40352 15856 40392 15896
rect 40434 15856 40474 15896
rect 40516 15856 40556 15896
rect 40598 15856 40638 15896
rect 40680 15856 40720 15896
rect 44352 15856 44392 15896
rect 44434 15856 44474 15896
rect 44516 15856 44556 15896
rect 44598 15856 44638 15896
rect 44680 15856 44720 15896
rect 48352 15856 48392 15896
rect 48434 15856 48474 15896
rect 48516 15856 48556 15896
rect 48598 15856 48638 15896
rect 48680 15856 48720 15896
rect 52352 15856 52392 15896
rect 52434 15856 52474 15896
rect 52516 15856 52556 15896
rect 52598 15856 52638 15896
rect 52680 15856 52720 15896
rect 56352 15856 56392 15896
rect 56434 15856 56474 15896
rect 56516 15856 56556 15896
rect 56598 15856 56638 15896
rect 56680 15856 56720 15896
rect 60352 15856 60392 15896
rect 60434 15856 60474 15896
rect 60516 15856 60556 15896
rect 60598 15856 60638 15896
rect 60680 15856 60720 15896
rect 64352 15856 64392 15896
rect 64434 15856 64474 15896
rect 64516 15856 64556 15896
rect 64598 15856 64638 15896
rect 64680 15856 64720 15896
rect 68352 15856 68392 15896
rect 68434 15856 68474 15896
rect 68516 15856 68556 15896
rect 68598 15856 68638 15896
rect 68680 15856 68720 15896
rect 72352 15856 72392 15896
rect 72434 15856 72474 15896
rect 72516 15856 72556 15896
rect 72598 15856 72638 15896
rect 72680 15856 72720 15896
rect 76352 15856 76392 15896
rect 76434 15856 76474 15896
rect 76516 15856 76556 15896
rect 76598 15856 76638 15896
rect 76680 15856 76720 15896
rect 80352 15856 80392 15896
rect 80434 15856 80474 15896
rect 80516 15856 80556 15896
rect 80598 15856 80638 15896
rect 80680 15856 80720 15896
rect 84352 15856 84392 15896
rect 84434 15856 84474 15896
rect 84516 15856 84556 15896
rect 84598 15856 84638 15896
rect 84680 15856 84720 15896
rect 88352 15856 88392 15896
rect 88434 15856 88474 15896
rect 88516 15856 88556 15896
rect 88598 15856 88638 15896
rect 88680 15856 88720 15896
rect 92352 15856 92392 15896
rect 92434 15856 92474 15896
rect 92516 15856 92556 15896
rect 92598 15856 92638 15896
rect 92680 15856 92720 15896
rect 96352 15856 96392 15896
rect 96434 15856 96474 15896
rect 96516 15856 96556 15896
rect 96598 15856 96638 15896
rect 96680 15856 96720 15896
rect 3112 15100 3152 15140
rect 3194 15100 3234 15140
rect 3276 15100 3316 15140
rect 3358 15100 3398 15140
rect 3440 15100 3480 15140
rect 7112 15100 7152 15140
rect 7194 15100 7234 15140
rect 7276 15100 7316 15140
rect 7358 15100 7398 15140
rect 7440 15100 7480 15140
rect 11112 15100 11152 15140
rect 11194 15100 11234 15140
rect 11276 15100 11316 15140
rect 11358 15100 11398 15140
rect 11440 15100 11480 15140
rect 15112 15100 15152 15140
rect 15194 15100 15234 15140
rect 15276 15100 15316 15140
rect 15358 15100 15398 15140
rect 15440 15100 15480 15140
rect 19112 15100 19152 15140
rect 19194 15100 19234 15140
rect 19276 15100 19316 15140
rect 19358 15100 19398 15140
rect 19440 15100 19480 15140
rect 23112 15100 23152 15140
rect 23194 15100 23234 15140
rect 23276 15100 23316 15140
rect 23358 15100 23398 15140
rect 23440 15100 23480 15140
rect 27112 15100 27152 15140
rect 27194 15100 27234 15140
rect 27276 15100 27316 15140
rect 27358 15100 27398 15140
rect 27440 15100 27480 15140
rect 31112 15100 31152 15140
rect 31194 15100 31234 15140
rect 31276 15100 31316 15140
rect 31358 15100 31398 15140
rect 31440 15100 31480 15140
rect 35112 15100 35152 15140
rect 35194 15100 35234 15140
rect 35276 15100 35316 15140
rect 35358 15100 35398 15140
rect 35440 15100 35480 15140
rect 39112 15100 39152 15140
rect 39194 15100 39234 15140
rect 39276 15100 39316 15140
rect 39358 15100 39398 15140
rect 39440 15100 39480 15140
rect 43112 15100 43152 15140
rect 43194 15100 43234 15140
rect 43276 15100 43316 15140
rect 43358 15100 43398 15140
rect 43440 15100 43480 15140
rect 47112 15100 47152 15140
rect 47194 15100 47234 15140
rect 47276 15100 47316 15140
rect 47358 15100 47398 15140
rect 47440 15100 47480 15140
rect 51112 15100 51152 15140
rect 51194 15100 51234 15140
rect 51276 15100 51316 15140
rect 51358 15100 51398 15140
rect 51440 15100 51480 15140
rect 55112 15100 55152 15140
rect 55194 15100 55234 15140
rect 55276 15100 55316 15140
rect 55358 15100 55398 15140
rect 55440 15100 55480 15140
rect 59112 15100 59152 15140
rect 59194 15100 59234 15140
rect 59276 15100 59316 15140
rect 59358 15100 59398 15140
rect 59440 15100 59480 15140
rect 63112 15100 63152 15140
rect 63194 15100 63234 15140
rect 63276 15100 63316 15140
rect 63358 15100 63398 15140
rect 63440 15100 63480 15140
rect 67112 15100 67152 15140
rect 67194 15100 67234 15140
rect 67276 15100 67316 15140
rect 67358 15100 67398 15140
rect 67440 15100 67480 15140
rect 4352 14344 4392 14384
rect 4434 14344 4474 14384
rect 4516 14344 4556 14384
rect 4598 14344 4638 14384
rect 4680 14344 4720 14384
rect 8352 14344 8392 14384
rect 8434 14344 8474 14384
rect 8516 14344 8556 14384
rect 8598 14344 8638 14384
rect 8680 14344 8720 14384
rect 12352 14344 12392 14384
rect 12434 14344 12474 14384
rect 12516 14344 12556 14384
rect 12598 14344 12638 14384
rect 12680 14344 12720 14384
rect 16352 14344 16392 14384
rect 16434 14344 16474 14384
rect 16516 14344 16556 14384
rect 16598 14344 16638 14384
rect 16680 14344 16720 14384
rect 20352 14344 20392 14384
rect 20434 14344 20474 14384
rect 20516 14344 20556 14384
rect 20598 14344 20638 14384
rect 20680 14344 20720 14384
rect 24352 14344 24392 14384
rect 24434 14344 24474 14384
rect 24516 14344 24556 14384
rect 24598 14344 24638 14384
rect 24680 14344 24720 14384
rect 28352 14344 28392 14384
rect 28434 14344 28474 14384
rect 28516 14344 28556 14384
rect 28598 14344 28638 14384
rect 28680 14344 28720 14384
rect 32352 14344 32392 14384
rect 32434 14344 32474 14384
rect 32516 14344 32556 14384
rect 32598 14344 32638 14384
rect 32680 14344 32720 14384
rect 36352 14344 36392 14384
rect 36434 14344 36474 14384
rect 36516 14344 36556 14384
rect 36598 14344 36638 14384
rect 36680 14344 36720 14384
rect 40352 14344 40392 14384
rect 40434 14344 40474 14384
rect 40516 14344 40556 14384
rect 40598 14344 40638 14384
rect 40680 14344 40720 14384
rect 44352 14344 44392 14384
rect 44434 14344 44474 14384
rect 44516 14344 44556 14384
rect 44598 14344 44638 14384
rect 44680 14344 44720 14384
rect 48352 14344 48392 14384
rect 48434 14344 48474 14384
rect 48516 14344 48556 14384
rect 48598 14344 48638 14384
rect 48680 14344 48720 14384
rect 52352 14344 52392 14384
rect 52434 14344 52474 14384
rect 52516 14344 52556 14384
rect 52598 14344 52638 14384
rect 52680 14344 52720 14384
rect 56352 14344 56392 14384
rect 56434 14344 56474 14384
rect 56516 14344 56556 14384
rect 56598 14344 56638 14384
rect 56680 14344 56720 14384
rect 60352 14344 60392 14384
rect 60434 14344 60474 14384
rect 60516 14344 60556 14384
rect 60598 14344 60638 14384
rect 60680 14344 60720 14384
rect 64352 14344 64392 14384
rect 64434 14344 64474 14384
rect 64516 14344 64556 14384
rect 64598 14344 64638 14384
rect 64680 14344 64720 14384
rect 68352 14344 68392 14384
rect 68434 14344 68474 14384
rect 68516 14344 68556 14384
rect 68598 14344 68638 14384
rect 68680 14344 68720 14384
rect 3112 13588 3152 13628
rect 3194 13588 3234 13628
rect 3276 13588 3316 13628
rect 3358 13588 3398 13628
rect 3440 13588 3480 13628
rect 7112 13588 7152 13628
rect 7194 13588 7234 13628
rect 7276 13588 7316 13628
rect 7358 13588 7398 13628
rect 7440 13588 7480 13628
rect 11112 13588 11152 13628
rect 11194 13588 11234 13628
rect 11276 13588 11316 13628
rect 11358 13588 11398 13628
rect 11440 13588 11480 13628
rect 15112 13588 15152 13628
rect 15194 13588 15234 13628
rect 15276 13588 15316 13628
rect 15358 13588 15398 13628
rect 15440 13588 15480 13628
rect 19112 13588 19152 13628
rect 19194 13588 19234 13628
rect 19276 13588 19316 13628
rect 19358 13588 19398 13628
rect 19440 13588 19480 13628
rect 23112 13588 23152 13628
rect 23194 13588 23234 13628
rect 23276 13588 23316 13628
rect 23358 13588 23398 13628
rect 23440 13588 23480 13628
rect 27112 13588 27152 13628
rect 27194 13588 27234 13628
rect 27276 13588 27316 13628
rect 27358 13588 27398 13628
rect 27440 13588 27480 13628
rect 31112 13588 31152 13628
rect 31194 13588 31234 13628
rect 31276 13588 31316 13628
rect 31358 13588 31398 13628
rect 31440 13588 31480 13628
rect 35112 13588 35152 13628
rect 35194 13588 35234 13628
rect 35276 13588 35316 13628
rect 35358 13588 35398 13628
rect 35440 13588 35480 13628
rect 39112 13588 39152 13628
rect 39194 13588 39234 13628
rect 39276 13588 39316 13628
rect 39358 13588 39398 13628
rect 39440 13588 39480 13628
rect 43112 13588 43152 13628
rect 43194 13588 43234 13628
rect 43276 13588 43316 13628
rect 43358 13588 43398 13628
rect 43440 13588 43480 13628
rect 47112 13588 47152 13628
rect 47194 13588 47234 13628
rect 47276 13588 47316 13628
rect 47358 13588 47398 13628
rect 47440 13588 47480 13628
rect 51112 13588 51152 13628
rect 51194 13588 51234 13628
rect 51276 13588 51316 13628
rect 51358 13588 51398 13628
rect 51440 13588 51480 13628
rect 55112 13588 55152 13628
rect 55194 13588 55234 13628
rect 55276 13588 55316 13628
rect 55358 13588 55398 13628
rect 55440 13588 55480 13628
rect 59112 13588 59152 13628
rect 59194 13588 59234 13628
rect 59276 13588 59316 13628
rect 59358 13588 59398 13628
rect 59440 13588 59480 13628
rect 63112 13588 63152 13628
rect 63194 13588 63234 13628
rect 63276 13588 63316 13628
rect 63358 13588 63398 13628
rect 63440 13588 63480 13628
rect 67112 13588 67152 13628
rect 67194 13588 67234 13628
rect 67276 13588 67316 13628
rect 67358 13588 67398 13628
rect 67440 13588 67480 13628
rect 4352 12832 4392 12872
rect 4434 12832 4474 12872
rect 4516 12832 4556 12872
rect 4598 12832 4638 12872
rect 4680 12832 4720 12872
rect 8352 12832 8392 12872
rect 8434 12832 8474 12872
rect 8516 12832 8556 12872
rect 8598 12832 8638 12872
rect 8680 12832 8720 12872
rect 12352 12832 12392 12872
rect 12434 12832 12474 12872
rect 12516 12832 12556 12872
rect 12598 12832 12638 12872
rect 12680 12832 12720 12872
rect 16352 12832 16392 12872
rect 16434 12832 16474 12872
rect 16516 12832 16556 12872
rect 16598 12832 16638 12872
rect 16680 12832 16720 12872
rect 20352 12832 20392 12872
rect 20434 12832 20474 12872
rect 20516 12832 20556 12872
rect 20598 12832 20638 12872
rect 20680 12832 20720 12872
rect 24352 12832 24392 12872
rect 24434 12832 24474 12872
rect 24516 12832 24556 12872
rect 24598 12832 24638 12872
rect 24680 12832 24720 12872
rect 28352 12832 28392 12872
rect 28434 12832 28474 12872
rect 28516 12832 28556 12872
rect 28598 12832 28638 12872
rect 28680 12832 28720 12872
rect 32352 12832 32392 12872
rect 32434 12832 32474 12872
rect 32516 12832 32556 12872
rect 32598 12832 32638 12872
rect 32680 12832 32720 12872
rect 36352 12832 36392 12872
rect 36434 12832 36474 12872
rect 36516 12832 36556 12872
rect 36598 12832 36638 12872
rect 36680 12832 36720 12872
rect 40352 12832 40392 12872
rect 40434 12832 40474 12872
rect 40516 12832 40556 12872
rect 40598 12832 40638 12872
rect 40680 12832 40720 12872
rect 44352 12832 44392 12872
rect 44434 12832 44474 12872
rect 44516 12832 44556 12872
rect 44598 12832 44638 12872
rect 44680 12832 44720 12872
rect 48352 12832 48392 12872
rect 48434 12832 48474 12872
rect 48516 12832 48556 12872
rect 48598 12832 48638 12872
rect 48680 12832 48720 12872
rect 52352 12832 52392 12872
rect 52434 12832 52474 12872
rect 52516 12832 52556 12872
rect 52598 12832 52638 12872
rect 52680 12832 52720 12872
rect 56352 12832 56392 12872
rect 56434 12832 56474 12872
rect 56516 12832 56556 12872
rect 56598 12832 56638 12872
rect 56680 12832 56720 12872
rect 60352 12832 60392 12872
rect 60434 12832 60474 12872
rect 60516 12832 60556 12872
rect 60598 12832 60638 12872
rect 60680 12832 60720 12872
rect 64352 12832 64392 12872
rect 64434 12832 64474 12872
rect 64516 12832 64556 12872
rect 64598 12832 64638 12872
rect 64680 12832 64720 12872
rect 68352 12832 68392 12872
rect 68434 12832 68474 12872
rect 68516 12832 68556 12872
rect 68598 12832 68638 12872
rect 68680 12832 68720 12872
rect 3112 12076 3152 12116
rect 3194 12076 3234 12116
rect 3276 12076 3316 12116
rect 3358 12076 3398 12116
rect 3440 12076 3480 12116
rect 7112 12076 7152 12116
rect 7194 12076 7234 12116
rect 7276 12076 7316 12116
rect 7358 12076 7398 12116
rect 7440 12076 7480 12116
rect 11112 12076 11152 12116
rect 11194 12076 11234 12116
rect 11276 12076 11316 12116
rect 11358 12076 11398 12116
rect 11440 12076 11480 12116
rect 15112 12076 15152 12116
rect 15194 12076 15234 12116
rect 15276 12076 15316 12116
rect 15358 12076 15398 12116
rect 15440 12076 15480 12116
rect 19112 12076 19152 12116
rect 19194 12076 19234 12116
rect 19276 12076 19316 12116
rect 19358 12076 19398 12116
rect 19440 12076 19480 12116
rect 23112 12076 23152 12116
rect 23194 12076 23234 12116
rect 23276 12076 23316 12116
rect 23358 12076 23398 12116
rect 23440 12076 23480 12116
rect 27112 12076 27152 12116
rect 27194 12076 27234 12116
rect 27276 12076 27316 12116
rect 27358 12076 27398 12116
rect 27440 12076 27480 12116
rect 31112 12076 31152 12116
rect 31194 12076 31234 12116
rect 31276 12076 31316 12116
rect 31358 12076 31398 12116
rect 31440 12076 31480 12116
rect 35112 12076 35152 12116
rect 35194 12076 35234 12116
rect 35276 12076 35316 12116
rect 35358 12076 35398 12116
rect 35440 12076 35480 12116
rect 39112 12076 39152 12116
rect 39194 12076 39234 12116
rect 39276 12076 39316 12116
rect 39358 12076 39398 12116
rect 39440 12076 39480 12116
rect 43112 12076 43152 12116
rect 43194 12076 43234 12116
rect 43276 12076 43316 12116
rect 43358 12076 43398 12116
rect 43440 12076 43480 12116
rect 47112 12076 47152 12116
rect 47194 12076 47234 12116
rect 47276 12076 47316 12116
rect 47358 12076 47398 12116
rect 47440 12076 47480 12116
rect 51112 12076 51152 12116
rect 51194 12076 51234 12116
rect 51276 12076 51316 12116
rect 51358 12076 51398 12116
rect 51440 12076 51480 12116
rect 55112 12076 55152 12116
rect 55194 12076 55234 12116
rect 55276 12076 55316 12116
rect 55358 12076 55398 12116
rect 55440 12076 55480 12116
rect 59112 12076 59152 12116
rect 59194 12076 59234 12116
rect 59276 12076 59316 12116
rect 59358 12076 59398 12116
rect 59440 12076 59480 12116
rect 63112 12076 63152 12116
rect 63194 12076 63234 12116
rect 63276 12076 63316 12116
rect 63358 12076 63398 12116
rect 63440 12076 63480 12116
rect 67112 12076 67152 12116
rect 67194 12076 67234 12116
rect 67276 12076 67316 12116
rect 67358 12076 67398 12116
rect 67440 12076 67480 12116
rect 4352 11320 4392 11360
rect 4434 11320 4474 11360
rect 4516 11320 4556 11360
rect 4598 11320 4638 11360
rect 4680 11320 4720 11360
rect 8352 11320 8392 11360
rect 8434 11320 8474 11360
rect 8516 11320 8556 11360
rect 8598 11320 8638 11360
rect 8680 11320 8720 11360
rect 12352 11320 12392 11360
rect 12434 11320 12474 11360
rect 12516 11320 12556 11360
rect 12598 11320 12638 11360
rect 12680 11320 12720 11360
rect 16352 11320 16392 11360
rect 16434 11320 16474 11360
rect 16516 11320 16556 11360
rect 16598 11320 16638 11360
rect 16680 11320 16720 11360
rect 20352 11320 20392 11360
rect 20434 11320 20474 11360
rect 20516 11320 20556 11360
rect 20598 11320 20638 11360
rect 20680 11320 20720 11360
rect 24352 11320 24392 11360
rect 24434 11320 24474 11360
rect 24516 11320 24556 11360
rect 24598 11320 24638 11360
rect 24680 11320 24720 11360
rect 28352 11320 28392 11360
rect 28434 11320 28474 11360
rect 28516 11320 28556 11360
rect 28598 11320 28638 11360
rect 28680 11320 28720 11360
rect 32352 11320 32392 11360
rect 32434 11320 32474 11360
rect 32516 11320 32556 11360
rect 32598 11320 32638 11360
rect 32680 11320 32720 11360
rect 36352 11320 36392 11360
rect 36434 11320 36474 11360
rect 36516 11320 36556 11360
rect 36598 11320 36638 11360
rect 36680 11320 36720 11360
rect 40352 11320 40392 11360
rect 40434 11320 40474 11360
rect 40516 11320 40556 11360
rect 40598 11320 40638 11360
rect 40680 11320 40720 11360
rect 44352 11320 44392 11360
rect 44434 11320 44474 11360
rect 44516 11320 44556 11360
rect 44598 11320 44638 11360
rect 44680 11320 44720 11360
rect 48352 11320 48392 11360
rect 48434 11320 48474 11360
rect 48516 11320 48556 11360
rect 48598 11320 48638 11360
rect 48680 11320 48720 11360
rect 52352 11320 52392 11360
rect 52434 11320 52474 11360
rect 52516 11320 52556 11360
rect 52598 11320 52638 11360
rect 52680 11320 52720 11360
rect 56352 11320 56392 11360
rect 56434 11320 56474 11360
rect 56516 11320 56556 11360
rect 56598 11320 56638 11360
rect 56680 11320 56720 11360
rect 60352 11320 60392 11360
rect 60434 11320 60474 11360
rect 60516 11320 60556 11360
rect 60598 11320 60638 11360
rect 60680 11320 60720 11360
rect 64352 11320 64392 11360
rect 64434 11320 64474 11360
rect 64516 11320 64556 11360
rect 64598 11320 64638 11360
rect 64680 11320 64720 11360
rect 68352 11320 68392 11360
rect 68434 11320 68474 11360
rect 68516 11320 68556 11360
rect 68598 11320 68638 11360
rect 68680 11320 68720 11360
rect 3112 10564 3152 10604
rect 3194 10564 3234 10604
rect 3276 10564 3316 10604
rect 3358 10564 3398 10604
rect 3440 10564 3480 10604
rect 7112 10564 7152 10604
rect 7194 10564 7234 10604
rect 7276 10564 7316 10604
rect 7358 10564 7398 10604
rect 7440 10564 7480 10604
rect 11112 10564 11152 10604
rect 11194 10564 11234 10604
rect 11276 10564 11316 10604
rect 11358 10564 11398 10604
rect 11440 10564 11480 10604
rect 15112 10564 15152 10604
rect 15194 10564 15234 10604
rect 15276 10564 15316 10604
rect 15358 10564 15398 10604
rect 15440 10564 15480 10604
rect 19112 10564 19152 10604
rect 19194 10564 19234 10604
rect 19276 10564 19316 10604
rect 19358 10564 19398 10604
rect 19440 10564 19480 10604
rect 23112 10564 23152 10604
rect 23194 10564 23234 10604
rect 23276 10564 23316 10604
rect 23358 10564 23398 10604
rect 23440 10564 23480 10604
rect 27112 10564 27152 10604
rect 27194 10564 27234 10604
rect 27276 10564 27316 10604
rect 27358 10564 27398 10604
rect 27440 10564 27480 10604
rect 31112 10564 31152 10604
rect 31194 10564 31234 10604
rect 31276 10564 31316 10604
rect 31358 10564 31398 10604
rect 31440 10564 31480 10604
rect 35112 10564 35152 10604
rect 35194 10564 35234 10604
rect 35276 10564 35316 10604
rect 35358 10564 35398 10604
rect 35440 10564 35480 10604
rect 39112 10564 39152 10604
rect 39194 10564 39234 10604
rect 39276 10564 39316 10604
rect 39358 10564 39398 10604
rect 39440 10564 39480 10604
rect 43112 10564 43152 10604
rect 43194 10564 43234 10604
rect 43276 10564 43316 10604
rect 43358 10564 43398 10604
rect 43440 10564 43480 10604
rect 47112 10564 47152 10604
rect 47194 10564 47234 10604
rect 47276 10564 47316 10604
rect 47358 10564 47398 10604
rect 47440 10564 47480 10604
rect 51112 10564 51152 10604
rect 51194 10564 51234 10604
rect 51276 10564 51316 10604
rect 51358 10564 51398 10604
rect 51440 10564 51480 10604
rect 55112 10564 55152 10604
rect 55194 10564 55234 10604
rect 55276 10564 55316 10604
rect 55358 10564 55398 10604
rect 55440 10564 55480 10604
rect 59112 10564 59152 10604
rect 59194 10564 59234 10604
rect 59276 10564 59316 10604
rect 59358 10564 59398 10604
rect 59440 10564 59480 10604
rect 63112 10564 63152 10604
rect 63194 10564 63234 10604
rect 63276 10564 63316 10604
rect 63358 10564 63398 10604
rect 63440 10564 63480 10604
rect 67112 10564 67152 10604
rect 67194 10564 67234 10604
rect 67276 10564 67316 10604
rect 67358 10564 67398 10604
rect 67440 10564 67480 10604
rect 4352 9808 4392 9848
rect 4434 9808 4474 9848
rect 4516 9808 4556 9848
rect 4598 9808 4638 9848
rect 4680 9808 4720 9848
rect 8352 9808 8392 9848
rect 8434 9808 8474 9848
rect 8516 9808 8556 9848
rect 8598 9808 8638 9848
rect 8680 9808 8720 9848
rect 12352 9808 12392 9848
rect 12434 9808 12474 9848
rect 12516 9808 12556 9848
rect 12598 9808 12638 9848
rect 12680 9808 12720 9848
rect 16352 9808 16392 9848
rect 16434 9808 16474 9848
rect 16516 9808 16556 9848
rect 16598 9808 16638 9848
rect 16680 9808 16720 9848
rect 20352 9808 20392 9848
rect 20434 9808 20474 9848
rect 20516 9808 20556 9848
rect 20598 9808 20638 9848
rect 20680 9808 20720 9848
rect 24352 9808 24392 9848
rect 24434 9808 24474 9848
rect 24516 9808 24556 9848
rect 24598 9808 24638 9848
rect 24680 9808 24720 9848
rect 28352 9808 28392 9848
rect 28434 9808 28474 9848
rect 28516 9808 28556 9848
rect 28598 9808 28638 9848
rect 28680 9808 28720 9848
rect 32352 9808 32392 9848
rect 32434 9808 32474 9848
rect 32516 9808 32556 9848
rect 32598 9808 32638 9848
rect 32680 9808 32720 9848
rect 36352 9808 36392 9848
rect 36434 9808 36474 9848
rect 36516 9808 36556 9848
rect 36598 9808 36638 9848
rect 36680 9808 36720 9848
rect 40352 9808 40392 9848
rect 40434 9808 40474 9848
rect 40516 9808 40556 9848
rect 40598 9808 40638 9848
rect 40680 9808 40720 9848
rect 44352 9808 44392 9848
rect 44434 9808 44474 9848
rect 44516 9808 44556 9848
rect 44598 9808 44638 9848
rect 44680 9808 44720 9848
rect 48352 9808 48392 9848
rect 48434 9808 48474 9848
rect 48516 9808 48556 9848
rect 48598 9808 48638 9848
rect 48680 9808 48720 9848
rect 52352 9808 52392 9848
rect 52434 9808 52474 9848
rect 52516 9808 52556 9848
rect 52598 9808 52638 9848
rect 52680 9808 52720 9848
rect 56352 9808 56392 9848
rect 56434 9808 56474 9848
rect 56516 9808 56556 9848
rect 56598 9808 56638 9848
rect 56680 9808 56720 9848
rect 60352 9808 60392 9848
rect 60434 9808 60474 9848
rect 60516 9808 60556 9848
rect 60598 9808 60638 9848
rect 60680 9808 60720 9848
rect 64352 9808 64392 9848
rect 64434 9808 64474 9848
rect 64516 9808 64556 9848
rect 64598 9808 64638 9848
rect 64680 9808 64720 9848
rect 68352 9808 68392 9848
rect 68434 9808 68474 9848
rect 68516 9808 68556 9848
rect 68598 9808 68638 9848
rect 68680 9808 68720 9848
rect 3112 9052 3152 9092
rect 3194 9052 3234 9092
rect 3276 9052 3316 9092
rect 3358 9052 3398 9092
rect 3440 9052 3480 9092
rect 7112 9052 7152 9092
rect 7194 9052 7234 9092
rect 7276 9052 7316 9092
rect 7358 9052 7398 9092
rect 7440 9052 7480 9092
rect 11112 9052 11152 9092
rect 11194 9052 11234 9092
rect 11276 9052 11316 9092
rect 11358 9052 11398 9092
rect 11440 9052 11480 9092
rect 15112 9052 15152 9092
rect 15194 9052 15234 9092
rect 15276 9052 15316 9092
rect 15358 9052 15398 9092
rect 15440 9052 15480 9092
rect 19112 9052 19152 9092
rect 19194 9052 19234 9092
rect 19276 9052 19316 9092
rect 19358 9052 19398 9092
rect 19440 9052 19480 9092
rect 23112 9052 23152 9092
rect 23194 9052 23234 9092
rect 23276 9052 23316 9092
rect 23358 9052 23398 9092
rect 23440 9052 23480 9092
rect 27112 9052 27152 9092
rect 27194 9052 27234 9092
rect 27276 9052 27316 9092
rect 27358 9052 27398 9092
rect 27440 9052 27480 9092
rect 31112 9052 31152 9092
rect 31194 9052 31234 9092
rect 31276 9052 31316 9092
rect 31358 9052 31398 9092
rect 31440 9052 31480 9092
rect 35112 9052 35152 9092
rect 35194 9052 35234 9092
rect 35276 9052 35316 9092
rect 35358 9052 35398 9092
rect 35440 9052 35480 9092
rect 39112 9052 39152 9092
rect 39194 9052 39234 9092
rect 39276 9052 39316 9092
rect 39358 9052 39398 9092
rect 39440 9052 39480 9092
rect 43112 9052 43152 9092
rect 43194 9052 43234 9092
rect 43276 9052 43316 9092
rect 43358 9052 43398 9092
rect 43440 9052 43480 9092
rect 47112 9052 47152 9092
rect 47194 9052 47234 9092
rect 47276 9052 47316 9092
rect 47358 9052 47398 9092
rect 47440 9052 47480 9092
rect 51112 9052 51152 9092
rect 51194 9052 51234 9092
rect 51276 9052 51316 9092
rect 51358 9052 51398 9092
rect 51440 9052 51480 9092
rect 55112 9052 55152 9092
rect 55194 9052 55234 9092
rect 55276 9052 55316 9092
rect 55358 9052 55398 9092
rect 55440 9052 55480 9092
rect 59112 9052 59152 9092
rect 59194 9052 59234 9092
rect 59276 9052 59316 9092
rect 59358 9052 59398 9092
rect 59440 9052 59480 9092
rect 63112 9052 63152 9092
rect 63194 9052 63234 9092
rect 63276 9052 63316 9092
rect 63358 9052 63398 9092
rect 63440 9052 63480 9092
rect 67112 9052 67152 9092
rect 67194 9052 67234 9092
rect 67276 9052 67316 9092
rect 67358 9052 67398 9092
rect 67440 9052 67480 9092
rect 4352 8296 4392 8336
rect 4434 8296 4474 8336
rect 4516 8296 4556 8336
rect 4598 8296 4638 8336
rect 4680 8296 4720 8336
rect 8352 8296 8392 8336
rect 8434 8296 8474 8336
rect 8516 8296 8556 8336
rect 8598 8296 8638 8336
rect 8680 8296 8720 8336
rect 12352 8296 12392 8336
rect 12434 8296 12474 8336
rect 12516 8296 12556 8336
rect 12598 8296 12638 8336
rect 12680 8296 12720 8336
rect 16352 8296 16392 8336
rect 16434 8296 16474 8336
rect 16516 8296 16556 8336
rect 16598 8296 16638 8336
rect 16680 8296 16720 8336
rect 20352 8296 20392 8336
rect 20434 8296 20474 8336
rect 20516 8296 20556 8336
rect 20598 8296 20638 8336
rect 20680 8296 20720 8336
rect 24352 8296 24392 8336
rect 24434 8296 24474 8336
rect 24516 8296 24556 8336
rect 24598 8296 24638 8336
rect 24680 8296 24720 8336
rect 28352 8296 28392 8336
rect 28434 8296 28474 8336
rect 28516 8296 28556 8336
rect 28598 8296 28638 8336
rect 28680 8296 28720 8336
rect 32352 8296 32392 8336
rect 32434 8296 32474 8336
rect 32516 8296 32556 8336
rect 32598 8296 32638 8336
rect 32680 8296 32720 8336
rect 36352 8296 36392 8336
rect 36434 8296 36474 8336
rect 36516 8296 36556 8336
rect 36598 8296 36638 8336
rect 36680 8296 36720 8336
rect 40352 8296 40392 8336
rect 40434 8296 40474 8336
rect 40516 8296 40556 8336
rect 40598 8296 40638 8336
rect 40680 8296 40720 8336
rect 44352 8296 44392 8336
rect 44434 8296 44474 8336
rect 44516 8296 44556 8336
rect 44598 8296 44638 8336
rect 44680 8296 44720 8336
rect 48352 8296 48392 8336
rect 48434 8296 48474 8336
rect 48516 8296 48556 8336
rect 48598 8296 48638 8336
rect 48680 8296 48720 8336
rect 52352 8296 52392 8336
rect 52434 8296 52474 8336
rect 52516 8296 52556 8336
rect 52598 8296 52638 8336
rect 52680 8296 52720 8336
rect 56352 8296 56392 8336
rect 56434 8296 56474 8336
rect 56516 8296 56556 8336
rect 56598 8296 56638 8336
rect 56680 8296 56720 8336
rect 60352 8296 60392 8336
rect 60434 8296 60474 8336
rect 60516 8296 60556 8336
rect 60598 8296 60638 8336
rect 60680 8296 60720 8336
rect 64352 8296 64392 8336
rect 64434 8296 64474 8336
rect 64516 8296 64556 8336
rect 64598 8296 64638 8336
rect 64680 8296 64720 8336
rect 68352 8296 68392 8336
rect 68434 8296 68474 8336
rect 68516 8296 68556 8336
rect 68598 8296 68638 8336
rect 68680 8296 68720 8336
rect 3112 7540 3152 7580
rect 3194 7540 3234 7580
rect 3276 7540 3316 7580
rect 3358 7540 3398 7580
rect 3440 7540 3480 7580
rect 7112 7540 7152 7580
rect 7194 7540 7234 7580
rect 7276 7540 7316 7580
rect 7358 7540 7398 7580
rect 7440 7540 7480 7580
rect 11112 7540 11152 7580
rect 11194 7540 11234 7580
rect 11276 7540 11316 7580
rect 11358 7540 11398 7580
rect 11440 7540 11480 7580
rect 15112 7540 15152 7580
rect 15194 7540 15234 7580
rect 15276 7540 15316 7580
rect 15358 7540 15398 7580
rect 15440 7540 15480 7580
rect 19112 7540 19152 7580
rect 19194 7540 19234 7580
rect 19276 7540 19316 7580
rect 19358 7540 19398 7580
rect 19440 7540 19480 7580
rect 23112 7540 23152 7580
rect 23194 7540 23234 7580
rect 23276 7540 23316 7580
rect 23358 7540 23398 7580
rect 23440 7540 23480 7580
rect 27112 7540 27152 7580
rect 27194 7540 27234 7580
rect 27276 7540 27316 7580
rect 27358 7540 27398 7580
rect 27440 7540 27480 7580
rect 31112 7540 31152 7580
rect 31194 7540 31234 7580
rect 31276 7540 31316 7580
rect 31358 7540 31398 7580
rect 31440 7540 31480 7580
rect 35112 7540 35152 7580
rect 35194 7540 35234 7580
rect 35276 7540 35316 7580
rect 35358 7540 35398 7580
rect 35440 7540 35480 7580
rect 39112 7540 39152 7580
rect 39194 7540 39234 7580
rect 39276 7540 39316 7580
rect 39358 7540 39398 7580
rect 39440 7540 39480 7580
rect 43112 7540 43152 7580
rect 43194 7540 43234 7580
rect 43276 7540 43316 7580
rect 43358 7540 43398 7580
rect 43440 7540 43480 7580
rect 47112 7540 47152 7580
rect 47194 7540 47234 7580
rect 47276 7540 47316 7580
rect 47358 7540 47398 7580
rect 47440 7540 47480 7580
rect 51112 7540 51152 7580
rect 51194 7540 51234 7580
rect 51276 7540 51316 7580
rect 51358 7540 51398 7580
rect 51440 7540 51480 7580
rect 55112 7540 55152 7580
rect 55194 7540 55234 7580
rect 55276 7540 55316 7580
rect 55358 7540 55398 7580
rect 55440 7540 55480 7580
rect 59112 7540 59152 7580
rect 59194 7540 59234 7580
rect 59276 7540 59316 7580
rect 59358 7540 59398 7580
rect 59440 7540 59480 7580
rect 63112 7540 63152 7580
rect 63194 7540 63234 7580
rect 63276 7540 63316 7580
rect 63358 7540 63398 7580
rect 63440 7540 63480 7580
rect 67112 7540 67152 7580
rect 67194 7540 67234 7580
rect 67276 7540 67316 7580
rect 67358 7540 67398 7580
rect 67440 7540 67480 7580
rect 86668 7456 86708 7496
rect 4352 6784 4392 6824
rect 4434 6784 4474 6824
rect 4516 6784 4556 6824
rect 4598 6784 4638 6824
rect 4680 6784 4720 6824
rect 8352 6784 8392 6824
rect 8434 6784 8474 6824
rect 8516 6784 8556 6824
rect 8598 6784 8638 6824
rect 8680 6784 8720 6824
rect 12352 6784 12392 6824
rect 12434 6784 12474 6824
rect 12516 6784 12556 6824
rect 12598 6784 12638 6824
rect 12680 6784 12720 6824
rect 16352 6784 16392 6824
rect 16434 6784 16474 6824
rect 16516 6784 16556 6824
rect 16598 6784 16638 6824
rect 16680 6784 16720 6824
rect 20352 6784 20392 6824
rect 20434 6784 20474 6824
rect 20516 6784 20556 6824
rect 20598 6784 20638 6824
rect 20680 6784 20720 6824
rect 24352 6784 24392 6824
rect 24434 6784 24474 6824
rect 24516 6784 24556 6824
rect 24598 6784 24638 6824
rect 24680 6784 24720 6824
rect 28352 6784 28392 6824
rect 28434 6784 28474 6824
rect 28516 6784 28556 6824
rect 28598 6784 28638 6824
rect 28680 6784 28720 6824
rect 32352 6784 32392 6824
rect 32434 6784 32474 6824
rect 32516 6784 32556 6824
rect 32598 6784 32638 6824
rect 32680 6784 32720 6824
rect 36352 6784 36392 6824
rect 36434 6784 36474 6824
rect 36516 6784 36556 6824
rect 36598 6784 36638 6824
rect 36680 6784 36720 6824
rect 40352 6784 40392 6824
rect 40434 6784 40474 6824
rect 40516 6784 40556 6824
rect 40598 6784 40638 6824
rect 40680 6784 40720 6824
rect 44352 6784 44392 6824
rect 44434 6784 44474 6824
rect 44516 6784 44556 6824
rect 44598 6784 44638 6824
rect 44680 6784 44720 6824
rect 48352 6784 48392 6824
rect 48434 6784 48474 6824
rect 48516 6784 48556 6824
rect 48598 6784 48638 6824
rect 48680 6784 48720 6824
rect 52352 6784 52392 6824
rect 52434 6784 52474 6824
rect 52516 6784 52556 6824
rect 52598 6784 52638 6824
rect 52680 6784 52720 6824
rect 56352 6784 56392 6824
rect 56434 6784 56474 6824
rect 56516 6784 56556 6824
rect 56598 6784 56638 6824
rect 56680 6784 56720 6824
rect 60352 6784 60392 6824
rect 60434 6784 60474 6824
rect 60516 6784 60556 6824
rect 60598 6784 60638 6824
rect 60680 6784 60720 6824
rect 64352 6784 64392 6824
rect 64434 6784 64474 6824
rect 64516 6784 64556 6824
rect 64598 6784 64638 6824
rect 64680 6784 64720 6824
rect 68352 6784 68392 6824
rect 68434 6784 68474 6824
rect 68516 6784 68556 6824
rect 68598 6784 68638 6824
rect 68680 6784 68720 6824
rect 3112 6028 3152 6068
rect 3194 6028 3234 6068
rect 3276 6028 3316 6068
rect 3358 6028 3398 6068
rect 3440 6028 3480 6068
rect 7112 6028 7152 6068
rect 7194 6028 7234 6068
rect 7276 6028 7316 6068
rect 7358 6028 7398 6068
rect 7440 6028 7480 6068
rect 11112 6028 11152 6068
rect 11194 6028 11234 6068
rect 11276 6028 11316 6068
rect 11358 6028 11398 6068
rect 11440 6028 11480 6068
rect 15112 6028 15152 6068
rect 15194 6028 15234 6068
rect 15276 6028 15316 6068
rect 15358 6028 15398 6068
rect 15440 6028 15480 6068
rect 19112 6028 19152 6068
rect 19194 6028 19234 6068
rect 19276 6028 19316 6068
rect 19358 6028 19398 6068
rect 19440 6028 19480 6068
rect 23112 6028 23152 6068
rect 23194 6028 23234 6068
rect 23276 6028 23316 6068
rect 23358 6028 23398 6068
rect 23440 6028 23480 6068
rect 27112 6028 27152 6068
rect 27194 6028 27234 6068
rect 27276 6028 27316 6068
rect 27358 6028 27398 6068
rect 27440 6028 27480 6068
rect 31112 6028 31152 6068
rect 31194 6028 31234 6068
rect 31276 6028 31316 6068
rect 31358 6028 31398 6068
rect 31440 6028 31480 6068
rect 35112 6028 35152 6068
rect 35194 6028 35234 6068
rect 35276 6028 35316 6068
rect 35358 6028 35398 6068
rect 35440 6028 35480 6068
rect 39112 6028 39152 6068
rect 39194 6028 39234 6068
rect 39276 6028 39316 6068
rect 39358 6028 39398 6068
rect 39440 6028 39480 6068
rect 43112 6028 43152 6068
rect 43194 6028 43234 6068
rect 43276 6028 43316 6068
rect 43358 6028 43398 6068
rect 43440 6028 43480 6068
rect 47112 6028 47152 6068
rect 47194 6028 47234 6068
rect 47276 6028 47316 6068
rect 47358 6028 47398 6068
rect 47440 6028 47480 6068
rect 51112 6028 51152 6068
rect 51194 6028 51234 6068
rect 51276 6028 51316 6068
rect 51358 6028 51398 6068
rect 51440 6028 51480 6068
rect 55112 6028 55152 6068
rect 55194 6028 55234 6068
rect 55276 6028 55316 6068
rect 55358 6028 55398 6068
rect 55440 6028 55480 6068
rect 59112 6028 59152 6068
rect 59194 6028 59234 6068
rect 59276 6028 59316 6068
rect 59358 6028 59398 6068
rect 59440 6028 59480 6068
rect 63112 6028 63152 6068
rect 63194 6028 63234 6068
rect 63276 6028 63316 6068
rect 63358 6028 63398 6068
rect 63440 6028 63480 6068
rect 67112 6028 67152 6068
rect 67194 6028 67234 6068
rect 67276 6028 67316 6068
rect 67358 6028 67398 6068
rect 67440 6028 67480 6068
rect 4352 5272 4392 5312
rect 4434 5272 4474 5312
rect 4516 5272 4556 5312
rect 4598 5272 4638 5312
rect 4680 5272 4720 5312
rect 8352 5272 8392 5312
rect 8434 5272 8474 5312
rect 8516 5272 8556 5312
rect 8598 5272 8638 5312
rect 8680 5272 8720 5312
rect 12352 5272 12392 5312
rect 12434 5272 12474 5312
rect 12516 5272 12556 5312
rect 12598 5272 12638 5312
rect 12680 5272 12720 5312
rect 16352 5272 16392 5312
rect 16434 5272 16474 5312
rect 16516 5272 16556 5312
rect 16598 5272 16638 5312
rect 16680 5272 16720 5312
rect 20352 5272 20392 5312
rect 20434 5272 20474 5312
rect 20516 5272 20556 5312
rect 20598 5272 20638 5312
rect 20680 5272 20720 5312
rect 24352 5272 24392 5312
rect 24434 5272 24474 5312
rect 24516 5272 24556 5312
rect 24598 5272 24638 5312
rect 24680 5272 24720 5312
rect 28352 5272 28392 5312
rect 28434 5272 28474 5312
rect 28516 5272 28556 5312
rect 28598 5272 28638 5312
rect 28680 5272 28720 5312
rect 32352 5272 32392 5312
rect 32434 5272 32474 5312
rect 32516 5272 32556 5312
rect 32598 5272 32638 5312
rect 32680 5272 32720 5312
rect 36352 5272 36392 5312
rect 36434 5272 36474 5312
rect 36516 5272 36556 5312
rect 36598 5272 36638 5312
rect 36680 5272 36720 5312
rect 40352 5272 40392 5312
rect 40434 5272 40474 5312
rect 40516 5272 40556 5312
rect 40598 5272 40638 5312
rect 40680 5272 40720 5312
rect 44352 5272 44392 5312
rect 44434 5272 44474 5312
rect 44516 5272 44556 5312
rect 44598 5272 44638 5312
rect 44680 5272 44720 5312
rect 48352 5272 48392 5312
rect 48434 5272 48474 5312
rect 48516 5272 48556 5312
rect 48598 5272 48638 5312
rect 48680 5272 48720 5312
rect 52352 5272 52392 5312
rect 52434 5272 52474 5312
rect 52516 5272 52556 5312
rect 52598 5272 52638 5312
rect 52680 5272 52720 5312
rect 56352 5272 56392 5312
rect 56434 5272 56474 5312
rect 56516 5272 56556 5312
rect 56598 5272 56638 5312
rect 56680 5272 56720 5312
rect 60352 5272 60392 5312
rect 60434 5272 60474 5312
rect 60516 5272 60556 5312
rect 60598 5272 60638 5312
rect 60680 5272 60720 5312
rect 64352 5272 64392 5312
rect 64434 5272 64474 5312
rect 64516 5272 64556 5312
rect 64598 5272 64638 5312
rect 64680 5272 64720 5312
rect 68352 5272 68392 5312
rect 68434 5272 68474 5312
rect 68516 5272 68556 5312
rect 68598 5272 68638 5312
rect 68680 5272 68720 5312
rect 72352 5272 72392 5312
rect 72434 5272 72474 5312
rect 72516 5272 72556 5312
rect 72598 5272 72638 5312
rect 72680 5272 72720 5312
rect 76352 5272 76392 5312
rect 76434 5272 76474 5312
rect 76516 5272 76556 5312
rect 76598 5272 76638 5312
rect 76680 5272 76720 5312
rect 80352 5272 80392 5312
rect 80434 5272 80474 5312
rect 80516 5272 80556 5312
rect 80598 5272 80638 5312
rect 80680 5272 80720 5312
rect 84352 5272 84392 5312
rect 84434 5272 84474 5312
rect 84516 5272 84556 5312
rect 84598 5272 84638 5312
rect 84680 5272 84720 5312
rect 88352 5272 88392 5312
rect 88434 5272 88474 5312
rect 88516 5272 88556 5312
rect 88598 5272 88638 5312
rect 88680 5272 88720 5312
rect 92352 5272 92392 5312
rect 92434 5272 92474 5312
rect 92516 5272 92556 5312
rect 92598 5272 92638 5312
rect 92680 5272 92720 5312
rect 96352 5272 96392 5312
rect 96434 5272 96474 5312
rect 96516 5272 96556 5312
rect 96598 5272 96638 5312
rect 96680 5272 96720 5312
rect 3112 4516 3152 4556
rect 3194 4516 3234 4556
rect 3276 4516 3316 4556
rect 3358 4516 3398 4556
rect 3440 4516 3480 4556
rect 7112 4516 7152 4556
rect 7194 4516 7234 4556
rect 7276 4516 7316 4556
rect 7358 4516 7398 4556
rect 7440 4516 7480 4556
rect 11112 4516 11152 4556
rect 11194 4516 11234 4556
rect 11276 4516 11316 4556
rect 11358 4516 11398 4556
rect 11440 4516 11480 4556
rect 15112 4516 15152 4556
rect 15194 4516 15234 4556
rect 15276 4516 15316 4556
rect 15358 4516 15398 4556
rect 15440 4516 15480 4556
rect 19112 4516 19152 4556
rect 19194 4516 19234 4556
rect 19276 4516 19316 4556
rect 19358 4516 19398 4556
rect 19440 4516 19480 4556
rect 23112 4516 23152 4556
rect 23194 4516 23234 4556
rect 23276 4516 23316 4556
rect 23358 4516 23398 4556
rect 23440 4516 23480 4556
rect 27112 4516 27152 4556
rect 27194 4516 27234 4556
rect 27276 4516 27316 4556
rect 27358 4516 27398 4556
rect 27440 4516 27480 4556
rect 31112 4516 31152 4556
rect 31194 4516 31234 4556
rect 31276 4516 31316 4556
rect 31358 4516 31398 4556
rect 31440 4516 31480 4556
rect 35112 4516 35152 4556
rect 35194 4516 35234 4556
rect 35276 4516 35316 4556
rect 35358 4516 35398 4556
rect 35440 4516 35480 4556
rect 39112 4516 39152 4556
rect 39194 4516 39234 4556
rect 39276 4516 39316 4556
rect 39358 4516 39398 4556
rect 39440 4516 39480 4556
rect 43112 4516 43152 4556
rect 43194 4516 43234 4556
rect 43276 4516 43316 4556
rect 43358 4516 43398 4556
rect 43440 4516 43480 4556
rect 47112 4516 47152 4556
rect 47194 4516 47234 4556
rect 47276 4516 47316 4556
rect 47358 4516 47398 4556
rect 47440 4516 47480 4556
rect 51112 4516 51152 4556
rect 51194 4516 51234 4556
rect 51276 4516 51316 4556
rect 51358 4516 51398 4556
rect 51440 4516 51480 4556
rect 55112 4516 55152 4556
rect 55194 4516 55234 4556
rect 55276 4516 55316 4556
rect 55358 4516 55398 4556
rect 55440 4516 55480 4556
rect 59112 4516 59152 4556
rect 59194 4516 59234 4556
rect 59276 4516 59316 4556
rect 59358 4516 59398 4556
rect 59440 4516 59480 4556
rect 63112 4516 63152 4556
rect 63194 4516 63234 4556
rect 63276 4516 63316 4556
rect 63358 4516 63398 4556
rect 63440 4516 63480 4556
rect 67112 4516 67152 4556
rect 67194 4516 67234 4556
rect 67276 4516 67316 4556
rect 67358 4516 67398 4556
rect 67440 4516 67480 4556
rect 71112 4516 71152 4556
rect 71194 4516 71234 4556
rect 71276 4516 71316 4556
rect 71358 4516 71398 4556
rect 71440 4516 71480 4556
rect 75112 4516 75152 4556
rect 75194 4516 75234 4556
rect 75276 4516 75316 4556
rect 75358 4516 75398 4556
rect 75440 4516 75480 4556
rect 79112 4516 79152 4556
rect 79194 4516 79234 4556
rect 79276 4516 79316 4556
rect 79358 4516 79398 4556
rect 79440 4516 79480 4556
rect 83112 4516 83152 4556
rect 83194 4516 83234 4556
rect 83276 4516 83316 4556
rect 83358 4516 83398 4556
rect 83440 4516 83480 4556
rect 87112 4516 87152 4556
rect 87194 4516 87234 4556
rect 87276 4516 87316 4556
rect 87358 4516 87398 4556
rect 87440 4516 87480 4556
rect 91112 4516 91152 4556
rect 91194 4516 91234 4556
rect 91276 4516 91316 4556
rect 91358 4516 91398 4556
rect 91440 4516 91480 4556
rect 95112 4516 95152 4556
rect 95194 4516 95234 4556
rect 95276 4516 95316 4556
rect 95358 4516 95398 4556
rect 95440 4516 95480 4556
rect 99112 4516 99152 4556
rect 99194 4516 99234 4556
rect 99276 4516 99316 4556
rect 99358 4516 99398 4556
rect 99440 4516 99480 4556
rect 4352 3760 4392 3800
rect 4434 3760 4474 3800
rect 4516 3760 4556 3800
rect 4598 3760 4638 3800
rect 4680 3760 4720 3800
rect 8352 3760 8392 3800
rect 8434 3760 8474 3800
rect 8516 3760 8556 3800
rect 8598 3760 8638 3800
rect 8680 3760 8720 3800
rect 12352 3760 12392 3800
rect 12434 3760 12474 3800
rect 12516 3760 12556 3800
rect 12598 3760 12638 3800
rect 12680 3760 12720 3800
rect 16352 3760 16392 3800
rect 16434 3760 16474 3800
rect 16516 3760 16556 3800
rect 16598 3760 16638 3800
rect 16680 3760 16720 3800
rect 20352 3760 20392 3800
rect 20434 3760 20474 3800
rect 20516 3760 20556 3800
rect 20598 3760 20638 3800
rect 20680 3760 20720 3800
rect 24352 3760 24392 3800
rect 24434 3760 24474 3800
rect 24516 3760 24556 3800
rect 24598 3760 24638 3800
rect 24680 3760 24720 3800
rect 28352 3760 28392 3800
rect 28434 3760 28474 3800
rect 28516 3760 28556 3800
rect 28598 3760 28638 3800
rect 28680 3760 28720 3800
rect 32352 3760 32392 3800
rect 32434 3760 32474 3800
rect 32516 3760 32556 3800
rect 32598 3760 32638 3800
rect 32680 3760 32720 3800
rect 36352 3760 36392 3800
rect 36434 3760 36474 3800
rect 36516 3760 36556 3800
rect 36598 3760 36638 3800
rect 36680 3760 36720 3800
rect 40352 3760 40392 3800
rect 40434 3760 40474 3800
rect 40516 3760 40556 3800
rect 40598 3760 40638 3800
rect 40680 3760 40720 3800
rect 44352 3760 44392 3800
rect 44434 3760 44474 3800
rect 44516 3760 44556 3800
rect 44598 3760 44638 3800
rect 44680 3760 44720 3800
rect 48352 3760 48392 3800
rect 48434 3760 48474 3800
rect 48516 3760 48556 3800
rect 48598 3760 48638 3800
rect 48680 3760 48720 3800
rect 52352 3760 52392 3800
rect 52434 3760 52474 3800
rect 52516 3760 52556 3800
rect 52598 3760 52638 3800
rect 52680 3760 52720 3800
rect 56352 3760 56392 3800
rect 56434 3760 56474 3800
rect 56516 3760 56556 3800
rect 56598 3760 56638 3800
rect 56680 3760 56720 3800
rect 60352 3760 60392 3800
rect 60434 3760 60474 3800
rect 60516 3760 60556 3800
rect 60598 3760 60638 3800
rect 60680 3760 60720 3800
rect 64352 3760 64392 3800
rect 64434 3760 64474 3800
rect 64516 3760 64556 3800
rect 64598 3760 64638 3800
rect 64680 3760 64720 3800
rect 68352 3760 68392 3800
rect 68434 3760 68474 3800
rect 68516 3760 68556 3800
rect 68598 3760 68638 3800
rect 68680 3760 68720 3800
rect 72352 3760 72392 3800
rect 72434 3760 72474 3800
rect 72516 3760 72556 3800
rect 72598 3760 72638 3800
rect 72680 3760 72720 3800
rect 76352 3760 76392 3800
rect 76434 3760 76474 3800
rect 76516 3760 76556 3800
rect 76598 3760 76638 3800
rect 76680 3760 76720 3800
rect 80352 3760 80392 3800
rect 80434 3760 80474 3800
rect 80516 3760 80556 3800
rect 80598 3760 80638 3800
rect 80680 3760 80720 3800
rect 84352 3760 84392 3800
rect 84434 3760 84474 3800
rect 84516 3760 84556 3800
rect 84598 3760 84638 3800
rect 84680 3760 84720 3800
rect 88352 3760 88392 3800
rect 88434 3760 88474 3800
rect 88516 3760 88556 3800
rect 88598 3760 88638 3800
rect 88680 3760 88720 3800
rect 92352 3760 92392 3800
rect 92434 3760 92474 3800
rect 92516 3760 92556 3800
rect 92598 3760 92638 3800
rect 92680 3760 92720 3800
rect 96352 3760 96392 3800
rect 96434 3760 96474 3800
rect 96516 3760 96556 3800
rect 96598 3760 96638 3800
rect 96680 3760 96720 3800
rect 3112 3004 3152 3044
rect 3194 3004 3234 3044
rect 3276 3004 3316 3044
rect 3358 3004 3398 3044
rect 3440 3004 3480 3044
rect 7112 3004 7152 3044
rect 7194 3004 7234 3044
rect 7276 3004 7316 3044
rect 7358 3004 7398 3044
rect 7440 3004 7480 3044
rect 11112 3004 11152 3044
rect 11194 3004 11234 3044
rect 11276 3004 11316 3044
rect 11358 3004 11398 3044
rect 11440 3004 11480 3044
rect 15112 3004 15152 3044
rect 15194 3004 15234 3044
rect 15276 3004 15316 3044
rect 15358 3004 15398 3044
rect 15440 3004 15480 3044
rect 19112 3004 19152 3044
rect 19194 3004 19234 3044
rect 19276 3004 19316 3044
rect 19358 3004 19398 3044
rect 19440 3004 19480 3044
rect 23112 3004 23152 3044
rect 23194 3004 23234 3044
rect 23276 3004 23316 3044
rect 23358 3004 23398 3044
rect 23440 3004 23480 3044
rect 27112 3004 27152 3044
rect 27194 3004 27234 3044
rect 27276 3004 27316 3044
rect 27358 3004 27398 3044
rect 27440 3004 27480 3044
rect 31112 3004 31152 3044
rect 31194 3004 31234 3044
rect 31276 3004 31316 3044
rect 31358 3004 31398 3044
rect 31440 3004 31480 3044
rect 35112 3004 35152 3044
rect 35194 3004 35234 3044
rect 35276 3004 35316 3044
rect 35358 3004 35398 3044
rect 35440 3004 35480 3044
rect 39112 3004 39152 3044
rect 39194 3004 39234 3044
rect 39276 3004 39316 3044
rect 39358 3004 39398 3044
rect 39440 3004 39480 3044
rect 43112 3004 43152 3044
rect 43194 3004 43234 3044
rect 43276 3004 43316 3044
rect 43358 3004 43398 3044
rect 43440 3004 43480 3044
rect 47112 3004 47152 3044
rect 47194 3004 47234 3044
rect 47276 3004 47316 3044
rect 47358 3004 47398 3044
rect 47440 3004 47480 3044
rect 51112 3004 51152 3044
rect 51194 3004 51234 3044
rect 51276 3004 51316 3044
rect 51358 3004 51398 3044
rect 51440 3004 51480 3044
rect 55112 3004 55152 3044
rect 55194 3004 55234 3044
rect 55276 3004 55316 3044
rect 55358 3004 55398 3044
rect 55440 3004 55480 3044
rect 59112 3004 59152 3044
rect 59194 3004 59234 3044
rect 59276 3004 59316 3044
rect 59358 3004 59398 3044
rect 59440 3004 59480 3044
rect 63112 3004 63152 3044
rect 63194 3004 63234 3044
rect 63276 3004 63316 3044
rect 63358 3004 63398 3044
rect 63440 3004 63480 3044
rect 67112 3004 67152 3044
rect 67194 3004 67234 3044
rect 67276 3004 67316 3044
rect 67358 3004 67398 3044
rect 67440 3004 67480 3044
rect 71112 3004 71152 3044
rect 71194 3004 71234 3044
rect 71276 3004 71316 3044
rect 71358 3004 71398 3044
rect 71440 3004 71480 3044
rect 75112 3004 75152 3044
rect 75194 3004 75234 3044
rect 75276 3004 75316 3044
rect 75358 3004 75398 3044
rect 75440 3004 75480 3044
rect 79112 3004 79152 3044
rect 79194 3004 79234 3044
rect 79276 3004 79316 3044
rect 79358 3004 79398 3044
rect 79440 3004 79480 3044
rect 83112 3004 83152 3044
rect 83194 3004 83234 3044
rect 83276 3004 83316 3044
rect 83358 3004 83398 3044
rect 83440 3004 83480 3044
rect 87112 3004 87152 3044
rect 87194 3004 87234 3044
rect 87276 3004 87316 3044
rect 87358 3004 87398 3044
rect 87440 3004 87480 3044
rect 91112 3004 91152 3044
rect 91194 3004 91234 3044
rect 91276 3004 91316 3044
rect 91358 3004 91398 3044
rect 91440 3004 91480 3044
rect 95112 3004 95152 3044
rect 95194 3004 95234 3044
rect 95276 3004 95316 3044
rect 95358 3004 95398 3044
rect 95440 3004 95480 3044
rect 99112 3004 99152 3044
rect 99194 3004 99234 3044
rect 99276 3004 99316 3044
rect 99358 3004 99398 3044
rect 99440 3004 99480 3044
rect 4352 2248 4392 2288
rect 4434 2248 4474 2288
rect 4516 2248 4556 2288
rect 4598 2248 4638 2288
rect 4680 2248 4720 2288
rect 8352 2248 8392 2288
rect 8434 2248 8474 2288
rect 8516 2248 8556 2288
rect 8598 2248 8638 2288
rect 8680 2248 8720 2288
rect 12352 2248 12392 2288
rect 12434 2248 12474 2288
rect 12516 2248 12556 2288
rect 12598 2248 12638 2288
rect 12680 2248 12720 2288
rect 16352 2248 16392 2288
rect 16434 2248 16474 2288
rect 16516 2248 16556 2288
rect 16598 2248 16638 2288
rect 16680 2248 16720 2288
rect 20352 2248 20392 2288
rect 20434 2248 20474 2288
rect 20516 2248 20556 2288
rect 20598 2248 20638 2288
rect 20680 2248 20720 2288
rect 24352 2248 24392 2288
rect 24434 2248 24474 2288
rect 24516 2248 24556 2288
rect 24598 2248 24638 2288
rect 24680 2248 24720 2288
rect 28352 2248 28392 2288
rect 28434 2248 28474 2288
rect 28516 2248 28556 2288
rect 28598 2248 28638 2288
rect 28680 2248 28720 2288
rect 32352 2248 32392 2288
rect 32434 2248 32474 2288
rect 32516 2248 32556 2288
rect 32598 2248 32638 2288
rect 32680 2248 32720 2288
rect 36352 2248 36392 2288
rect 36434 2248 36474 2288
rect 36516 2248 36556 2288
rect 36598 2248 36638 2288
rect 36680 2248 36720 2288
rect 40352 2248 40392 2288
rect 40434 2248 40474 2288
rect 40516 2248 40556 2288
rect 40598 2248 40638 2288
rect 40680 2248 40720 2288
rect 44352 2248 44392 2288
rect 44434 2248 44474 2288
rect 44516 2248 44556 2288
rect 44598 2248 44638 2288
rect 44680 2248 44720 2288
rect 48352 2248 48392 2288
rect 48434 2248 48474 2288
rect 48516 2248 48556 2288
rect 48598 2248 48638 2288
rect 48680 2248 48720 2288
rect 52352 2248 52392 2288
rect 52434 2248 52474 2288
rect 52516 2248 52556 2288
rect 52598 2248 52638 2288
rect 52680 2248 52720 2288
rect 56352 2248 56392 2288
rect 56434 2248 56474 2288
rect 56516 2248 56556 2288
rect 56598 2248 56638 2288
rect 56680 2248 56720 2288
rect 60352 2248 60392 2288
rect 60434 2248 60474 2288
rect 60516 2248 60556 2288
rect 60598 2248 60638 2288
rect 60680 2248 60720 2288
rect 64352 2248 64392 2288
rect 64434 2248 64474 2288
rect 64516 2248 64556 2288
rect 64598 2248 64638 2288
rect 64680 2248 64720 2288
rect 68352 2248 68392 2288
rect 68434 2248 68474 2288
rect 68516 2248 68556 2288
rect 68598 2248 68638 2288
rect 68680 2248 68720 2288
rect 72352 2248 72392 2288
rect 72434 2248 72474 2288
rect 72516 2248 72556 2288
rect 72598 2248 72638 2288
rect 72680 2248 72720 2288
rect 76352 2248 76392 2288
rect 76434 2248 76474 2288
rect 76516 2248 76556 2288
rect 76598 2248 76638 2288
rect 76680 2248 76720 2288
rect 80352 2248 80392 2288
rect 80434 2248 80474 2288
rect 80516 2248 80556 2288
rect 80598 2248 80638 2288
rect 80680 2248 80720 2288
rect 84352 2248 84392 2288
rect 84434 2248 84474 2288
rect 84516 2248 84556 2288
rect 84598 2248 84638 2288
rect 84680 2248 84720 2288
rect 88352 2248 88392 2288
rect 88434 2248 88474 2288
rect 88516 2248 88556 2288
rect 88598 2248 88638 2288
rect 88680 2248 88720 2288
rect 92352 2248 92392 2288
rect 92434 2248 92474 2288
rect 92516 2248 92556 2288
rect 92598 2248 92638 2288
rect 92680 2248 92720 2288
rect 96352 2248 96392 2288
rect 96434 2248 96474 2288
rect 96516 2248 96556 2288
rect 96598 2248 96638 2288
rect 96680 2248 96720 2288
rect 3112 1492 3152 1532
rect 3194 1492 3234 1532
rect 3276 1492 3316 1532
rect 3358 1492 3398 1532
rect 3440 1492 3480 1532
rect 7112 1492 7152 1532
rect 7194 1492 7234 1532
rect 7276 1492 7316 1532
rect 7358 1492 7398 1532
rect 7440 1492 7480 1532
rect 11112 1492 11152 1532
rect 11194 1492 11234 1532
rect 11276 1492 11316 1532
rect 11358 1492 11398 1532
rect 11440 1492 11480 1532
rect 15112 1492 15152 1532
rect 15194 1492 15234 1532
rect 15276 1492 15316 1532
rect 15358 1492 15398 1532
rect 15440 1492 15480 1532
rect 19112 1492 19152 1532
rect 19194 1492 19234 1532
rect 19276 1492 19316 1532
rect 19358 1492 19398 1532
rect 19440 1492 19480 1532
rect 23112 1492 23152 1532
rect 23194 1492 23234 1532
rect 23276 1492 23316 1532
rect 23358 1492 23398 1532
rect 23440 1492 23480 1532
rect 27112 1492 27152 1532
rect 27194 1492 27234 1532
rect 27276 1492 27316 1532
rect 27358 1492 27398 1532
rect 27440 1492 27480 1532
rect 31112 1492 31152 1532
rect 31194 1492 31234 1532
rect 31276 1492 31316 1532
rect 31358 1492 31398 1532
rect 31440 1492 31480 1532
rect 35112 1492 35152 1532
rect 35194 1492 35234 1532
rect 35276 1492 35316 1532
rect 35358 1492 35398 1532
rect 35440 1492 35480 1532
rect 39112 1492 39152 1532
rect 39194 1492 39234 1532
rect 39276 1492 39316 1532
rect 39358 1492 39398 1532
rect 39440 1492 39480 1532
rect 43112 1492 43152 1532
rect 43194 1492 43234 1532
rect 43276 1492 43316 1532
rect 43358 1492 43398 1532
rect 43440 1492 43480 1532
rect 47112 1492 47152 1532
rect 47194 1492 47234 1532
rect 47276 1492 47316 1532
rect 47358 1492 47398 1532
rect 47440 1492 47480 1532
rect 51112 1492 51152 1532
rect 51194 1492 51234 1532
rect 51276 1492 51316 1532
rect 51358 1492 51398 1532
rect 51440 1492 51480 1532
rect 55112 1492 55152 1532
rect 55194 1492 55234 1532
rect 55276 1492 55316 1532
rect 55358 1492 55398 1532
rect 55440 1492 55480 1532
rect 59112 1492 59152 1532
rect 59194 1492 59234 1532
rect 59276 1492 59316 1532
rect 59358 1492 59398 1532
rect 59440 1492 59480 1532
rect 63112 1492 63152 1532
rect 63194 1492 63234 1532
rect 63276 1492 63316 1532
rect 63358 1492 63398 1532
rect 63440 1492 63480 1532
rect 67112 1492 67152 1532
rect 67194 1492 67234 1532
rect 67276 1492 67316 1532
rect 67358 1492 67398 1532
rect 67440 1492 67480 1532
rect 71112 1492 71152 1532
rect 71194 1492 71234 1532
rect 71276 1492 71316 1532
rect 71358 1492 71398 1532
rect 71440 1492 71480 1532
rect 75112 1492 75152 1532
rect 75194 1492 75234 1532
rect 75276 1492 75316 1532
rect 75358 1492 75398 1532
rect 75440 1492 75480 1532
rect 79112 1492 79152 1532
rect 79194 1492 79234 1532
rect 79276 1492 79316 1532
rect 79358 1492 79398 1532
rect 79440 1492 79480 1532
rect 83112 1492 83152 1532
rect 83194 1492 83234 1532
rect 83276 1492 83316 1532
rect 83358 1492 83398 1532
rect 83440 1492 83480 1532
rect 87112 1492 87152 1532
rect 87194 1492 87234 1532
rect 87276 1492 87316 1532
rect 87358 1492 87398 1532
rect 87440 1492 87480 1532
rect 91112 1492 91152 1532
rect 91194 1492 91234 1532
rect 91276 1492 91316 1532
rect 91358 1492 91398 1532
rect 91440 1492 91480 1532
rect 95112 1492 95152 1532
rect 95194 1492 95234 1532
rect 95276 1492 95316 1532
rect 95358 1492 95398 1532
rect 95440 1492 95480 1532
rect 99112 1492 99152 1532
rect 99194 1492 99234 1532
rect 99276 1492 99316 1532
rect 99358 1492 99398 1532
rect 99440 1492 99480 1532
rect 4352 736 4392 776
rect 4434 736 4474 776
rect 4516 736 4556 776
rect 4598 736 4638 776
rect 4680 736 4720 776
rect 8352 736 8392 776
rect 8434 736 8474 776
rect 8516 736 8556 776
rect 8598 736 8638 776
rect 8680 736 8720 776
rect 12352 736 12392 776
rect 12434 736 12474 776
rect 12516 736 12556 776
rect 12598 736 12638 776
rect 12680 736 12720 776
rect 16352 736 16392 776
rect 16434 736 16474 776
rect 16516 736 16556 776
rect 16598 736 16638 776
rect 16680 736 16720 776
rect 20352 736 20392 776
rect 20434 736 20474 776
rect 20516 736 20556 776
rect 20598 736 20638 776
rect 20680 736 20720 776
rect 24352 736 24392 776
rect 24434 736 24474 776
rect 24516 736 24556 776
rect 24598 736 24638 776
rect 24680 736 24720 776
rect 28352 736 28392 776
rect 28434 736 28474 776
rect 28516 736 28556 776
rect 28598 736 28638 776
rect 28680 736 28720 776
rect 32352 736 32392 776
rect 32434 736 32474 776
rect 32516 736 32556 776
rect 32598 736 32638 776
rect 32680 736 32720 776
rect 36352 736 36392 776
rect 36434 736 36474 776
rect 36516 736 36556 776
rect 36598 736 36638 776
rect 36680 736 36720 776
rect 40352 736 40392 776
rect 40434 736 40474 776
rect 40516 736 40556 776
rect 40598 736 40638 776
rect 40680 736 40720 776
rect 44352 736 44392 776
rect 44434 736 44474 776
rect 44516 736 44556 776
rect 44598 736 44638 776
rect 44680 736 44720 776
rect 48352 736 48392 776
rect 48434 736 48474 776
rect 48516 736 48556 776
rect 48598 736 48638 776
rect 48680 736 48720 776
rect 52352 736 52392 776
rect 52434 736 52474 776
rect 52516 736 52556 776
rect 52598 736 52638 776
rect 52680 736 52720 776
rect 56352 736 56392 776
rect 56434 736 56474 776
rect 56516 736 56556 776
rect 56598 736 56638 776
rect 56680 736 56720 776
rect 60352 736 60392 776
rect 60434 736 60474 776
rect 60516 736 60556 776
rect 60598 736 60638 776
rect 60680 736 60720 776
rect 64352 736 64392 776
rect 64434 736 64474 776
rect 64516 736 64556 776
rect 64598 736 64638 776
rect 64680 736 64720 776
rect 68352 736 68392 776
rect 68434 736 68474 776
rect 68516 736 68556 776
rect 68598 736 68638 776
rect 68680 736 68720 776
rect 72352 736 72392 776
rect 72434 736 72474 776
rect 72516 736 72556 776
rect 72598 736 72638 776
rect 72680 736 72720 776
rect 76352 736 76392 776
rect 76434 736 76474 776
rect 76516 736 76556 776
rect 76598 736 76638 776
rect 76680 736 76720 776
rect 80352 736 80392 776
rect 80434 736 80474 776
rect 80516 736 80556 776
rect 80598 736 80638 776
rect 80680 736 80720 776
rect 84352 736 84392 776
rect 84434 736 84474 776
rect 84516 736 84556 776
rect 84598 736 84638 776
rect 84680 736 84720 776
rect 88352 736 88392 776
rect 88434 736 88474 776
rect 88516 736 88556 776
rect 88598 736 88638 776
rect 88680 736 88720 776
rect 92352 736 92392 776
rect 92434 736 92474 776
rect 92516 736 92556 776
rect 92598 736 92638 776
rect 92680 736 92720 776
rect 96352 736 96392 776
rect 96434 736 96474 776
rect 96516 736 96556 776
rect 96598 736 96638 776
rect 96680 736 96720 776
<< metal5 >>
rect 4343 38599 4729 38618
rect 4343 38576 4409 38599
rect 4495 38576 4577 38599
rect 4663 38576 4729 38599
rect 4343 38536 4352 38576
rect 4392 38536 4409 38576
rect 4495 38536 4516 38576
rect 4556 38536 4577 38576
rect 4663 38536 4680 38576
rect 4720 38536 4729 38576
rect 4343 38513 4409 38536
rect 4495 38513 4577 38536
rect 4663 38513 4729 38536
rect 4343 38494 4729 38513
rect 8343 38599 8729 38618
rect 8343 38576 8409 38599
rect 8495 38576 8577 38599
rect 8663 38576 8729 38599
rect 8343 38536 8352 38576
rect 8392 38536 8409 38576
rect 8495 38536 8516 38576
rect 8556 38536 8577 38576
rect 8663 38536 8680 38576
rect 8720 38536 8729 38576
rect 8343 38513 8409 38536
rect 8495 38513 8577 38536
rect 8663 38513 8729 38536
rect 8343 38494 8729 38513
rect 12343 38599 12729 38618
rect 12343 38576 12409 38599
rect 12495 38576 12577 38599
rect 12663 38576 12729 38599
rect 12343 38536 12352 38576
rect 12392 38536 12409 38576
rect 12495 38536 12516 38576
rect 12556 38536 12577 38576
rect 12663 38536 12680 38576
rect 12720 38536 12729 38576
rect 12343 38513 12409 38536
rect 12495 38513 12577 38536
rect 12663 38513 12729 38536
rect 12343 38494 12729 38513
rect 16343 38599 16729 38618
rect 16343 38576 16409 38599
rect 16495 38576 16577 38599
rect 16663 38576 16729 38599
rect 16343 38536 16352 38576
rect 16392 38536 16409 38576
rect 16495 38536 16516 38576
rect 16556 38536 16577 38576
rect 16663 38536 16680 38576
rect 16720 38536 16729 38576
rect 16343 38513 16409 38536
rect 16495 38513 16577 38536
rect 16663 38513 16729 38536
rect 16343 38494 16729 38513
rect 20343 38599 20729 38618
rect 20343 38576 20409 38599
rect 20495 38576 20577 38599
rect 20663 38576 20729 38599
rect 20343 38536 20352 38576
rect 20392 38536 20409 38576
rect 20495 38536 20516 38576
rect 20556 38536 20577 38576
rect 20663 38536 20680 38576
rect 20720 38536 20729 38576
rect 20343 38513 20409 38536
rect 20495 38513 20577 38536
rect 20663 38513 20729 38536
rect 20343 38494 20729 38513
rect 24343 38599 24729 38618
rect 24343 38576 24409 38599
rect 24495 38576 24577 38599
rect 24663 38576 24729 38599
rect 24343 38536 24352 38576
rect 24392 38536 24409 38576
rect 24495 38536 24516 38576
rect 24556 38536 24577 38576
rect 24663 38536 24680 38576
rect 24720 38536 24729 38576
rect 24343 38513 24409 38536
rect 24495 38513 24577 38536
rect 24663 38513 24729 38536
rect 24343 38494 24729 38513
rect 28343 38599 28729 38618
rect 28343 38576 28409 38599
rect 28495 38576 28577 38599
rect 28663 38576 28729 38599
rect 28343 38536 28352 38576
rect 28392 38536 28409 38576
rect 28495 38536 28516 38576
rect 28556 38536 28577 38576
rect 28663 38536 28680 38576
rect 28720 38536 28729 38576
rect 28343 38513 28409 38536
rect 28495 38513 28577 38536
rect 28663 38513 28729 38536
rect 28343 38494 28729 38513
rect 32343 38599 32729 38618
rect 32343 38576 32409 38599
rect 32495 38576 32577 38599
rect 32663 38576 32729 38599
rect 32343 38536 32352 38576
rect 32392 38536 32409 38576
rect 32495 38536 32516 38576
rect 32556 38536 32577 38576
rect 32663 38536 32680 38576
rect 32720 38536 32729 38576
rect 32343 38513 32409 38536
rect 32495 38513 32577 38536
rect 32663 38513 32729 38536
rect 32343 38494 32729 38513
rect 36343 38599 36729 38618
rect 36343 38576 36409 38599
rect 36495 38576 36577 38599
rect 36663 38576 36729 38599
rect 36343 38536 36352 38576
rect 36392 38536 36409 38576
rect 36495 38536 36516 38576
rect 36556 38536 36577 38576
rect 36663 38536 36680 38576
rect 36720 38536 36729 38576
rect 36343 38513 36409 38536
rect 36495 38513 36577 38536
rect 36663 38513 36729 38536
rect 36343 38494 36729 38513
rect 40343 38599 40729 38618
rect 40343 38576 40409 38599
rect 40495 38576 40577 38599
rect 40663 38576 40729 38599
rect 40343 38536 40352 38576
rect 40392 38536 40409 38576
rect 40495 38536 40516 38576
rect 40556 38536 40577 38576
rect 40663 38536 40680 38576
rect 40720 38536 40729 38576
rect 40343 38513 40409 38536
rect 40495 38513 40577 38536
rect 40663 38513 40729 38536
rect 40343 38494 40729 38513
rect 44343 38599 44729 38618
rect 44343 38576 44409 38599
rect 44495 38576 44577 38599
rect 44663 38576 44729 38599
rect 44343 38536 44352 38576
rect 44392 38536 44409 38576
rect 44495 38536 44516 38576
rect 44556 38536 44577 38576
rect 44663 38536 44680 38576
rect 44720 38536 44729 38576
rect 44343 38513 44409 38536
rect 44495 38513 44577 38536
rect 44663 38513 44729 38536
rect 44343 38494 44729 38513
rect 48343 38599 48729 38618
rect 48343 38576 48409 38599
rect 48495 38576 48577 38599
rect 48663 38576 48729 38599
rect 48343 38536 48352 38576
rect 48392 38536 48409 38576
rect 48495 38536 48516 38576
rect 48556 38536 48577 38576
rect 48663 38536 48680 38576
rect 48720 38536 48729 38576
rect 48343 38513 48409 38536
rect 48495 38513 48577 38536
rect 48663 38513 48729 38536
rect 48343 38494 48729 38513
rect 52343 38599 52729 38618
rect 52343 38576 52409 38599
rect 52495 38576 52577 38599
rect 52663 38576 52729 38599
rect 52343 38536 52352 38576
rect 52392 38536 52409 38576
rect 52495 38536 52516 38576
rect 52556 38536 52577 38576
rect 52663 38536 52680 38576
rect 52720 38536 52729 38576
rect 52343 38513 52409 38536
rect 52495 38513 52577 38536
rect 52663 38513 52729 38536
rect 52343 38494 52729 38513
rect 56343 38599 56729 38618
rect 56343 38576 56409 38599
rect 56495 38576 56577 38599
rect 56663 38576 56729 38599
rect 56343 38536 56352 38576
rect 56392 38536 56409 38576
rect 56495 38536 56516 38576
rect 56556 38536 56577 38576
rect 56663 38536 56680 38576
rect 56720 38536 56729 38576
rect 56343 38513 56409 38536
rect 56495 38513 56577 38536
rect 56663 38513 56729 38536
rect 56343 38494 56729 38513
rect 60343 38599 60729 38618
rect 60343 38576 60409 38599
rect 60495 38576 60577 38599
rect 60663 38576 60729 38599
rect 60343 38536 60352 38576
rect 60392 38536 60409 38576
rect 60495 38536 60516 38576
rect 60556 38536 60577 38576
rect 60663 38536 60680 38576
rect 60720 38536 60729 38576
rect 60343 38513 60409 38536
rect 60495 38513 60577 38536
rect 60663 38513 60729 38536
rect 60343 38494 60729 38513
rect 64343 38599 64729 38618
rect 64343 38576 64409 38599
rect 64495 38576 64577 38599
rect 64663 38576 64729 38599
rect 64343 38536 64352 38576
rect 64392 38536 64409 38576
rect 64495 38536 64516 38576
rect 64556 38536 64577 38576
rect 64663 38536 64680 38576
rect 64720 38536 64729 38576
rect 64343 38513 64409 38536
rect 64495 38513 64577 38536
rect 64663 38513 64729 38536
rect 64343 38494 64729 38513
rect 68343 38599 68729 38618
rect 68343 38576 68409 38599
rect 68495 38576 68577 38599
rect 68663 38576 68729 38599
rect 68343 38536 68352 38576
rect 68392 38536 68409 38576
rect 68495 38536 68516 38576
rect 68556 38536 68577 38576
rect 68663 38536 68680 38576
rect 68720 38536 68729 38576
rect 68343 38513 68409 38536
rect 68495 38513 68577 38536
rect 68663 38513 68729 38536
rect 68343 38494 68729 38513
rect 72343 38599 72729 38618
rect 72343 38576 72409 38599
rect 72495 38576 72577 38599
rect 72663 38576 72729 38599
rect 72343 38536 72352 38576
rect 72392 38536 72409 38576
rect 72495 38536 72516 38576
rect 72556 38536 72577 38576
rect 72663 38536 72680 38576
rect 72720 38536 72729 38576
rect 72343 38513 72409 38536
rect 72495 38513 72577 38536
rect 72663 38513 72729 38536
rect 72343 38494 72729 38513
rect 76343 38599 76729 38618
rect 76343 38576 76409 38599
rect 76495 38576 76577 38599
rect 76663 38576 76729 38599
rect 76343 38536 76352 38576
rect 76392 38536 76409 38576
rect 76495 38536 76516 38576
rect 76556 38536 76577 38576
rect 76663 38536 76680 38576
rect 76720 38536 76729 38576
rect 76343 38513 76409 38536
rect 76495 38513 76577 38536
rect 76663 38513 76729 38536
rect 76343 38494 76729 38513
rect 80343 38599 80729 38618
rect 80343 38576 80409 38599
rect 80495 38576 80577 38599
rect 80663 38576 80729 38599
rect 80343 38536 80352 38576
rect 80392 38536 80409 38576
rect 80495 38536 80516 38576
rect 80556 38536 80577 38576
rect 80663 38536 80680 38576
rect 80720 38536 80729 38576
rect 80343 38513 80409 38536
rect 80495 38513 80577 38536
rect 80663 38513 80729 38536
rect 80343 38494 80729 38513
rect 84343 38599 84729 38618
rect 84343 38576 84409 38599
rect 84495 38576 84577 38599
rect 84663 38576 84729 38599
rect 84343 38536 84352 38576
rect 84392 38536 84409 38576
rect 84495 38536 84516 38576
rect 84556 38536 84577 38576
rect 84663 38536 84680 38576
rect 84720 38536 84729 38576
rect 84343 38513 84409 38536
rect 84495 38513 84577 38536
rect 84663 38513 84729 38536
rect 84343 38494 84729 38513
rect 88343 38599 88729 38618
rect 88343 38576 88409 38599
rect 88495 38576 88577 38599
rect 88663 38576 88729 38599
rect 88343 38536 88352 38576
rect 88392 38536 88409 38576
rect 88495 38536 88516 38576
rect 88556 38536 88577 38576
rect 88663 38536 88680 38576
rect 88720 38536 88729 38576
rect 88343 38513 88409 38536
rect 88495 38513 88577 38536
rect 88663 38513 88729 38536
rect 88343 38494 88729 38513
rect 92343 38599 92729 38618
rect 92343 38576 92409 38599
rect 92495 38576 92577 38599
rect 92663 38576 92729 38599
rect 92343 38536 92352 38576
rect 92392 38536 92409 38576
rect 92495 38536 92516 38576
rect 92556 38536 92577 38576
rect 92663 38536 92680 38576
rect 92720 38536 92729 38576
rect 92343 38513 92409 38536
rect 92495 38513 92577 38536
rect 92663 38513 92729 38536
rect 92343 38494 92729 38513
rect 96343 38599 96729 38618
rect 96343 38576 96409 38599
rect 96495 38576 96577 38599
rect 96663 38576 96729 38599
rect 96343 38536 96352 38576
rect 96392 38536 96409 38576
rect 96495 38536 96516 38576
rect 96556 38536 96577 38576
rect 96663 38536 96680 38576
rect 96720 38536 96729 38576
rect 96343 38513 96409 38536
rect 96495 38513 96577 38536
rect 96663 38513 96729 38536
rect 96343 38494 96729 38513
rect 3103 37843 3489 37862
rect 3103 37820 3169 37843
rect 3255 37820 3337 37843
rect 3423 37820 3489 37843
rect 3103 37780 3112 37820
rect 3152 37780 3169 37820
rect 3255 37780 3276 37820
rect 3316 37780 3337 37820
rect 3423 37780 3440 37820
rect 3480 37780 3489 37820
rect 3103 37757 3169 37780
rect 3255 37757 3337 37780
rect 3423 37757 3489 37780
rect 3103 37738 3489 37757
rect 7103 37843 7489 37862
rect 7103 37820 7169 37843
rect 7255 37820 7337 37843
rect 7423 37820 7489 37843
rect 7103 37780 7112 37820
rect 7152 37780 7169 37820
rect 7255 37780 7276 37820
rect 7316 37780 7337 37820
rect 7423 37780 7440 37820
rect 7480 37780 7489 37820
rect 7103 37757 7169 37780
rect 7255 37757 7337 37780
rect 7423 37757 7489 37780
rect 7103 37738 7489 37757
rect 11103 37843 11489 37862
rect 11103 37820 11169 37843
rect 11255 37820 11337 37843
rect 11423 37820 11489 37843
rect 11103 37780 11112 37820
rect 11152 37780 11169 37820
rect 11255 37780 11276 37820
rect 11316 37780 11337 37820
rect 11423 37780 11440 37820
rect 11480 37780 11489 37820
rect 11103 37757 11169 37780
rect 11255 37757 11337 37780
rect 11423 37757 11489 37780
rect 11103 37738 11489 37757
rect 15103 37843 15489 37862
rect 15103 37820 15169 37843
rect 15255 37820 15337 37843
rect 15423 37820 15489 37843
rect 15103 37780 15112 37820
rect 15152 37780 15169 37820
rect 15255 37780 15276 37820
rect 15316 37780 15337 37820
rect 15423 37780 15440 37820
rect 15480 37780 15489 37820
rect 15103 37757 15169 37780
rect 15255 37757 15337 37780
rect 15423 37757 15489 37780
rect 15103 37738 15489 37757
rect 19103 37843 19489 37862
rect 19103 37820 19169 37843
rect 19255 37820 19337 37843
rect 19423 37820 19489 37843
rect 19103 37780 19112 37820
rect 19152 37780 19169 37820
rect 19255 37780 19276 37820
rect 19316 37780 19337 37820
rect 19423 37780 19440 37820
rect 19480 37780 19489 37820
rect 19103 37757 19169 37780
rect 19255 37757 19337 37780
rect 19423 37757 19489 37780
rect 19103 37738 19489 37757
rect 23103 37843 23489 37862
rect 23103 37820 23169 37843
rect 23255 37820 23337 37843
rect 23423 37820 23489 37843
rect 23103 37780 23112 37820
rect 23152 37780 23169 37820
rect 23255 37780 23276 37820
rect 23316 37780 23337 37820
rect 23423 37780 23440 37820
rect 23480 37780 23489 37820
rect 23103 37757 23169 37780
rect 23255 37757 23337 37780
rect 23423 37757 23489 37780
rect 23103 37738 23489 37757
rect 27103 37843 27489 37862
rect 27103 37820 27169 37843
rect 27255 37820 27337 37843
rect 27423 37820 27489 37843
rect 27103 37780 27112 37820
rect 27152 37780 27169 37820
rect 27255 37780 27276 37820
rect 27316 37780 27337 37820
rect 27423 37780 27440 37820
rect 27480 37780 27489 37820
rect 27103 37757 27169 37780
rect 27255 37757 27337 37780
rect 27423 37757 27489 37780
rect 27103 37738 27489 37757
rect 31103 37843 31489 37862
rect 31103 37820 31169 37843
rect 31255 37820 31337 37843
rect 31423 37820 31489 37843
rect 31103 37780 31112 37820
rect 31152 37780 31169 37820
rect 31255 37780 31276 37820
rect 31316 37780 31337 37820
rect 31423 37780 31440 37820
rect 31480 37780 31489 37820
rect 31103 37757 31169 37780
rect 31255 37757 31337 37780
rect 31423 37757 31489 37780
rect 31103 37738 31489 37757
rect 35103 37843 35489 37862
rect 35103 37820 35169 37843
rect 35255 37820 35337 37843
rect 35423 37820 35489 37843
rect 35103 37780 35112 37820
rect 35152 37780 35169 37820
rect 35255 37780 35276 37820
rect 35316 37780 35337 37820
rect 35423 37780 35440 37820
rect 35480 37780 35489 37820
rect 35103 37757 35169 37780
rect 35255 37757 35337 37780
rect 35423 37757 35489 37780
rect 35103 37738 35489 37757
rect 39103 37843 39489 37862
rect 39103 37820 39169 37843
rect 39255 37820 39337 37843
rect 39423 37820 39489 37843
rect 39103 37780 39112 37820
rect 39152 37780 39169 37820
rect 39255 37780 39276 37820
rect 39316 37780 39337 37820
rect 39423 37780 39440 37820
rect 39480 37780 39489 37820
rect 39103 37757 39169 37780
rect 39255 37757 39337 37780
rect 39423 37757 39489 37780
rect 39103 37738 39489 37757
rect 43103 37843 43489 37862
rect 43103 37820 43169 37843
rect 43255 37820 43337 37843
rect 43423 37820 43489 37843
rect 43103 37780 43112 37820
rect 43152 37780 43169 37820
rect 43255 37780 43276 37820
rect 43316 37780 43337 37820
rect 43423 37780 43440 37820
rect 43480 37780 43489 37820
rect 43103 37757 43169 37780
rect 43255 37757 43337 37780
rect 43423 37757 43489 37780
rect 43103 37738 43489 37757
rect 47103 37843 47489 37862
rect 47103 37820 47169 37843
rect 47255 37820 47337 37843
rect 47423 37820 47489 37843
rect 47103 37780 47112 37820
rect 47152 37780 47169 37820
rect 47255 37780 47276 37820
rect 47316 37780 47337 37820
rect 47423 37780 47440 37820
rect 47480 37780 47489 37820
rect 47103 37757 47169 37780
rect 47255 37757 47337 37780
rect 47423 37757 47489 37780
rect 47103 37738 47489 37757
rect 51103 37843 51489 37862
rect 51103 37820 51169 37843
rect 51255 37820 51337 37843
rect 51423 37820 51489 37843
rect 51103 37780 51112 37820
rect 51152 37780 51169 37820
rect 51255 37780 51276 37820
rect 51316 37780 51337 37820
rect 51423 37780 51440 37820
rect 51480 37780 51489 37820
rect 51103 37757 51169 37780
rect 51255 37757 51337 37780
rect 51423 37757 51489 37780
rect 51103 37738 51489 37757
rect 55103 37843 55489 37862
rect 55103 37820 55169 37843
rect 55255 37820 55337 37843
rect 55423 37820 55489 37843
rect 55103 37780 55112 37820
rect 55152 37780 55169 37820
rect 55255 37780 55276 37820
rect 55316 37780 55337 37820
rect 55423 37780 55440 37820
rect 55480 37780 55489 37820
rect 55103 37757 55169 37780
rect 55255 37757 55337 37780
rect 55423 37757 55489 37780
rect 55103 37738 55489 37757
rect 59103 37843 59489 37862
rect 59103 37820 59169 37843
rect 59255 37820 59337 37843
rect 59423 37820 59489 37843
rect 59103 37780 59112 37820
rect 59152 37780 59169 37820
rect 59255 37780 59276 37820
rect 59316 37780 59337 37820
rect 59423 37780 59440 37820
rect 59480 37780 59489 37820
rect 59103 37757 59169 37780
rect 59255 37757 59337 37780
rect 59423 37757 59489 37780
rect 59103 37738 59489 37757
rect 63103 37843 63489 37862
rect 63103 37820 63169 37843
rect 63255 37820 63337 37843
rect 63423 37820 63489 37843
rect 63103 37780 63112 37820
rect 63152 37780 63169 37820
rect 63255 37780 63276 37820
rect 63316 37780 63337 37820
rect 63423 37780 63440 37820
rect 63480 37780 63489 37820
rect 63103 37757 63169 37780
rect 63255 37757 63337 37780
rect 63423 37757 63489 37780
rect 63103 37738 63489 37757
rect 67103 37843 67489 37862
rect 67103 37820 67169 37843
rect 67255 37820 67337 37843
rect 67423 37820 67489 37843
rect 67103 37780 67112 37820
rect 67152 37780 67169 37820
rect 67255 37780 67276 37820
rect 67316 37780 67337 37820
rect 67423 37780 67440 37820
rect 67480 37780 67489 37820
rect 67103 37757 67169 37780
rect 67255 37757 67337 37780
rect 67423 37757 67489 37780
rect 67103 37738 67489 37757
rect 71103 37843 71489 37862
rect 71103 37820 71169 37843
rect 71255 37820 71337 37843
rect 71423 37820 71489 37843
rect 71103 37780 71112 37820
rect 71152 37780 71169 37820
rect 71255 37780 71276 37820
rect 71316 37780 71337 37820
rect 71423 37780 71440 37820
rect 71480 37780 71489 37820
rect 71103 37757 71169 37780
rect 71255 37757 71337 37780
rect 71423 37757 71489 37780
rect 71103 37738 71489 37757
rect 75103 37843 75489 37862
rect 75103 37820 75169 37843
rect 75255 37820 75337 37843
rect 75423 37820 75489 37843
rect 75103 37780 75112 37820
rect 75152 37780 75169 37820
rect 75255 37780 75276 37820
rect 75316 37780 75337 37820
rect 75423 37780 75440 37820
rect 75480 37780 75489 37820
rect 75103 37757 75169 37780
rect 75255 37757 75337 37780
rect 75423 37757 75489 37780
rect 75103 37738 75489 37757
rect 79103 37843 79489 37862
rect 79103 37820 79169 37843
rect 79255 37820 79337 37843
rect 79423 37820 79489 37843
rect 79103 37780 79112 37820
rect 79152 37780 79169 37820
rect 79255 37780 79276 37820
rect 79316 37780 79337 37820
rect 79423 37780 79440 37820
rect 79480 37780 79489 37820
rect 79103 37757 79169 37780
rect 79255 37757 79337 37780
rect 79423 37757 79489 37780
rect 79103 37738 79489 37757
rect 83103 37843 83489 37862
rect 83103 37820 83169 37843
rect 83255 37820 83337 37843
rect 83423 37820 83489 37843
rect 83103 37780 83112 37820
rect 83152 37780 83169 37820
rect 83255 37780 83276 37820
rect 83316 37780 83337 37820
rect 83423 37780 83440 37820
rect 83480 37780 83489 37820
rect 83103 37757 83169 37780
rect 83255 37757 83337 37780
rect 83423 37757 83489 37780
rect 83103 37738 83489 37757
rect 87103 37843 87489 37862
rect 87103 37820 87169 37843
rect 87255 37820 87337 37843
rect 87423 37820 87489 37843
rect 87103 37780 87112 37820
rect 87152 37780 87169 37820
rect 87255 37780 87276 37820
rect 87316 37780 87337 37820
rect 87423 37780 87440 37820
rect 87480 37780 87489 37820
rect 87103 37757 87169 37780
rect 87255 37757 87337 37780
rect 87423 37757 87489 37780
rect 87103 37738 87489 37757
rect 91103 37843 91489 37862
rect 91103 37820 91169 37843
rect 91255 37820 91337 37843
rect 91423 37820 91489 37843
rect 91103 37780 91112 37820
rect 91152 37780 91169 37820
rect 91255 37780 91276 37820
rect 91316 37780 91337 37820
rect 91423 37780 91440 37820
rect 91480 37780 91489 37820
rect 91103 37757 91169 37780
rect 91255 37757 91337 37780
rect 91423 37757 91489 37780
rect 91103 37738 91489 37757
rect 95103 37843 95489 37862
rect 95103 37820 95169 37843
rect 95255 37820 95337 37843
rect 95423 37820 95489 37843
rect 95103 37780 95112 37820
rect 95152 37780 95169 37820
rect 95255 37780 95276 37820
rect 95316 37780 95337 37820
rect 95423 37780 95440 37820
rect 95480 37780 95489 37820
rect 95103 37757 95169 37780
rect 95255 37757 95337 37780
rect 95423 37757 95489 37780
rect 95103 37738 95489 37757
rect 99103 37843 99489 37862
rect 99103 37820 99169 37843
rect 99255 37820 99337 37843
rect 99423 37820 99489 37843
rect 99103 37780 99112 37820
rect 99152 37780 99169 37820
rect 99255 37780 99276 37820
rect 99316 37780 99337 37820
rect 99423 37780 99440 37820
rect 99480 37780 99489 37820
rect 99103 37757 99169 37780
rect 99255 37757 99337 37780
rect 99423 37757 99489 37780
rect 99103 37738 99489 37757
rect 4343 37087 4729 37106
rect 4343 37064 4409 37087
rect 4495 37064 4577 37087
rect 4663 37064 4729 37087
rect 4343 37024 4352 37064
rect 4392 37024 4409 37064
rect 4495 37024 4516 37064
rect 4556 37024 4577 37064
rect 4663 37024 4680 37064
rect 4720 37024 4729 37064
rect 4343 37001 4409 37024
rect 4495 37001 4577 37024
rect 4663 37001 4729 37024
rect 4343 36982 4729 37001
rect 8343 37087 8729 37106
rect 8343 37064 8409 37087
rect 8495 37064 8577 37087
rect 8663 37064 8729 37087
rect 8343 37024 8352 37064
rect 8392 37024 8409 37064
rect 8495 37024 8516 37064
rect 8556 37024 8577 37064
rect 8663 37024 8680 37064
rect 8720 37024 8729 37064
rect 8343 37001 8409 37024
rect 8495 37001 8577 37024
rect 8663 37001 8729 37024
rect 8343 36982 8729 37001
rect 12343 37087 12729 37106
rect 12343 37064 12409 37087
rect 12495 37064 12577 37087
rect 12663 37064 12729 37087
rect 12343 37024 12352 37064
rect 12392 37024 12409 37064
rect 12495 37024 12516 37064
rect 12556 37024 12577 37064
rect 12663 37024 12680 37064
rect 12720 37024 12729 37064
rect 12343 37001 12409 37024
rect 12495 37001 12577 37024
rect 12663 37001 12729 37024
rect 12343 36982 12729 37001
rect 16343 37087 16729 37106
rect 16343 37064 16409 37087
rect 16495 37064 16577 37087
rect 16663 37064 16729 37087
rect 16343 37024 16352 37064
rect 16392 37024 16409 37064
rect 16495 37024 16516 37064
rect 16556 37024 16577 37064
rect 16663 37024 16680 37064
rect 16720 37024 16729 37064
rect 16343 37001 16409 37024
rect 16495 37001 16577 37024
rect 16663 37001 16729 37024
rect 16343 36982 16729 37001
rect 20343 37087 20729 37106
rect 20343 37064 20409 37087
rect 20495 37064 20577 37087
rect 20663 37064 20729 37087
rect 20343 37024 20352 37064
rect 20392 37024 20409 37064
rect 20495 37024 20516 37064
rect 20556 37024 20577 37064
rect 20663 37024 20680 37064
rect 20720 37024 20729 37064
rect 20343 37001 20409 37024
rect 20495 37001 20577 37024
rect 20663 37001 20729 37024
rect 20343 36982 20729 37001
rect 24343 37087 24729 37106
rect 24343 37064 24409 37087
rect 24495 37064 24577 37087
rect 24663 37064 24729 37087
rect 24343 37024 24352 37064
rect 24392 37024 24409 37064
rect 24495 37024 24516 37064
rect 24556 37024 24577 37064
rect 24663 37024 24680 37064
rect 24720 37024 24729 37064
rect 24343 37001 24409 37024
rect 24495 37001 24577 37024
rect 24663 37001 24729 37024
rect 24343 36982 24729 37001
rect 28343 37087 28729 37106
rect 28343 37064 28409 37087
rect 28495 37064 28577 37087
rect 28663 37064 28729 37087
rect 28343 37024 28352 37064
rect 28392 37024 28409 37064
rect 28495 37024 28516 37064
rect 28556 37024 28577 37064
rect 28663 37024 28680 37064
rect 28720 37024 28729 37064
rect 28343 37001 28409 37024
rect 28495 37001 28577 37024
rect 28663 37001 28729 37024
rect 28343 36982 28729 37001
rect 32343 37087 32729 37106
rect 32343 37064 32409 37087
rect 32495 37064 32577 37087
rect 32663 37064 32729 37087
rect 32343 37024 32352 37064
rect 32392 37024 32409 37064
rect 32495 37024 32516 37064
rect 32556 37024 32577 37064
rect 32663 37024 32680 37064
rect 32720 37024 32729 37064
rect 32343 37001 32409 37024
rect 32495 37001 32577 37024
rect 32663 37001 32729 37024
rect 32343 36982 32729 37001
rect 36343 37087 36729 37106
rect 36343 37064 36409 37087
rect 36495 37064 36577 37087
rect 36663 37064 36729 37087
rect 36343 37024 36352 37064
rect 36392 37024 36409 37064
rect 36495 37024 36516 37064
rect 36556 37024 36577 37064
rect 36663 37024 36680 37064
rect 36720 37024 36729 37064
rect 36343 37001 36409 37024
rect 36495 37001 36577 37024
rect 36663 37001 36729 37024
rect 36343 36982 36729 37001
rect 40343 37087 40729 37106
rect 40343 37064 40409 37087
rect 40495 37064 40577 37087
rect 40663 37064 40729 37087
rect 40343 37024 40352 37064
rect 40392 37024 40409 37064
rect 40495 37024 40516 37064
rect 40556 37024 40577 37064
rect 40663 37024 40680 37064
rect 40720 37024 40729 37064
rect 40343 37001 40409 37024
rect 40495 37001 40577 37024
rect 40663 37001 40729 37024
rect 40343 36982 40729 37001
rect 44343 37087 44729 37106
rect 44343 37064 44409 37087
rect 44495 37064 44577 37087
rect 44663 37064 44729 37087
rect 44343 37024 44352 37064
rect 44392 37024 44409 37064
rect 44495 37024 44516 37064
rect 44556 37024 44577 37064
rect 44663 37024 44680 37064
rect 44720 37024 44729 37064
rect 44343 37001 44409 37024
rect 44495 37001 44577 37024
rect 44663 37001 44729 37024
rect 44343 36982 44729 37001
rect 48343 37087 48729 37106
rect 48343 37064 48409 37087
rect 48495 37064 48577 37087
rect 48663 37064 48729 37087
rect 48343 37024 48352 37064
rect 48392 37024 48409 37064
rect 48495 37024 48516 37064
rect 48556 37024 48577 37064
rect 48663 37024 48680 37064
rect 48720 37024 48729 37064
rect 48343 37001 48409 37024
rect 48495 37001 48577 37024
rect 48663 37001 48729 37024
rect 48343 36982 48729 37001
rect 52343 37087 52729 37106
rect 52343 37064 52409 37087
rect 52495 37064 52577 37087
rect 52663 37064 52729 37087
rect 52343 37024 52352 37064
rect 52392 37024 52409 37064
rect 52495 37024 52516 37064
rect 52556 37024 52577 37064
rect 52663 37024 52680 37064
rect 52720 37024 52729 37064
rect 52343 37001 52409 37024
rect 52495 37001 52577 37024
rect 52663 37001 52729 37024
rect 52343 36982 52729 37001
rect 56343 37087 56729 37106
rect 56343 37064 56409 37087
rect 56495 37064 56577 37087
rect 56663 37064 56729 37087
rect 56343 37024 56352 37064
rect 56392 37024 56409 37064
rect 56495 37024 56516 37064
rect 56556 37024 56577 37064
rect 56663 37024 56680 37064
rect 56720 37024 56729 37064
rect 56343 37001 56409 37024
rect 56495 37001 56577 37024
rect 56663 37001 56729 37024
rect 56343 36982 56729 37001
rect 60343 37087 60729 37106
rect 60343 37064 60409 37087
rect 60495 37064 60577 37087
rect 60663 37064 60729 37087
rect 60343 37024 60352 37064
rect 60392 37024 60409 37064
rect 60495 37024 60516 37064
rect 60556 37024 60577 37064
rect 60663 37024 60680 37064
rect 60720 37024 60729 37064
rect 60343 37001 60409 37024
rect 60495 37001 60577 37024
rect 60663 37001 60729 37024
rect 60343 36982 60729 37001
rect 64343 37087 64729 37106
rect 64343 37064 64409 37087
rect 64495 37064 64577 37087
rect 64663 37064 64729 37087
rect 64343 37024 64352 37064
rect 64392 37024 64409 37064
rect 64495 37024 64516 37064
rect 64556 37024 64577 37064
rect 64663 37024 64680 37064
rect 64720 37024 64729 37064
rect 64343 37001 64409 37024
rect 64495 37001 64577 37024
rect 64663 37001 64729 37024
rect 64343 36982 64729 37001
rect 68343 37087 68729 37106
rect 68343 37064 68409 37087
rect 68495 37064 68577 37087
rect 68663 37064 68729 37087
rect 68343 37024 68352 37064
rect 68392 37024 68409 37064
rect 68495 37024 68516 37064
rect 68556 37024 68577 37064
rect 68663 37024 68680 37064
rect 68720 37024 68729 37064
rect 68343 37001 68409 37024
rect 68495 37001 68577 37024
rect 68663 37001 68729 37024
rect 68343 36982 68729 37001
rect 72343 37087 72729 37106
rect 72343 37064 72409 37087
rect 72495 37064 72577 37087
rect 72663 37064 72729 37087
rect 72343 37024 72352 37064
rect 72392 37024 72409 37064
rect 72495 37024 72516 37064
rect 72556 37024 72577 37064
rect 72663 37024 72680 37064
rect 72720 37024 72729 37064
rect 72343 37001 72409 37024
rect 72495 37001 72577 37024
rect 72663 37001 72729 37024
rect 72343 36982 72729 37001
rect 76343 37087 76729 37106
rect 76343 37064 76409 37087
rect 76495 37064 76577 37087
rect 76663 37064 76729 37087
rect 76343 37024 76352 37064
rect 76392 37024 76409 37064
rect 76495 37024 76516 37064
rect 76556 37024 76577 37064
rect 76663 37024 76680 37064
rect 76720 37024 76729 37064
rect 76343 37001 76409 37024
rect 76495 37001 76577 37024
rect 76663 37001 76729 37024
rect 76343 36982 76729 37001
rect 80343 37087 80729 37106
rect 80343 37064 80409 37087
rect 80495 37064 80577 37087
rect 80663 37064 80729 37087
rect 80343 37024 80352 37064
rect 80392 37024 80409 37064
rect 80495 37024 80516 37064
rect 80556 37024 80577 37064
rect 80663 37024 80680 37064
rect 80720 37024 80729 37064
rect 80343 37001 80409 37024
rect 80495 37001 80577 37024
rect 80663 37001 80729 37024
rect 80343 36982 80729 37001
rect 84343 37087 84729 37106
rect 84343 37064 84409 37087
rect 84495 37064 84577 37087
rect 84663 37064 84729 37087
rect 84343 37024 84352 37064
rect 84392 37024 84409 37064
rect 84495 37024 84516 37064
rect 84556 37024 84577 37064
rect 84663 37024 84680 37064
rect 84720 37024 84729 37064
rect 84343 37001 84409 37024
rect 84495 37001 84577 37024
rect 84663 37001 84729 37024
rect 84343 36982 84729 37001
rect 88343 37087 88729 37106
rect 88343 37064 88409 37087
rect 88495 37064 88577 37087
rect 88663 37064 88729 37087
rect 88343 37024 88352 37064
rect 88392 37024 88409 37064
rect 88495 37024 88516 37064
rect 88556 37024 88577 37064
rect 88663 37024 88680 37064
rect 88720 37024 88729 37064
rect 88343 37001 88409 37024
rect 88495 37001 88577 37024
rect 88663 37001 88729 37024
rect 88343 36982 88729 37001
rect 92343 37087 92729 37106
rect 92343 37064 92409 37087
rect 92495 37064 92577 37087
rect 92663 37064 92729 37087
rect 92343 37024 92352 37064
rect 92392 37024 92409 37064
rect 92495 37024 92516 37064
rect 92556 37024 92577 37064
rect 92663 37024 92680 37064
rect 92720 37024 92729 37064
rect 92343 37001 92409 37024
rect 92495 37001 92577 37024
rect 92663 37001 92729 37024
rect 92343 36982 92729 37001
rect 96343 37087 96729 37106
rect 96343 37064 96409 37087
rect 96495 37064 96577 37087
rect 96663 37064 96729 37087
rect 96343 37024 96352 37064
rect 96392 37024 96409 37064
rect 96495 37024 96516 37064
rect 96556 37024 96577 37064
rect 96663 37024 96680 37064
rect 96720 37024 96729 37064
rect 96343 37001 96409 37024
rect 96495 37001 96577 37024
rect 96663 37001 96729 37024
rect 96343 36982 96729 37001
rect 3103 36331 3489 36350
rect 3103 36308 3169 36331
rect 3255 36308 3337 36331
rect 3423 36308 3489 36331
rect 3103 36268 3112 36308
rect 3152 36268 3169 36308
rect 3255 36268 3276 36308
rect 3316 36268 3337 36308
rect 3423 36268 3440 36308
rect 3480 36268 3489 36308
rect 3103 36245 3169 36268
rect 3255 36245 3337 36268
rect 3423 36245 3489 36268
rect 3103 36226 3489 36245
rect 7103 36331 7489 36350
rect 7103 36308 7169 36331
rect 7255 36308 7337 36331
rect 7423 36308 7489 36331
rect 7103 36268 7112 36308
rect 7152 36268 7169 36308
rect 7255 36268 7276 36308
rect 7316 36268 7337 36308
rect 7423 36268 7440 36308
rect 7480 36268 7489 36308
rect 7103 36245 7169 36268
rect 7255 36245 7337 36268
rect 7423 36245 7489 36268
rect 7103 36226 7489 36245
rect 11103 36331 11489 36350
rect 11103 36308 11169 36331
rect 11255 36308 11337 36331
rect 11423 36308 11489 36331
rect 11103 36268 11112 36308
rect 11152 36268 11169 36308
rect 11255 36268 11276 36308
rect 11316 36268 11337 36308
rect 11423 36268 11440 36308
rect 11480 36268 11489 36308
rect 11103 36245 11169 36268
rect 11255 36245 11337 36268
rect 11423 36245 11489 36268
rect 11103 36226 11489 36245
rect 15103 36331 15489 36350
rect 15103 36308 15169 36331
rect 15255 36308 15337 36331
rect 15423 36308 15489 36331
rect 15103 36268 15112 36308
rect 15152 36268 15169 36308
rect 15255 36268 15276 36308
rect 15316 36268 15337 36308
rect 15423 36268 15440 36308
rect 15480 36268 15489 36308
rect 15103 36245 15169 36268
rect 15255 36245 15337 36268
rect 15423 36245 15489 36268
rect 15103 36226 15489 36245
rect 19103 36331 19489 36350
rect 19103 36308 19169 36331
rect 19255 36308 19337 36331
rect 19423 36308 19489 36331
rect 19103 36268 19112 36308
rect 19152 36268 19169 36308
rect 19255 36268 19276 36308
rect 19316 36268 19337 36308
rect 19423 36268 19440 36308
rect 19480 36268 19489 36308
rect 19103 36245 19169 36268
rect 19255 36245 19337 36268
rect 19423 36245 19489 36268
rect 19103 36226 19489 36245
rect 23103 36331 23489 36350
rect 23103 36308 23169 36331
rect 23255 36308 23337 36331
rect 23423 36308 23489 36331
rect 23103 36268 23112 36308
rect 23152 36268 23169 36308
rect 23255 36268 23276 36308
rect 23316 36268 23337 36308
rect 23423 36268 23440 36308
rect 23480 36268 23489 36308
rect 23103 36245 23169 36268
rect 23255 36245 23337 36268
rect 23423 36245 23489 36268
rect 23103 36226 23489 36245
rect 27103 36331 27489 36350
rect 27103 36308 27169 36331
rect 27255 36308 27337 36331
rect 27423 36308 27489 36331
rect 27103 36268 27112 36308
rect 27152 36268 27169 36308
rect 27255 36268 27276 36308
rect 27316 36268 27337 36308
rect 27423 36268 27440 36308
rect 27480 36268 27489 36308
rect 27103 36245 27169 36268
rect 27255 36245 27337 36268
rect 27423 36245 27489 36268
rect 27103 36226 27489 36245
rect 31103 36331 31489 36350
rect 31103 36308 31169 36331
rect 31255 36308 31337 36331
rect 31423 36308 31489 36331
rect 31103 36268 31112 36308
rect 31152 36268 31169 36308
rect 31255 36268 31276 36308
rect 31316 36268 31337 36308
rect 31423 36268 31440 36308
rect 31480 36268 31489 36308
rect 31103 36245 31169 36268
rect 31255 36245 31337 36268
rect 31423 36245 31489 36268
rect 31103 36226 31489 36245
rect 35103 36331 35489 36350
rect 35103 36308 35169 36331
rect 35255 36308 35337 36331
rect 35423 36308 35489 36331
rect 35103 36268 35112 36308
rect 35152 36268 35169 36308
rect 35255 36268 35276 36308
rect 35316 36268 35337 36308
rect 35423 36268 35440 36308
rect 35480 36268 35489 36308
rect 35103 36245 35169 36268
rect 35255 36245 35337 36268
rect 35423 36245 35489 36268
rect 35103 36226 35489 36245
rect 39103 36331 39489 36350
rect 39103 36308 39169 36331
rect 39255 36308 39337 36331
rect 39423 36308 39489 36331
rect 39103 36268 39112 36308
rect 39152 36268 39169 36308
rect 39255 36268 39276 36308
rect 39316 36268 39337 36308
rect 39423 36268 39440 36308
rect 39480 36268 39489 36308
rect 39103 36245 39169 36268
rect 39255 36245 39337 36268
rect 39423 36245 39489 36268
rect 39103 36226 39489 36245
rect 43103 36331 43489 36350
rect 43103 36308 43169 36331
rect 43255 36308 43337 36331
rect 43423 36308 43489 36331
rect 43103 36268 43112 36308
rect 43152 36268 43169 36308
rect 43255 36268 43276 36308
rect 43316 36268 43337 36308
rect 43423 36268 43440 36308
rect 43480 36268 43489 36308
rect 43103 36245 43169 36268
rect 43255 36245 43337 36268
rect 43423 36245 43489 36268
rect 43103 36226 43489 36245
rect 47103 36331 47489 36350
rect 47103 36308 47169 36331
rect 47255 36308 47337 36331
rect 47423 36308 47489 36331
rect 47103 36268 47112 36308
rect 47152 36268 47169 36308
rect 47255 36268 47276 36308
rect 47316 36268 47337 36308
rect 47423 36268 47440 36308
rect 47480 36268 47489 36308
rect 47103 36245 47169 36268
rect 47255 36245 47337 36268
rect 47423 36245 47489 36268
rect 47103 36226 47489 36245
rect 51103 36331 51489 36350
rect 51103 36308 51169 36331
rect 51255 36308 51337 36331
rect 51423 36308 51489 36331
rect 51103 36268 51112 36308
rect 51152 36268 51169 36308
rect 51255 36268 51276 36308
rect 51316 36268 51337 36308
rect 51423 36268 51440 36308
rect 51480 36268 51489 36308
rect 51103 36245 51169 36268
rect 51255 36245 51337 36268
rect 51423 36245 51489 36268
rect 51103 36226 51489 36245
rect 55103 36331 55489 36350
rect 55103 36308 55169 36331
rect 55255 36308 55337 36331
rect 55423 36308 55489 36331
rect 55103 36268 55112 36308
rect 55152 36268 55169 36308
rect 55255 36268 55276 36308
rect 55316 36268 55337 36308
rect 55423 36268 55440 36308
rect 55480 36268 55489 36308
rect 55103 36245 55169 36268
rect 55255 36245 55337 36268
rect 55423 36245 55489 36268
rect 55103 36226 55489 36245
rect 59103 36331 59489 36350
rect 59103 36308 59169 36331
rect 59255 36308 59337 36331
rect 59423 36308 59489 36331
rect 59103 36268 59112 36308
rect 59152 36268 59169 36308
rect 59255 36268 59276 36308
rect 59316 36268 59337 36308
rect 59423 36268 59440 36308
rect 59480 36268 59489 36308
rect 59103 36245 59169 36268
rect 59255 36245 59337 36268
rect 59423 36245 59489 36268
rect 59103 36226 59489 36245
rect 63103 36331 63489 36350
rect 63103 36308 63169 36331
rect 63255 36308 63337 36331
rect 63423 36308 63489 36331
rect 63103 36268 63112 36308
rect 63152 36268 63169 36308
rect 63255 36268 63276 36308
rect 63316 36268 63337 36308
rect 63423 36268 63440 36308
rect 63480 36268 63489 36308
rect 63103 36245 63169 36268
rect 63255 36245 63337 36268
rect 63423 36245 63489 36268
rect 63103 36226 63489 36245
rect 67103 36331 67489 36350
rect 67103 36308 67169 36331
rect 67255 36308 67337 36331
rect 67423 36308 67489 36331
rect 67103 36268 67112 36308
rect 67152 36268 67169 36308
rect 67255 36268 67276 36308
rect 67316 36268 67337 36308
rect 67423 36268 67440 36308
rect 67480 36268 67489 36308
rect 67103 36245 67169 36268
rect 67255 36245 67337 36268
rect 67423 36245 67489 36268
rect 67103 36226 67489 36245
rect 71103 36331 71489 36350
rect 71103 36308 71169 36331
rect 71255 36308 71337 36331
rect 71423 36308 71489 36331
rect 71103 36268 71112 36308
rect 71152 36268 71169 36308
rect 71255 36268 71276 36308
rect 71316 36268 71337 36308
rect 71423 36268 71440 36308
rect 71480 36268 71489 36308
rect 71103 36245 71169 36268
rect 71255 36245 71337 36268
rect 71423 36245 71489 36268
rect 71103 36226 71489 36245
rect 75103 36331 75489 36350
rect 75103 36308 75169 36331
rect 75255 36308 75337 36331
rect 75423 36308 75489 36331
rect 75103 36268 75112 36308
rect 75152 36268 75169 36308
rect 75255 36268 75276 36308
rect 75316 36268 75337 36308
rect 75423 36268 75440 36308
rect 75480 36268 75489 36308
rect 75103 36245 75169 36268
rect 75255 36245 75337 36268
rect 75423 36245 75489 36268
rect 75103 36226 75489 36245
rect 79103 36331 79489 36350
rect 79103 36308 79169 36331
rect 79255 36308 79337 36331
rect 79423 36308 79489 36331
rect 79103 36268 79112 36308
rect 79152 36268 79169 36308
rect 79255 36268 79276 36308
rect 79316 36268 79337 36308
rect 79423 36268 79440 36308
rect 79480 36268 79489 36308
rect 79103 36245 79169 36268
rect 79255 36245 79337 36268
rect 79423 36245 79489 36268
rect 79103 36226 79489 36245
rect 83103 36331 83489 36350
rect 83103 36308 83169 36331
rect 83255 36308 83337 36331
rect 83423 36308 83489 36331
rect 83103 36268 83112 36308
rect 83152 36268 83169 36308
rect 83255 36268 83276 36308
rect 83316 36268 83337 36308
rect 83423 36268 83440 36308
rect 83480 36268 83489 36308
rect 83103 36245 83169 36268
rect 83255 36245 83337 36268
rect 83423 36245 83489 36268
rect 83103 36226 83489 36245
rect 87103 36331 87489 36350
rect 87103 36308 87169 36331
rect 87255 36308 87337 36331
rect 87423 36308 87489 36331
rect 87103 36268 87112 36308
rect 87152 36268 87169 36308
rect 87255 36268 87276 36308
rect 87316 36268 87337 36308
rect 87423 36268 87440 36308
rect 87480 36268 87489 36308
rect 87103 36245 87169 36268
rect 87255 36245 87337 36268
rect 87423 36245 87489 36268
rect 87103 36226 87489 36245
rect 91103 36331 91489 36350
rect 91103 36308 91169 36331
rect 91255 36308 91337 36331
rect 91423 36308 91489 36331
rect 91103 36268 91112 36308
rect 91152 36268 91169 36308
rect 91255 36268 91276 36308
rect 91316 36268 91337 36308
rect 91423 36268 91440 36308
rect 91480 36268 91489 36308
rect 91103 36245 91169 36268
rect 91255 36245 91337 36268
rect 91423 36245 91489 36268
rect 91103 36226 91489 36245
rect 95103 36331 95489 36350
rect 95103 36308 95169 36331
rect 95255 36308 95337 36331
rect 95423 36308 95489 36331
rect 95103 36268 95112 36308
rect 95152 36268 95169 36308
rect 95255 36268 95276 36308
rect 95316 36268 95337 36308
rect 95423 36268 95440 36308
rect 95480 36268 95489 36308
rect 95103 36245 95169 36268
rect 95255 36245 95337 36268
rect 95423 36245 95489 36268
rect 95103 36226 95489 36245
rect 99103 36331 99489 36350
rect 99103 36308 99169 36331
rect 99255 36308 99337 36331
rect 99423 36308 99489 36331
rect 99103 36268 99112 36308
rect 99152 36268 99169 36308
rect 99255 36268 99276 36308
rect 99316 36268 99337 36308
rect 99423 36268 99440 36308
rect 99480 36268 99489 36308
rect 99103 36245 99169 36268
rect 99255 36245 99337 36268
rect 99423 36245 99489 36268
rect 99103 36226 99489 36245
rect 4343 35575 4729 35594
rect 4343 35552 4409 35575
rect 4495 35552 4577 35575
rect 4663 35552 4729 35575
rect 4343 35512 4352 35552
rect 4392 35512 4409 35552
rect 4495 35512 4516 35552
rect 4556 35512 4577 35552
rect 4663 35512 4680 35552
rect 4720 35512 4729 35552
rect 4343 35489 4409 35512
rect 4495 35489 4577 35512
rect 4663 35489 4729 35512
rect 4343 35470 4729 35489
rect 8343 35575 8729 35594
rect 8343 35552 8409 35575
rect 8495 35552 8577 35575
rect 8663 35552 8729 35575
rect 8343 35512 8352 35552
rect 8392 35512 8409 35552
rect 8495 35512 8516 35552
rect 8556 35512 8577 35552
rect 8663 35512 8680 35552
rect 8720 35512 8729 35552
rect 8343 35489 8409 35512
rect 8495 35489 8577 35512
rect 8663 35489 8729 35512
rect 8343 35470 8729 35489
rect 12343 35575 12729 35594
rect 12343 35552 12409 35575
rect 12495 35552 12577 35575
rect 12663 35552 12729 35575
rect 12343 35512 12352 35552
rect 12392 35512 12409 35552
rect 12495 35512 12516 35552
rect 12556 35512 12577 35552
rect 12663 35512 12680 35552
rect 12720 35512 12729 35552
rect 12343 35489 12409 35512
rect 12495 35489 12577 35512
rect 12663 35489 12729 35512
rect 12343 35470 12729 35489
rect 16343 35575 16729 35594
rect 16343 35552 16409 35575
rect 16495 35552 16577 35575
rect 16663 35552 16729 35575
rect 16343 35512 16352 35552
rect 16392 35512 16409 35552
rect 16495 35512 16516 35552
rect 16556 35512 16577 35552
rect 16663 35512 16680 35552
rect 16720 35512 16729 35552
rect 16343 35489 16409 35512
rect 16495 35489 16577 35512
rect 16663 35489 16729 35512
rect 16343 35470 16729 35489
rect 20343 35575 20729 35594
rect 20343 35552 20409 35575
rect 20495 35552 20577 35575
rect 20663 35552 20729 35575
rect 20343 35512 20352 35552
rect 20392 35512 20409 35552
rect 20495 35512 20516 35552
rect 20556 35512 20577 35552
rect 20663 35512 20680 35552
rect 20720 35512 20729 35552
rect 20343 35489 20409 35512
rect 20495 35489 20577 35512
rect 20663 35489 20729 35512
rect 20343 35470 20729 35489
rect 24343 35575 24729 35594
rect 24343 35552 24409 35575
rect 24495 35552 24577 35575
rect 24663 35552 24729 35575
rect 24343 35512 24352 35552
rect 24392 35512 24409 35552
rect 24495 35512 24516 35552
rect 24556 35512 24577 35552
rect 24663 35512 24680 35552
rect 24720 35512 24729 35552
rect 24343 35489 24409 35512
rect 24495 35489 24577 35512
rect 24663 35489 24729 35512
rect 24343 35470 24729 35489
rect 28343 35575 28729 35594
rect 28343 35552 28409 35575
rect 28495 35552 28577 35575
rect 28663 35552 28729 35575
rect 28343 35512 28352 35552
rect 28392 35512 28409 35552
rect 28495 35512 28516 35552
rect 28556 35512 28577 35552
rect 28663 35512 28680 35552
rect 28720 35512 28729 35552
rect 28343 35489 28409 35512
rect 28495 35489 28577 35512
rect 28663 35489 28729 35512
rect 28343 35470 28729 35489
rect 32343 35575 32729 35594
rect 32343 35552 32409 35575
rect 32495 35552 32577 35575
rect 32663 35552 32729 35575
rect 32343 35512 32352 35552
rect 32392 35512 32409 35552
rect 32495 35512 32516 35552
rect 32556 35512 32577 35552
rect 32663 35512 32680 35552
rect 32720 35512 32729 35552
rect 32343 35489 32409 35512
rect 32495 35489 32577 35512
rect 32663 35489 32729 35512
rect 32343 35470 32729 35489
rect 36343 35575 36729 35594
rect 36343 35552 36409 35575
rect 36495 35552 36577 35575
rect 36663 35552 36729 35575
rect 36343 35512 36352 35552
rect 36392 35512 36409 35552
rect 36495 35512 36516 35552
rect 36556 35512 36577 35552
rect 36663 35512 36680 35552
rect 36720 35512 36729 35552
rect 36343 35489 36409 35512
rect 36495 35489 36577 35512
rect 36663 35489 36729 35512
rect 36343 35470 36729 35489
rect 40343 35575 40729 35594
rect 40343 35552 40409 35575
rect 40495 35552 40577 35575
rect 40663 35552 40729 35575
rect 40343 35512 40352 35552
rect 40392 35512 40409 35552
rect 40495 35512 40516 35552
rect 40556 35512 40577 35552
rect 40663 35512 40680 35552
rect 40720 35512 40729 35552
rect 40343 35489 40409 35512
rect 40495 35489 40577 35512
rect 40663 35489 40729 35512
rect 40343 35470 40729 35489
rect 44343 35575 44729 35594
rect 44343 35552 44409 35575
rect 44495 35552 44577 35575
rect 44663 35552 44729 35575
rect 44343 35512 44352 35552
rect 44392 35512 44409 35552
rect 44495 35512 44516 35552
rect 44556 35512 44577 35552
rect 44663 35512 44680 35552
rect 44720 35512 44729 35552
rect 44343 35489 44409 35512
rect 44495 35489 44577 35512
rect 44663 35489 44729 35512
rect 44343 35470 44729 35489
rect 48343 35575 48729 35594
rect 48343 35552 48409 35575
rect 48495 35552 48577 35575
rect 48663 35552 48729 35575
rect 48343 35512 48352 35552
rect 48392 35512 48409 35552
rect 48495 35512 48516 35552
rect 48556 35512 48577 35552
rect 48663 35512 48680 35552
rect 48720 35512 48729 35552
rect 48343 35489 48409 35512
rect 48495 35489 48577 35512
rect 48663 35489 48729 35512
rect 48343 35470 48729 35489
rect 52343 35575 52729 35594
rect 52343 35552 52409 35575
rect 52495 35552 52577 35575
rect 52663 35552 52729 35575
rect 52343 35512 52352 35552
rect 52392 35512 52409 35552
rect 52495 35512 52516 35552
rect 52556 35512 52577 35552
rect 52663 35512 52680 35552
rect 52720 35512 52729 35552
rect 52343 35489 52409 35512
rect 52495 35489 52577 35512
rect 52663 35489 52729 35512
rect 52343 35470 52729 35489
rect 56343 35575 56729 35594
rect 56343 35552 56409 35575
rect 56495 35552 56577 35575
rect 56663 35552 56729 35575
rect 56343 35512 56352 35552
rect 56392 35512 56409 35552
rect 56495 35512 56516 35552
rect 56556 35512 56577 35552
rect 56663 35512 56680 35552
rect 56720 35512 56729 35552
rect 56343 35489 56409 35512
rect 56495 35489 56577 35512
rect 56663 35489 56729 35512
rect 56343 35470 56729 35489
rect 60343 35575 60729 35594
rect 60343 35552 60409 35575
rect 60495 35552 60577 35575
rect 60663 35552 60729 35575
rect 60343 35512 60352 35552
rect 60392 35512 60409 35552
rect 60495 35512 60516 35552
rect 60556 35512 60577 35552
rect 60663 35512 60680 35552
rect 60720 35512 60729 35552
rect 60343 35489 60409 35512
rect 60495 35489 60577 35512
rect 60663 35489 60729 35512
rect 60343 35470 60729 35489
rect 64343 35575 64729 35594
rect 64343 35552 64409 35575
rect 64495 35552 64577 35575
rect 64663 35552 64729 35575
rect 64343 35512 64352 35552
rect 64392 35512 64409 35552
rect 64495 35512 64516 35552
rect 64556 35512 64577 35552
rect 64663 35512 64680 35552
rect 64720 35512 64729 35552
rect 64343 35489 64409 35512
rect 64495 35489 64577 35512
rect 64663 35489 64729 35512
rect 64343 35470 64729 35489
rect 68343 35575 68729 35594
rect 68343 35552 68409 35575
rect 68495 35552 68577 35575
rect 68663 35552 68729 35575
rect 68343 35512 68352 35552
rect 68392 35512 68409 35552
rect 68495 35512 68516 35552
rect 68556 35512 68577 35552
rect 68663 35512 68680 35552
rect 68720 35512 68729 35552
rect 68343 35489 68409 35512
rect 68495 35489 68577 35512
rect 68663 35489 68729 35512
rect 68343 35470 68729 35489
rect 72343 35575 72729 35594
rect 72343 35552 72409 35575
rect 72495 35552 72577 35575
rect 72663 35552 72729 35575
rect 72343 35512 72352 35552
rect 72392 35512 72409 35552
rect 72495 35512 72516 35552
rect 72556 35512 72577 35552
rect 72663 35512 72680 35552
rect 72720 35512 72729 35552
rect 72343 35489 72409 35512
rect 72495 35489 72577 35512
rect 72663 35489 72729 35512
rect 72343 35470 72729 35489
rect 76343 35575 76729 35594
rect 76343 35552 76409 35575
rect 76495 35552 76577 35575
rect 76663 35552 76729 35575
rect 76343 35512 76352 35552
rect 76392 35512 76409 35552
rect 76495 35512 76516 35552
rect 76556 35512 76577 35552
rect 76663 35512 76680 35552
rect 76720 35512 76729 35552
rect 76343 35489 76409 35512
rect 76495 35489 76577 35512
rect 76663 35489 76729 35512
rect 76343 35470 76729 35489
rect 80343 35575 80729 35594
rect 80343 35552 80409 35575
rect 80495 35552 80577 35575
rect 80663 35552 80729 35575
rect 80343 35512 80352 35552
rect 80392 35512 80409 35552
rect 80495 35512 80516 35552
rect 80556 35512 80577 35552
rect 80663 35512 80680 35552
rect 80720 35512 80729 35552
rect 80343 35489 80409 35512
rect 80495 35489 80577 35512
rect 80663 35489 80729 35512
rect 80343 35470 80729 35489
rect 84343 35575 84729 35594
rect 84343 35552 84409 35575
rect 84495 35552 84577 35575
rect 84663 35552 84729 35575
rect 84343 35512 84352 35552
rect 84392 35512 84409 35552
rect 84495 35512 84516 35552
rect 84556 35512 84577 35552
rect 84663 35512 84680 35552
rect 84720 35512 84729 35552
rect 84343 35489 84409 35512
rect 84495 35489 84577 35512
rect 84663 35489 84729 35512
rect 84343 35470 84729 35489
rect 88343 35575 88729 35594
rect 88343 35552 88409 35575
rect 88495 35552 88577 35575
rect 88663 35552 88729 35575
rect 88343 35512 88352 35552
rect 88392 35512 88409 35552
rect 88495 35512 88516 35552
rect 88556 35512 88577 35552
rect 88663 35512 88680 35552
rect 88720 35512 88729 35552
rect 88343 35489 88409 35512
rect 88495 35489 88577 35512
rect 88663 35489 88729 35512
rect 88343 35470 88729 35489
rect 92343 35575 92729 35594
rect 92343 35552 92409 35575
rect 92495 35552 92577 35575
rect 92663 35552 92729 35575
rect 92343 35512 92352 35552
rect 92392 35512 92409 35552
rect 92495 35512 92516 35552
rect 92556 35512 92577 35552
rect 92663 35512 92680 35552
rect 92720 35512 92729 35552
rect 92343 35489 92409 35512
rect 92495 35489 92577 35512
rect 92663 35489 92729 35512
rect 92343 35470 92729 35489
rect 96343 35575 96729 35594
rect 96343 35552 96409 35575
rect 96495 35552 96577 35575
rect 96663 35552 96729 35575
rect 96343 35512 96352 35552
rect 96392 35512 96409 35552
rect 96495 35512 96516 35552
rect 96556 35512 96577 35552
rect 96663 35512 96680 35552
rect 96720 35512 96729 35552
rect 96343 35489 96409 35512
rect 96495 35489 96577 35512
rect 96663 35489 96729 35512
rect 96343 35470 96729 35489
rect 3103 34819 3489 34838
rect 3103 34796 3169 34819
rect 3255 34796 3337 34819
rect 3423 34796 3489 34819
rect 3103 34756 3112 34796
rect 3152 34756 3169 34796
rect 3255 34756 3276 34796
rect 3316 34756 3337 34796
rect 3423 34756 3440 34796
rect 3480 34756 3489 34796
rect 3103 34733 3169 34756
rect 3255 34733 3337 34756
rect 3423 34733 3489 34756
rect 3103 34714 3489 34733
rect 7103 34819 7489 34838
rect 7103 34796 7169 34819
rect 7255 34796 7337 34819
rect 7423 34796 7489 34819
rect 7103 34756 7112 34796
rect 7152 34756 7169 34796
rect 7255 34756 7276 34796
rect 7316 34756 7337 34796
rect 7423 34756 7440 34796
rect 7480 34756 7489 34796
rect 7103 34733 7169 34756
rect 7255 34733 7337 34756
rect 7423 34733 7489 34756
rect 7103 34714 7489 34733
rect 11103 34819 11489 34838
rect 11103 34796 11169 34819
rect 11255 34796 11337 34819
rect 11423 34796 11489 34819
rect 11103 34756 11112 34796
rect 11152 34756 11169 34796
rect 11255 34756 11276 34796
rect 11316 34756 11337 34796
rect 11423 34756 11440 34796
rect 11480 34756 11489 34796
rect 11103 34733 11169 34756
rect 11255 34733 11337 34756
rect 11423 34733 11489 34756
rect 11103 34714 11489 34733
rect 15103 34819 15489 34838
rect 15103 34796 15169 34819
rect 15255 34796 15337 34819
rect 15423 34796 15489 34819
rect 15103 34756 15112 34796
rect 15152 34756 15169 34796
rect 15255 34756 15276 34796
rect 15316 34756 15337 34796
rect 15423 34756 15440 34796
rect 15480 34756 15489 34796
rect 15103 34733 15169 34756
rect 15255 34733 15337 34756
rect 15423 34733 15489 34756
rect 15103 34714 15489 34733
rect 19103 34819 19489 34838
rect 19103 34796 19169 34819
rect 19255 34796 19337 34819
rect 19423 34796 19489 34819
rect 19103 34756 19112 34796
rect 19152 34756 19169 34796
rect 19255 34756 19276 34796
rect 19316 34756 19337 34796
rect 19423 34756 19440 34796
rect 19480 34756 19489 34796
rect 19103 34733 19169 34756
rect 19255 34733 19337 34756
rect 19423 34733 19489 34756
rect 19103 34714 19489 34733
rect 23103 34819 23489 34838
rect 23103 34796 23169 34819
rect 23255 34796 23337 34819
rect 23423 34796 23489 34819
rect 23103 34756 23112 34796
rect 23152 34756 23169 34796
rect 23255 34756 23276 34796
rect 23316 34756 23337 34796
rect 23423 34756 23440 34796
rect 23480 34756 23489 34796
rect 23103 34733 23169 34756
rect 23255 34733 23337 34756
rect 23423 34733 23489 34756
rect 23103 34714 23489 34733
rect 27103 34819 27489 34838
rect 27103 34796 27169 34819
rect 27255 34796 27337 34819
rect 27423 34796 27489 34819
rect 27103 34756 27112 34796
rect 27152 34756 27169 34796
rect 27255 34756 27276 34796
rect 27316 34756 27337 34796
rect 27423 34756 27440 34796
rect 27480 34756 27489 34796
rect 27103 34733 27169 34756
rect 27255 34733 27337 34756
rect 27423 34733 27489 34756
rect 27103 34714 27489 34733
rect 31103 34819 31489 34838
rect 31103 34796 31169 34819
rect 31255 34796 31337 34819
rect 31423 34796 31489 34819
rect 31103 34756 31112 34796
rect 31152 34756 31169 34796
rect 31255 34756 31276 34796
rect 31316 34756 31337 34796
rect 31423 34756 31440 34796
rect 31480 34756 31489 34796
rect 31103 34733 31169 34756
rect 31255 34733 31337 34756
rect 31423 34733 31489 34756
rect 31103 34714 31489 34733
rect 35103 34819 35489 34838
rect 35103 34796 35169 34819
rect 35255 34796 35337 34819
rect 35423 34796 35489 34819
rect 35103 34756 35112 34796
rect 35152 34756 35169 34796
rect 35255 34756 35276 34796
rect 35316 34756 35337 34796
rect 35423 34756 35440 34796
rect 35480 34756 35489 34796
rect 35103 34733 35169 34756
rect 35255 34733 35337 34756
rect 35423 34733 35489 34756
rect 35103 34714 35489 34733
rect 39103 34819 39489 34838
rect 39103 34796 39169 34819
rect 39255 34796 39337 34819
rect 39423 34796 39489 34819
rect 39103 34756 39112 34796
rect 39152 34756 39169 34796
rect 39255 34756 39276 34796
rect 39316 34756 39337 34796
rect 39423 34756 39440 34796
rect 39480 34756 39489 34796
rect 39103 34733 39169 34756
rect 39255 34733 39337 34756
rect 39423 34733 39489 34756
rect 39103 34714 39489 34733
rect 43103 34819 43489 34838
rect 43103 34796 43169 34819
rect 43255 34796 43337 34819
rect 43423 34796 43489 34819
rect 43103 34756 43112 34796
rect 43152 34756 43169 34796
rect 43255 34756 43276 34796
rect 43316 34756 43337 34796
rect 43423 34756 43440 34796
rect 43480 34756 43489 34796
rect 43103 34733 43169 34756
rect 43255 34733 43337 34756
rect 43423 34733 43489 34756
rect 43103 34714 43489 34733
rect 47103 34819 47489 34838
rect 47103 34796 47169 34819
rect 47255 34796 47337 34819
rect 47423 34796 47489 34819
rect 47103 34756 47112 34796
rect 47152 34756 47169 34796
rect 47255 34756 47276 34796
rect 47316 34756 47337 34796
rect 47423 34756 47440 34796
rect 47480 34756 47489 34796
rect 47103 34733 47169 34756
rect 47255 34733 47337 34756
rect 47423 34733 47489 34756
rect 47103 34714 47489 34733
rect 51103 34819 51489 34838
rect 51103 34796 51169 34819
rect 51255 34796 51337 34819
rect 51423 34796 51489 34819
rect 51103 34756 51112 34796
rect 51152 34756 51169 34796
rect 51255 34756 51276 34796
rect 51316 34756 51337 34796
rect 51423 34756 51440 34796
rect 51480 34756 51489 34796
rect 51103 34733 51169 34756
rect 51255 34733 51337 34756
rect 51423 34733 51489 34756
rect 51103 34714 51489 34733
rect 55103 34819 55489 34838
rect 55103 34796 55169 34819
rect 55255 34796 55337 34819
rect 55423 34796 55489 34819
rect 55103 34756 55112 34796
rect 55152 34756 55169 34796
rect 55255 34756 55276 34796
rect 55316 34756 55337 34796
rect 55423 34756 55440 34796
rect 55480 34756 55489 34796
rect 55103 34733 55169 34756
rect 55255 34733 55337 34756
rect 55423 34733 55489 34756
rect 55103 34714 55489 34733
rect 59103 34819 59489 34838
rect 59103 34796 59169 34819
rect 59255 34796 59337 34819
rect 59423 34796 59489 34819
rect 59103 34756 59112 34796
rect 59152 34756 59169 34796
rect 59255 34756 59276 34796
rect 59316 34756 59337 34796
rect 59423 34756 59440 34796
rect 59480 34756 59489 34796
rect 59103 34733 59169 34756
rect 59255 34733 59337 34756
rect 59423 34733 59489 34756
rect 59103 34714 59489 34733
rect 63103 34819 63489 34838
rect 63103 34796 63169 34819
rect 63255 34796 63337 34819
rect 63423 34796 63489 34819
rect 63103 34756 63112 34796
rect 63152 34756 63169 34796
rect 63255 34756 63276 34796
rect 63316 34756 63337 34796
rect 63423 34756 63440 34796
rect 63480 34756 63489 34796
rect 63103 34733 63169 34756
rect 63255 34733 63337 34756
rect 63423 34733 63489 34756
rect 63103 34714 63489 34733
rect 67103 34819 67489 34838
rect 67103 34796 67169 34819
rect 67255 34796 67337 34819
rect 67423 34796 67489 34819
rect 67103 34756 67112 34796
rect 67152 34756 67169 34796
rect 67255 34756 67276 34796
rect 67316 34756 67337 34796
rect 67423 34756 67440 34796
rect 67480 34756 67489 34796
rect 67103 34733 67169 34756
rect 67255 34733 67337 34756
rect 67423 34733 67489 34756
rect 67103 34714 67489 34733
rect 71103 34819 71489 34838
rect 71103 34796 71169 34819
rect 71255 34796 71337 34819
rect 71423 34796 71489 34819
rect 71103 34756 71112 34796
rect 71152 34756 71169 34796
rect 71255 34756 71276 34796
rect 71316 34756 71337 34796
rect 71423 34756 71440 34796
rect 71480 34756 71489 34796
rect 71103 34733 71169 34756
rect 71255 34733 71337 34756
rect 71423 34733 71489 34756
rect 71103 34714 71489 34733
rect 75103 34819 75489 34838
rect 75103 34796 75169 34819
rect 75255 34796 75337 34819
rect 75423 34796 75489 34819
rect 75103 34756 75112 34796
rect 75152 34756 75169 34796
rect 75255 34756 75276 34796
rect 75316 34756 75337 34796
rect 75423 34756 75440 34796
rect 75480 34756 75489 34796
rect 75103 34733 75169 34756
rect 75255 34733 75337 34756
rect 75423 34733 75489 34756
rect 75103 34714 75489 34733
rect 79103 34819 79489 34838
rect 79103 34796 79169 34819
rect 79255 34796 79337 34819
rect 79423 34796 79489 34819
rect 79103 34756 79112 34796
rect 79152 34756 79169 34796
rect 79255 34756 79276 34796
rect 79316 34756 79337 34796
rect 79423 34756 79440 34796
rect 79480 34756 79489 34796
rect 79103 34733 79169 34756
rect 79255 34733 79337 34756
rect 79423 34733 79489 34756
rect 79103 34714 79489 34733
rect 83103 34819 83489 34838
rect 83103 34796 83169 34819
rect 83255 34796 83337 34819
rect 83423 34796 83489 34819
rect 83103 34756 83112 34796
rect 83152 34756 83169 34796
rect 83255 34756 83276 34796
rect 83316 34756 83337 34796
rect 83423 34756 83440 34796
rect 83480 34756 83489 34796
rect 83103 34733 83169 34756
rect 83255 34733 83337 34756
rect 83423 34733 83489 34756
rect 83103 34714 83489 34733
rect 87103 34819 87489 34838
rect 87103 34796 87169 34819
rect 87255 34796 87337 34819
rect 87423 34796 87489 34819
rect 87103 34756 87112 34796
rect 87152 34756 87169 34796
rect 87255 34756 87276 34796
rect 87316 34756 87337 34796
rect 87423 34756 87440 34796
rect 87480 34756 87489 34796
rect 87103 34733 87169 34756
rect 87255 34733 87337 34756
rect 87423 34733 87489 34756
rect 87103 34714 87489 34733
rect 91103 34819 91489 34838
rect 91103 34796 91169 34819
rect 91255 34796 91337 34819
rect 91423 34796 91489 34819
rect 91103 34756 91112 34796
rect 91152 34756 91169 34796
rect 91255 34756 91276 34796
rect 91316 34756 91337 34796
rect 91423 34756 91440 34796
rect 91480 34756 91489 34796
rect 91103 34733 91169 34756
rect 91255 34733 91337 34756
rect 91423 34733 91489 34756
rect 91103 34714 91489 34733
rect 95103 34819 95489 34838
rect 95103 34796 95169 34819
rect 95255 34796 95337 34819
rect 95423 34796 95489 34819
rect 95103 34756 95112 34796
rect 95152 34756 95169 34796
rect 95255 34756 95276 34796
rect 95316 34756 95337 34796
rect 95423 34756 95440 34796
rect 95480 34756 95489 34796
rect 95103 34733 95169 34756
rect 95255 34733 95337 34756
rect 95423 34733 95489 34756
rect 95103 34714 95489 34733
rect 99103 34819 99489 34838
rect 99103 34796 99169 34819
rect 99255 34796 99337 34819
rect 99423 34796 99489 34819
rect 99103 34756 99112 34796
rect 99152 34756 99169 34796
rect 99255 34756 99276 34796
rect 99316 34756 99337 34796
rect 99423 34756 99440 34796
rect 99480 34756 99489 34796
rect 99103 34733 99169 34756
rect 99255 34733 99337 34756
rect 99423 34733 99489 34756
rect 99103 34714 99489 34733
rect 4343 34063 4729 34082
rect 4343 34040 4409 34063
rect 4495 34040 4577 34063
rect 4663 34040 4729 34063
rect 4343 34000 4352 34040
rect 4392 34000 4409 34040
rect 4495 34000 4516 34040
rect 4556 34000 4577 34040
rect 4663 34000 4680 34040
rect 4720 34000 4729 34040
rect 4343 33977 4409 34000
rect 4495 33977 4577 34000
rect 4663 33977 4729 34000
rect 4343 33958 4729 33977
rect 8343 34063 8729 34082
rect 8343 34040 8409 34063
rect 8495 34040 8577 34063
rect 8663 34040 8729 34063
rect 8343 34000 8352 34040
rect 8392 34000 8409 34040
rect 8495 34000 8516 34040
rect 8556 34000 8577 34040
rect 8663 34000 8680 34040
rect 8720 34000 8729 34040
rect 8343 33977 8409 34000
rect 8495 33977 8577 34000
rect 8663 33977 8729 34000
rect 8343 33958 8729 33977
rect 12343 34063 12729 34082
rect 12343 34040 12409 34063
rect 12495 34040 12577 34063
rect 12663 34040 12729 34063
rect 12343 34000 12352 34040
rect 12392 34000 12409 34040
rect 12495 34000 12516 34040
rect 12556 34000 12577 34040
rect 12663 34000 12680 34040
rect 12720 34000 12729 34040
rect 12343 33977 12409 34000
rect 12495 33977 12577 34000
rect 12663 33977 12729 34000
rect 12343 33958 12729 33977
rect 16343 34063 16729 34082
rect 16343 34040 16409 34063
rect 16495 34040 16577 34063
rect 16663 34040 16729 34063
rect 16343 34000 16352 34040
rect 16392 34000 16409 34040
rect 16495 34000 16516 34040
rect 16556 34000 16577 34040
rect 16663 34000 16680 34040
rect 16720 34000 16729 34040
rect 16343 33977 16409 34000
rect 16495 33977 16577 34000
rect 16663 33977 16729 34000
rect 16343 33958 16729 33977
rect 20343 34063 20729 34082
rect 20343 34040 20409 34063
rect 20495 34040 20577 34063
rect 20663 34040 20729 34063
rect 20343 34000 20352 34040
rect 20392 34000 20409 34040
rect 20495 34000 20516 34040
rect 20556 34000 20577 34040
rect 20663 34000 20680 34040
rect 20720 34000 20729 34040
rect 20343 33977 20409 34000
rect 20495 33977 20577 34000
rect 20663 33977 20729 34000
rect 20343 33958 20729 33977
rect 24343 34063 24729 34082
rect 24343 34040 24409 34063
rect 24495 34040 24577 34063
rect 24663 34040 24729 34063
rect 24343 34000 24352 34040
rect 24392 34000 24409 34040
rect 24495 34000 24516 34040
rect 24556 34000 24577 34040
rect 24663 34000 24680 34040
rect 24720 34000 24729 34040
rect 24343 33977 24409 34000
rect 24495 33977 24577 34000
rect 24663 33977 24729 34000
rect 24343 33958 24729 33977
rect 28343 34063 28729 34082
rect 28343 34040 28409 34063
rect 28495 34040 28577 34063
rect 28663 34040 28729 34063
rect 28343 34000 28352 34040
rect 28392 34000 28409 34040
rect 28495 34000 28516 34040
rect 28556 34000 28577 34040
rect 28663 34000 28680 34040
rect 28720 34000 28729 34040
rect 28343 33977 28409 34000
rect 28495 33977 28577 34000
rect 28663 33977 28729 34000
rect 28343 33958 28729 33977
rect 32343 34063 32729 34082
rect 32343 34040 32409 34063
rect 32495 34040 32577 34063
rect 32663 34040 32729 34063
rect 32343 34000 32352 34040
rect 32392 34000 32409 34040
rect 32495 34000 32516 34040
rect 32556 34000 32577 34040
rect 32663 34000 32680 34040
rect 32720 34000 32729 34040
rect 32343 33977 32409 34000
rect 32495 33977 32577 34000
rect 32663 33977 32729 34000
rect 32343 33958 32729 33977
rect 36343 34063 36729 34082
rect 36343 34040 36409 34063
rect 36495 34040 36577 34063
rect 36663 34040 36729 34063
rect 36343 34000 36352 34040
rect 36392 34000 36409 34040
rect 36495 34000 36516 34040
rect 36556 34000 36577 34040
rect 36663 34000 36680 34040
rect 36720 34000 36729 34040
rect 36343 33977 36409 34000
rect 36495 33977 36577 34000
rect 36663 33977 36729 34000
rect 36343 33958 36729 33977
rect 40343 34063 40729 34082
rect 40343 34040 40409 34063
rect 40495 34040 40577 34063
rect 40663 34040 40729 34063
rect 40343 34000 40352 34040
rect 40392 34000 40409 34040
rect 40495 34000 40516 34040
rect 40556 34000 40577 34040
rect 40663 34000 40680 34040
rect 40720 34000 40729 34040
rect 40343 33977 40409 34000
rect 40495 33977 40577 34000
rect 40663 33977 40729 34000
rect 40343 33958 40729 33977
rect 44343 34063 44729 34082
rect 44343 34040 44409 34063
rect 44495 34040 44577 34063
rect 44663 34040 44729 34063
rect 44343 34000 44352 34040
rect 44392 34000 44409 34040
rect 44495 34000 44516 34040
rect 44556 34000 44577 34040
rect 44663 34000 44680 34040
rect 44720 34000 44729 34040
rect 44343 33977 44409 34000
rect 44495 33977 44577 34000
rect 44663 33977 44729 34000
rect 44343 33958 44729 33977
rect 48343 34063 48729 34082
rect 48343 34040 48409 34063
rect 48495 34040 48577 34063
rect 48663 34040 48729 34063
rect 48343 34000 48352 34040
rect 48392 34000 48409 34040
rect 48495 34000 48516 34040
rect 48556 34000 48577 34040
rect 48663 34000 48680 34040
rect 48720 34000 48729 34040
rect 48343 33977 48409 34000
rect 48495 33977 48577 34000
rect 48663 33977 48729 34000
rect 48343 33958 48729 33977
rect 52343 34063 52729 34082
rect 52343 34040 52409 34063
rect 52495 34040 52577 34063
rect 52663 34040 52729 34063
rect 52343 34000 52352 34040
rect 52392 34000 52409 34040
rect 52495 34000 52516 34040
rect 52556 34000 52577 34040
rect 52663 34000 52680 34040
rect 52720 34000 52729 34040
rect 52343 33977 52409 34000
rect 52495 33977 52577 34000
rect 52663 33977 52729 34000
rect 52343 33958 52729 33977
rect 56343 34063 56729 34082
rect 56343 34040 56409 34063
rect 56495 34040 56577 34063
rect 56663 34040 56729 34063
rect 56343 34000 56352 34040
rect 56392 34000 56409 34040
rect 56495 34000 56516 34040
rect 56556 34000 56577 34040
rect 56663 34000 56680 34040
rect 56720 34000 56729 34040
rect 56343 33977 56409 34000
rect 56495 33977 56577 34000
rect 56663 33977 56729 34000
rect 56343 33958 56729 33977
rect 60343 34063 60729 34082
rect 60343 34040 60409 34063
rect 60495 34040 60577 34063
rect 60663 34040 60729 34063
rect 60343 34000 60352 34040
rect 60392 34000 60409 34040
rect 60495 34000 60516 34040
rect 60556 34000 60577 34040
rect 60663 34000 60680 34040
rect 60720 34000 60729 34040
rect 60343 33977 60409 34000
rect 60495 33977 60577 34000
rect 60663 33977 60729 34000
rect 60343 33958 60729 33977
rect 64343 34063 64729 34082
rect 64343 34040 64409 34063
rect 64495 34040 64577 34063
rect 64663 34040 64729 34063
rect 64343 34000 64352 34040
rect 64392 34000 64409 34040
rect 64495 34000 64516 34040
rect 64556 34000 64577 34040
rect 64663 34000 64680 34040
rect 64720 34000 64729 34040
rect 64343 33977 64409 34000
rect 64495 33977 64577 34000
rect 64663 33977 64729 34000
rect 64343 33958 64729 33977
rect 68343 34063 68729 34082
rect 68343 34040 68409 34063
rect 68495 34040 68577 34063
rect 68663 34040 68729 34063
rect 68343 34000 68352 34040
rect 68392 34000 68409 34040
rect 68495 34000 68516 34040
rect 68556 34000 68577 34040
rect 68663 34000 68680 34040
rect 68720 34000 68729 34040
rect 68343 33977 68409 34000
rect 68495 33977 68577 34000
rect 68663 33977 68729 34000
rect 68343 33958 68729 33977
rect 86450 33475 86574 33494
rect 86450 33389 86469 33475
rect 86555 33452 86574 33475
rect 86555 33412 87052 33452
rect 87092 33412 87101 33452
rect 86555 33389 86574 33412
rect 86450 33370 86574 33389
rect 3103 33307 3489 33326
rect 3103 33284 3169 33307
rect 3255 33284 3337 33307
rect 3423 33284 3489 33307
rect 3103 33244 3112 33284
rect 3152 33244 3169 33284
rect 3255 33244 3276 33284
rect 3316 33244 3337 33284
rect 3423 33244 3440 33284
rect 3480 33244 3489 33284
rect 3103 33221 3169 33244
rect 3255 33221 3337 33244
rect 3423 33221 3489 33244
rect 3103 33202 3489 33221
rect 7103 33307 7489 33326
rect 7103 33284 7169 33307
rect 7255 33284 7337 33307
rect 7423 33284 7489 33307
rect 7103 33244 7112 33284
rect 7152 33244 7169 33284
rect 7255 33244 7276 33284
rect 7316 33244 7337 33284
rect 7423 33244 7440 33284
rect 7480 33244 7489 33284
rect 7103 33221 7169 33244
rect 7255 33221 7337 33244
rect 7423 33221 7489 33244
rect 7103 33202 7489 33221
rect 11103 33307 11489 33326
rect 11103 33284 11169 33307
rect 11255 33284 11337 33307
rect 11423 33284 11489 33307
rect 11103 33244 11112 33284
rect 11152 33244 11169 33284
rect 11255 33244 11276 33284
rect 11316 33244 11337 33284
rect 11423 33244 11440 33284
rect 11480 33244 11489 33284
rect 11103 33221 11169 33244
rect 11255 33221 11337 33244
rect 11423 33221 11489 33244
rect 11103 33202 11489 33221
rect 15103 33307 15489 33326
rect 15103 33284 15169 33307
rect 15255 33284 15337 33307
rect 15423 33284 15489 33307
rect 15103 33244 15112 33284
rect 15152 33244 15169 33284
rect 15255 33244 15276 33284
rect 15316 33244 15337 33284
rect 15423 33244 15440 33284
rect 15480 33244 15489 33284
rect 15103 33221 15169 33244
rect 15255 33221 15337 33244
rect 15423 33221 15489 33244
rect 15103 33202 15489 33221
rect 19103 33307 19489 33326
rect 19103 33284 19169 33307
rect 19255 33284 19337 33307
rect 19423 33284 19489 33307
rect 19103 33244 19112 33284
rect 19152 33244 19169 33284
rect 19255 33244 19276 33284
rect 19316 33244 19337 33284
rect 19423 33244 19440 33284
rect 19480 33244 19489 33284
rect 19103 33221 19169 33244
rect 19255 33221 19337 33244
rect 19423 33221 19489 33244
rect 19103 33202 19489 33221
rect 23103 33307 23489 33326
rect 23103 33284 23169 33307
rect 23255 33284 23337 33307
rect 23423 33284 23489 33307
rect 23103 33244 23112 33284
rect 23152 33244 23169 33284
rect 23255 33244 23276 33284
rect 23316 33244 23337 33284
rect 23423 33244 23440 33284
rect 23480 33244 23489 33284
rect 23103 33221 23169 33244
rect 23255 33221 23337 33244
rect 23423 33221 23489 33244
rect 23103 33202 23489 33221
rect 27103 33307 27489 33326
rect 27103 33284 27169 33307
rect 27255 33284 27337 33307
rect 27423 33284 27489 33307
rect 27103 33244 27112 33284
rect 27152 33244 27169 33284
rect 27255 33244 27276 33284
rect 27316 33244 27337 33284
rect 27423 33244 27440 33284
rect 27480 33244 27489 33284
rect 27103 33221 27169 33244
rect 27255 33221 27337 33244
rect 27423 33221 27489 33244
rect 27103 33202 27489 33221
rect 31103 33307 31489 33326
rect 31103 33284 31169 33307
rect 31255 33284 31337 33307
rect 31423 33284 31489 33307
rect 31103 33244 31112 33284
rect 31152 33244 31169 33284
rect 31255 33244 31276 33284
rect 31316 33244 31337 33284
rect 31423 33244 31440 33284
rect 31480 33244 31489 33284
rect 31103 33221 31169 33244
rect 31255 33221 31337 33244
rect 31423 33221 31489 33244
rect 31103 33202 31489 33221
rect 35103 33307 35489 33326
rect 35103 33284 35169 33307
rect 35255 33284 35337 33307
rect 35423 33284 35489 33307
rect 35103 33244 35112 33284
rect 35152 33244 35169 33284
rect 35255 33244 35276 33284
rect 35316 33244 35337 33284
rect 35423 33244 35440 33284
rect 35480 33244 35489 33284
rect 35103 33221 35169 33244
rect 35255 33221 35337 33244
rect 35423 33221 35489 33244
rect 35103 33202 35489 33221
rect 39103 33307 39489 33326
rect 39103 33284 39169 33307
rect 39255 33284 39337 33307
rect 39423 33284 39489 33307
rect 39103 33244 39112 33284
rect 39152 33244 39169 33284
rect 39255 33244 39276 33284
rect 39316 33244 39337 33284
rect 39423 33244 39440 33284
rect 39480 33244 39489 33284
rect 39103 33221 39169 33244
rect 39255 33221 39337 33244
rect 39423 33221 39489 33244
rect 39103 33202 39489 33221
rect 43103 33307 43489 33326
rect 43103 33284 43169 33307
rect 43255 33284 43337 33307
rect 43423 33284 43489 33307
rect 43103 33244 43112 33284
rect 43152 33244 43169 33284
rect 43255 33244 43276 33284
rect 43316 33244 43337 33284
rect 43423 33244 43440 33284
rect 43480 33244 43489 33284
rect 43103 33221 43169 33244
rect 43255 33221 43337 33244
rect 43423 33221 43489 33244
rect 43103 33202 43489 33221
rect 47103 33307 47489 33326
rect 47103 33284 47169 33307
rect 47255 33284 47337 33307
rect 47423 33284 47489 33307
rect 47103 33244 47112 33284
rect 47152 33244 47169 33284
rect 47255 33244 47276 33284
rect 47316 33244 47337 33284
rect 47423 33244 47440 33284
rect 47480 33244 47489 33284
rect 47103 33221 47169 33244
rect 47255 33221 47337 33244
rect 47423 33221 47489 33244
rect 47103 33202 47489 33221
rect 51103 33307 51489 33326
rect 51103 33284 51169 33307
rect 51255 33284 51337 33307
rect 51423 33284 51489 33307
rect 51103 33244 51112 33284
rect 51152 33244 51169 33284
rect 51255 33244 51276 33284
rect 51316 33244 51337 33284
rect 51423 33244 51440 33284
rect 51480 33244 51489 33284
rect 51103 33221 51169 33244
rect 51255 33221 51337 33244
rect 51423 33221 51489 33244
rect 51103 33202 51489 33221
rect 55103 33307 55489 33326
rect 55103 33284 55169 33307
rect 55255 33284 55337 33307
rect 55423 33284 55489 33307
rect 55103 33244 55112 33284
rect 55152 33244 55169 33284
rect 55255 33244 55276 33284
rect 55316 33244 55337 33284
rect 55423 33244 55440 33284
rect 55480 33244 55489 33284
rect 55103 33221 55169 33244
rect 55255 33221 55337 33244
rect 55423 33221 55489 33244
rect 55103 33202 55489 33221
rect 59103 33307 59489 33326
rect 59103 33284 59169 33307
rect 59255 33284 59337 33307
rect 59423 33284 59489 33307
rect 59103 33244 59112 33284
rect 59152 33244 59169 33284
rect 59255 33244 59276 33284
rect 59316 33244 59337 33284
rect 59423 33244 59440 33284
rect 59480 33244 59489 33284
rect 59103 33221 59169 33244
rect 59255 33221 59337 33244
rect 59423 33221 59489 33244
rect 59103 33202 59489 33221
rect 63103 33307 63489 33326
rect 63103 33284 63169 33307
rect 63255 33284 63337 33307
rect 63423 33284 63489 33307
rect 63103 33244 63112 33284
rect 63152 33244 63169 33284
rect 63255 33244 63276 33284
rect 63316 33244 63337 33284
rect 63423 33244 63440 33284
rect 63480 33244 63489 33284
rect 63103 33221 63169 33244
rect 63255 33221 63337 33244
rect 63423 33221 63489 33244
rect 63103 33202 63489 33221
rect 67103 33307 67489 33326
rect 67103 33284 67169 33307
rect 67255 33284 67337 33307
rect 67423 33284 67489 33307
rect 67103 33244 67112 33284
rect 67152 33244 67169 33284
rect 67255 33244 67276 33284
rect 67316 33244 67337 33284
rect 67423 33244 67440 33284
rect 67480 33244 67489 33284
rect 67103 33221 67169 33244
rect 67255 33221 67337 33244
rect 67423 33221 67489 33244
rect 67103 33202 67489 33221
rect 73226 32887 73350 32906
rect 73226 32801 73245 32887
rect 73331 32864 73350 32887
rect 73331 32824 73612 32864
rect 73652 32824 73661 32864
rect 73331 32801 73350 32824
rect 73226 32782 73350 32801
rect 4343 32551 4729 32570
rect 4343 32528 4409 32551
rect 4495 32528 4577 32551
rect 4663 32528 4729 32551
rect 4343 32488 4352 32528
rect 4392 32488 4409 32528
rect 4495 32488 4516 32528
rect 4556 32488 4577 32528
rect 4663 32488 4680 32528
rect 4720 32488 4729 32528
rect 4343 32465 4409 32488
rect 4495 32465 4577 32488
rect 4663 32465 4729 32488
rect 4343 32446 4729 32465
rect 8343 32551 8729 32570
rect 8343 32528 8409 32551
rect 8495 32528 8577 32551
rect 8663 32528 8729 32551
rect 8343 32488 8352 32528
rect 8392 32488 8409 32528
rect 8495 32488 8516 32528
rect 8556 32488 8577 32528
rect 8663 32488 8680 32528
rect 8720 32488 8729 32528
rect 8343 32465 8409 32488
rect 8495 32465 8577 32488
rect 8663 32465 8729 32488
rect 8343 32446 8729 32465
rect 12343 32551 12729 32570
rect 12343 32528 12409 32551
rect 12495 32528 12577 32551
rect 12663 32528 12729 32551
rect 12343 32488 12352 32528
rect 12392 32488 12409 32528
rect 12495 32488 12516 32528
rect 12556 32488 12577 32528
rect 12663 32488 12680 32528
rect 12720 32488 12729 32528
rect 12343 32465 12409 32488
rect 12495 32465 12577 32488
rect 12663 32465 12729 32488
rect 12343 32446 12729 32465
rect 16343 32551 16729 32570
rect 16343 32528 16409 32551
rect 16495 32528 16577 32551
rect 16663 32528 16729 32551
rect 16343 32488 16352 32528
rect 16392 32488 16409 32528
rect 16495 32488 16516 32528
rect 16556 32488 16577 32528
rect 16663 32488 16680 32528
rect 16720 32488 16729 32528
rect 16343 32465 16409 32488
rect 16495 32465 16577 32488
rect 16663 32465 16729 32488
rect 16343 32446 16729 32465
rect 20343 32551 20729 32570
rect 20343 32528 20409 32551
rect 20495 32528 20577 32551
rect 20663 32528 20729 32551
rect 20343 32488 20352 32528
rect 20392 32488 20409 32528
rect 20495 32488 20516 32528
rect 20556 32488 20577 32528
rect 20663 32488 20680 32528
rect 20720 32488 20729 32528
rect 20343 32465 20409 32488
rect 20495 32465 20577 32488
rect 20663 32465 20729 32488
rect 20343 32446 20729 32465
rect 24343 32551 24729 32570
rect 24343 32528 24409 32551
rect 24495 32528 24577 32551
rect 24663 32528 24729 32551
rect 24343 32488 24352 32528
rect 24392 32488 24409 32528
rect 24495 32488 24516 32528
rect 24556 32488 24577 32528
rect 24663 32488 24680 32528
rect 24720 32488 24729 32528
rect 24343 32465 24409 32488
rect 24495 32465 24577 32488
rect 24663 32465 24729 32488
rect 24343 32446 24729 32465
rect 28343 32551 28729 32570
rect 28343 32528 28409 32551
rect 28495 32528 28577 32551
rect 28663 32528 28729 32551
rect 28343 32488 28352 32528
rect 28392 32488 28409 32528
rect 28495 32488 28516 32528
rect 28556 32488 28577 32528
rect 28663 32488 28680 32528
rect 28720 32488 28729 32528
rect 28343 32465 28409 32488
rect 28495 32465 28577 32488
rect 28663 32465 28729 32488
rect 28343 32446 28729 32465
rect 32343 32551 32729 32570
rect 32343 32528 32409 32551
rect 32495 32528 32577 32551
rect 32663 32528 32729 32551
rect 32343 32488 32352 32528
rect 32392 32488 32409 32528
rect 32495 32488 32516 32528
rect 32556 32488 32577 32528
rect 32663 32488 32680 32528
rect 32720 32488 32729 32528
rect 32343 32465 32409 32488
rect 32495 32465 32577 32488
rect 32663 32465 32729 32488
rect 32343 32446 32729 32465
rect 36343 32551 36729 32570
rect 36343 32528 36409 32551
rect 36495 32528 36577 32551
rect 36663 32528 36729 32551
rect 36343 32488 36352 32528
rect 36392 32488 36409 32528
rect 36495 32488 36516 32528
rect 36556 32488 36577 32528
rect 36663 32488 36680 32528
rect 36720 32488 36729 32528
rect 36343 32465 36409 32488
rect 36495 32465 36577 32488
rect 36663 32465 36729 32488
rect 36343 32446 36729 32465
rect 40343 32551 40729 32570
rect 40343 32528 40409 32551
rect 40495 32528 40577 32551
rect 40663 32528 40729 32551
rect 40343 32488 40352 32528
rect 40392 32488 40409 32528
rect 40495 32488 40516 32528
rect 40556 32488 40577 32528
rect 40663 32488 40680 32528
rect 40720 32488 40729 32528
rect 40343 32465 40409 32488
rect 40495 32465 40577 32488
rect 40663 32465 40729 32488
rect 40343 32446 40729 32465
rect 44343 32551 44729 32570
rect 44343 32528 44409 32551
rect 44495 32528 44577 32551
rect 44663 32528 44729 32551
rect 44343 32488 44352 32528
rect 44392 32488 44409 32528
rect 44495 32488 44516 32528
rect 44556 32488 44577 32528
rect 44663 32488 44680 32528
rect 44720 32488 44729 32528
rect 44343 32465 44409 32488
rect 44495 32465 44577 32488
rect 44663 32465 44729 32488
rect 44343 32446 44729 32465
rect 48343 32551 48729 32570
rect 48343 32528 48409 32551
rect 48495 32528 48577 32551
rect 48663 32528 48729 32551
rect 48343 32488 48352 32528
rect 48392 32488 48409 32528
rect 48495 32488 48516 32528
rect 48556 32488 48577 32528
rect 48663 32488 48680 32528
rect 48720 32488 48729 32528
rect 48343 32465 48409 32488
rect 48495 32465 48577 32488
rect 48663 32465 48729 32488
rect 48343 32446 48729 32465
rect 52343 32551 52729 32570
rect 52343 32528 52409 32551
rect 52495 32528 52577 32551
rect 52663 32528 52729 32551
rect 52343 32488 52352 32528
rect 52392 32488 52409 32528
rect 52495 32488 52516 32528
rect 52556 32488 52577 32528
rect 52663 32488 52680 32528
rect 52720 32488 52729 32528
rect 52343 32465 52409 32488
rect 52495 32465 52577 32488
rect 52663 32465 52729 32488
rect 52343 32446 52729 32465
rect 56343 32551 56729 32570
rect 56343 32528 56409 32551
rect 56495 32528 56577 32551
rect 56663 32528 56729 32551
rect 56343 32488 56352 32528
rect 56392 32488 56409 32528
rect 56495 32488 56516 32528
rect 56556 32488 56577 32528
rect 56663 32488 56680 32528
rect 56720 32488 56729 32528
rect 56343 32465 56409 32488
rect 56495 32465 56577 32488
rect 56663 32465 56729 32488
rect 56343 32446 56729 32465
rect 60343 32551 60729 32570
rect 60343 32528 60409 32551
rect 60495 32528 60577 32551
rect 60663 32528 60729 32551
rect 60343 32488 60352 32528
rect 60392 32488 60409 32528
rect 60495 32488 60516 32528
rect 60556 32488 60577 32528
rect 60663 32488 60680 32528
rect 60720 32488 60729 32528
rect 60343 32465 60409 32488
rect 60495 32465 60577 32488
rect 60663 32465 60729 32488
rect 60343 32446 60729 32465
rect 64343 32551 64729 32570
rect 64343 32528 64409 32551
rect 64495 32528 64577 32551
rect 64663 32528 64729 32551
rect 64343 32488 64352 32528
rect 64392 32488 64409 32528
rect 64495 32488 64516 32528
rect 64556 32488 64577 32528
rect 64663 32488 64680 32528
rect 64720 32488 64729 32528
rect 64343 32465 64409 32488
rect 64495 32465 64577 32488
rect 64663 32465 64729 32488
rect 64343 32446 64729 32465
rect 68343 32551 68729 32570
rect 68343 32528 68409 32551
rect 68495 32528 68577 32551
rect 68663 32528 68729 32551
rect 68343 32488 68352 32528
rect 68392 32488 68409 32528
rect 68495 32488 68516 32528
rect 68556 32488 68577 32528
rect 68663 32488 68680 32528
rect 68720 32488 68729 32528
rect 68343 32465 68409 32488
rect 68495 32465 68577 32488
rect 68663 32465 68729 32488
rect 68343 32446 68729 32465
rect 72316 31856 72756 31986
rect 3103 31795 3489 31814
rect 3103 31772 3169 31795
rect 3255 31772 3337 31795
rect 3423 31772 3489 31795
rect 3103 31732 3112 31772
rect 3152 31732 3169 31772
rect 3255 31732 3276 31772
rect 3316 31732 3337 31772
rect 3423 31732 3440 31772
rect 3480 31732 3489 31772
rect 3103 31709 3169 31732
rect 3255 31709 3337 31732
rect 3423 31709 3489 31732
rect 3103 31690 3489 31709
rect 7103 31795 7489 31814
rect 7103 31772 7169 31795
rect 7255 31772 7337 31795
rect 7423 31772 7489 31795
rect 7103 31732 7112 31772
rect 7152 31732 7169 31772
rect 7255 31732 7276 31772
rect 7316 31732 7337 31772
rect 7423 31732 7440 31772
rect 7480 31732 7489 31772
rect 7103 31709 7169 31732
rect 7255 31709 7337 31732
rect 7423 31709 7489 31732
rect 7103 31690 7489 31709
rect 11103 31795 11489 31814
rect 11103 31772 11169 31795
rect 11255 31772 11337 31795
rect 11423 31772 11489 31795
rect 11103 31732 11112 31772
rect 11152 31732 11169 31772
rect 11255 31732 11276 31772
rect 11316 31732 11337 31772
rect 11423 31732 11440 31772
rect 11480 31732 11489 31772
rect 11103 31709 11169 31732
rect 11255 31709 11337 31732
rect 11423 31709 11489 31732
rect 11103 31690 11489 31709
rect 15103 31795 15489 31814
rect 15103 31772 15169 31795
rect 15255 31772 15337 31795
rect 15423 31772 15489 31795
rect 15103 31732 15112 31772
rect 15152 31732 15169 31772
rect 15255 31732 15276 31772
rect 15316 31732 15337 31772
rect 15423 31732 15440 31772
rect 15480 31732 15489 31772
rect 15103 31709 15169 31732
rect 15255 31709 15337 31732
rect 15423 31709 15489 31732
rect 15103 31690 15489 31709
rect 19103 31795 19489 31814
rect 19103 31772 19169 31795
rect 19255 31772 19337 31795
rect 19423 31772 19489 31795
rect 19103 31732 19112 31772
rect 19152 31732 19169 31772
rect 19255 31732 19276 31772
rect 19316 31732 19337 31772
rect 19423 31732 19440 31772
rect 19480 31732 19489 31772
rect 19103 31709 19169 31732
rect 19255 31709 19337 31732
rect 19423 31709 19489 31732
rect 19103 31690 19489 31709
rect 23103 31795 23489 31814
rect 23103 31772 23169 31795
rect 23255 31772 23337 31795
rect 23423 31772 23489 31795
rect 23103 31732 23112 31772
rect 23152 31732 23169 31772
rect 23255 31732 23276 31772
rect 23316 31732 23337 31772
rect 23423 31732 23440 31772
rect 23480 31732 23489 31772
rect 23103 31709 23169 31732
rect 23255 31709 23337 31732
rect 23423 31709 23489 31732
rect 23103 31690 23489 31709
rect 27103 31795 27489 31814
rect 27103 31772 27169 31795
rect 27255 31772 27337 31795
rect 27423 31772 27489 31795
rect 27103 31732 27112 31772
rect 27152 31732 27169 31772
rect 27255 31732 27276 31772
rect 27316 31732 27337 31772
rect 27423 31732 27440 31772
rect 27480 31732 27489 31772
rect 27103 31709 27169 31732
rect 27255 31709 27337 31732
rect 27423 31709 27489 31732
rect 27103 31690 27489 31709
rect 31103 31795 31489 31814
rect 31103 31772 31169 31795
rect 31255 31772 31337 31795
rect 31423 31772 31489 31795
rect 31103 31732 31112 31772
rect 31152 31732 31169 31772
rect 31255 31732 31276 31772
rect 31316 31732 31337 31772
rect 31423 31732 31440 31772
rect 31480 31732 31489 31772
rect 31103 31709 31169 31732
rect 31255 31709 31337 31732
rect 31423 31709 31489 31732
rect 31103 31690 31489 31709
rect 35103 31795 35489 31814
rect 35103 31772 35169 31795
rect 35255 31772 35337 31795
rect 35423 31772 35489 31795
rect 35103 31732 35112 31772
rect 35152 31732 35169 31772
rect 35255 31732 35276 31772
rect 35316 31732 35337 31772
rect 35423 31732 35440 31772
rect 35480 31732 35489 31772
rect 35103 31709 35169 31732
rect 35255 31709 35337 31732
rect 35423 31709 35489 31732
rect 35103 31690 35489 31709
rect 39103 31795 39489 31814
rect 39103 31772 39169 31795
rect 39255 31772 39337 31795
rect 39423 31772 39489 31795
rect 39103 31732 39112 31772
rect 39152 31732 39169 31772
rect 39255 31732 39276 31772
rect 39316 31732 39337 31772
rect 39423 31732 39440 31772
rect 39480 31732 39489 31772
rect 39103 31709 39169 31732
rect 39255 31709 39337 31732
rect 39423 31709 39489 31732
rect 39103 31690 39489 31709
rect 43103 31795 43489 31814
rect 43103 31772 43169 31795
rect 43255 31772 43337 31795
rect 43423 31772 43489 31795
rect 43103 31732 43112 31772
rect 43152 31732 43169 31772
rect 43255 31732 43276 31772
rect 43316 31732 43337 31772
rect 43423 31732 43440 31772
rect 43480 31732 43489 31772
rect 43103 31709 43169 31732
rect 43255 31709 43337 31732
rect 43423 31709 43489 31732
rect 43103 31690 43489 31709
rect 47103 31795 47489 31814
rect 47103 31772 47169 31795
rect 47255 31772 47337 31795
rect 47423 31772 47489 31795
rect 47103 31732 47112 31772
rect 47152 31732 47169 31772
rect 47255 31732 47276 31772
rect 47316 31732 47337 31772
rect 47423 31732 47440 31772
rect 47480 31732 47489 31772
rect 47103 31709 47169 31732
rect 47255 31709 47337 31732
rect 47423 31709 47489 31732
rect 47103 31690 47489 31709
rect 51103 31795 51489 31814
rect 51103 31772 51169 31795
rect 51255 31772 51337 31795
rect 51423 31772 51489 31795
rect 51103 31732 51112 31772
rect 51152 31732 51169 31772
rect 51255 31732 51276 31772
rect 51316 31732 51337 31772
rect 51423 31732 51440 31772
rect 51480 31732 51489 31772
rect 51103 31709 51169 31732
rect 51255 31709 51337 31732
rect 51423 31709 51489 31732
rect 51103 31690 51489 31709
rect 55103 31795 55489 31814
rect 55103 31772 55169 31795
rect 55255 31772 55337 31795
rect 55423 31772 55489 31795
rect 55103 31732 55112 31772
rect 55152 31732 55169 31772
rect 55255 31732 55276 31772
rect 55316 31732 55337 31772
rect 55423 31732 55440 31772
rect 55480 31732 55489 31772
rect 55103 31709 55169 31732
rect 55255 31709 55337 31732
rect 55423 31709 55489 31732
rect 55103 31690 55489 31709
rect 59103 31795 59489 31814
rect 59103 31772 59169 31795
rect 59255 31772 59337 31795
rect 59423 31772 59489 31795
rect 59103 31732 59112 31772
rect 59152 31732 59169 31772
rect 59255 31732 59276 31772
rect 59316 31732 59337 31772
rect 59423 31732 59440 31772
rect 59480 31732 59489 31772
rect 59103 31709 59169 31732
rect 59255 31709 59337 31732
rect 59423 31709 59489 31732
rect 59103 31690 59489 31709
rect 63103 31795 63489 31814
rect 63103 31772 63169 31795
rect 63255 31772 63337 31795
rect 63423 31772 63489 31795
rect 63103 31732 63112 31772
rect 63152 31732 63169 31772
rect 63255 31732 63276 31772
rect 63316 31732 63337 31772
rect 63423 31732 63440 31772
rect 63480 31732 63489 31772
rect 63103 31709 63169 31732
rect 63255 31709 63337 31732
rect 63423 31709 63489 31732
rect 63103 31690 63489 31709
rect 67103 31795 67489 31814
rect 67103 31772 67169 31795
rect 67255 31772 67337 31795
rect 67423 31772 67489 31795
rect 67103 31732 67112 31772
rect 67152 31732 67169 31772
rect 67255 31732 67276 31772
rect 67316 31732 67337 31772
rect 67423 31732 67440 31772
rect 67480 31732 67489 31772
rect 67103 31709 67169 31732
rect 67255 31709 67337 31732
rect 67423 31709 67489 31732
rect 67103 31690 67489 31709
rect 72316 31770 72409 31856
rect 72495 31770 72577 31856
rect 72663 31770 72756 31856
rect 72316 31688 72756 31770
rect 72316 31602 72409 31688
rect 72495 31602 72577 31688
rect 72663 31602 72756 31688
rect 72316 31520 72756 31602
rect 72316 31434 72409 31520
rect 72495 31434 72577 31520
rect 72663 31434 72756 31520
rect 72316 31352 72756 31434
rect 72316 31266 72409 31352
rect 72495 31266 72577 31352
rect 72663 31266 72756 31352
rect 72316 31184 72756 31266
rect 72316 31098 72409 31184
rect 72495 31098 72577 31184
rect 72663 31098 72756 31184
rect 4343 31039 4729 31058
rect 4343 31016 4409 31039
rect 4495 31016 4577 31039
rect 4663 31016 4729 31039
rect 4343 30976 4352 31016
rect 4392 30976 4409 31016
rect 4495 30976 4516 31016
rect 4556 30976 4577 31016
rect 4663 30976 4680 31016
rect 4720 30976 4729 31016
rect 4343 30953 4409 30976
rect 4495 30953 4577 30976
rect 4663 30953 4729 30976
rect 4343 30934 4729 30953
rect 8343 31039 8729 31058
rect 8343 31016 8409 31039
rect 8495 31016 8577 31039
rect 8663 31016 8729 31039
rect 8343 30976 8352 31016
rect 8392 30976 8409 31016
rect 8495 30976 8516 31016
rect 8556 30976 8577 31016
rect 8663 30976 8680 31016
rect 8720 30976 8729 31016
rect 8343 30953 8409 30976
rect 8495 30953 8577 30976
rect 8663 30953 8729 30976
rect 8343 30934 8729 30953
rect 12343 31039 12729 31058
rect 12343 31016 12409 31039
rect 12495 31016 12577 31039
rect 12663 31016 12729 31039
rect 12343 30976 12352 31016
rect 12392 30976 12409 31016
rect 12495 30976 12516 31016
rect 12556 30976 12577 31016
rect 12663 30976 12680 31016
rect 12720 30976 12729 31016
rect 12343 30953 12409 30976
rect 12495 30953 12577 30976
rect 12663 30953 12729 30976
rect 12343 30934 12729 30953
rect 16343 31039 16729 31058
rect 16343 31016 16409 31039
rect 16495 31016 16577 31039
rect 16663 31016 16729 31039
rect 16343 30976 16352 31016
rect 16392 30976 16409 31016
rect 16495 30976 16516 31016
rect 16556 30976 16577 31016
rect 16663 30976 16680 31016
rect 16720 30976 16729 31016
rect 16343 30953 16409 30976
rect 16495 30953 16577 30976
rect 16663 30953 16729 30976
rect 16343 30934 16729 30953
rect 20343 31039 20729 31058
rect 20343 31016 20409 31039
rect 20495 31016 20577 31039
rect 20663 31016 20729 31039
rect 20343 30976 20352 31016
rect 20392 30976 20409 31016
rect 20495 30976 20516 31016
rect 20556 30976 20577 31016
rect 20663 30976 20680 31016
rect 20720 30976 20729 31016
rect 20343 30953 20409 30976
rect 20495 30953 20577 30976
rect 20663 30953 20729 30976
rect 20343 30934 20729 30953
rect 24343 31039 24729 31058
rect 24343 31016 24409 31039
rect 24495 31016 24577 31039
rect 24663 31016 24729 31039
rect 24343 30976 24352 31016
rect 24392 30976 24409 31016
rect 24495 30976 24516 31016
rect 24556 30976 24577 31016
rect 24663 30976 24680 31016
rect 24720 30976 24729 31016
rect 24343 30953 24409 30976
rect 24495 30953 24577 30976
rect 24663 30953 24729 30976
rect 24343 30934 24729 30953
rect 28343 31039 28729 31058
rect 28343 31016 28409 31039
rect 28495 31016 28577 31039
rect 28663 31016 28729 31039
rect 28343 30976 28352 31016
rect 28392 30976 28409 31016
rect 28495 30976 28516 31016
rect 28556 30976 28577 31016
rect 28663 30976 28680 31016
rect 28720 30976 28729 31016
rect 28343 30953 28409 30976
rect 28495 30953 28577 30976
rect 28663 30953 28729 30976
rect 28343 30934 28729 30953
rect 32343 31039 32729 31058
rect 32343 31016 32409 31039
rect 32495 31016 32577 31039
rect 32663 31016 32729 31039
rect 32343 30976 32352 31016
rect 32392 30976 32409 31016
rect 32495 30976 32516 31016
rect 32556 30976 32577 31016
rect 32663 30976 32680 31016
rect 32720 30976 32729 31016
rect 32343 30953 32409 30976
rect 32495 30953 32577 30976
rect 32663 30953 32729 30976
rect 32343 30934 32729 30953
rect 36343 31039 36729 31058
rect 36343 31016 36409 31039
rect 36495 31016 36577 31039
rect 36663 31016 36729 31039
rect 36343 30976 36352 31016
rect 36392 30976 36409 31016
rect 36495 30976 36516 31016
rect 36556 30976 36577 31016
rect 36663 30976 36680 31016
rect 36720 30976 36729 31016
rect 36343 30953 36409 30976
rect 36495 30953 36577 30976
rect 36663 30953 36729 30976
rect 36343 30934 36729 30953
rect 40343 31039 40729 31058
rect 40343 31016 40409 31039
rect 40495 31016 40577 31039
rect 40663 31016 40729 31039
rect 40343 30976 40352 31016
rect 40392 30976 40409 31016
rect 40495 30976 40516 31016
rect 40556 30976 40577 31016
rect 40663 30976 40680 31016
rect 40720 30976 40729 31016
rect 40343 30953 40409 30976
rect 40495 30953 40577 30976
rect 40663 30953 40729 30976
rect 40343 30934 40729 30953
rect 44343 31039 44729 31058
rect 44343 31016 44409 31039
rect 44495 31016 44577 31039
rect 44663 31016 44729 31039
rect 44343 30976 44352 31016
rect 44392 30976 44409 31016
rect 44495 30976 44516 31016
rect 44556 30976 44577 31016
rect 44663 30976 44680 31016
rect 44720 30976 44729 31016
rect 44343 30953 44409 30976
rect 44495 30953 44577 30976
rect 44663 30953 44729 30976
rect 44343 30934 44729 30953
rect 48343 31039 48729 31058
rect 48343 31016 48409 31039
rect 48495 31016 48577 31039
rect 48663 31016 48729 31039
rect 48343 30976 48352 31016
rect 48392 30976 48409 31016
rect 48495 30976 48516 31016
rect 48556 30976 48577 31016
rect 48663 30976 48680 31016
rect 48720 30976 48729 31016
rect 48343 30953 48409 30976
rect 48495 30953 48577 30976
rect 48663 30953 48729 30976
rect 48343 30934 48729 30953
rect 52343 31039 52729 31058
rect 52343 31016 52409 31039
rect 52495 31016 52577 31039
rect 52663 31016 52729 31039
rect 52343 30976 52352 31016
rect 52392 30976 52409 31016
rect 52495 30976 52516 31016
rect 52556 30976 52577 31016
rect 52663 30976 52680 31016
rect 52720 30976 52729 31016
rect 52343 30953 52409 30976
rect 52495 30953 52577 30976
rect 52663 30953 52729 30976
rect 52343 30934 52729 30953
rect 56343 31039 56729 31058
rect 56343 31016 56409 31039
rect 56495 31016 56577 31039
rect 56663 31016 56729 31039
rect 56343 30976 56352 31016
rect 56392 30976 56409 31016
rect 56495 30976 56516 31016
rect 56556 30976 56577 31016
rect 56663 30976 56680 31016
rect 56720 30976 56729 31016
rect 56343 30953 56409 30976
rect 56495 30953 56577 30976
rect 56663 30953 56729 30976
rect 56343 30934 56729 30953
rect 60343 31039 60729 31058
rect 60343 31016 60409 31039
rect 60495 31016 60577 31039
rect 60663 31016 60729 31039
rect 60343 30976 60352 31016
rect 60392 30976 60409 31016
rect 60495 30976 60516 31016
rect 60556 30976 60577 31016
rect 60663 30976 60680 31016
rect 60720 30976 60729 31016
rect 60343 30953 60409 30976
rect 60495 30953 60577 30976
rect 60663 30953 60729 30976
rect 60343 30934 60729 30953
rect 64343 31039 64729 31058
rect 64343 31016 64409 31039
rect 64495 31016 64577 31039
rect 64663 31016 64729 31039
rect 64343 30976 64352 31016
rect 64392 30976 64409 31016
rect 64495 30976 64516 31016
rect 64556 30976 64577 31016
rect 64663 30976 64680 31016
rect 64720 30976 64729 31016
rect 64343 30953 64409 30976
rect 64495 30953 64577 30976
rect 64663 30953 64729 30976
rect 64343 30934 64729 30953
rect 68343 31039 68729 31058
rect 68343 31016 68409 31039
rect 68495 31016 68577 31039
rect 68663 31016 68729 31039
rect 68343 30976 68352 31016
rect 68392 30976 68409 31016
rect 68495 30976 68516 31016
rect 68556 30976 68577 31016
rect 68663 30976 68680 31016
rect 68720 30976 68729 31016
rect 68343 30953 68409 30976
rect 68495 30953 68577 30976
rect 68663 30953 68729 30976
rect 68343 30934 68729 30953
rect 72316 31016 72756 31098
rect 72316 30930 72409 31016
rect 72495 30930 72577 31016
rect 72663 30930 72756 31016
rect 72316 30848 72756 30930
rect 72316 30762 72409 30848
rect 72495 30762 72577 30848
rect 72663 30762 72756 30848
rect 72316 30680 72756 30762
rect 72316 30594 72409 30680
rect 72495 30594 72577 30680
rect 72663 30594 72756 30680
rect 72316 30512 72756 30594
rect 72316 30426 72409 30512
rect 72495 30426 72577 30512
rect 72663 30426 72756 30512
rect 72316 30344 72756 30426
rect 3103 30283 3489 30302
rect 3103 30260 3169 30283
rect 3255 30260 3337 30283
rect 3423 30260 3489 30283
rect 3103 30220 3112 30260
rect 3152 30220 3169 30260
rect 3255 30220 3276 30260
rect 3316 30220 3337 30260
rect 3423 30220 3440 30260
rect 3480 30220 3489 30260
rect 3103 30197 3169 30220
rect 3255 30197 3337 30220
rect 3423 30197 3489 30220
rect 3103 30178 3489 30197
rect 7103 30283 7489 30302
rect 7103 30260 7169 30283
rect 7255 30260 7337 30283
rect 7423 30260 7489 30283
rect 7103 30220 7112 30260
rect 7152 30220 7169 30260
rect 7255 30220 7276 30260
rect 7316 30220 7337 30260
rect 7423 30220 7440 30260
rect 7480 30220 7489 30260
rect 7103 30197 7169 30220
rect 7255 30197 7337 30220
rect 7423 30197 7489 30220
rect 7103 30178 7489 30197
rect 11103 30283 11489 30302
rect 11103 30260 11169 30283
rect 11255 30260 11337 30283
rect 11423 30260 11489 30283
rect 11103 30220 11112 30260
rect 11152 30220 11169 30260
rect 11255 30220 11276 30260
rect 11316 30220 11337 30260
rect 11423 30220 11440 30260
rect 11480 30220 11489 30260
rect 11103 30197 11169 30220
rect 11255 30197 11337 30220
rect 11423 30197 11489 30220
rect 11103 30178 11489 30197
rect 15103 30283 15489 30302
rect 15103 30260 15169 30283
rect 15255 30260 15337 30283
rect 15423 30260 15489 30283
rect 15103 30220 15112 30260
rect 15152 30220 15169 30260
rect 15255 30220 15276 30260
rect 15316 30220 15337 30260
rect 15423 30220 15440 30260
rect 15480 30220 15489 30260
rect 15103 30197 15169 30220
rect 15255 30197 15337 30220
rect 15423 30197 15489 30220
rect 15103 30178 15489 30197
rect 19103 30283 19489 30302
rect 19103 30260 19169 30283
rect 19255 30260 19337 30283
rect 19423 30260 19489 30283
rect 19103 30220 19112 30260
rect 19152 30220 19169 30260
rect 19255 30220 19276 30260
rect 19316 30220 19337 30260
rect 19423 30220 19440 30260
rect 19480 30220 19489 30260
rect 19103 30197 19169 30220
rect 19255 30197 19337 30220
rect 19423 30197 19489 30220
rect 19103 30178 19489 30197
rect 23103 30283 23489 30302
rect 23103 30260 23169 30283
rect 23255 30260 23337 30283
rect 23423 30260 23489 30283
rect 23103 30220 23112 30260
rect 23152 30220 23169 30260
rect 23255 30220 23276 30260
rect 23316 30220 23337 30260
rect 23423 30220 23440 30260
rect 23480 30220 23489 30260
rect 23103 30197 23169 30220
rect 23255 30197 23337 30220
rect 23423 30197 23489 30220
rect 23103 30178 23489 30197
rect 27103 30283 27489 30302
rect 27103 30260 27169 30283
rect 27255 30260 27337 30283
rect 27423 30260 27489 30283
rect 27103 30220 27112 30260
rect 27152 30220 27169 30260
rect 27255 30220 27276 30260
rect 27316 30220 27337 30260
rect 27423 30220 27440 30260
rect 27480 30220 27489 30260
rect 27103 30197 27169 30220
rect 27255 30197 27337 30220
rect 27423 30197 27489 30220
rect 27103 30178 27489 30197
rect 31103 30283 31489 30302
rect 31103 30260 31169 30283
rect 31255 30260 31337 30283
rect 31423 30260 31489 30283
rect 31103 30220 31112 30260
rect 31152 30220 31169 30260
rect 31255 30220 31276 30260
rect 31316 30220 31337 30260
rect 31423 30220 31440 30260
rect 31480 30220 31489 30260
rect 31103 30197 31169 30220
rect 31255 30197 31337 30220
rect 31423 30197 31489 30220
rect 31103 30178 31489 30197
rect 35103 30283 35489 30302
rect 35103 30260 35169 30283
rect 35255 30260 35337 30283
rect 35423 30260 35489 30283
rect 35103 30220 35112 30260
rect 35152 30220 35169 30260
rect 35255 30220 35276 30260
rect 35316 30220 35337 30260
rect 35423 30220 35440 30260
rect 35480 30220 35489 30260
rect 35103 30197 35169 30220
rect 35255 30197 35337 30220
rect 35423 30197 35489 30220
rect 35103 30178 35489 30197
rect 39103 30283 39489 30302
rect 39103 30260 39169 30283
rect 39255 30260 39337 30283
rect 39423 30260 39489 30283
rect 39103 30220 39112 30260
rect 39152 30220 39169 30260
rect 39255 30220 39276 30260
rect 39316 30220 39337 30260
rect 39423 30220 39440 30260
rect 39480 30220 39489 30260
rect 39103 30197 39169 30220
rect 39255 30197 39337 30220
rect 39423 30197 39489 30220
rect 39103 30178 39489 30197
rect 43103 30283 43489 30302
rect 43103 30260 43169 30283
rect 43255 30260 43337 30283
rect 43423 30260 43489 30283
rect 43103 30220 43112 30260
rect 43152 30220 43169 30260
rect 43255 30220 43276 30260
rect 43316 30220 43337 30260
rect 43423 30220 43440 30260
rect 43480 30220 43489 30260
rect 43103 30197 43169 30220
rect 43255 30197 43337 30220
rect 43423 30197 43489 30220
rect 43103 30178 43489 30197
rect 47103 30283 47489 30302
rect 47103 30260 47169 30283
rect 47255 30260 47337 30283
rect 47423 30260 47489 30283
rect 47103 30220 47112 30260
rect 47152 30220 47169 30260
rect 47255 30220 47276 30260
rect 47316 30220 47337 30260
rect 47423 30220 47440 30260
rect 47480 30220 47489 30260
rect 47103 30197 47169 30220
rect 47255 30197 47337 30220
rect 47423 30197 47489 30220
rect 47103 30178 47489 30197
rect 51103 30283 51489 30302
rect 51103 30260 51169 30283
rect 51255 30260 51337 30283
rect 51423 30260 51489 30283
rect 51103 30220 51112 30260
rect 51152 30220 51169 30260
rect 51255 30220 51276 30260
rect 51316 30220 51337 30260
rect 51423 30220 51440 30260
rect 51480 30220 51489 30260
rect 51103 30197 51169 30220
rect 51255 30197 51337 30220
rect 51423 30197 51489 30220
rect 51103 30178 51489 30197
rect 55103 30283 55489 30302
rect 55103 30260 55169 30283
rect 55255 30260 55337 30283
rect 55423 30260 55489 30283
rect 55103 30220 55112 30260
rect 55152 30220 55169 30260
rect 55255 30220 55276 30260
rect 55316 30220 55337 30260
rect 55423 30220 55440 30260
rect 55480 30220 55489 30260
rect 55103 30197 55169 30220
rect 55255 30197 55337 30220
rect 55423 30197 55489 30220
rect 55103 30178 55489 30197
rect 59103 30283 59489 30302
rect 59103 30260 59169 30283
rect 59255 30260 59337 30283
rect 59423 30260 59489 30283
rect 59103 30220 59112 30260
rect 59152 30220 59169 30260
rect 59255 30220 59276 30260
rect 59316 30220 59337 30260
rect 59423 30220 59440 30260
rect 59480 30220 59489 30260
rect 59103 30197 59169 30220
rect 59255 30197 59337 30220
rect 59423 30197 59489 30220
rect 59103 30178 59489 30197
rect 63103 30283 63489 30302
rect 63103 30260 63169 30283
rect 63255 30260 63337 30283
rect 63423 30260 63489 30283
rect 63103 30220 63112 30260
rect 63152 30220 63169 30260
rect 63255 30220 63276 30260
rect 63316 30220 63337 30260
rect 63423 30220 63440 30260
rect 63480 30220 63489 30260
rect 63103 30197 63169 30220
rect 63255 30197 63337 30220
rect 63423 30197 63489 30220
rect 63103 30178 63489 30197
rect 67103 30283 67489 30302
rect 67103 30260 67169 30283
rect 67255 30260 67337 30283
rect 67423 30260 67489 30283
rect 67103 30220 67112 30260
rect 67152 30220 67169 30260
rect 67255 30220 67276 30260
rect 67316 30220 67337 30260
rect 67423 30220 67440 30260
rect 67480 30220 67489 30260
rect 67103 30197 67169 30220
rect 67255 30197 67337 30220
rect 67423 30197 67489 30220
rect 67103 30178 67489 30197
rect 72316 30258 72409 30344
rect 72495 30258 72577 30344
rect 72663 30258 72756 30344
rect 72316 30176 72756 30258
rect 72316 30090 72409 30176
rect 72495 30090 72577 30176
rect 72663 30090 72756 30176
rect 72316 30008 72756 30090
rect 72316 29922 72409 30008
rect 72495 29922 72577 30008
rect 72663 29922 72756 30008
rect 72316 29840 72756 29922
rect 72316 29754 72409 29840
rect 72495 29754 72577 29840
rect 72663 29754 72756 29840
rect 72316 29624 72756 29754
rect 76316 31856 76756 31986
rect 76316 31770 76409 31856
rect 76495 31770 76577 31856
rect 76663 31770 76756 31856
rect 76316 31688 76756 31770
rect 76316 31602 76409 31688
rect 76495 31602 76577 31688
rect 76663 31602 76756 31688
rect 76316 31520 76756 31602
rect 76316 31434 76409 31520
rect 76495 31434 76577 31520
rect 76663 31434 76756 31520
rect 76316 31352 76756 31434
rect 76316 31266 76409 31352
rect 76495 31266 76577 31352
rect 76663 31266 76756 31352
rect 76316 31184 76756 31266
rect 76316 31098 76409 31184
rect 76495 31098 76577 31184
rect 76663 31098 76756 31184
rect 76316 31016 76756 31098
rect 76316 30930 76409 31016
rect 76495 30930 76577 31016
rect 76663 30930 76756 31016
rect 76316 30848 76756 30930
rect 76316 30762 76409 30848
rect 76495 30762 76577 30848
rect 76663 30762 76756 30848
rect 76316 30680 76756 30762
rect 76316 30594 76409 30680
rect 76495 30594 76577 30680
rect 76663 30594 76756 30680
rect 76316 30512 76756 30594
rect 76316 30426 76409 30512
rect 76495 30426 76577 30512
rect 76663 30426 76756 30512
rect 76316 30344 76756 30426
rect 76316 30258 76409 30344
rect 76495 30258 76577 30344
rect 76663 30258 76756 30344
rect 76316 30176 76756 30258
rect 76316 30090 76409 30176
rect 76495 30090 76577 30176
rect 76663 30090 76756 30176
rect 76316 30008 76756 30090
rect 76316 29922 76409 30008
rect 76495 29922 76577 30008
rect 76663 29922 76756 30008
rect 76316 29840 76756 29922
rect 76316 29754 76409 29840
rect 76495 29754 76577 29840
rect 76663 29754 76756 29840
rect 76316 29624 76756 29754
rect 80316 31856 80756 31986
rect 80316 31770 80409 31856
rect 80495 31770 80577 31856
rect 80663 31770 80756 31856
rect 80316 31688 80756 31770
rect 80316 31602 80409 31688
rect 80495 31602 80577 31688
rect 80663 31602 80756 31688
rect 80316 31520 80756 31602
rect 80316 31434 80409 31520
rect 80495 31434 80577 31520
rect 80663 31434 80756 31520
rect 80316 31352 80756 31434
rect 80316 31266 80409 31352
rect 80495 31266 80577 31352
rect 80663 31266 80756 31352
rect 80316 31184 80756 31266
rect 80316 31098 80409 31184
rect 80495 31098 80577 31184
rect 80663 31098 80756 31184
rect 80316 31016 80756 31098
rect 80316 30930 80409 31016
rect 80495 30930 80577 31016
rect 80663 30930 80756 31016
rect 80316 30848 80756 30930
rect 80316 30762 80409 30848
rect 80495 30762 80577 30848
rect 80663 30762 80756 30848
rect 80316 30680 80756 30762
rect 80316 30594 80409 30680
rect 80495 30594 80577 30680
rect 80663 30594 80756 30680
rect 80316 30512 80756 30594
rect 80316 30426 80409 30512
rect 80495 30426 80577 30512
rect 80663 30426 80756 30512
rect 80316 30344 80756 30426
rect 80316 30258 80409 30344
rect 80495 30258 80577 30344
rect 80663 30258 80756 30344
rect 80316 30176 80756 30258
rect 80316 30090 80409 30176
rect 80495 30090 80577 30176
rect 80663 30090 80756 30176
rect 80316 30008 80756 30090
rect 80316 29922 80409 30008
rect 80495 29922 80577 30008
rect 80663 29922 80756 30008
rect 80316 29840 80756 29922
rect 80316 29754 80409 29840
rect 80495 29754 80577 29840
rect 80663 29754 80756 29840
rect 80316 29624 80756 29754
rect 84316 31856 84756 31986
rect 84316 31770 84409 31856
rect 84495 31770 84577 31856
rect 84663 31770 84756 31856
rect 84316 31688 84756 31770
rect 84316 31602 84409 31688
rect 84495 31602 84577 31688
rect 84663 31602 84756 31688
rect 84316 31520 84756 31602
rect 84316 31434 84409 31520
rect 84495 31434 84577 31520
rect 84663 31434 84756 31520
rect 84316 31352 84756 31434
rect 84316 31266 84409 31352
rect 84495 31266 84577 31352
rect 84663 31266 84756 31352
rect 84316 31184 84756 31266
rect 84316 31098 84409 31184
rect 84495 31098 84577 31184
rect 84663 31098 84756 31184
rect 84316 31016 84756 31098
rect 84316 30930 84409 31016
rect 84495 30930 84577 31016
rect 84663 30930 84756 31016
rect 84316 30848 84756 30930
rect 84316 30762 84409 30848
rect 84495 30762 84577 30848
rect 84663 30762 84756 30848
rect 84316 30680 84756 30762
rect 84316 30594 84409 30680
rect 84495 30594 84577 30680
rect 84663 30594 84756 30680
rect 84316 30512 84756 30594
rect 84316 30426 84409 30512
rect 84495 30426 84577 30512
rect 84663 30426 84756 30512
rect 84316 30344 84756 30426
rect 84316 30258 84409 30344
rect 84495 30258 84577 30344
rect 84663 30258 84756 30344
rect 84316 30176 84756 30258
rect 84316 30090 84409 30176
rect 84495 30090 84577 30176
rect 84663 30090 84756 30176
rect 84316 30008 84756 30090
rect 84316 29922 84409 30008
rect 84495 29922 84577 30008
rect 84663 29922 84756 30008
rect 84316 29840 84756 29922
rect 84316 29754 84409 29840
rect 84495 29754 84577 29840
rect 84663 29754 84756 29840
rect 84316 29624 84756 29754
rect 88316 31856 88756 31986
rect 88316 31770 88409 31856
rect 88495 31770 88577 31856
rect 88663 31770 88756 31856
rect 88316 31688 88756 31770
rect 88316 31602 88409 31688
rect 88495 31602 88577 31688
rect 88663 31602 88756 31688
rect 88316 31520 88756 31602
rect 88316 31434 88409 31520
rect 88495 31434 88577 31520
rect 88663 31434 88756 31520
rect 88316 31352 88756 31434
rect 88316 31266 88409 31352
rect 88495 31266 88577 31352
rect 88663 31266 88756 31352
rect 88316 31184 88756 31266
rect 88316 31098 88409 31184
rect 88495 31098 88577 31184
rect 88663 31098 88756 31184
rect 88316 31016 88756 31098
rect 88316 30930 88409 31016
rect 88495 30930 88577 31016
rect 88663 30930 88756 31016
rect 88316 30848 88756 30930
rect 88316 30762 88409 30848
rect 88495 30762 88577 30848
rect 88663 30762 88756 30848
rect 88316 30680 88756 30762
rect 88316 30594 88409 30680
rect 88495 30594 88577 30680
rect 88663 30594 88756 30680
rect 88316 30512 88756 30594
rect 88316 30426 88409 30512
rect 88495 30426 88577 30512
rect 88663 30426 88756 30512
rect 88316 30344 88756 30426
rect 88316 30258 88409 30344
rect 88495 30258 88577 30344
rect 88663 30258 88756 30344
rect 88316 30176 88756 30258
rect 88316 30090 88409 30176
rect 88495 30090 88577 30176
rect 88663 30090 88756 30176
rect 88316 30008 88756 30090
rect 88316 29922 88409 30008
rect 88495 29922 88577 30008
rect 88663 29922 88756 30008
rect 88316 29840 88756 29922
rect 88316 29754 88409 29840
rect 88495 29754 88577 29840
rect 88663 29754 88756 29840
rect 88316 29624 88756 29754
rect 92316 31856 92756 31986
rect 92316 31770 92409 31856
rect 92495 31770 92577 31856
rect 92663 31770 92756 31856
rect 92316 31688 92756 31770
rect 92316 31602 92409 31688
rect 92495 31602 92577 31688
rect 92663 31602 92756 31688
rect 92316 31520 92756 31602
rect 92316 31434 92409 31520
rect 92495 31434 92577 31520
rect 92663 31434 92756 31520
rect 92316 31352 92756 31434
rect 92316 31266 92409 31352
rect 92495 31266 92577 31352
rect 92663 31266 92756 31352
rect 92316 31184 92756 31266
rect 92316 31098 92409 31184
rect 92495 31098 92577 31184
rect 92663 31098 92756 31184
rect 92316 31016 92756 31098
rect 92316 30930 92409 31016
rect 92495 30930 92577 31016
rect 92663 30930 92756 31016
rect 92316 30848 92756 30930
rect 92316 30762 92409 30848
rect 92495 30762 92577 30848
rect 92663 30762 92756 30848
rect 92316 30680 92756 30762
rect 92316 30594 92409 30680
rect 92495 30594 92577 30680
rect 92663 30594 92756 30680
rect 92316 30512 92756 30594
rect 92316 30426 92409 30512
rect 92495 30426 92577 30512
rect 92663 30426 92756 30512
rect 92316 30344 92756 30426
rect 92316 30258 92409 30344
rect 92495 30258 92577 30344
rect 92663 30258 92756 30344
rect 92316 30176 92756 30258
rect 92316 30090 92409 30176
rect 92495 30090 92577 30176
rect 92663 30090 92756 30176
rect 92316 30008 92756 30090
rect 92316 29922 92409 30008
rect 92495 29922 92577 30008
rect 92663 29922 92756 30008
rect 92316 29840 92756 29922
rect 92316 29754 92409 29840
rect 92495 29754 92577 29840
rect 92663 29754 92756 29840
rect 92316 29624 92756 29754
rect 96316 31856 96756 31986
rect 96316 31770 96409 31856
rect 96495 31770 96577 31856
rect 96663 31770 96756 31856
rect 96316 31688 96756 31770
rect 96316 31602 96409 31688
rect 96495 31602 96577 31688
rect 96663 31602 96756 31688
rect 96316 31520 96756 31602
rect 96316 31434 96409 31520
rect 96495 31434 96577 31520
rect 96663 31434 96756 31520
rect 96316 31352 96756 31434
rect 96316 31266 96409 31352
rect 96495 31266 96577 31352
rect 96663 31266 96756 31352
rect 96316 31184 96756 31266
rect 96316 31098 96409 31184
rect 96495 31098 96577 31184
rect 96663 31098 96756 31184
rect 96316 31016 96756 31098
rect 96316 30930 96409 31016
rect 96495 30930 96577 31016
rect 96663 30930 96756 31016
rect 96316 30848 96756 30930
rect 96316 30762 96409 30848
rect 96495 30762 96577 30848
rect 96663 30762 96756 30848
rect 96316 30680 96756 30762
rect 96316 30594 96409 30680
rect 96495 30594 96577 30680
rect 96663 30594 96756 30680
rect 96316 30512 96756 30594
rect 96316 30426 96409 30512
rect 96495 30426 96577 30512
rect 96663 30426 96756 30512
rect 96316 30344 96756 30426
rect 96316 30258 96409 30344
rect 96495 30258 96577 30344
rect 96663 30258 96756 30344
rect 96316 30176 96756 30258
rect 96316 30090 96409 30176
rect 96495 30090 96577 30176
rect 96663 30090 96756 30176
rect 96316 30008 96756 30090
rect 96316 29922 96409 30008
rect 96495 29922 96577 30008
rect 96663 29922 96756 30008
rect 96316 29840 96756 29922
rect 96316 29754 96409 29840
rect 96495 29754 96577 29840
rect 96663 29754 96756 29840
rect 96316 29624 96756 29754
rect 4343 29527 4729 29546
rect 4343 29504 4409 29527
rect 4495 29504 4577 29527
rect 4663 29504 4729 29527
rect 4343 29464 4352 29504
rect 4392 29464 4409 29504
rect 4495 29464 4516 29504
rect 4556 29464 4577 29504
rect 4663 29464 4680 29504
rect 4720 29464 4729 29504
rect 4343 29441 4409 29464
rect 4495 29441 4577 29464
rect 4663 29441 4729 29464
rect 4343 29422 4729 29441
rect 8343 29527 8729 29546
rect 8343 29504 8409 29527
rect 8495 29504 8577 29527
rect 8663 29504 8729 29527
rect 8343 29464 8352 29504
rect 8392 29464 8409 29504
rect 8495 29464 8516 29504
rect 8556 29464 8577 29504
rect 8663 29464 8680 29504
rect 8720 29464 8729 29504
rect 8343 29441 8409 29464
rect 8495 29441 8577 29464
rect 8663 29441 8729 29464
rect 8343 29422 8729 29441
rect 12343 29527 12729 29546
rect 12343 29504 12409 29527
rect 12495 29504 12577 29527
rect 12663 29504 12729 29527
rect 12343 29464 12352 29504
rect 12392 29464 12409 29504
rect 12495 29464 12516 29504
rect 12556 29464 12577 29504
rect 12663 29464 12680 29504
rect 12720 29464 12729 29504
rect 12343 29441 12409 29464
rect 12495 29441 12577 29464
rect 12663 29441 12729 29464
rect 12343 29422 12729 29441
rect 16343 29527 16729 29546
rect 16343 29504 16409 29527
rect 16495 29504 16577 29527
rect 16663 29504 16729 29527
rect 16343 29464 16352 29504
rect 16392 29464 16409 29504
rect 16495 29464 16516 29504
rect 16556 29464 16577 29504
rect 16663 29464 16680 29504
rect 16720 29464 16729 29504
rect 16343 29441 16409 29464
rect 16495 29441 16577 29464
rect 16663 29441 16729 29464
rect 16343 29422 16729 29441
rect 20343 29527 20729 29546
rect 20343 29504 20409 29527
rect 20495 29504 20577 29527
rect 20663 29504 20729 29527
rect 20343 29464 20352 29504
rect 20392 29464 20409 29504
rect 20495 29464 20516 29504
rect 20556 29464 20577 29504
rect 20663 29464 20680 29504
rect 20720 29464 20729 29504
rect 20343 29441 20409 29464
rect 20495 29441 20577 29464
rect 20663 29441 20729 29464
rect 20343 29422 20729 29441
rect 24343 29527 24729 29546
rect 24343 29504 24409 29527
rect 24495 29504 24577 29527
rect 24663 29504 24729 29527
rect 24343 29464 24352 29504
rect 24392 29464 24409 29504
rect 24495 29464 24516 29504
rect 24556 29464 24577 29504
rect 24663 29464 24680 29504
rect 24720 29464 24729 29504
rect 24343 29441 24409 29464
rect 24495 29441 24577 29464
rect 24663 29441 24729 29464
rect 24343 29422 24729 29441
rect 28343 29527 28729 29546
rect 28343 29504 28409 29527
rect 28495 29504 28577 29527
rect 28663 29504 28729 29527
rect 28343 29464 28352 29504
rect 28392 29464 28409 29504
rect 28495 29464 28516 29504
rect 28556 29464 28577 29504
rect 28663 29464 28680 29504
rect 28720 29464 28729 29504
rect 28343 29441 28409 29464
rect 28495 29441 28577 29464
rect 28663 29441 28729 29464
rect 28343 29422 28729 29441
rect 32343 29527 32729 29546
rect 32343 29504 32409 29527
rect 32495 29504 32577 29527
rect 32663 29504 32729 29527
rect 32343 29464 32352 29504
rect 32392 29464 32409 29504
rect 32495 29464 32516 29504
rect 32556 29464 32577 29504
rect 32663 29464 32680 29504
rect 32720 29464 32729 29504
rect 32343 29441 32409 29464
rect 32495 29441 32577 29464
rect 32663 29441 32729 29464
rect 32343 29422 32729 29441
rect 36343 29527 36729 29546
rect 36343 29504 36409 29527
rect 36495 29504 36577 29527
rect 36663 29504 36729 29527
rect 36343 29464 36352 29504
rect 36392 29464 36409 29504
rect 36495 29464 36516 29504
rect 36556 29464 36577 29504
rect 36663 29464 36680 29504
rect 36720 29464 36729 29504
rect 36343 29441 36409 29464
rect 36495 29441 36577 29464
rect 36663 29441 36729 29464
rect 36343 29422 36729 29441
rect 40343 29527 40729 29546
rect 40343 29504 40409 29527
rect 40495 29504 40577 29527
rect 40663 29504 40729 29527
rect 40343 29464 40352 29504
rect 40392 29464 40409 29504
rect 40495 29464 40516 29504
rect 40556 29464 40577 29504
rect 40663 29464 40680 29504
rect 40720 29464 40729 29504
rect 40343 29441 40409 29464
rect 40495 29441 40577 29464
rect 40663 29441 40729 29464
rect 40343 29422 40729 29441
rect 44343 29527 44729 29546
rect 44343 29504 44409 29527
rect 44495 29504 44577 29527
rect 44663 29504 44729 29527
rect 44343 29464 44352 29504
rect 44392 29464 44409 29504
rect 44495 29464 44516 29504
rect 44556 29464 44577 29504
rect 44663 29464 44680 29504
rect 44720 29464 44729 29504
rect 44343 29441 44409 29464
rect 44495 29441 44577 29464
rect 44663 29441 44729 29464
rect 44343 29422 44729 29441
rect 48343 29527 48729 29546
rect 48343 29504 48409 29527
rect 48495 29504 48577 29527
rect 48663 29504 48729 29527
rect 48343 29464 48352 29504
rect 48392 29464 48409 29504
rect 48495 29464 48516 29504
rect 48556 29464 48577 29504
rect 48663 29464 48680 29504
rect 48720 29464 48729 29504
rect 48343 29441 48409 29464
rect 48495 29441 48577 29464
rect 48663 29441 48729 29464
rect 48343 29422 48729 29441
rect 52343 29527 52729 29546
rect 52343 29504 52409 29527
rect 52495 29504 52577 29527
rect 52663 29504 52729 29527
rect 52343 29464 52352 29504
rect 52392 29464 52409 29504
rect 52495 29464 52516 29504
rect 52556 29464 52577 29504
rect 52663 29464 52680 29504
rect 52720 29464 52729 29504
rect 52343 29441 52409 29464
rect 52495 29441 52577 29464
rect 52663 29441 52729 29464
rect 52343 29422 52729 29441
rect 56343 29527 56729 29546
rect 56343 29504 56409 29527
rect 56495 29504 56577 29527
rect 56663 29504 56729 29527
rect 56343 29464 56352 29504
rect 56392 29464 56409 29504
rect 56495 29464 56516 29504
rect 56556 29464 56577 29504
rect 56663 29464 56680 29504
rect 56720 29464 56729 29504
rect 56343 29441 56409 29464
rect 56495 29441 56577 29464
rect 56663 29441 56729 29464
rect 56343 29422 56729 29441
rect 60343 29527 60729 29546
rect 60343 29504 60409 29527
rect 60495 29504 60577 29527
rect 60663 29504 60729 29527
rect 60343 29464 60352 29504
rect 60392 29464 60409 29504
rect 60495 29464 60516 29504
rect 60556 29464 60577 29504
rect 60663 29464 60680 29504
rect 60720 29464 60729 29504
rect 60343 29441 60409 29464
rect 60495 29441 60577 29464
rect 60663 29441 60729 29464
rect 60343 29422 60729 29441
rect 64343 29527 64729 29546
rect 64343 29504 64409 29527
rect 64495 29504 64577 29527
rect 64663 29504 64729 29527
rect 64343 29464 64352 29504
rect 64392 29464 64409 29504
rect 64495 29464 64516 29504
rect 64556 29464 64577 29504
rect 64663 29464 64680 29504
rect 64720 29464 64729 29504
rect 64343 29441 64409 29464
rect 64495 29441 64577 29464
rect 64663 29441 64729 29464
rect 64343 29422 64729 29441
rect 68343 29527 68729 29546
rect 68343 29504 68409 29527
rect 68495 29504 68577 29527
rect 68663 29504 68729 29527
rect 68343 29464 68352 29504
rect 68392 29464 68409 29504
rect 68495 29464 68516 29504
rect 68556 29464 68577 29504
rect 68663 29464 68680 29504
rect 68720 29464 68729 29504
rect 68343 29441 68409 29464
rect 68495 29441 68577 29464
rect 68663 29441 68729 29464
rect 68343 29422 68729 29441
rect 75076 28980 75516 29110
rect 75076 28894 75169 28980
rect 75255 28894 75337 28980
rect 75423 28894 75516 28980
rect 75076 28812 75516 28894
rect 3103 28771 3489 28790
rect 3103 28748 3169 28771
rect 3255 28748 3337 28771
rect 3423 28748 3489 28771
rect 3103 28708 3112 28748
rect 3152 28708 3169 28748
rect 3255 28708 3276 28748
rect 3316 28708 3337 28748
rect 3423 28708 3440 28748
rect 3480 28708 3489 28748
rect 3103 28685 3169 28708
rect 3255 28685 3337 28708
rect 3423 28685 3489 28708
rect 3103 28666 3489 28685
rect 7103 28771 7489 28790
rect 7103 28748 7169 28771
rect 7255 28748 7337 28771
rect 7423 28748 7489 28771
rect 7103 28708 7112 28748
rect 7152 28708 7169 28748
rect 7255 28708 7276 28748
rect 7316 28708 7337 28748
rect 7423 28708 7440 28748
rect 7480 28708 7489 28748
rect 7103 28685 7169 28708
rect 7255 28685 7337 28708
rect 7423 28685 7489 28708
rect 7103 28666 7489 28685
rect 11103 28771 11489 28790
rect 11103 28748 11169 28771
rect 11255 28748 11337 28771
rect 11423 28748 11489 28771
rect 11103 28708 11112 28748
rect 11152 28708 11169 28748
rect 11255 28708 11276 28748
rect 11316 28708 11337 28748
rect 11423 28708 11440 28748
rect 11480 28708 11489 28748
rect 11103 28685 11169 28708
rect 11255 28685 11337 28708
rect 11423 28685 11489 28708
rect 11103 28666 11489 28685
rect 15103 28771 15489 28790
rect 15103 28748 15169 28771
rect 15255 28748 15337 28771
rect 15423 28748 15489 28771
rect 15103 28708 15112 28748
rect 15152 28708 15169 28748
rect 15255 28708 15276 28748
rect 15316 28708 15337 28748
rect 15423 28708 15440 28748
rect 15480 28708 15489 28748
rect 15103 28685 15169 28708
rect 15255 28685 15337 28708
rect 15423 28685 15489 28708
rect 15103 28666 15489 28685
rect 19103 28771 19489 28790
rect 19103 28748 19169 28771
rect 19255 28748 19337 28771
rect 19423 28748 19489 28771
rect 19103 28708 19112 28748
rect 19152 28708 19169 28748
rect 19255 28708 19276 28748
rect 19316 28708 19337 28748
rect 19423 28708 19440 28748
rect 19480 28708 19489 28748
rect 19103 28685 19169 28708
rect 19255 28685 19337 28708
rect 19423 28685 19489 28708
rect 19103 28666 19489 28685
rect 23103 28771 23489 28790
rect 23103 28748 23169 28771
rect 23255 28748 23337 28771
rect 23423 28748 23489 28771
rect 23103 28708 23112 28748
rect 23152 28708 23169 28748
rect 23255 28708 23276 28748
rect 23316 28708 23337 28748
rect 23423 28708 23440 28748
rect 23480 28708 23489 28748
rect 23103 28685 23169 28708
rect 23255 28685 23337 28708
rect 23423 28685 23489 28708
rect 23103 28666 23489 28685
rect 27103 28771 27489 28790
rect 27103 28748 27169 28771
rect 27255 28748 27337 28771
rect 27423 28748 27489 28771
rect 27103 28708 27112 28748
rect 27152 28708 27169 28748
rect 27255 28708 27276 28748
rect 27316 28708 27337 28748
rect 27423 28708 27440 28748
rect 27480 28708 27489 28748
rect 27103 28685 27169 28708
rect 27255 28685 27337 28708
rect 27423 28685 27489 28708
rect 27103 28666 27489 28685
rect 31103 28771 31489 28790
rect 31103 28748 31169 28771
rect 31255 28748 31337 28771
rect 31423 28748 31489 28771
rect 31103 28708 31112 28748
rect 31152 28708 31169 28748
rect 31255 28708 31276 28748
rect 31316 28708 31337 28748
rect 31423 28708 31440 28748
rect 31480 28708 31489 28748
rect 31103 28685 31169 28708
rect 31255 28685 31337 28708
rect 31423 28685 31489 28708
rect 31103 28666 31489 28685
rect 35103 28771 35489 28790
rect 35103 28748 35169 28771
rect 35255 28748 35337 28771
rect 35423 28748 35489 28771
rect 35103 28708 35112 28748
rect 35152 28708 35169 28748
rect 35255 28708 35276 28748
rect 35316 28708 35337 28748
rect 35423 28708 35440 28748
rect 35480 28708 35489 28748
rect 35103 28685 35169 28708
rect 35255 28685 35337 28708
rect 35423 28685 35489 28708
rect 35103 28666 35489 28685
rect 39103 28771 39489 28790
rect 39103 28748 39169 28771
rect 39255 28748 39337 28771
rect 39423 28748 39489 28771
rect 39103 28708 39112 28748
rect 39152 28708 39169 28748
rect 39255 28708 39276 28748
rect 39316 28708 39337 28748
rect 39423 28708 39440 28748
rect 39480 28708 39489 28748
rect 39103 28685 39169 28708
rect 39255 28685 39337 28708
rect 39423 28685 39489 28708
rect 39103 28666 39489 28685
rect 43103 28771 43489 28790
rect 43103 28748 43169 28771
rect 43255 28748 43337 28771
rect 43423 28748 43489 28771
rect 43103 28708 43112 28748
rect 43152 28708 43169 28748
rect 43255 28708 43276 28748
rect 43316 28708 43337 28748
rect 43423 28708 43440 28748
rect 43480 28708 43489 28748
rect 43103 28685 43169 28708
rect 43255 28685 43337 28708
rect 43423 28685 43489 28708
rect 43103 28666 43489 28685
rect 47103 28771 47489 28790
rect 47103 28748 47169 28771
rect 47255 28748 47337 28771
rect 47423 28748 47489 28771
rect 47103 28708 47112 28748
rect 47152 28708 47169 28748
rect 47255 28708 47276 28748
rect 47316 28708 47337 28748
rect 47423 28708 47440 28748
rect 47480 28708 47489 28748
rect 47103 28685 47169 28708
rect 47255 28685 47337 28708
rect 47423 28685 47489 28708
rect 47103 28666 47489 28685
rect 51103 28771 51489 28790
rect 51103 28748 51169 28771
rect 51255 28748 51337 28771
rect 51423 28748 51489 28771
rect 51103 28708 51112 28748
rect 51152 28708 51169 28748
rect 51255 28708 51276 28748
rect 51316 28708 51337 28748
rect 51423 28708 51440 28748
rect 51480 28708 51489 28748
rect 51103 28685 51169 28708
rect 51255 28685 51337 28708
rect 51423 28685 51489 28708
rect 51103 28666 51489 28685
rect 55103 28771 55489 28790
rect 55103 28748 55169 28771
rect 55255 28748 55337 28771
rect 55423 28748 55489 28771
rect 55103 28708 55112 28748
rect 55152 28708 55169 28748
rect 55255 28708 55276 28748
rect 55316 28708 55337 28748
rect 55423 28708 55440 28748
rect 55480 28708 55489 28748
rect 55103 28685 55169 28708
rect 55255 28685 55337 28708
rect 55423 28685 55489 28708
rect 55103 28666 55489 28685
rect 59103 28771 59489 28790
rect 59103 28748 59169 28771
rect 59255 28748 59337 28771
rect 59423 28748 59489 28771
rect 59103 28708 59112 28748
rect 59152 28708 59169 28748
rect 59255 28708 59276 28748
rect 59316 28708 59337 28748
rect 59423 28708 59440 28748
rect 59480 28708 59489 28748
rect 59103 28685 59169 28708
rect 59255 28685 59337 28708
rect 59423 28685 59489 28708
rect 59103 28666 59489 28685
rect 63103 28771 63489 28790
rect 63103 28748 63169 28771
rect 63255 28748 63337 28771
rect 63423 28748 63489 28771
rect 63103 28708 63112 28748
rect 63152 28708 63169 28748
rect 63255 28708 63276 28748
rect 63316 28708 63337 28748
rect 63423 28708 63440 28748
rect 63480 28708 63489 28748
rect 63103 28685 63169 28708
rect 63255 28685 63337 28708
rect 63423 28685 63489 28708
rect 63103 28666 63489 28685
rect 67103 28771 67489 28790
rect 67103 28748 67169 28771
rect 67255 28748 67337 28771
rect 67423 28748 67489 28771
rect 67103 28708 67112 28748
rect 67152 28708 67169 28748
rect 67255 28708 67276 28748
rect 67316 28708 67337 28748
rect 67423 28708 67440 28748
rect 67480 28708 67489 28748
rect 67103 28685 67169 28708
rect 67255 28685 67337 28708
rect 67423 28685 67489 28708
rect 67103 28666 67489 28685
rect 75076 28726 75169 28812
rect 75255 28726 75337 28812
rect 75423 28726 75516 28812
rect 75076 28644 75516 28726
rect 75076 28558 75169 28644
rect 75255 28558 75337 28644
rect 75423 28558 75516 28644
rect 75076 28476 75516 28558
rect 75076 28390 75169 28476
rect 75255 28390 75337 28476
rect 75423 28390 75516 28476
rect 75076 28308 75516 28390
rect 75076 28222 75169 28308
rect 75255 28222 75337 28308
rect 75423 28222 75516 28308
rect 75076 28140 75516 28222
rect 75076 28054 75169 28140
rect 75255 28054 75337 28140
rect 75423 28054 75516 28140
rect 4343 28015 4729 28034
rect 4343 27992 4409 28015
rect 4495 27992 4577 28015
rect 4663 27992 4729 28015
rect 4343 27952 4352 27992
rect 4392 27952 4409 27992
rect 4495 27952 4516 27992
rect 4556 27952 4577 27992
rect 4663 27952 4680 27992
rect 4720 27952 4729 27992
rect 4343 27929 4409 27952
rect 4495 27929 4577 27952
rect 4663 27929 4729 27952
rect 4343 27910 4729 27929
rect 8343 28015 8729 28034
rect 8343 27992 8409 28015
rect 8495 27992 8577 28015
rect 8663 27992 8729 28015
rect 8343 27952 8352 27992
rect 8392 27952 8409 27992
rect 8495 27952 8516 27992
rect 8556 27952 8577 27992
rect 8663 27952 8680 27992
rect 8720 27952 8729 27992
rect 8343 27929 8409 27952
rect 8495 27929 8577 27952
rect 8663 27929 8729 27952
rect 8343 27910 8729 27929
rect 12343 28015 12729 28034
rect 12343 27992 12409 28015
rect 12495 27992 12577 28015
rect 12663 27992 12729 28015
rect 12343 27952 12352 27992
rect 12392 27952 12409 27992
rect 12495 27952 12516 27992
rect 12556 27952 12577 27992
rect 12663 27952 12680 27992
rect 12720 27952 12729 27992
rect 12343 27929 12409 27952
rect 12495 27929 12577 27952
rect 12663 27929 12729 27952
rect 12343 27910 12729 27929
rect 16343 28015 16729 28034
rect 16343 27992 16409 28015
rect 16495 27992 16577 28015
rect 16663 27992 16729 28015
rect 16343 27952 16352 27992
rect 16392 27952 16409 27992
rect 16495 27952 16516 27992
rect 16556 27952 16577 27992
rect 16663 27952 16680 27992
rect 16720 27952 16729 27992
rect 16343 27929 16409 27952
rect 16495 27929 16577 27952
rect 16663 27929 16729 27952
rect 16343 27910 16729 27929
rect 20343 28015 20729 28034
rect 20343 27992 20409 28015
rect 20495 27992 20577 28015
rect 20663 27992 20729 28015
rect 20343 27952 20352 27992
rect 20392 27952 20409 27992
rect 20495 27952 20516 27992
rect 20556 27952 20577 27992
rect 20663 27952 20680 27992
rect 20720 27952 20729 27992
rect 20343 27929 20409 27952
rect 20495 27929 20577 27952
rect 20663 27929 20729 27952
rect 20343 27910 20729 27929
rect 24343 28015 24729 28034
rect 24343 27992 24409 28015
rect 24495 27992 24577 28015
rect 24663 27992 24729 28015
rect 24343 27952 24352 27992
rect 24392 27952 24409 27992
rect 24495 27952 24516 27992
rect 24556 27952 24577 27992
rect 24663 27952 24680 27992
rect 24720 27952 24729 27992
rect 24343 27929 24409 27952
rect 24495 27929 24577 27952
rect 24663 27929 24729 27952
rect 24343 27910 24729 27929
rect 28343 28015 28729 28034
rect 28343 27992 28409 28015
rect 28495 27992 28577 28015
rect 28663 27992 28729 28015
rect 28343 27952 28352 27992
rect 28392 27952 28409 27992
rect 28495 27952 28516 27992
rect 28556 27952 28577 27992
rect 28663 27952 28680 27992
rect 28720 27952 28729 27992
rect 28343 27929 28409 27952
rect 28495 27929 28577 27952
rect 28663 27929 28729 27952
rect 28343 27910 28729 27929
rect 32343 28015 32729 28034
rect 32343 27992 32409 28015
rect 32495 27992 32577 28015
rect 32663 27992 32729 28015
rect 32343 27952 32352 27992
rect 32392 27952 32409 27992
rect 32495 27952 32516 27992
rect 32556 27952 32577 27992
rect 32663 27952 32680 27992
rect 32720 27952 32729 27992
rect 32343 27929 32409 27952
rect 32495 27929 32577 27952
rect 32663 27929 32729 27952
rect 32343 27910 32729 27929
rect 36343 28015 36729 28034
rect 36343 27992 36409 28015
rect 36495 27992 36577 28015
rect 36663 27992 36729 28015
rect 36343 27952 36352 27992
rect 36392 27952 36409 27992
rect 36495 27952 36516 27992
rect 36556 27952 36577 27992
rect 36663 27952 36680 27992
rect 36720 27952 36729 27992
rect 36343 27929 36409 27952
rect 36495 27929 36577 27952
rect 36663 27929 36729 27952
rect 36343 27910 36729 27929
rect 40343 28015 40729 28034
rect 40343 27992 40409 28015
rect 40495 27992 40577 28015
rect 40663 27992 40729 28015
rect 40343 27952 40352 27992
rect 40392 27952 40409 27992
rect 40495 27952 40516 27992
rect 40556 27952 40577 27992
rect 40663 27952 40680 27992
rect 40720 27952 40729 27992
rect 40343 27929 40409 27952
rect 40495 27929 40577 27952
rect 40663 27929 40729 27952
rect 40343 27910 40729 27929
rect 44343 28015 44729 28034
rect 44343 27992 44409 28015
rect 44495 27992 44577 28015
rect 44663 27992 44729 28015
rect 44343 27952 44352 27992
rect 44392 27952 44409 27992
rect 44495 27952 44516 27992
rect 44556 27952 44577 27992
rect 44663 27952 44680 27992
rect 44720 27952 44729 27992
rect 44343 27929 44409 27952
rect 44495 27929 44577 27952
rect 44663 27929 44729 27952
rect 44343 27910 44729 27929
rect 48343 28015 48729 28034
rect 48343 27992 48409 28015
rect 48495 27992 48577 28015
rect 48663 27992 48729 28015
rect 48343 27952 48352 27992
rect 48392 27952 48409 27992
rect 48495 27952 48516 27992
rect 48556 27952 48577 27992
rect 48663 27952 48680 27992
rect 48720 27952 48729 27992
rect 48343 27929 48409 27952
rect 48495 27929 48577 27952
rect 48663 27929 48729 27952
rect 48343 27910 48729 27929
rect 52343 28015 52729 28034
rect 52343 27992 52409 28015
rect 52495 27992 52577 28015
rect 52663 27992 52729 28015
rect 52343 27952 52352 27992
rect 52392 27952 52409 27992
rect 52495 27952 52516 27992
rect 52556 27952 52577 27992
rect 52663 27952 52680 27992
rect 52720 27952 52729 27992
rect 52343 27929 52409 27952
rect 52495 27929 52577 27952
rect 52663 27929 52729 27952
rect 52343 27910 52729 27929
rect 56343 28015 56729 28034
rect 56343 27992 56409 28015
rect 56495 27992 56577 28015
rect 56663 27992 56729 28015
rect 56343 27952 56352 27992
rect 56392 27952 56409 27992
rect 56495 27952 56516 27992
rect 56556 27952 56577 27992
rect 56663 27952 56680 27992
rect 56720 27952 56729 27992
rect 56343 27929 56409 27952
rect 56495 27929 56577 27952
rect 56663 27929 56729 27952
rect 56343 27910 56729 27929
rect 60343 28015 60729 28034
rect 60343 27992 60409 28015
rect 60495 27992 60577 28015
rect 60663 27992 60729 28015
rect 60343 27952 60352 27992
rect 60392 27952 60409 27992
rect 60495 27952 60516 27992
rect 60556 27952 60577 27992
rect 60663 27952 60680 27992
rect 60720 27952 60729 27992
rect 60343 27929 60409 27952
rect 60495 27929 60577 27952
rect 60663 27929 60729 27952
rect 60343 27910 60729 27929
rect 64343 28015 64729 28034
rect 64343 27992 64409 28015
rect 64495 27992 64577 28015
rect 64663 27992 64729 28015
rect 64343 27952 64352 27992
rect 64392 27952 64409 27992
rect 64495 27952 64516 27992
rect 64556 27952 64577 27992
rect 64663 27952 64680 27992
rect 64720 27952 64729 27992
rect 64343 27929 64409 27952
rect 64495 27929 64577 27952
rect 64663 27929 64729 27952
rect 64343 27910 64729 27929
rect 68343 28015 68729 28034
rect 68343 27992 68409 28015
rect 68495 27992 68577 28015
rect 68663 27992 68729 28015
rect 68343 27952 68352 27992
rect 68392 27952 68409 27992
rect 68495 27952 68516 27992
rect 68556 27952 68577 27992
rect 68663 27952 68680 27992
rect 68720 27952 68729 27992
rect 68343 27929 68409 27952
rect 68495 27929 68577 27952
rect 68663 27929 68729 27952
rect 68343 27910 68729 27929
rect 75076 27972 75516 28054
rect 75076 27886 75169 27972
rect 75255 27886 75337 27972
rect 75423 27886 75516 27972
rect 75076 27804 75516 27886
rect 75076 27718 75169 27804
rect 75255 27718 75337 27804
rect 75423 27718 75516 27804
rect 75076 27636 75516 27718
rect 75076 27550 75169 27636
rect 75255 27550 75337 27636
rect 75423 27550 75516 27636
rect 75076 27468 75516 27550
rect 75076 27382 75169 27468
rect 75255 27382 75337 27468
rect 75423 27382 75516 27468
rect 75076 27300 75516 27382
rect 3103 27259 3489 27278
rect 3103 27236 3169 27259
rect 3255 27236 3337 27259
rect 3423 27236 3489 27259
rect 3103 27196 3112 27236
rect 3152 27196 3169 27236
rect 3255 27196 3276 27236
rect 3316 27196 3337 27236
rect 3423 27196 3440 27236
rect 3480 27196 3489 27236
rect 3103 27173 3169 27196
rect 3255 27173 3337 27196
rect 3423 27173 3489 27196
rect 3103 27154 3489 27173
rect 7103 27259 7489 27278
rect 7103 27236 7169 27259
rect 7255 27236 7337 27259
rect 7423 27236 7489 27259
rect 7103 27196 7112 27236
rect 7152 27196 7169 27236
rect 7255 27196 7276 27236
rect 7316 27196 7337 27236
rect 7423 27196 7440 27236
rect 7480 27196 7489 27236
rect 7103 27173 7169 27196
rect 7255 27173 7337 27196
rect 7423 27173 7489 27196
rect 7103 27154 7489 27173
rect 11103 27259 11489 27278
rect 11103 27236 11169 27259
rect 11255 27236 11337 27259
rect 11423 27236 11489 27259
rect 11103 27196 11112 27236
rect 11152 27196 11169 27236
rect 11255 27196 11276 27236
rect 11316 27196 11337 27236
rect 11423 27196 11440 27236
rect 11480 27196 11489 27236
rect 11103 27173 11169 27196
rect 11255 27173 11337 27196
rect 11423 27173 11489 27196
rect 11103 27154 11489 27173
rect 15103 27259 15489 27278
rect 15103 27236 15169 27259
rect 15255 27236 15337 27259
rect 15423 27236 15489 27259
rect 15103 27196 15112 27236
rect 15152 27196 15169 27236
rect 15255 27196 15276 27236
rect 15316 27196 15337 27236
rect 15423 27196 15440 27236
rect 15480 27196 15489 27236
rect 15103 27173 15169 27196
rect 15255 27173 15337 27196
rect 15423 27173 15489 27196
rect 15103 27154 15489 27173
rect 19103 27259 19489 27278
rect 19103 27236 19169 27259
rect 19255 27236 19337 27259
rect 19423 27236 19489 27259
rect 19103 27196 19112 27236
rect 19152 27196 19169 27236
rect 19255 27196 19276 27236
rect 19316 27196 19337 27236
rect 19423 27196 19440 27236
rect 19480 27196 19489 27236
rect 19103 27173 19169 27196
rect 19255 27173 19337 27196
rect 19423 27173 19489 27196
rect 19103 27154 19489 27173
rect 23103 27259 23489 27278
rect 23103 27236 23169 27259
rect 23255 27236 23337 27259
rect 23423 27236 23489 27259
rect 23103 27196 23112 27236
rect 23152 27196 23169 27236
rect 23255 27196 23276 27236
rect 23316 27196 23337 27236
rect 23423 27196 23440 27236
rect 23480 27196 23489 27236
rect 23103 27173 23169 27196
rect 23255 27173 23337 27196
rect 23423 27173 23489 27196
rect 23103 27154 23489 27173
rect 27103 27259 27489 27278
rect 27103 27236 27169 27259
rect 27255 27236 27337 27259
rect 27423 27236 27489 27259
rect 27103 27196 27112 27236
rect 27152 27196 27169 27236
rect 27255 27196 27276 27236
rect 27316 27196 27337 27236
rect 27423 27196 27440 27236
rect 27480 27196 27489 27236
rect 27103 27173 27169 27196
rect 27255 27173 27337 27196
rect 27423 27173 27489 27196
rect 27103 27154 27489 27173
rect 31103 27259 31489 27278
rect 31103 27236 31169 27259
rect 31255 27236 31337 27259
rect 31423 27236 31489 27259
rect 31103 27196 31112 27236
rect 31152 27196 31169 27236
rect 31255 27196 31276 27236
rect 31316 27196 31337 27236
rect 31423 27196 31440 27236
rect 31480 27196 31489 27236
rect 31103 27173 31169 27196
rect 31255 27173 31337 27196
rect 31423 27173 31489 27196
rect 31103 27154 31489 27173
rect 35103 27259 35489 27278
rect 35103 27236 35169 27259
rect 35255 27236 35337 27259
rect 35423 27236 35489 27259
rect 35103 27196 35112 27236
rect 35152 27196 35169 27236
rect 35255 27196 35276 27236
rect 35316 27196 35337 27236
rect 35423 27196 35440 27236
rect 35480 27196 35489 27236
rect 35103 27173 35169 27196
rect 35255 27173 35337 27196
rect 35423 27173 35489 27196
rect 35103 27154 35489 27173
rect 39103 27259 39489 27278
rect 39103 27236 39169 27259
rect 39255 27236 39337 27259
rect 39423 27236 39489 27259
rect 39103 27196 39112 27236
rect 39152 27196 39169 27236
rect 39255 27196 39276 27236
rect 39316 27196 39337 27236
rect 39423 27196 39440 27236
rect 39480 27196 39489 27236
rect 39103 27173 39169 27196
rect 39255 27173 39337 27196
rect 39423 27173 39489 27196
rect 39103 27154 39489 27173
rect 43103 27259 43489 27278
rect 43103 27236 43169 27259
rect 43255 27236 43337 27259
rect 43423 27236 43489 27259
rect 43103 27196 43112 27236
rect 43152 27196 43169 27236
rect 43255 27196 43276 27236
rect 43316 27196 43337 27236
rect 43423 27196 43440 27236
rect 43480 27196 43489 27236
rect 43103 27173 43169 27196
rect 43255 27173 43337 27196
rect 43423 27173 43489 27196
rect 43103 27154 43489 27173
rect 47103 27259 47489 27278
rect 47103 27236 47169 27259
rect 47255 27236 47337 27259
rect 47423 27236 47489 27259
rect 47103 27196 47112 27236
rect 47152 27196 47169 27236
rect 47255 27196 47276 27236
rect 47316 27196 47337 27236
rect 47423 27196 47440 27236
rect 47480 27196 47489 27236
rect 47103 27173 47169 27196
rect 47255 27173 47337 27196
rect 47423 27173 47489 27196
rect 47103 27154 47489 27173
rect 51103 27259 51489 27278
rect 51103 27236 51169 27259
rect 51255 27236 51337 27259
rect 51423 27236 51489 27259
rect 51103 27196 51112 27236
rect 51152 27196 51169 27236
rect 51255 27196 51276 27236
rect 51316 27196 51337 27236
rect 51423 27196 51440 27236
rect 51480 27196 51489 27236
rect 51103 27173 51169 27196
rect 51255 27173 51337 27196
rect 51423 27173 51489 27196
rect 51103 27154 51489 27173
rect 55103 27259 55489 27278
rect 55103 27236 55169 27259
rect 55255 27236 55337 27259
rect 55423 27236 55489 27259
rect 55103 27196 55112 27236
rect 55152 27196 55169 27236
rect 55255 27196 55276 27236
rect 55316 27196 55337 27236
rect 55423 27196 55440 27236
rect 55480 27196 55489 27236
rect 55103 27173 55169 27196
rect 55255 27173 55337 27196
rect 55423 27173 55489 27196
rect 55103 27154 55489 27173
rect 59103 27259 59489 27278
rect 59103 27236 59169 27259
rect 59255 27236 59337 27259
rect 59423 27236 59489 27259
rect 59103 27196 59112 27236
rect 59152 27196 59169 27236
rect 59255 27196 59276 27236
rect 59316 27196 59337 27236
rect 59423 27196 59440 27236
rect 59480 27196 59489 27236
rect 59103 27173 59169 27196
rect 59255 27173 59337 27196
rect 59423 27173 59489 27196
rect 59103 27154 59489 27173
rect 63103 27259 63489 27278
rect 63103 27236 63169 27259
rect 63255 27236 63337 27259
rect 63423 27236 63489 27259
rect 63103 27196 63112 27236
rect 63152 27196 63169 27236
rect 63255 27196 63276 27236
rect 63316 27196 63337 27236
rect 63423 27196 63440 27236
rect 63480 27196 63489 27236
rect 63103 27173 63169 27196
rect 63255 27173 63337 27196
rect 63423 27173 63489 27196
rect 63103 27154 63489 27173
rect 67103 27259 67489 27278
rect 67103 27236 67169 27259
rect 67255 27236 67337 27259
rect 67423 27236 67489 27259
rect 67103 27196 67112 27236
rect 67152 27196 67169 27236
rect 67255 27196 67276 27236
rect 67316 27196 67337 27236
rect 67423 27196 67440 27236
rect 67480 27196 67489 27236
rect 67103 27173 67169 27196
rect 67255 27173 67337 27196
rect 67423 27173 67489 27196
rect 67103 27154 67489 27173
rect 75076 27214 75169 27300
rect 75255 27214 75337 27300
rect 75423 27214 75516 27300
rect 75076 27132 75516 27214
rect 75076 27046 75169 27132
rect 75255 27046 75337 27132
rect 75423 27046 75516 27132
rect 75076 26964 75516 27046
rect 75076 26878 75169 26964
rect 75255 26878 75337 26964
rect 75423 26878 75516 26964
rect 75076 26748 75516 26878
rect 79076 28980 79516 29110
rect 79076 28894 79169 28980
rect 79255 28894 79337 28980
rect 79423 28894 79516 28980
rect 79076 28812 79516 28894
rect 79076 28726 79169 28812
rect 79255 28726 79337 28812
rect 79423 28726 79516 28812
rect 79076 28644 79516 28726
rect 79076 28558 79169 28644
rect 79255 28558 79337 28644
rect 79423 28558 79516 28644
rect 79076 28476 79516 28558
rect 79076 28390 79169 28476
rect 79255 28390 79337 28476
rect 79423 28390 79516 28476
rect 79076 28308 79516 28390
rect 79076 28222 79169 28308
rect 79255 28222 79337 28308
rect 79423 28222 79516 28308
rect 79076 28140 79516 28222
rect 79076 28054 79169 28140
rect 79255 28054 79337 28140
rect 79423 28054 79516 28140
rect 79076 27972 79516 28054
rect 79076 27886 79169 27972
rect 79255 27886 79337 27972
rect 79423 27886 79516 27972
rect 79076 27804 79516 27886
rect 79076 27718 79169 27804
rect 79255 27718 79337 27804
rect 79423 27718 79516 27804
rect 79076 27636 79516 27718
rect 79076 27550 79169 27636
rect 79255 27550 79337 27636
rect 79423 27550 79516 27636
rect 79076 27468 79516 27550
rect 79076 27382 79169 27468
rect 79255 27382 79337 27468
rect 79423 27382 79516 27468
rect 79076 27300 79516 27382
rect 79076 27214 79169 27300
rect 79255 27214 79337 27300
rect 79423 27214 79516 27300
rect 79076 27132 79516 27214
rect 79076 27046 79169 27132
rect 79255 27046 79337 27132
rect 79423 27046 79516 27132
rect 79076 26964 79516 27046
rect 79076 26878 79169 26964
rect 79255 26878 79337 26964
rect 79423 26878 79516 26964
rect 79076 26748 79516 26878
rect 83076 28980 83516 29110
rect 83076 28894 83169 28980
rect 83255 28894 83337 28980
rect 83423 28894 83516 28980
rect 83076 28812 83516 28894
rect 83076 28726 83169 28812
rect 83255 28726 83337 28812
rect 83423 28726 83516 28812
rect 83076 28644 83516 28726
rect 83076 28558 83169 28644
rect 83255 28558 83337 28644
rect 83423 28558 83516 28644
rect 83076 28476 83516 28558
rect 83076 28390 83169 28476
rect 83255 28390 83337 28476
rect 83423 28390 83516 28476
rect 83076 28308 83516 28390
rect 83076 28222 83169 28308
rect 83255 28222 83337 28308
rect 83423 28222 83516 28308
rect 83076 28140 83516 28222
rect 83076 28054 83169 28140
rect 83255 28054 83337 28140
rect 83423 28054 83516 28140
rect 83076 27972 83516 28054
rect 83076 27886 83169 27972
rect 83255 27886 83337 27972
rect 83423 27886 83516 27972
rect 83076 27804 83516 27886
rect 83076 27718 83169 27804
rect 83255 27718 83337 27804
rect 83423 27718 83516 27804
rect 83076 27636 83516 27718
rect 83076 27550 83169 27636
rect 83255 27550 83337 27636
rect 83423 27550 83516 27636
rect 83076 27468 83516 27550
rect 83076 27382 83169 27468
rect 83255 27382 83337 27468
rect 83423 27382 83516 27468
rect 83076 27300 83516 27382
rect 83076 27214 83169 27300
rect 83255 27214 83337 27300
rect 83423 27214 83516 27300
rect 83076 27132 83516 27214
rect 83076 27046 83169 27132
rect 83255 27046 83337 27132
rect 83423 27046 83516 27132
rect 83076 26964 83516 27046
rect 83076 26878 83169 26964
rect 83255 26878 83337 26964
rect 83423 26878 83516 26964
rect 83076 26748 83516 26878
rect 87076 28980 87516 29110
rect 87076 28894 87169 28980
rect 87255 28894 87337 28980
rect 87423 28894 87516 28980
rect 87076 28812 87516 28894
rect 87076 28726 87169 28812
rect 87255 28726 87337 28812
rect 87423 28726 87516 28812
rect 87076 28644 87516 28726
rect 87076 28558 87169 28644
rect 87255 28558 87337 28644
rect 87423 28558 87516 28644
rect 87076 28476 87516 28558
rect 87076 28390 87169 28476
rect 87255 28390 87337 28476
rect 87423 28390 87516 28476
rect 87076 28308 87516 28390
rect 87076 28222 87169 28308
rect 87255 28222 87337 28308
rect 87423 28222 87516 28308
rect 87076 28140 87516 28222
rect 87076 28054 87169 28140
rect 87255 28054 87337 28140
rect 87423 28054 87516 28140
rect 87076 27972 87516 28054
rect 87076 27886 87169 27972
rect 87255 27886 87337 27972
rect 87423 27886 87516 27972
rect 87076 27804 87516 27886
rect 87076 27718 87169 27804
rect 87255 27718 87337 27804
rect 87423 27718 87516 27804
rect 87076 27636 87516 27718
rect 87076 27550 87169 27636
rect 87255 27550 87337 27636
rect 87423 27550 87516 27636
rect 87076 27468 87516 27550
rect 87076 27382 87169 27468
rect 87255 27382 87337 27468
rect 87423 27382 87516 27468
rect 87076 27300 87516 27382
rect 87076 27214 87169 27300
rect 87255 27214 87337 27300
rect 87423 27214 87516 27300
rect 87076 27132 87516 27214
rect 87076 27046 87169 27132
rect 87255 27046 87337 27132
rect 87423 27046 87516 27132
rect 87076 26964 87516 27046
rect 87076 26878 87169 26964
rect 87255 26878 87337 26964
rect 87423 26878 87516 26964
rect 87076 26748 87516 26878
rect 91076 28980 91516 29110
rect 91076 28894 91169 28980
rect 91255 28894 91337 28980
rect 91423 28894 91516 28980
rect 91076 28812 91516 28894
rect 91076 28726 91169 28812
rect 91255 28726 91337 28812
rect 91423 28726 91516 28812
rect 91076 28644 91516 28726
rect 91076 28558 91169 28644
rect 91255 28558 91337 28644
rect 91423 28558 91516 28644
rect 91076 28476 91516 28558
rect 91076 28390 91169 28476
rect 91255 28390 91337 28476
rect 91423 28390 91516 28476
rect 91076 28308 91516 28390
rect 91076 28222 91169 28308
rect 91255 28222 91337 28308
rect 91423 28222 91516 28308
rect 91076 28140 91516 28222
rect 91076 28054 91169 28140
rect 91255 28054 91337 28140
rect 91423 28054 91516 28140
rect 91076 27972 91516 28054
rect 91076 27886 91169 27972
rect 91255 27886 91337 27972
rect 91423 27886 91516 27972
rect 91076 27804 91516 27886
rect 91076 27718 91169 27804
rect 91255 27718 91337 27804
rect 91423 27718 91516 27804
rect 91076 27636 91516 27718
rect 91076 27550 91169 27636
rect 91255 27550 91337 27636
rect 91423 27550 91516 27636
rect 91076 27468 91516 27550
rect 91076 27382 91169 27468
rect 91255 27382 91337 27468
rect 91423 27382 91516 27468
rect 91076 27300 91516 27382
rect 91076 27214 91169 27300
rect 91255 27214 91337 27300
rect 91423 27214 91516 27300
rect 91076 27132 91516 27214
rect 91076 27046 91169 27132
rect 91255 27046 91337 27132
rect 91423 27046 91516 27132
rect 91076 26964 91516 27046
rect 91076 26878 91169 26964
rect 91255 26878 91337 26964
rect 91423 26878 91516 26964
rect 91076 26748 91516 26878
rect 95076 28980 95516 29110
rect 95076 28894 95169 28980
rect 95255 28894 95337 28980
rect 95423 28894 95516 28980
rect 95076 28812 95516 28894
rect 95076 28726 95169 28812
rect 95255 28726 95337 28812
rect 95423 28726 95516 28812
rect 95076 28644 95516 28726
rect 95076 28558 95169 28644
rect 95255 28558 95337 28644
rect 95423 28558 95516 28644
rect 95076 28476 95516 28558
rect 95076 28390 95169 28476
rect 95255 28390 95337 28476
rect 95423 28390 95516 28476
rect 95076 28308 95516 28390
rect 95076 28222 95169 28308
rect 95255 28222 95337 28308
rect 95423 28222 95516 28308
rect 95076 28140 95516 28222
rect 95076 28054 95169 28140
rect 95255 28054 95337 28140
rect 95423 28054 95516 28140
rect 95076 27972 95516 28054
rect 95076 27886 95169 27972
rect 95255 27886 95337 27972
rect 95423 27886 95516 27972
rect 95076 27804 95516 27886
rect 95076 27718 95169 27804
rect 95255 27718 95337 27804
rect 95423 27718 95516 27804
rect 95076 27636 95516 27718
rect 95076 27550 95169 27636
rect 95255 27550 95337 27636
rect 95423 27550 95516 27636
rect 95076 27468 95516 27550
rect 95076 27382 95169 27468
rect 95255 27382 95337 27468
rect 95423 27382 95516 27468
rect 95076 27300 95516 27382
rect 95076 27214 95169 27300
rect 95255 27214 95337 27300
rect 95423 27214 95516 27300
rect 95076 27132 95516 27214
rect 95076 27046 95169 27132
rect 95255 27046 95337 27132
rect 95423 27046 95516 27132
rect 95076 26964 95516 27046
rect 95076 26878 95169 26964
rect 95255 26878 95337 26964
rect 95423 26878 95516 26964
rect 95076 26748 95516 26878
rect 73226 26587 73350 26606
rect 73226 26564 73245 26587
rect 71875 26524 71884 26564
rect 71924 26524 73228 26564
rect 4343 26503 4729 26522
rect 4343 26480 4409 26503
rect 4495 26480 4577 26503
rect 4663 26480 4729 26503
rect 4343 26440 4352 26480
rect 4392 26440 4409 26480
rect 4495 26440 4516 26480
rect 4556 26440 4577 26480
rect 4663 26440 4680 26480
rect 4720 26440 4729 26480
rect 4343 26417 4409 26440
rect 4495 26417 4577 26440
rect 4663 26417 4729 26440
rect 4343 26398 4729 26417
rect 8343 26503 8729 26522
rect 8343 26480 8409 26503
rect 8495 26480 8577 26503
rect 8663 26480 8729 26503
rect 8343 26440 8352 26480
rect 8392 26440 8409 26480
rect 8495 26440 8516 26480
rect 8556 26440 8577 26480
rect 8663 26440 8680 26480
rect 8720 26440 8729 26480
rect 8343 26417 8409 26440
rect 8495 26417 8577 26440
rect 8663 26417 8729 26440
rect 8343 26398 8729 26417
rect 12343 26503 12729 26522
rect 12343 26480 12409 26503
rect 12495 26480 12577 26503
rect 12663 26480 12729 26503
rect 12343 26440 12352 26480
rect 12392 26440 12409 26480
rect 12495 26440 12516 26480
rect 12556 26440 12577 26480
rect 12663 26440 12680 26480
rect 12720 26440 12729 26480
rect 12343 26417 12409 26440
rect 12495 26417 12577 26440
rect 12663 26417 12729 26440
rect 12343 26398 12729 26417
rect 16343 26503 16729 26522
rect 16343 26480 16409 26503
rect 16495 26480 16577 26503
rect 16663 26480 16729 26503
rect 16343 26440 16352 26480
rect 16392 26440 16409 26480
rect 16495 26440 16516 26480
rect 16556 26440 16577 26480
rect 16663 26440 16680 26480
rect 16720 26440 16729 26480
rect 16343 26417 16409 26440
rect 16495 26417 16577 26440
rect 16663 26417 16729 26440
rect 16343 26398 16729 26417
rect 20343 26503 20729 26522
rect 20343 26480 20409 26503
rect 20495 26480 20577 26503
rect 20663 26480 20729 26503
rect 20343 26440 20352 26480
rect 20392 26440 20409 26480
rect 20495 26440 20516 26480
rect 20556 26440 20577 26480
rect 20663 26440 20680 26480
rect 20720 26440 20729 26480
rect 20343 26417 20409 26440
rect 20495 26417 20577 26440
rect 20663 26417 20729 26440
rect 20343 26398 20729 26417
rect 24343 26503 24729 26522
rect 24343 26480 24409 26503
rect 24495 26480 24577 26503
rect 24663 26480 24729 26503
rect 24343 26440 24352 26480
rect 24392 26440 24409 26480
rect 24495 26440 24516 26480
rect 24556 26440 24577 26480
rect 24663 26440 24680 26480
rect 24720 26440 24729 26480
rect 24343 26417 24409 26440
rect 24495 26417 24577 26440
rect 24663 26417 24729 26440
rect 24343 26398 24729 26417
rect 28343 26503 28729 26522
rect 28343 26480 28409 26503
rect 28495 26480 28577 26503
rect 28663 26480 28729 26503
rect 28343 26440 28352 26480
rect 28392 26440 28409 26480
rect 28495 26440 28516 26480
rect 28556 26440 28577 26480
rect 28663 26440 28680 26480
rect 28720 26440 28729 26480
rect 28343 26417 28409 26440
rect 28495 26417 28577 26440
rect 28663 26417 28729 26440
rect 28343 26398 28729 26417
rect 32343 26503 32729 26522
rect 32343 26480 32409 26503
rect 32495 26480 32577 26503
rect 32663 26480 32729 26503
rect 32343 26440 32352 26480
rect 32392 26440 32409 26480
rect 32495 26440 32516 26480
rect 32556 26440 32577 26480
rect 32663 26440 32680 26480
rect 32720 26440 32729 26480
rect 32343 26417 32409 26440
rect 32495 26417 32577 26440
rect 32663 26417 32729 26440
rect 32343 26398 32729 26417
rect 36343 26503 36729 26522
rect 36343 26480 36409 26503
rect 36495 26480 36577 26503
rect 36663 26480 36729 26503
rect 36343 26440 36352 26480
rect 36392 26440 36409 26480
rect 36495 26440 36516 26480
rect 36556 26440 36577 26480
rect 36663 26440 36680 26480
rect 36720 26440 36729 26480
rect 36343 26417 36409 26440
rect 36495 26417 36577 26440
rect 36663 26417 36729 26440
rect 36343 26398 36729 26417
rect 40343 26503 40729 26522
rect 40343 26480 40409 26503
rect 40495 26480 40577 26503
rect 40663 26480 40729 26503
rect 40343 26440 40352 26480
rect 40392 26440 40409 26480
rect 40495 26440 40516 26480
rect 40556 26440 40577 26480
rect 40663 26440 40680 26480
rect 40720 26440 40729 26480
rect 40343 26417 40409 26440
rect 40495 26417 40577 26440
rect 40663 26417 40729 26440
rect 40343 26398 40729 26417
rect 44343 26503 44729 26522
rect 44343 26480 44409 26503
rect 44495 26480 44577 26503
rect 44663 26480 44729 26503
rect 44343 26440 44352 26480
rect 44392 26440 44409 26480
rect 44495 26440 44516 26480
rect 44556 26440 44577 26480
rect 44663 26440 44680 26480
rect 44720 26440 44729 26480
rect 44343 26417 44409 26440
rect 44495 26417 44577 26440
rect 44663 26417 44729 26440
rect 44343 26398 44729 26417
rect 48343 26503 48729 26522
rect 48343 26480 48409 26503
rect 48495 26480 48577 26503
rect 48663 26480 48729 26503
rect 48343 26440 48352 26480
rect 48392 26440 48409 26480
rect 48495 26440 48516 26480
rect 48556 26440 48577 26480
rect 48663 26440 48680 26480
rect 48720 26440 48729 26480
rect 48343 26417 48409 26440
rect 48495 26417 48577 26440
rect 48663 26417 48729 26440
rect 48343 26398 48729 26417
rect 52343 26503 52729 26522
rect 52343 26480 52409 26503
rect 52495 26480 52577 26503
rect 52663 26480 52729 26503
rect 52343 26440 52352 26480
rect 52392 26440 52409 26480
rect 52495 26440 52516 26480
rect 52556 26440 52577 26480
rect 52663 26440 52680 26480
rect 52720 26440 52729 26480
rect 52343 26417 52409 26440
rect 52495 26417 52577 26440
rect 52663 26417 52729 26440
rect 52343 26398 52729 26417
rect 56343 26503 56729 26522
rect 56343 26480 56409 26503
rect 56495 26480 56577 26503
rect 56663 26480 56729 26503
rect 56343 26440 56352 26480
rect 56392 26440 56409 26480
rect 56495 26440 56516 26480
rect 56556 26440 56577 26480
rect 56663 26440 56680 26480
rect 56720 26440 56729 26480
rect 56343 26417 56409 26440
rect 56495 26417 56577 26440
rect 56663 26417 56729 26440
rect 56343 26398 56729 26417
rect 60343 26503 60729 26522
rect 60343 26480 60409 26503
rect 60495 26480 60577 26503
rect 60663 26480 60729 26503
rect 60343 26440 60352 26480
rect 60392 26440 60409 26480
rect 60495 26440 60516 26480
rect 60556 26440 60577 26480
rect 60663 26440 60680 26480
rect 60720 26440 60729 26480
rect 60343 26417 60409 26440
rect 60495 26417 60577 26440
rect 60663 26417 60729 26440
rect 60343 26398 60729 26417
rect 64343 26503 64729 26522
rect 64343 26480 64409 26503
rect 64495 26480 64577 26503
rect 64663 26480 64729 26503
rect 64343 26440 64352 26480
rect 64392 26440 64409 26480
rect 64495 26440 64516 26480
rect 64556 26440 64577 26480
rect 64663 26440 64680 26480
rect 64720 26440 64729 26480
rect 64343 26417 64409 26440
rect 64495 26417 64577 26440
rect 64663 26417 64729 26440
rect 64343 26398 64729 26417
rect 68343 26503 68729 26522
rect 68343 26480 68409 26503
rect 68495 26480 68577 26503
rect 68663 26480 68729 26503
rect 73226 26501 73245 26524
rect 73331 26501 73350 26587
rect 73226 26482 73350 26501
rect 68343 26440 68352 26480
rect 68392 26440 68409 26480
rect 68495 26440 68516 26480
rect 68556 26440 68577 26480
rect 68663 26440 68680 26480
rect 68720 26440 68729 26480
rect 68343 26417 68409 26440
rect 68495 26417 68577 26440
rect 68663 26417 68729 26440
rect 68343 26398 68729 26417
rect 3103 25747 3489 25766
rect 3103 25724 3169 25747
rect 3255 25724 3337 25747
rect 3423 25724 3489 25747
rect 3103 25684 3112 25724
rect 3152 25684 3169 25724
rect 3255 25684 3276 25724
rect 3316 25684 3337 25724
rect 3423 25684 3440 25724
rect 3480 25684 3489 25724
rect 3103 25661 3169 25684
rect 3255 25661 3337 25684
rect 3423 25661 3489 25684
rect 3103 25642 3489 25661
rect 7103 25747 7489 25766
rect 7103 25724 7169 25747
rect 7255 25724 7337 25747
rect 7423 25724 7489 25747
rect 7103 25684 7112 25724
rect 7152 25684 7169 25724
rect 7255 25684 7276 25724
rect 7316 25684 7337 25724
rect 7423 25684 7440 25724
rect 7480 25684 7489 25724
rect 7103 25661 7169 25684
rect 7255 25661 7337 25684
rect 7423 25661 7489 25684
rect 7103 25642 7489 25661
rect 11103 25747 11489 25766
rect 11103 25724 11169 25747
rect 11255 25724 11337 25747
rect 11423 25724 11489 25747
rect 11103 25684 11112 25724
rect 11152 25684 11169 25724
rect 11255 25684 11276 25724
rect 11316 25684 11337 25724
rect 11423 25684 11440 25724
rect 11480 25684 11489 25724
rect 11103 25661 11169 25684
rect 11255 25661 11337 25684
rect 11423 25661 11489 25684
rect 11103 25642 11489 25661
rect 15103 25747 15489 25766
rect 15103 25724 15169 25747
rect 15255 25724 15337 25747
rect 15423 25724 15489 25747
rect 15103 25684 15112 25724
rect 15152 25684 15169 25724
rect 15255 25684 15276 25724
rect 15316 25684 15337 25724
rect 15423 25684 15440 25724
rect 15480 25684 15489 25724
rect 15103 25661 15169 25684
rect 15255 25661 15337 25684
rect 15423 25661 15489 25684
rect 15103 25642 15489 25661
rect 19103 25747 19489 25766
rect 19103 25724 19169 25747
rect 19255 25724 19337 25747
rect 19423 25724 19489 25747
rect 19103 25684 19112 25724
rect 19152 25684 19169 25724
rect 19255 25684 19276 25724
rect 19316 25684 19337 25724
rect 19423 25684 19440 25724
rect 19480 25684 19489 25724
rect 19103 25661 19169 25684
rect 19255 25661 19337 25684
rect 19423 25661 19489 25684
rect 19103 25642 19489 25661
rect 23103 25747 23489 25766
rect 23103 25724 23169 25747
rect 23255 25724 23337 25747
rect 23423 25724 23489 25747
rect 23103 25684 23112 25724
rect 23152 25684 23169 25724
rect 23255 25684 23276 25724
rect 23316 25684 23337 25724
rect 23423 25684 23440 25724
rect 23480 25684 23489 25724
rect 23103 25661 23169 25684
rect 23255 25661 23337 25684
rect 23423 25661 23489 25684
rect 23103 25642 23489 25661
rect 27103 25747 27489 25766
rect 27103 25724 27169 25747
rect 27255 25724 27337 25747
rect 27423 25724 27489 25747
rect 27103 25684 27112 25724
rect 27152 25684 27169 25724
rect 27255 25684 27276 25724
rect 27316 25684 27337 25724
rect 27423 25684 27440 25724
rect 27480 25684 27489 25724
rect 27103 25661 27169 25684
rect 27255 25661 27337 25684
rect 27423 25661 27489 25684
rect 27103 25642 27489 25661
rect 31103 25747 31489 25766
rect 31103 25724 31169 25747
rect 31255 25724 31337 25747
rect 31423 25724 31489 25747
rect 31103 25684 31112 25724
rect 31152 25684 31169 25724
rect 31255 25684 31276 25724
rect 31316 25684 31337 25724
rect 31423 25684 31440 25724
rect 31480 25684 31489 25724
rect 31103 25661 31169 25684
rect 31255 25661 31337 25684
rect 31423 25661 31489 25684
rect 31103 25642 31489 25661
rect 35103 25747 35489 25766
rect 35103 25724 35169 25747
rect 35255 25724 35337 25747
rect 35423 25724 35489 25747
rect 35103 25684 35112 25724
rect 35152 25684 35169 25724
rect 35255 25684 35276 25724
rect 35316 25684 35337 25724
rect 35423 25684 35440 25724
rect 35480 25684 35489 25724
rect 35103 25661 35169 25684
rect 35255 25661 35337 25684
rect 35423 25661 35489 25684
rect 35103 25642 35489 25661
rect 39103 25747 39489 25766
rect 39103 25724 39169 25747
rect 39255 25724 39337 25747
rect 39423 25724 39489 25747
rect 39103 25684 39112 25724
rect 39152 25684 39169 25724
rect 39255 25684 39276 25724
rect 39316 25684 39337 25724
rect 39423 25684 39440 25724
rect 39480 25684 39489 25724
rect 39103 25661 39169 25684
rect 39255 25661 39337 25684
rect 39423 25661 39489 25684
rect 39103 25642 39489 25661
rect 43103 25747 43489 25766
rect 43103 25724 43169 25747
rect 43255 25724 43337 25747
rect 43423 25724 43489 25747
rect 43103 25684 43112 25724
rect 43152 25684 43169 25724
rect 43255 25684 43276 25724
rect 43316 25684 43337 25724
rect 43423 25684 43440 25724
rect 43480 25684 43489 25724
rect 43103 25661 43169 25684
rect 43255 25661 43337 25684
rect 43423 25661 43489 25684
rect 43103 25642 43489 25661
rect 47103 25747 47489 25766
rect 47103 25724 47169 25747
rect 47255 25724 47337 25747
rect 47423 25724 47489 25747
rect 47103 25684 47112 25724
rect 47152 25684 47169 25724
rect 47255 25684 47276 25724
rect 47316 25684 47337 25724
rect 47423 25684 47440 25724
rect 47480 25684 47489 25724
rect 47103 25661 47169 25684
rect 47255 25661 47337 25684
rect 47423 25661 47489 25684
rect 47103 25642 47489 25661
rect 51103 25747 51489 25766
rect 51103 25724 51169 25747
rect 51255 25724 51337 25747
rect 51423 25724 51489 25747
rect 51103 25684 51112 25724
rect 51152 25684 51169 25724
rect 51255 25684 51276 25724
rect 51316 25684 51337 25724
rect 51423 25684 51440 25724
rect 51480 25684 51489 25724
rect 51103 25661 51169 25684
rect 51255 25661 51337 25684
rect 51423 25661 51489 25684
rect 51103 25642 51489 25661
rect 55103 25747 55489 25766
rect 55103 25724 55169 25747
rect 55255 25724 55337 25747
rect 55423 25724 55489 25747
rect 55103 25684 55112 25724
rect 55152 25684 55169 25724
rect 55255 25684 55276 25724
rect 55316 25684 55337 25724
rect 55423 25684 55440 25724
rect 55480 25684 55489 25724
rect 55103 25661 55169 25684
rect 55255 25661 55337 25684
rect 55423 25661 55489 25684
rect 55103 25642 55489 25661
rect 59103 25747 59489 25766
rect 59103 25724 59169 25747
rect 59255 25724 59337 25747
rect 59423 25724 59489 25747
rect 59103 25684 59112 25724
rect 59152 25684 59169 25724
rect 59255 25684 59276 25724
rect 59316 25684 59337 25724
rect 59423 25684 59440 25724
rect 59480 25684 59489 25724
rect 59103 25661 59169 25684
rect 59255 25661 59337 25684
rect 59423 25661 59489 25684
rect 59103 25642 59489 25661
rect 63103 25747 63489 25766
rect 63103 25724 63169 25747
rect 63255 25724 63337 25747
rect 63423 25724 63489 25747
rect 63103 25684 63112 25724
rect 63152 25684 63169 25724
rect 63255 25684 63276 25724
rect 63316 25684 63337 25724
rect 63423 25684 63440 25724
rect 63480 25684 63489 25724
rect 63103 25661 63169 25684
rect 63255 25661 63337 25684
rect 63423 25661 63489 25684
rect 63103 25642 63489 25661
rect 67103 25747 67489 25766
rect 67103 25724 67169 25747
rect 67255 25724 67337 25747
rect 67423 25724 67489 25747
rect 67103 25684 67112 25724
rect 67152 25684 67169 25724
rect 67255 25684 67276 25724
rect 67316 25684 67337 25724
rect 67423 25684 67440 25724
rect 67480 25684 67489 25724
rect 67103 25661 67169 25684
rect 67255 25661 67337 25684
rect 67423 25661 67489 25684
rect 67103 25642 67489 25661
rect 86450 25411 86574 25430
rect 86450 25388 86469 25411
rect 85699 25348 85708 25388
rect 85748 25348 86469 25388
rect 86450 25325 86469 25348
rect 86555 25388 86574 25411
rect 86555 25348 86860 25388
rect 86900 25348 86909 25388
rect 86555 25325 86574 25348
rect 86450 25306 86574 25325
rect 4343 24991 4729 25010
rect 4343 24968 4409 24991
rect 4495 24968 4577 24991
rect 4663 24968 4729 24991
rect 4343 24928 4352 24968
rect 4392 24928 4409 24968
rect 4495 24928 4516 24968
rect 4556 24928 4577 24968
rect 4663 24928 4680 24968
rect 4720 24928 4729 24968
rect 4343 24905 4409 24928
rect 4495 24905 4577 24928
rect 4663 24905 4729 24928
rect 4343 24886 4729 24905
rect 8343 24991 8729 25010
rect 8343 24968 8409 24991
rect 8495 24968 8577 24991
rect 8663 24968 8729 24991
rect 8343 24928 8352 24968
rect 8392 24928 8409 24968
rect 8495 24928 8516 24968
rect 8556 24928 8577 24968
rect 8663 24928 8680 24968
rect 8720 24928 8729 24968
rect 8343 24905 8409 24928
rect 8495 24905 8577 24928
rect 8663 24905 8729 24928
rect 8343 24886 8729 24905
rect 12343 24991 12729 25010
rect 12343 24968 12409 24991
rect 12495 24968 12577 24991
rect 12663 24968 12729 24991
rect 12343 24928 12352 24968
rect 12392 24928 12409 24968
rect 12495 24928 12516 24968
rect 12556 24928 12577 24968
rect 12663 24928 12680 24968
rect 12720 24928 12729 24968
rect 12343 24905 12409 24928
rect 12495 24905 12577 24928
rect 12663 24905 12729 24928
rect 12343 24886 12729 24905
rect 16343 24991 16729 25010
rect 16343 24968 16409 24991
rect 16495 24968 16577 24991
rect 16663 24968 16729 24991
rect 16343 24928 16352 24968
rect 16392 24928 16409 24968
rect 16495 24928 16516 24968
rect 16556 24928 16577 24968
rect 16663 24928 16680 24968
rect 16720 24928 16729 24968
rect 16343 24905 16409 24928
rect 16495 24905 16577 24928
rect 16663 24905 16729 24928
rect 16343 24886 16729 24905
rect 20343 24991 20729 25010
rect 20343 24968 20409 24991
rect 20495 24968 20577 24991
rect 20663 24968 20729 24991
rect 20343 24928 20352 24968
rect 20392 24928 20409 24968
rect 20495 24928 20516 24968
rect 20556 24928 20577 24968
rect 20663 24928 20680 24968
rect 20720 24928 20729 24968
rect 20343 24905 20409 24928
rect 20495 24905 20577 24928
rect 20663 24905 20729 24928
rect 20343 24886 20729 24905
rect 24343 24991 24729 25010
rect 24343 24968 24409 24991
rect 24495 24968 24577 24991
rect 24663 24968 24729 24991
rect 24343 24928 24352 24968
rect 24392 24928 24409 24968
rect 24495 24928 24516 24968
rect 24556 24928 24577 24968
rect 24663 24928 24680 24968
rect 24720 24928 24729 24968
rect 24343 24905 24409 24928
rect 24495 24905 24577 24928
rect 24663 24905 24729 24928
rect 24343 24886 24729 24905
rect 28343 24991 28729 25010
rect 28343 24968 28409 24991
rect 28495 24968 28577 24991
rect 28663 24968 28729 24991
rect 28343 24928 28352 24968
rect 28392 24928 28409 24968
rect 28495 24928 28516 24968
rect 28556 24928 28577 24968
rect 28663 24928 28680 24968
rect 28720 24928 28729 24968
rect 28343 24905 28409 24928
rect 28495 24905 28577 24928
rect 28663 24905 28729 24928
rect 28343 24886 28729 24905
rect 32343 24991 32729 25010
rect 32343 24968 32409 24991
rect 32495 24968 32577 24991
rect 32663 24968 32729 24991
rect 32343 24928 32352 24968
rect 32392 24928 32409 24968
rect 32495 24928 32516 24968
rect 32556 24928 32577 24968
rect 32663 24928 32680 24968
rect 32720 24928 32729 24968
rect 32343 24905 32409 24928
rect 32495 24905 32577 24928
rect 32663 24905 32729 24928
rect 32343 24886 32729 24905
rect 36343 24991 36729 25010
rect 36343 24968 36409 24991
rect 36495 24968 36577 24991
rect 36663 24968 36729 24991
rect 36343 24928 36352 24968
rect 36392 24928 36409 24968
rect 36495 24928 36516 24968
rect 36556 24928 36577 24968
rect 36663 24928 36680 24968
rect 36720 24928 36729 24968
rect 36343 24905 36409 24928
rect 36495 24905 36577 24928
rect 36663 24905 36729 24928
rect 36343 24886 36729 24905
rect 40343 24991 40729 25010
rect 40343 24968 40409 24991
rect 40495 24968 40577 24991
rect 40663 24968 40729 24991
rect 40343 24928 40352 24968
rect 40392 24928 40409 24968
rect 40495 24928 40516 24968
rect 40556 24928 40577 24968
rect 40663 24928 40680 24968
rect 40720 24928 40729 24968
rect 40343 24905 40409 24928
rect 40495 24905 40577 24928
rect 40663 24905 40729 24928
rect 40343 24886 40729 24905
rect 44343 24991 44729 25010
rect 44343 24968 44409 24991
rect 44495 24968 44577 24991
rect 44663 24968 44729 24991
rect 44343 24928 44352 24968
rect 44392 24928 44409 24968
rect 44495 24928 44516 24968
rect 44556 24928 44577 24968
rect 44663 24928 44680 24968
rect 44720 24928 44729 24968
rect 44343 24905 44409 24928
rect 44495 24905 44577 24928
rect 44663 24905 44729 24928
rect 44343 24886 44729 24905
rect 48343 24991 48729 25010
rect 48343 24968 48409 24991
rect 48495 24968 48577 24991
rect 48663 24968 48729 24991
rect 48343 24928 48352 24968
rect 48392 24928 48409 24968
rect 48495 24928 48516 24968
rect 48556 24928 48577 24968
rect 48663 24928 48680 24968
rect 48720 24928 48729 24968
rect 48343 24905 48409 24928
rect 48495 24905 48577 24928
rect 48663 24905 48729 24928
rect 48343 24886 48729 24905
rect 52343 24991 52729 25010
rect 52343 24968 52409 24991
rect 52495 24968 52577 24991
rect 52663 24968 52729 24991
rect 52343 24928 52352 24968
rect 52392 24928 52409 24968
rect 52495 24928 52516 24968
rect 52556 24928 52577 24968
rect 52663 24928 52680 24968
rect 52720 24928 52729 24968
rect 52343 24905 52409 24928
rect 52495 24905 52577 24928
rect 52663 24905 52729 24928
rect 52343 24886 52729 24905
rect 56343 24991 56729 25010
rect 56343 24968 56409 24991
rect 56495 24968 56577 24991
rect 56663 24968 56729 24991
rect 56343 24928 56352 24968
rect 56392 24928 56409 24968
rect 56495 24928 56516 24968
rect 56556 24928 56577 24968
rect 56663 24928 56680 24968
rect 56720 24928 56729 24968
rect 56343 24905 56409 24928
rect 56495 24905 56577 24928
rect 56663 24905 56729 24928
rect 56343 24886 56729 24905
rect 60343 24991 60729 25010
rect 60343 24968 60409 24991
rect 60495 24968 60577 24991
rect 60663 24968 60729 24991
rect 60343 24928 60352 24968
rect 60392 24928 60409 24968
rect 60495 24928 60516 24968
rect 60556 24928 60577 24968
rect 60663 24928 60680 24968
rect 60720 24928 60729 24968
rect 60343 24905 60409 24928
rect 60495 24905 60577 24928
rect 60663 24905 60729 24928
rect 60343 24886 60729 24905
rect 64343 24991 64729 25010
rect 64343 24968 64409 24991
rect 64495 24968 64577 24991
rect 64663 24968 64729 24991
rect 64343 24928 64352 24968
rect 64392 24928 64409 24968
rect 64495 24928 64516 24968
rect 64556 24928 64577 24968
rect 64663 24928 64680 24968
rect 64720 24928 64729 24968
rect 64343 24905 64409 24928
rect 64495 24905 64577 24928
rect 64663 24905 64729 24928
rect 64343 24886 64729 24905
rect 68343 24991 68729 25010
rect 68343 24968 68409 24991
rect 68495 24968 68577 24991
rect 68663 24968 68729 24991
rect 68343 24928 68352 24968
rect 68392 24928 68409 24968
rect 68495 24928 68516 24968
rect 68556 24928 68577 24968
rect 68663 24928 68680 24968
rect 68720 24928 68729 24968
rect 68343 24905 68409 24928
rect 68495 24905 68577 24928
rect 68663 24905 68729 24928
rect 68343 24886 68729 24905
rect 3103 24235 3489 24254
rect 3103 24212 3169 24235
rect 3255 24212 3337 24235
rect 3423 24212 3489 24235
rect 3103 24172 3112 24212
rect 3152 24172 3169 24212
rect 3255 24172 3276 24212
rect 3316 24172 3337 24212
rect 3423 24172 3440 24212
rect 3480 24172 3489 24212
rect 3103 24149 3169 24172
rect 3255 24149 3337 24172
rect 3423 24149 3489 24172
rect 3103 24130 3489 24149
rect 7103 24235 7489 24254
rect 7103 24212 7169 24235
rect 7255 24212 7337 24235
rect 7423 24212 7489 24235
rect 7103 24172 7112 24212
rect 7152 24172 7169 24212
rect 7255 24172 7276 24212
rect 7316 24172 7337 24212
rect 7423 24172 7440 24212
rect 7480 24172 7489 24212
rect 7103 24149 7169 24172
rect 7255 24149 7337 24172
rect 7423 24149 7489 24172
rect 7103 24130 7489 24149
rect 11103 24235 11489 24254
rect 11103 24212 11169 24235
rect 11255 24212 11337 24235
rect 11423 24212 11489 24235
rect 11103 24172 11112 24212
rect 11152 24172 11169 24212
rect 11255 24172 11276 24212
rect 11316 24172 11337 24212
rect 11423 24172 11440 24212
rect 11480 24172 11489 24212
rect 11103 24149 11169 24172
rect 11255 24149 11337 24172
rect 11423 24149 11489 24172
rect 11103 24130 11489 24149
rect 15103 24235 15489 24254
rect 15103 24212 15169 24235
rect 15255 24212 15337 24235
rect 15423 24212 15489 24235
rect 15103 24172 15112 24212
rect 15152 24172 15169 24212
rect 15255 24172 15276 24212
rect 15316 24172 15337 24212
rect 15423 24172 15440 24212
rect 15480 24172 15489 24212
rect 15103 24149 15169 24172
rect 15255 24149 15337 24172
rect 15423 24149 15489 24172
rect 15103 24130 15489 24149
rect 19103 24235 19489 24254
rect 19103 24212 19169 24235
rect 19255 24212 19337 24235
rect 19423 24212 19489 24235
rect 19103 24172 19112 24212
rect 19152 24172 19169 24212
rect 19255 24172 19276 24212
rect 19316 24172 19337 24212
rect 19423 24172 19440 24212
rect 19480 24172 19489 24212
rect 19103 24149 19169 24172
rect 19255 24149 19337 24172
rect 19423 24149 19489 24172
rect 19103 24130 19489 24149
rect 23103 24235 23489 24254
rect 23103 24212 23169 24235
rect 23255 24212 23337 24235
rect 23423 24212 23489 24235
rect 23103 24172 23112 24212
rect 23152 24172 23169 24212
rect 23255 24172 23276 24212
rect 23316 24172 23337 24212
rect 23423 24172 23440 24212
rect 23480 24172 23489 24212
rect 23103 24149 23169 24172
rect 23255 24149 23337 24172
rect 23423 24149 23489 24172
rect 23103 24130 23489 24149
rect 27103 24235 27489 24254
rect 27103 24212 27169 24235
rect 27255 24212 27337 24235
rect 27423 24212 27489 24235
rect 27103 24172 27112 24212
rect 27152 24172 27169 24212
rect 27255 24172 27276 24212
rect 27316 24172 27337 24212
rect 27423 24172 27440 24212
rect 27480 24172 27489 24212
rect 27103 24149 27169 24172
rect 27255 24149 27337 24172
rect 27423 24149 27489 24172
rect 27103 24130 27489 24149
rect 31103 24235 31489 24254
rect 31103 24212 31169 24235
rect 31255 24212 31337 24235
rect 31423 24212 31489 24235
rect 31103 24172 31112 24212
rect 31152 24172 31169 24212
rect 31255 24172 31276 24212
rect 31316 24172 31337 24212
rect 31423 24172 31440 24212
rect 31480 24172 31489 24212
rect 31103 24149 31169 24172
rect 31255 24149 31337 24172
rect 31423 24149 31489 24172
rect 31103 24130 31489 24149
rect 35103 24235 35489 24254
rect 35103 24212 35169 24235
rect 35255 24212 35337 24235
rect 35423 24212 35489 24235
rect 35103 24172 35112 24212
rect 35152 24172 35169 24212
rect 35255 24172 35276 24212
rect 35316 24172 35337 24212
rect 35423 24172 35440 24212
rect 35480 24172 35489 24212
rect 35103 24149 35169 24172
rect 35255 24149 35337 24172
rect 35423 24149 35489 24172
rect 35103 24130 35489 24149
rect 39103 24235 39489 24254
rect 39103 24212 39169 24235
rect 39255 24212 39337 24235
rect 39423 24212 39489 24235
rect 39103 24172 39112 24212
rect 39152 24172 39169 24212
rect 39255 24172 39276 24212
rect 39316 24172 39337 24212
rect 39423 24172 39440 24212
rect 39480 24172 39489 24212
rect 39103 24149 39169 24172
rect 39255 24149 39337 24172
rect 39423 24149 39489 24172
rect 39103 24130 39489 24149
rect 43103 24235 43489 24254
rect 43103 24212 43169 24235
rect 43255 24212 43337 24235
rect 43423 24212 43489 24235
rect 43103 24172 43112 24212
rect 43152 24172 43169 24212
rect 43255 24172 43276 24212
rect 43316 24172 43337 24212
rect 43423 24172 43440 24212
rect 43480 24172 43489 24212
rect 43103 24149 43169 24172
rect 43255 24149 43337 24172
rect 43423 24149 43489 24172
rect 43103 24130 43489 24149
rect 47103 24235 47489 24254
rect 47103 24212 47169 24235
rect 47255 24212 47337 24235
rect 47423 24212 47489 24235
rect 47103 24172 47112 24212
rect 47152 24172 47169 24212
rect 47255 24172 47276 24212
rect 47316 24172 47337 24212
rect 47423 24172 47440 24212
rect 47480 24172 47489 24212
rect 47103 24149 47169 24172
rect 47255 24149 47337 24172
rect 47423 24149 47489 24172
rect 47103 24130 47489 24149
rect 51103 24235 51489 24254
rect 51103 24212 51169 24235
rect 51255 24212 51337 24235
rect 51423 24212 51489 24235
rect 51103 24172 51112 24212
rect 51152 24172 51169 24212
rect 51255 24172 51276 24212
rect 51316 24172 51337 24212
rect 51423 24172 51440 24212
rect 51480 24172 51489 24212
rect 51103 24149 51169 24172
rect 51255 24149 51337 24172
rect 51423 24149 51489 24172
rect 51103 24130 51489 24149
rect 55103 24235 55489 24254
rect 55103 24212 55169 24235
rect 55255 24212 55337 24235
rect 55423 24212 55489 24235
rect 55103 24172 55112 24212
rect 55152 24172 55169 24212
rect 55255 24172 55276 24212
rect 55316 24172 55337 24212
rect 55423 24172 55440 24212
rect 55480 24172 55489 24212
rect 55103 24149 55169 24172
rect 55255 24149 55337 24172
rect 55423 24149 55489 24172
rect 55103 24130 55489 24149
rect 59103 24235 59489 24254
rect 59103 24212 59169 24235
rect 59255 24212 59337 24235
rect 59423 24212 59489 24235
rect 59103 24172 59112 24212
rect 59152 24172 59169 24212
rect 59255 24172 59276 24212
rect 59316 24172 59337 24212
rect 59423 24172 59440 24212
rect 59480 24172 59489 24212
rect 59103 24149 59169 24172
rect 59255 24149 59337 24172
rect 59423 24149 59489 24172
rect 59103 24130 59489 24149
rect 63103 24235 63489 24254
rect 63103 24212 63169 24235
rect 63255 24212 63337 24235
rect 63423 24212 63489 24235
rect 63103 24172 63112 24212
rect 63152 24172 63169 24212
rect 63255 24172 63276 24212
rect 63316 24172 63337 24212
rect 63423 24172 63440 24212
rect 63480 24172 63489 24212
rect 63103 24149 63169 24172
rect 63255 24149 63337 24172
rect 63423 24149 63489 24172
rect 63103 24130 63489 24149
rect 67103 24235 67489 24254
rect 67103 24212 67169 24235
rect 67255 24212 67337 24235
rect 67423 24212 67489 24235
rect 67103 24172 67112 24212
rect 67152 24172 67169 24212
rect 67255 24172 67276 24212
rect 67316 24172 67337 24212
rect 67423 24172 67440 24212
rect 67480 24172 67489 24212
rect 67103 24149 67169 24172
rect 67255 24149 67337 24172
rect 67423 24149 67489 24172
rect 67103 24130 67489 24149
rect 71103 24235 71489 24254
rect 71103 24212 71169 24235
rect 71255 24212 71337 24235
rect 71423 24212 71489 24235
rect 71103 24172 71112 24212
rect 71152 24172 71169 24212
rect 71255 24172 71276 24212
rect 71316 24172 71337 24212
rect 71423 24172 71440 24212
rect 71480 24172 71489 24212
rect 71103 24149 71169 24172
rect 71255 24149 71337 24172
rect 71423 24149 71489 24172
rect 71103 24130 71489 24149
rect 75103 24235 75489 24254
rect 75103 24212 75169 24235
rect 75255 24212 75337 24235
rect 75423 24212 75489 24235
rect 75103 24172 75112 24212
rect 75152 24172 75169 24212
rect 75255 24172 75276 24212
rect 75316 24172 75337 24212
rect 75423 24172 75440 24212
rect 75480 24172 75489 24212
rect 75103 24149 75169 24172
rect 75255 24149 75337 24172
rect 75423 24149 75489 24172
rect 75103 24130 75489 24149
rect 79103 24235 79489 24254
rect 79103 24212 79169 24235
rect 79255 24212 79337 24235
rect 79423 24212 79489 24235
rect 79103 24172 79112 24212
rect 79152 24172 79169 24212
rect 79255 24172 79276 24212
rect 79316 24172 79337 24212
rect 79423 24172 79440 24212
rect 79480 24172 79489 24212
rect 79103 24149 79169 24172
rect 79255 24149 79337 24172
rect 79423 24149 79489 24172
rect 79103 24130 79489 24149
rect 83103 24235 83489 24254
rect 83103 24212 83169 24235
rect 83255 24212 83337 24235
rect 83423 24212 83489 24235
rect 83103 24172 83112 24212
rect 83152 24172 83169 24212
rect 83255 24172 83276 24212
rect 83316 24172 83337 24212
rect 83423 24172 83440 24212
rect 83480 24172 83489 24212
rect 83103 24149 83169 24172
rect 83255 24149 83337 24172
rect 83423 24149 83489 24172
rect 83103 24130 83489 24149
rect 87103 24235 87489 24254
rect 87103 24212 87169 24235
rect 87255 24212 87337 24235
rect 87423 24212 87489 24235
rect 87103 24172 87112 24212
rect 87152 24172 87169 24212
rect 87255 24172 87276 24212
rect 87316 24172 87337 24212
rect 87423 24172 87440 24212
rect 87480 24172 87489 24212
rect 87103 24149 87169 24172
rect 87255 24149 87337 24172
rect 87423 24149 87489 24172
rect 87103 24130 87489 24149
rect 91103 24235 91489 24254
rect 91103 24212 91169 24235
rect 91255 24212 91337 24235
rect 91423 24212 91489 24235
rect 91103 24172 91112 24212
rect 91152 24172 91169 24212
rect 91255 24172 91276 24212
rect 91316 24172 91337 24212
rect 91423 24172 91440 24212
rect 91480 24172 91489 24212
rect 91103 24149 91169 24172
rect 91255 24149 91337 24172
rect 91423 24149 91489 24172
rect 91103 24130 91489 24149
rect 95103 24235 95489 24254
rect 95103 24212 95169 24235
rect 95255 24212 95337 24235
rect 95423 24212 95489 24235
rect 95103 24172 95112 24212
rect 95152 24172 95169 24212
rect 95255 24172 95276 24212
rect 95316 24172 95337 24212
rect 95423 24172 95440 24212
rect 95480 24172 95489 24212
rect 95103 24149 95169 24172
rect 95255 24149 95337 24172
rect 95423 24149 95489 24172
rect 95103 24130 95489 24149
rect 99103 24235 99489 24254
rect 99103 24212 99169 24235
rect 99255 24212 99337 24235
rect 99423 24212 99489 24235
rect 99103 24172 99112 24212
rect 99152 24172 99169 24212
rect 99255 24172 99276 24212
rect 99316 24172 99337 24212
rect 99423 24172 99440 24212
rect 99480 24172 99489 24212
rect 99103 24149 99169 24172
rect 99255 24149 99337 24172
rect 99423 24149 99489 24172
rect 99103 24130 99489 24149
rect 4343 23479 4729 23498
rect 4343 23456 4409 23479
rect 4495 23456 4577 23479
rect 4663 23456 4729 23479
rect 4343 23416 4352 23456
rect 4392 23416 4409 23456
rect 4495 23416 4516 23456
rect 4556 23416 4577 23456
rect 4663 23416 4680 23456
rect 4720 23416 4729 23456
rect 4343 23393 4409 23416
rect 4495 23393 4577 23416
rect 4663 23393 4729 23416
rect 4343 23374 4729 23393
rect 8343 23479 8729 23498
rect 8343 23456 8409 23479
rect 8495 23456 8577 23479
rect 8663 23456 8729 23479
rect 8343 23416 8352 23456
rect 8392 23416 8409 23456
rect 8495 23416 8516 23456
rect 8556 23416 8577 23456
rect 8663 23416 8680 23456
rect 8720 23416 8729 23456
rect 8343 23393 8409 23416
rect 8495 23393 8577 23416
rect 8663 23393 8729 23416
rect 8343 23374 8729 23393
rect 12343 23479 12729 23498
rect 12343 23456 12409 23479
rect 12495 23456 12577 23479
rect 12663 23456 12729 23479
rect 12343 23416 12352 23456
rect 12392 23416 12409 23456
rect 12495 23416 12516 23456
rect 12556 23416 12577 23456
rect 12663 23416 12680 23456
rect 12720 23416 12729 23456
rect 12343 23393 12409 23416
rect 12495 23393 12577 23416
rect 12663 23393 12729 23416
rect 12343 23374 12729 23393
rect 16343 23479 16729 23498
rect 16343 23456 16409 23479
rect 16495 23456 16577 23479
rect 16663 23456 16729 23479
rect 16343 23416 16352 23456
rect 16392 23416 16409 23456
rect 16495 23416 16516 23456
rect 16556 23416 16577 23456
rect 16663 23416 16680 23456
rect 16720 23416 16729 23456
rect 16343 23393 16409 23416
rect 16495 23393 16577 23416
rect 16663 23393 16729 23416
rect 16343 23374 16729 23393
rect 20343 23479 20729 23498
rect 20343 23456 20409 23479
rect 20495 23456 20577 23479
rect 20663 23456 20729 23479
rect 20343 23416 20352 23456
rect 20392 23416 20409 23456
rect 20495 23416 20516 23456
rect 20556 23416 20577 23456
rect 20663 23416 20680 23456
rect 20720 23416 20729 23456
rect 20343 23393 20409 23416
rect 20495 23393 20577 23416
rect 20663 23393 20729 23416
rect 20343 23374 20729 23393
rect 24343 23479 24729 23498
rect 24343 23456 24409 23479
rect 24495 23456 24577 23479
rect 24663 23456 24729 23479
rect 24343 23416 24352 23456
rect 24392 23416 24409 23456
rect 24495 23416 24516 23456
rect 24556 23416 24577 23456
rect 24663 23416 24680 23456
rect 24720 23416 24729 23456
rect 24343 23393 24409 23416
rect 24495 23393 24577 23416
rect 24663 23393 24729 23416
rect 24343 23374 24729 23393
rect 28343 23479 28729 23498
rect 28343 23456 28409 23479
rect 28495 23456 28577 23479
rect 28663 23456 28729 23479
rect 28343 23416 28352 23456
rect 28392 23416 28409 23456
rect 28495 23416 28516 23456
rect 28556 23416 28577 23456
rect 28663 23416 28680 23456
rect 28720 23416 28729 23456
rect 28343 23393 28409 23416
rect 28495 23393 28577 23416
rect 28663 23393 28729 23416
rect 28343 23374 28729 23393
rect 32343 23479 32729 23498
rect 32343 23456 32409 23479
rect 32495 23456 32577 23479
rect 32663 23456 32729 23479
rect 32343 23416 32352 23456
rect 32392 23416 32409 23456
rect 32495 23416 32516 23456
rect 32556 23416 32577 23456
rect 32663 23416 32680 23456
rect 32720 23416 32729 23456
rect 32343 23393 32409 23416
rect 32495 23393 32577 23416
rect 32663 23393 32729 23416
rect 32343 23374 32729 23393
rect 36343 23479 36729 23498
rect 36343 23456 36409 23479
rect 36495 23456 36577 23479
rect 36663 23456 36729 23479
rect 36343 23416 36352 23456
rect 36392 23416 36409 23456
rect 36495 23416 36516 23456
rect 36556 23416 36577 23456
rect 36663 23416 36680 23456
rect 36720 23416 36729 23456
rect 36343 23393 36409 23416
rect 36495 23393 36577 23416
rect 36663 23393 36729 23416
rect 36343 23374 36729 23393
rect 40343 23479 40729 23498
rect 40343 23456 40409 23479
rect 40495 23456 40577 23479
rect 40663 23456 40729 23479
rect 40343 23416 40352 23456
rect 40392 23416 40409 23456
rect 40495 23416 40516 23456
rect 40556 23416 40577 23456
rect 40663 23416 40680 23456
rect 40720 23416 40729 23456
rect 40343 23393 40409 23416
rect 40495 23393 40577 23416
rect 40663 23393 40729 23416
rect 40343 23374 40729 23393
rect 44343 23479 44729 23498
rect 44343 23456 44409 23479
rect 44495 23456 44577 23479
rect 44663 23456 44729 23479
rect 44343 23416 44352 23456
rect 44392 23416 44409 23456
rect 44495 23416 44516 23456
rect 44556 23416 44577 23456
rect 44663 23416 44680 23456
rect 44720 23416 44729 23456
rect 44343 23393 44409 23416
rect 44495 23393 44577 23416
rect 44663 23393 44729 23416
rect 44343 23374 44729 23393
rect 48343 23479 48729 23498
rect 48343 23456 48409 23479
rect 48495 23456 48577 23479
rect 48663 23456 48729 23479
rect 48343 23416 48352 23456
rect 48392 23416 48409 23456
rect 48495 23416 48516 23456
rect 48556 23416 48577 23456
rect 48663 23416 48680 23456
rect 48720 23416 48729 23456
rect 48343 23393 48409 23416
rect 48495 23393 48577 23416
rect 48663 23393 48729 23416
rect 48343 23374 48729 23393
rect 52343 23479 52729 23498
rect 52343 23456 52409 23479
rect 52495 23456 52577 23479
rect 52663 23456 52729 23479
rect 52343 23416 52352 23456
rect 52392 23416 52409 23456
rect 52495 23416 52516 23456
rect 52556 23416 52577 23456
rect 52663 23416 52680 23456
rect 52720 23416 52729 23456
rect 52343 23393 52409 23416
rect 52495 23393 52577 23416
rect 52663 23393 52729 23416
rect 52343 23374 52729 23393
rect 56343 23479 56729 23498
rect 56343 23456 56409 23479
rect 56495 23456 56577 23479
rect 56663 23456 56729 23479
rect 56343 23416 56352 23456
rect 56392 23416 56409 23456
rect 56495 23416 56516 23456
rect 56556 23416 56577 23456
rect 56663 23416 56680 23456
rect 56720 23416 56729 23456
rect 56343 23393 56409 23416
rect 56495 23393 56577 23416
rect 56663 23393 56729 23416
rect 56343 23374 56729 23393
rect 60343 23479 60729 23498
rect 60343 23456 60409 23479
rect 60495 23456 60577 23479
rect 60663 23456 60729 23479
rect 60343 23416 60352 23456
rect 60392 23416 60409 23456
rect 60495 23416 60516 23456
rect 60556 23416 60577 23456
rect 60663 23416 60680 23456
rect 60720 23416 60729 23456
rect 60343 23393 60409 23416
rect 60495 23393 60577 23416
rect 60663 23393 60729 23416
rect 60343 23374 60729 23393
rect 64343 23479 64729 23498
rect 64343 23456 64409 23479
rect 64495 23456 64577 23479
rect 64663 23456 64729 23479
rect 64343 23416 64352 23456
rect 64392 23416 64409 23456
rect 64495 23416 64516 23456
rect 64556 23416 64577 23456
rect 64663 23416 64680 23456
rect 64720 23416 64729 23456
rect 64343 23393 64409 23416
rect 64495 23393 64577 23416
rect 64663 23393 64729 23416
rect 64343 23374 64729 23393
rect 68343 23479 68729 23498
rect 68343 23456 68409 23479
rect 68495 23456 68577 23479
rect 68663 23456 68729 23479
rect 68343 23416 68352 23456
rect 68392 23416 68409 23456
rect 68495 23416 68516 23456
rect 68556 23416 68577 23456
rect 68663 23416 68680 23456
rect 68720 23416 68729 23456
rect 68343 23393 68409 23416
rect 68495 23393 68577 23416
rect 68663 23393 68729 23416
rect 68343 23374 68729 23393
rect 72343 23479 72729 23498
rect 72343 23456 72409 23479
rect 72495 23456 72577 23479
rect 72663 23456 72729 23479
rect 72343 23416 72352 23456
rect 72392 23416 72409 23456
rect 72495 23416 72516 23456
rect 72556 23416 72577 23456
rect 72663 23416 72680 23456
rect 72720 23416 72729 23456
rect 72343 23393 72409 23416
rect 72495 23393 72577 23416
rect 72663 23393 72729 23416
rect 72343 23374 72729 23393
rect 76343 23479 76729 23498
rect 76343 23456 76409 23479
rect 76495 23456 76577 23479
rect 76663 23456 76729 23479
rect 76343 23416 76352 23456
rect 76392 23416 76409 23456
rect 76495 23416 76516 23456
rect 76556 23416 76577 23456
rect 76663 23416 76680 23456
rect 76720 23416 76729 23456
rect 76343 23393 76409 23416
rect 76495 23393 76577 23416
rect 76663 23393 76729 23416
rect 76343 23374 76729 23393
rect 80343 23479 80729 23498
rect 80343 23456 80409 23479
rect 80495 23456 80577 23479
rect 80663 23456 80729 23479
rect 80343 23416 80352 23456
rect 80392 23416 80409 23456
rect 80495 23416 80516 23456
rect 80556 23416 80577 23456
rect 80663 23416 80680 23456
rect 80720 23416 80729 23456
rect 80343 23393 80409 23416
rect 80495 23393 80577 23416
rect 80663 23393 80729 23416
rect 80343 23374 80729 23393
rect 84343 23479 84729 23498
rect 84343 23456 84409 23479
rect 84495 23456 84577 23479
rect 84663 23456 84729 23479
rect 84343 23416 84352 23456
rect 84392 23416 84409 23456
rect 84495 23416 84516 23456
rect 84556 23416 84577 23456
rect 84663 23416 84680 23456
rect 84720 23416 84729 23456
rect 84343 23393 84409 23416
rect 84495 23393 84577 23416
rect 84663 23393 84729 23416
rect 84343 23374 84729 23393
rect 88343 23479 88729 23498
rect 88343 23456 88409 23479
rect 88495 23456 88577 23479
rect 88663 23456 88729 23479
rect 88343 23416 88352 23456
rect 88392 23416 88409 23456
rect 88495 23416 88516 23456
rect 88556 23416 88577 23456
rect 88663 23416 88680 23456
rect 88720 23416 88729 23456
rect 88343 23393 88409 23416
rect 88495 23393 88577 23416
rect 88663 23393 88729 23416
rect 88343 23374 88729 23393
rect 92343 23479 92729 23498
rect 92343 23456 92409 23479
rect 92495 23456 92577 23479
rect 92663 23456 92729 23479
rect 92343 23416 92352 23456
rect 92392 23416 92409 23456
rect 92495 23416 92516 23456
rect 92556 23416 92577 23456
rect 92663 23416 92680 23456
rect 92720 23416 92729 23456
rect 92343 23393 92409 23416
rect 92495 23393 92577 23416
rect 92663 23393 92729 23416
rect 92343 23374 92729 23393
rect 96343 23479 96729 23498
rect 96343 23456 96409 23479
rect 96495 23456 96577 23479
rect 96663 23456 96729 23479
rect 96343 23416 96352 23456
rect 96392 23416 96409 23456
rect 96495 23416 96516 23456
rect 96556 23416 96577 23456
rect 96663 23416 96680 23456
rect 96720 23416 96729 23456
rect 96343 23393 96409 23416
rect 96495 23393 96577 23416
rect 96663 23393 96729 23416
rect 96343 23374 96729 23393
rect 3103 22723 3489 22742
rect 3103 22700 3169 22723
rect 3255 22700 3337 22723
rect 3423 22700 3489 22723
rect 3103 22660 3112 22700
rect 3152 22660 3169 22700
rect 3255 22660 3276 22700
rect 3316 22660 3337 22700
rect 3423 22660 3440 22700
rect 3480 22660 3489 22700
rect 3103 22637 3169 22660
rect 3255 22637 3337 22660
rect 3423 22637 3489 22660
rect 3103 22618 3489 22637
rect 7103 22723 7489 22742
rect 7103 22700 7169 22723
rect 7255 22700 7337 22723
rect 7423 22700 7489 22723
rect 7103 22660 7112 22700
rect 7152 22660 7169 22700
rect 7255 22660 7276 22700
rect 7316 22660 7337 22700
rect 7423 22660 7440 22700
rect 7480 22660 7489 22700
rect 7103 22637 7169 22660
rect 7255 22637 7337 22660
rect 7423 22637 7489 22660
rect 7103 22618 7489 22637
rect 11103 22723 11489 22742
rect 11103 22700 11169 22723
rect 11255 22700 11337 22723
rect 11423 22700 11489 22723
rect 11103 22660 11112 22700
rect 11152 22660 11169 22700
rect 11255 22660 11276 22700
rect 11316 22660 11337 22700
rect 11423 22660 11440 22700
rect 11480 22660 11489 22700
rect 11103 22637 11169 22660
rect 11255 22637 11337 22660
rect 11423 22637 11489 22660
rect 11103 22618 11489 22637
rect 15103 22723 15489 22742
rect 15103 22700 15169 22723
rect 15255 22700 15337 22723
rect 15423 22700 15489 22723
rect 15103 22660 15112 22700
rect 15152 22660 15169 22700
rect 15255 22660 15276 22700
rect 15316 22660 15337 22700
rect 15423 22660 15440 22700
rect 15480 22660 15489 22700
rect 15103 22637 15169 22660
rect 15255 22637 15337 22660
rect 15423 22637 15489 22660
rect 15103 22618 15489 22637
rect 19103 22723 19489 22742
rect 19103 22700 19169 22723
rect 19255 22700 19337 22723
rect 19423 22700 19489 22723
rect 19103 22660 19112 22700
rect 19152 22660 19169 22700
rect 19255 22660 19276 22700
rect 19316 22660 19337 22700
rect 19423 22660 19440 22700
rect 19480 22660 19489 22700
rect 19103 22637 19169 22660
rect 19255 22637 19337 22660
rect 19423 22637 19489 22660
rect 19103 22618 19489 22637
rect 23103 22723 23489 22742
rect 23103 22700 23169 22723
rect 23255 22700 23337 22723
rect 23423 22700 23489 22723
rect 23103 22660 23112 22700
rect 23152 22660 23169 22700
rect 23255 22660 23276 22700
rect 23316 22660 23337 22700
rect 23423 22660 23440 22700
rect 23480 22660 23489 22700
rect 23103 22637 23169 22660
rect 23255 22637 23337 22660
rect 23423 22637 23489 22660
rect 23103 22618 23489 22637
rect 27103 22723 27489 22742
rect 27103 22700 27169 22723
rect 27255 22700 27337 22723
rect 27423 22700 27489 22723
rect 27103 22660 27112 22700
rect 27152 22660 27169 22700
rect 27255 22660 27276 22700
rect 27316 22660 27337 22700
rect 27423 22660 27440 22700
rect 27480 22660 27489 22700
rect 27103 22637 27169 22660
rect 27255 22637 27337 22660
rect 27423 22637 27489 22660
rect 27103 22618 27489 22637
rect 31103 22723 31489 22742
rect 31103 22700 31169 22723
rect 31255 22700 31337 22723
rect 31423 22700 31489 22723
rect 31103 22660 31112 22700
rect 31152 22660 31169 22700
rect 31255 22660 31276 22700
rect 31316 22660 31337 22700
rect 31423 22660 31440 22700
rect 31480 22660 31489 22700
rect 31103 22637 31169 22660
rect 31255 22637 31337 22660
rect 31423 22637 31489 22660
rect 31103 22618 31489 22637
rect 35103 22723 35489 22742
rect 35103 22700 35169 22723
rect 35255 22700 35337 22723
rect 35423 22700 35489 22723
rect 35103 22660 35112 22700
rect 35152 22660 35169 22700
rect 35255 22660 35276 22700
rect 35316 22660 35337 22700
rect 35423 22660 35440 22700
rect 35480 22660 35489 22700
rect 35103 22637 35169 22660
rect 35255 22637 35337 22660
rect 35423 22637 35489 22660
rect 35103 22618 35489 22637
rect 39103 22723 39489 22742
rect 39103 22700 39169 22723
rect 39255 22700 39337 22723
rect 39423 22700 39489 22723
rect 39103 22660 39112 22700
rect 39152 22660 39169 22700
rect 39255 22660 39276 22700
rect 39316 22660 39337 22700
rect 39423 22660 39440 22700
rect 39480 22660 39489 22700
rect 39103 22637 39169 22660
rect 39255 22637 39337 22660
rect 39423 22637 39489 22660
rect 39103 22618 39489 22637
rect 43103 22723 43489 22742
rect 43103 22700 43169 22723
rect 43255 22700 43337 22723
rect 43423 22700 43489 22723
rect 43103 22660 43112 22700
rect 43152 22660 43169 22700
rect 43255 22660 43276 22700
rect 43316 22660 43337 22700
rect 43423 22660 43440 22700
rect 43480 22660 43489 22700
rect 43103 22637 43169 22660
rect 43255 22637 43337 22660
rect 43423 22637 43489 22660
rect 43103 22618 43489 22637
rect 47103 22723 47489 22742
rect 47103 22700 47169 22723
rect 47255 22700 47337 22723
rect 47423 22700 47489 22723
rect 47103 22660 47112 22700
rect 47152 22660 47169 22700
rect 47255 22660 47276 22700
rect 47316 22660 47337 22700
rect 47423 22660 47440 22700
rect 47480 22660 47489 22700
rect 47103 22637 47169 22660
rect 47255 22637 47337 22660
rect 47423 22637 47489 22660
rect 47103 22618 47489 22637
rect 51103 22723 51489 22742
rect 51103 22700 51169 22723
rect 51255 22700 51337 22723
rect 51423 22700 51489 22723
rect 51103 22660 51112 22700
rect 51152 22660 51169 22700
rect 51255 22660 51276 22700
rect 51316 22660 51337 22700
rect 51423 22660 51440 22700
rect 51480 22660 51489 22700
rect 51103 22637 51169 22660
rect 51255 22637 51337 22660
rect 51423 22637 51489 22660
rect 51103 22618 51489 22637
rect 55103 22723 55489 22742
rect 55103 22700 55169 22723
rect 55255 22700 55337 22723
rect 55423 22700 55489 22723
rect 55103 22660 55112 22700
rect 55152 22660 55169 22700
rect 55255 22660 55276 22700
rect 55316 22660 55337 22700
rect 55423 22660 55440 22700
rect 55480 22660 55489 22700
rect 55103 22637 55169 22660
rect 55255 22637 55337 22660
rect 55423 22637 55489 22660
rect 55103 22618 55489 22637
rect 59103 22723 59489 22742
rect 59103 22700 59169 22723
rect 59255 22700 59337 22723
rect 59423 22700 59489 22723
rect 59103 22660 59112 22700
rect 59152 22660 59169 22700
rect 59255 22660 59276 22700
rect 59316 22660 59337 22700
rect 59423 22660 59440 22700
rect 59480 22660 59489 22700
rect 59103 22637 59169 22660
rect 59255 22637 59337 22660
rect 59423 22637 59489 22660
rect 59103 22618 59489 22637
rect 63103 22723 63489 22742
rect 63103 22700 63169 22723
rect 63255 22700 63337 22723
rect 63423 22700 63489 22723
rect 63103 22660 63112 22700
rect 63152 22660 63169 22700
rect 63255 22660 63276 22700
rect 63316 22660 63337 22700
rect 63423 22660 63440 22700
rect 63480 22660 63489 22700
rect 63103 22637 63169 22660
rect 63255 22637 63337 22660
rect 63423 22637 63489 22660
rect 63103 22618 63489 22637
rect 67103 22723 67489 22742
rect 67103 22700 67169 22723
rect 67255 22700 67337 22723
rect 67423 22700 67489 22723
rect 67103 22660 67112 22700
rect 67152 22660 67169 22700
rect 67255 22660 67276 22700
rect 67316 22660 67337 22700
rect 67423 22660 67440 22700
rect 67480 22660 67489 22700
rect 67103 22637 67169 22660
rect 67255 22637 67337 22660
rect 67423 22637 67489 22660
rect 67103 22618 67489 22637
rect 71103 22723 71489 22742
rect 71103 22700 71169 22723
rect 71255 22700 71337 22723
rect 71423 22700 71489 22723
rect 71103 22660 71112 22700
rect 71152 22660 71169 22700
rect 71255 22660 71276 22700
rect 71316 22660 71337 22700
rect 71423 22660 71440 22700
rect 71480 22660 71489 22700
rect 71103 22637 71169 22660
rect 71255 22637 71337 22660
rect 71423 22637 71489 22660
rect 71103 22618 71489 22637
rect 75103 22723 75489 22742
rect 75103 22700 75169 22723
rect 75255 22700 75337 22723
rect 75423 22700 75489 22723
rect 75103 22660 75112 22700
rect 75152 22660 75169 22700
rect 75255 22660 75276 22700
rect 75316 22660 75337 22700
rect 75423 22660 75440 22700
rect 75480 22660 75489 22700
rect 75103 22637 75169 22660
rect 75255 22637 75337 22660
rect 75423 22637 75489 22660
rect 75103 22618 75489 22637
rect 79103 22723 79489 22742
rect 79103 22700 79169 22723
rect 79255 22700 79337 22723
rect 79423 22700 79489 22723
rect 79103 22660 79112 22700
rect 79152 22660 79169 22700
rect 79255 22660 79276 22700
rect 79316 22660 79337 22700
rect 79423 22660 79440 22700
rect 79480 22660 79489 22700
rect 79103 22637 79169 22660
rect 79255 22637 79337 22660
rect 79423 22637 79489 22660
rect 79103 22618 79489 22637
rect 83103 22723 83489 22742
rect 83103 22700 83169 22723
rect 83255 22700 83337 22723
rect 83423 22700 83489 22723
rect 83103 22660 83112 22700
rect 83152 22660 83169 22700
rect 83255 22660 83276 22700
rect 83316 22660 83337 22700
rect 83423 22660 83440 22700
rect 83480 22660 83489 22700
rect 83103 22637 83169 22660
rect 83255 22637 83337 22660
rect 83423 22637 83489 22660
rect 83103 22618 83489 22637
rect 87103 22723 87489 22742
rect 87103 22700 87169 22723
rect 87255 22700 87337 22723
rect 87423 22700 87489 22723
rect 87103 22660 87112 22700
rect 87152 22660 87169 22700
rect 87255 22660 87276 22700
rect 87316 22660 87337 22700
rect 87423 22660 87440 22700
rect 87480 22660 87489 22700
rect 87103 22637 87169 22660
rect 87255 22637 87337 22660
rect 87423 22637 87489 22660
rect 87103 22618 87489 22637
rect 91103 22723 91489 22742
rect 91103 22700 91169 22723
rect 91255 22700 91337 22723
rect 91423 22700 91489 22723
rect 91103 22660 91112 22700
rect 91152 22660 91169 22700
rect 91255 22660 91276 22700
rect 91316 22660 91337 22700
rect 91423 22660 91440 22700
rect 91480 22660 91489 22700
rect 91103 22637 91169 22660
rect 91255 22637 91337 22660
rect 91423 22637 91489 22660
rect 91103 22618 91489 22637
rect 95103 22723 95489 22742
rect 95103 22700 95169 22723
rect 95255 22700 95337 22723
rect 95423 22700 95489 22723
rect 95103 22660 95112 22700
rect 95152 22660 95169 22700
rect 95255 22660 95276 22700
rect 95316 22660 95337 22700
rect 95423 22660 95440 22700
rect 95480 22660 95489 22700
rect 95103 22637 95169 22660
rect 95255 22637 95337 22660
rect 95423 22637 95489 22660
rect 95103 22618 95489 22637
rect 99103 22723 99489 22742
rect 99103 22700 99169 22723
rect 99255 22700 99337 22723
rect 99423 22700 99489 22723
rect 99103 22660 99112 22700
rect 99152 22660 99169 22700
rect 99255 22660 99276 22700
rect 99316 22660 99337 22700
rect 99423 22660 99440 22700
rect 99480 22660 99489 22700
rect 99103 22637 99169 22660
rect 99255 22637 99337 22660
rect 99423 22637 99489 22660
rect 99103 22618 99489 22637
rect 4343 21967 4729 21986
rect 4343 21944 4409 21967
rect 4495 21944 4577 21967
rect 4663 21944 4729 21967
rect 4343 21904 4352 21944
rect 4392 21904 4409 21944
rect 4495 21904 4516 21944
rect 4556 21904 4577 21944
rect 4663 21904 4680 21944
rect 4720 21904 4729 21944
rect 4343 21881 4409 21904
rect 4495 21881 4577 21904
rect 4663 21881 4729 21904
rect 4343 21862 4729 21881
rect 8343 21967 8729 21986
rect 8343 21944 8409 21967
rect 8495 21944 8577 21967
rect 8663 21944 8729 21967
rect 8343 21904 8352 21944
rect 8392 21904 8409 21944
rect 8495 21904 8516 21944
rect 8556 21904 8577 21944
rect 8663 21904 8680 21944
rect 8720 21904 8729 21944
rect 8343 21881 8409 21904
rect 8495 21881 8577 21904
rect 8663 21881 8729 21904
rect 8343 21862 8729 21881
rect 12343 21967 12729 21986
rect 12343 21944 12409 21967
rect 12495 21944 12577 21967
rect 12663 21944 12729 21967
rect 12343 21904 12352 21944
rect 12392 21904 12409 21944
rect 12495 21904 12516 21944
rect 12556 21904 12577 21944
rect 12663 21904 12680 21944
rect 12720 21904 12729 21944
rect 12343 21881 12409 21904
rect 12495 21881 12577 21904
rect 12663 21881 12729 21904
rect 12343 21862 12729 21881
rect 16343 21967 16729 21986
rect 16343 21944 16409 21967
rect 16495 21944 16577 21967
rect 16663 21944 16729 21967
rect 16343 21904 16352 21944
rect 16392 21904 16409 21944
rect 16495 21904 16516 21944
rect 16556 21904 16577 21944
rect 16663 21904 16680 21944
rect 16720 21904 16729 21944
rect 16343 21881 16409 21904
rect 16495 21881 16577 21904
rect 16663 21881 16729 21904
rect 16343 21862 16729 21881
rect 20343 21967 20729 21986
rect 20343 21944 20409 21967
rect 20495 21944 20577 21967
rect 20663 21944 20729 21967
rect 20343 21904 20352 21944
rect 20392 21904 20409 21944
rect 20495 21904 20516 21944
rect 20556 21904 20577 21944
rect 20663 21904 20680 21944
rect 20720 21904 20729 21944
rect 20343 21881 20409 21904
rect 20495 21881 20577 21904
rect 20663 21881 20729 21904
rect 20343 21862 20729 21881
rect 24343 21967 24729 21986
rect 24343 21944 24409 21967
rect 24495 21944 24577 21967
rect 24663 21944 24729 21967
rect 24343 21904 24352 21944
rect 24392 21904 24409 21944
rect 24495 21904 24516 21944
rect 24556 21904 24577 21944
rect 24663 21904 24680 21944
rect 24720 21904 24729 21944
rect 24343 21881 24409 21904
rect 24495 21881 24577 21904
rect 24663 21881 24729 21904
rect 24343 21862 24729 21881
rect 28343 21967 28729 21986
rect 28343 21944 28409 21967
rect 28495 21944 28577 21967
rect 28663 21944 28729 21967
rect 28343 21904 28352 21944
rect 28392 21904 28409 21944
rect 28495 21904 28516 21944
rect 28556 21904 28577 21944
rect 28663 21904 28680 21944
rect 28720 21904 28729 21944
rect 28343 21881 28409 21904
rect 28495 21881 28577 21904
rect 28663 21881 28729 21904
rect 28343 21862 28729 21881
rect 32343 21967 32729 21986
rect 32343 21944 32409 21967
rect 32495 21944 32577 21967
rect 32663 21944 32729 21967
rect 32343 21904 32352 21944
rect 32392 21904 32409 21944
rect 32495 21904 32516 21944
rect 32556 21904 32577 21944
rect 32663 21904 32680 21944
rect 32720 21904 32729 21944
rect 32343 21881 32409 21904
rect 32495 21881 32577 21904
rect 32663 21881 32729 21904
rect 32343 21862 32729 21881
rect 36343 21967 36729 21986
rect 36343 21944 36409 21967
rect 36495 21944 36577 21967
rect 36663 21944 36729 21967
rect 36343 21904 36352 21944
rect 36392 21904 36409 21944
rect 36495 21904 36516 21944
rect 36556 21904 36577 21944
rect 36663 21904 36680 21944
rect 36720 21904 36729 21944
rect 36343 21881 36409 21904
rect 36495 21881 36577 21904
rect 36663 21881 36729 21904
rect 36343 21862 36729 21881
rect 40343 21967 40729 21986
rect 40343 21944 40409 21967
rect 40495 21944 40577 21967
rect 40663 21944 40729 21967
rect 40343 21904 40352 21944
rect 40392 21904 40409 21944
rect 40495 21904 40516 21944
rect 40556 21904 40577 21944
rect 40663 21904 40680 21944
rect 40720 21904 40729 21944
rect 40343 21881 40409 21904
rect 40495 21881 40577 21904
rect 40663 21881 40729 21904
rect 40343 21862 40729 21881
rect 44343 21967 44729 21986
rect 44343 21944 44409 21967
rect 44495 21944 44577 21967
rect 44663 21944 44729 21967
rect 44343 21904 44352 21944
rect 44392 21904 44409 21944
rect 44495 21904 44516 21944
rect 44556 21904 44577 21944
rect 44663 21904 44680 21944
rect 44720 21904 44729 21944
rect 44343 21881 44409 21904
rect 44495 21881 44577 21904
rect 44663 21881 44729 21904
rect 44343 21862 44729 21881
rect 48343 21967 48729 21986
rect 48343 21944 48409 21967
rect 48495 21944 48577 21967
rect 48663 21944 48729 21967
rect 48343 21904 48352 21944
rect 48392 21904 48409 21944
rect 48495 21904 48516 21944
rect 48556 21904 48577 21944
rect 48663 21904 48680 21944
rect 48720 21904 48729 21944
rect 48343 21881 48409 21904
rect 48495 21881 48577 21904
rect 48663 21881 48729 21904
rect 48343 21862 48729 21881
rect 52343 21967 52729 21986
rect 52343 21944 52409 21967
rect 52495 21944 52577 21967
rect 52663 21944 52729 21967
rect 52343 21904 52352 21944
rect 52392 21904 52409 21944
rect 52495 21904 52516 21944
rect 52556 21904 52577 21944
rect 52663 21904 52680 21944
rect 52720 21904 52729 21944
rect 52343 21881 52409 21904
rect 52495 21881 52577 21904
rect 52663 21881 52729 21904
rect 52343 21862 52729 21881
rect 56343 21967 56729 21986
rect 56343 21944 56409 21967
rect 56495 21944 56577 21967
rect 56663 21944 56729 21967
rect 56343 21904 56352 21944
rect 56392 21904 56409 21944
rect 56495 21904 56516 21944
rect 56556 21904 56577 21944
rect 56663 21904 56680 21944
rect 56720 21904 56729 21944
rect 56343 21881 56409 21904
rect 56495 21881 56577 21904
rect 56663 21881 56729 21904
rect 56343 21862 56729 21881
rect 60343 21967 60729 21986
rect 60343 21944 60409 21967
rect 60495 21944 60577 21967
rect 60663 21944 60729 21967
rect 60343 21904 60352 21944
rect 60392 21904 60409 21944
rect 60495 21904 60516 21944
rect 60556 21904 60577 21944
rect 60663 21904 60680 21944
rect 60720 21904 60729 21944
rect 60343 21881 60409 21904
rect 60495 21881 60577 21904
rect 60663 21881 60729 21904
rect 60343 21862 60729 21881
rect 64343 21967 64729 21986
rect 64343 21944 64409 21967
rect 64495 21944 64577 21967
rect 64663 21944 64729 21967
rect 64343 21904 64352 21944
rect 64392 21904 64409 21944
rect 64495 21904 64516 21944
rect 64556 21904 64577 21944
rect 64663 21904 64680 21944
rect 64720 21904 64729 21944
rect 64343 21881 64409 21904
rect 64495 21881 64577 21904
rect 64663 21881 64729 21904
rect 64343 21862 64729 21881
rect 68343 21967 68729 21986
rect 68343 21944 68409 21967
rect 68495 21944 68577 21967
rect 68663 21944 68729 21967
rect 68343 21904 68352 21944
rect 68392 21904 68409 21944
rect 68495 21904 68516 21944
rect 68556 21904 68577 21944
rect 68663 21904 68680 21944
rect 68720 21904 68729 21944
rect 68343 21881 68409 21904
rect 68495 21881 68577 21904
rect 68663 21881 68729 21904
rect 68343 21862 68729 21881
rect 72343 21967 72729 21986
rect 72343 21944 72409 21967
rect 72495 21944 72577 21967
rect 72663 21944 72729 21967
rect 72343 21904 72352 21944
rect 72392 21904 72409 21944
rect 72495 21904 72516 21944
rect 72556 21904 72577 21944
rect 72663 21904 72680 21944
rect 72720 21904 72729 21944
rect 72343 21881 72409 21904
rect 72495 21881 72577 21904
rect 72663 21881 72729 21904
rect 72343 21862 72729 21881
rect 76343 21967 76729 21986
rect 76343 21944 76409 21967
rect 76495 21944 76577 21967
rect 76663 21944 76729 21967
rect 76343 21904 76352 21944
rect 76392 21904 76409 21944
rect 76495 21904 76516 21944
rect 76556 21904 76577 21944
rect 76663 21904 76680 21944
rect 76720 21904 76729 21944
rect 76343 21881 76409 21904
rect 76495 21881 76577 21904
rect 76663 21881 76729 21904
rect 76343 21862 76729 21881
rect 80343 21967 80729 21986
rect 80343 21944 80409 21967
rect 80495 21944 80577 21967
rect 80663 21944 80729 21967
rect 80343 21904 80352 21944
rect 80392 21904 80409 21944
rect 80495 21904 80516 21944
rect 80556 21904 80577 21944
rect 80663 21904 80680 21944
rect 80720 21904 80729 21944
rect 80343 21881 80409 21904
rect 80495 21881 80577 21904
rect 80663 21881 80729 21904
rect 80343 21862 80729 21881
rect 84343 21967 84729 21986
rect 84343 21944 84409 21967
rect 84495 21944 84577 21967
rect 84663 21944 84729 21967
rect 84343 21904 84352 21944
rect 84392 21904 84409 21944
rect 84495 21904 84516 21944
rect 84556 21904 84577 21944
rect 84663 21904 84680 21944
rect 84720 21904 84729 21944
rect 84343 21881 84409 21904
rect 84495 21881 84577 21904
rect 84663 21881 84729 21904
rect 84343 21862 84729 21881
rect 88343 21967 88729 21986
rect 88343 21944 88409 21967
rect 88495 21944 88577 21967
rect 88663 21944 88729 21967
rect 88343 21904 88352 21944
rect 88392 21904 88409 21944
rect 88495 21904 88516 21944
rect 88556 21904 88577 21944
rect 88663 21904 88680 21944
rect 88720 21904 88729 21944
rect 88343 21881 88409 21904
rect 88495 21881 88577 21904
rect 88663 21881 88729 21904
rect 88343 21862 88729 21881
rect 92343 21967 92729 21986
rect 92343 21944 92409 21967
rect 92495 21944 92577 21967
rect 92663 21944 92729 21967
rect 92343 21904 92352 21944
rect 92392 21904 92409 21944
rect 92495 21904 92516 21944
rect 92556 21904 92577 21944
rect 92663 21904 92680 21944
rect 92720 21904 92729 21944
rect 92343 21881 92409 21904
rect 92495 21881 92577 21904
rect 92663 21881 92729 21904
rect 92343 21862 92729 21881
rect 96343 21967 96729 21986
rect 96343 21944 96409 21967
rect 96495 21944 96577 21967
rect 96663 21944 96729 21967
rect 96343 21904 96352 21944
rect 96392 21904 96409 21944
rect 96495 21904 96516 21944
rect 96556 21904 96577 21944
rect 96663 21904 96680 21944
rect 96720 21904 96729 21944
rect 96343 21881 96409 21904
rect 96495 21881 96577 21904
rect 96663 21881 96729 21904
rect 96343 21862 96729 21881
rect 3103 21211 3489 21230
rect 3103 21188 3169 21211
rect 3255 21188 3337 21211
rect 3423 21188 3489 21211
rect 3103 21148 3112 21188
rect 3152 21148 3169 21188
rect 3255 21148 3276 21188
rect 3316 21148 3337 21188
rect 3423 21148 3440 21188
rect 3480 21148 3489 21188
rect 3103 21125 3169 21148
rect 3255 21125 3337 21148
rect 3423 21125 3489 21148
rect 3103 21106 3489 21125
rect 7103 21211 7489 21230
rect 7103 21188 7169 21211
rect 7255 21188 7337 21211
rect 7423 21188 7489 21211
rect 7103 21148 7112 21188
rect 7152 21148 7169 21188
rect 7255 21148 7276 21188
rect 7316 21148 7337 21188
rect 7423 21148 7440 21188
rect 7480 21148 7489 21188
rect 7103 21125 7169 21148
rect 7255 21125 7337 21148
rect 7423 21125 7489 21148
rect 7103 21106 7489 21125
rect 11103 21211 11489 21230
rect 11103 21188 11169 21211
rect 11255 21188 11337 21211
rect 11423 21188 11489 21211
rect 11103 21148 11112 21188
rect 11152 21148 11169 21188
rect 11255 21148 11276 21188
rect 11316 21148 11337 21188
rect 11423 21148 11440 21188
rect 11480 21148 11489 21188
rect 11103 21125 11169 21148
rect 11255 21125 11337 21148
rect 11423 21125 11489 21148
rect 11103 21106 11489 21125
rect 15103 21211 15489 21230
rect 15103 21188 15169 21211
rect 15255 21188 15337 21211
rect 15423 21188 15489 21211
rect 15103 21148 15112 21188
rect 15152 21148 15169 21188
rect 15255 21148 15276 21188
rect 15316 21148 15337 21188
rect 15423 21148 15440 21188
rect 15480 21148 15489 21188
rect 15103 21125 15169 21148
rect 15255 21125 15337 21148
rect 15423 21125 15489 21148
rect 15103 21106 15489 21125
rect 19103 21211 19489 21230
rect 19103 21188 19169 21211
rect 19255 21188 19337 21211
rect 19423 21188 19489 21211
rect 19103 21148 19112 21188
rect 19152 21148 19169 21188
rect 19255 21148 19276 21188
rect 19316 21148 19337 21188
rect 19423 21148 19440 21188
rect 19480 21148 19489 21188
rect 19103 21125 19169 21148
rect 19255 21125 19337 21148
rect 19423 21125 19489 21148
rect 19103 21106 19489 21125
rect 23103 21211 23489 21230
rect 23103 21188 23169 21211
rect 23255 21188 23337 21211
rect 23423 21188 23489 21211
rect 23103 21148 23112 21188
rect 23152 21148 23169 21188
rect 23255 21148 23276 21188
rect 23316 21148 23337 21188
rect 23423 21148 23440 21188
rect 23480 21148 23489 21188
rect 23103 21125 23169 21148
rect 23255 21125 23337 21148
rect 23423 21125 23489 21148
rect 23103 21106 23489 21125
rect 27103 21211 27489 21230
rect 27103 21188 27169 21211
rect 27255 21188 27337 21211
rect 27423 21188 27489 21211
rect 27103 21148 27112 21188
rect 27152 21148 27169 21188
rect 27255 21148 27276 21188
rect 27316 21148 27337 21188
rect 27423 21148 27440 21188
rect 27480 21148 27489 21188
rect 27103 21125 27169 21148
rect 27255 21125 27337 21148
rect 27423 21125 27489 21148
rect 27103 21106 27489 21125
rect 31103 21211 31489 21230
rect 31103 21188 31169 21211
rect 31255 21188 31337 21211
rect 31423 21188 31489 21211
rect 31103 21148 31112 21188
rect 31152 21148 31169 21188
rect 31255 21148 31276 21188
rect 31316 21148 31337 21188
rect 31423 21148 31440 21188
rect 31480 21148 31489 21188
rect 31103 21125 31169 21148
rect 31255 21125 31337 21148
rect 31423 21125 31489 21148
rect 31103 21106 31489 21125
rect 35103 21211 35489 21230
rect 35103 21188 35169 21211
rect 35255 21188 35337 21211
rect 35423 21188 35489 21211
rect 35103 21148 35112 21188
rect 35152 21148 35169 21188
rect 35255 21148 35276 21188
rect 35316 21148 35337 21188
rect 35423 21148 35440 21188
rect 35480 21148 35489 21188
rect 35103 21125 35169 21148
rect 35255 21125 35337 21148
rect 35423 21125 35489 21148
rect 35103 21106 35489 21125
rect 39103 21211 39489 21230
rect 39103 21188 39169 21211
rect 39255 21188 39337 21211
rect 39423 21188 39489 21211
rect 39103 21148 39112 21188
rect 39152 21148 39169 21188
rect 39255 21148 39276 21188
rect 39316 21148 39337 21188
rect 39423 21148 39440 21188
rect 39480 21148 39489 21188
rect 39103 21125 39169 21148
rect 39255 21125 39337 21148
rect 39423 21125 39489 21148
rect 39103 21106 39489 21125
rect 43103 21211 43489 21230
rect 43103 21188 43169 21211
rect 43255 21188 43337 21211
rect 43423 21188 43489 21211
rect 43103 21148 43112 21188
rect 43152 21148 43169 21188
rect 43255 21148 43276 21188
rect 43316 21148 43337 21188
rect 43423 21148 43440 21188
rect 43480 21148 43489 21188
rect 43103 21125 43169 21148
rect 43255 21125 43337 21148
rect 43423 21125 43489 21148
rect 43103 21106 43489 21125
rect 47103 21211 47489 21230
rect 47103 21188 47169 21211
rect 47255 21188 47337 21211
rect 47423 21188 47489 21211
rect 47103 21148 47112 21188
rect 47152 21148 47169 21188
rect 47255 21148 47276 21188
rect 47316 21148 47337 21188
rect 47423 21148 47440 21188
rect 47480 21148 47489 21188
rect 47103 21125 47169 21148
rect 47255 21125 47337 21148
rect 47423 21125 47489 21148
rect 47103 21106 47489 21125
rect 51103 21211 51489 21230
rect 51103 21188 51169 21211
rect 51255 21188 51337 21211
rect 51423 21188 51489 21211
rect 51103 21148 51112 21188
rect 51152 21148 51169 21188
rect 51255 21148 51276 21188
rect 51316 21148 51337 21188
rect 51423 21148 51440 21188
rect 51480 21148 51489 21188
rect 51103 21125 51169 21148
rect 51255 21125 51337 21148
rect 51423 21125 51489 21148
rect 51103 21106 51489 21125
rect 55103 21211 55489 21230
rect 55103 21188 55169 21211
rect 55255 21188 55337 21211
rect 55423 21188 55489 21211
rect 55103 21148 55112 21188
rect 55152 21148 55169 21188
rect 55255 21148 55276 21188
rect 55316 21148 55337 21188
rect 55423 21148 55440 21188
rect 55480 21148 55489 21188
rect 55103 21125 55169 21148
rect 55255 21125 55337 21148
rect 55423 21125 55489 21148
rect 55103 21106 55489 21125
rect 59103 21211 59489 21230
rect 59103 21188 59169 21211
rect 59255 21188 59337 21211
rect 59423 21188 59489 21211
rect 59103 21148 59112 21188
rect 59152 21148 59169 21188
rect 59255 21148 59276 21188
rect 59316 21148 59337 21188
rect 59423 21148 59440 21188
rect 59480 21148 59489 21188
rect 59103 21125 59169 21148
rect 59255 21125 59337 21148
rect 59423 21125 59489 21148
rect 59103 21106 59489 21125
rect 63103 21211 63489 21230
rect 63103 21188 63169 21211
rect 63255 21188 63337 21211
rect 63423 21188 63489 21211
rect 63103 21148 63112 21188
rect 63152 21148 63169 21188
rect 63255 21148 63276 21188
rect 63316 21148 63337 21188
rect 63423 21148 63440 21188
rect 63480 21148 63489 21188
rect 63103 21125 63169 21148
rect 63255 21125 63337 21148
rect 63423 21125 63489 21148
rect 63103 21106 63489 21125
rect 67103 21211 67489 21230
rect 67103 21188 67169 21211
rect 67255 21188 67337 21211
rect 67423 21188 67489 21211
rect 67103 21148 67112 21188
rect 67152 21148 67169 21188
rect 67255 21148 67276 21188
rect 67316 21148 67337 21188
rect 67423 21148 67440 21188
rect 67480 21148 67489 21188
rect 67103 21125 67169 21148
rect 67255 21125 67337 21148
rect 67423 21125 67489 21148
rect 67103 21106 67489 21125
rect 71103 21211 71489 21230
rect 71103 21188 71169 21211
rect 71255 21188 71337 21211
rect 71423 21188 71489 21211
rect 71103 21148 71112 21188
rect 71152 21148 71169 21188
rect 71255 21148 71276 21188
rect 71316 21148 71337 21188
rect 71423 21148 71440 21188
rect 71480 21148 71489 21188
rect 71103 21125 71169 21148
rect 71255 21125 71337 21148
rect 71423 21125 71489 21148
rect 71103 21106 71489 21125
rect 75103 21211 75489 21230
rect 75103 21188 75169 21211
rect 75255 21188 75337 21211
rect 75423 21188 75489 21211
rect 75103 21148 75112 21188
rect 75152 21148 75169 21188
rect 75255 21148 75276 21188
rect 75316 21148 75337 21188
rect 75423 21148 75440 21188
rect 75480 21148 75489 21188
rect 75103 21125 75169 21148
rect 75255 21125 75337 21148
rect 75423 21125 75489 21148
rect 75103 21106 75489 21125
rect 79103 21211 79489 21230
rect 79103 21188 79169 21211
rect 79255 21188 79337 21211
rect 79423 21188 79489 21211
rect 79103 21148 79112 21188
rect 79152 21148 79169 21188
rect 79255 21148 79276 21188
rect 79316 21148 79337 21188
rect 79423 21148 79440 21188
rect 79480 21148 79489 21188
rect 79103 21125 79169 21148
rect 79255 21125 79337 21148
rect 79423 21125 79489 21148
rect 79103 21106 79489 21125
rect 83103 21211 83489 21230
rect 83103 21188 83169 21211
rect 83255 21188 83337 21211
rect 83423 21188 83489 21211
rect 83103 21148 83112 21188
rect 83152 21148 83169 21188
rect 83255 21148 83276 21188
rect 83316 21148 83337 21188
rect 83423 21148 83440 21188
rect 83480 21148 83489 21188
rect 83103 21125 83169 21148
rect 83255 21125 83337 21148
rect 83423 21125 83489 21148
rect 83103 21106 83489 21125
rect 87103 21211 87489 21230
rect 87103 21188 87169 21211
rect 87255 21188 87337 21211
rect 87423 21188 87489 21211
rect 87103 21148 87112 21188
rect 87152 21148 87169 21188
rect 87255 21148 87276 21188
rect 87316 21148 87337 21188
rect 87423 21148 87440 21188
rect 87480 21148 87489 21188
rect 87103 21125 87169 21148
rect 87255 21125 87337 21148
rect 87423 21125 87489 21148
rect 87103 21106 87489 21125
rect 91103 21211 91489 21230
rect 91103 21188 91169 21211
rect 91255 21188 91337 21211
rect 91423 21188 91489 21211
rect 91103 21148 91112 21188
rect 91152 21148 91169 21188
rect 91255 21148 91276 21188
rect 91316 21148 91337 21188
rect 91423 21148 91440 21188
rect 91480 21148 91489 21188
rect 91103 21125 91169 21148
rect 91255 21125 91337 21148
rect 91423 21125 91489 21148
rect 91103 21106 91489 21125
rect 95103 21211 95489 21230
rect 95103 21188 95169 21211
rect 95255 21188 95337 21211
rect 95423 21188 95489 21211
rect 95103 21148 95112 21188
rect 95152 21148 95169 21188
rect 95255 21148 95276 21188
rect 95316 21148 95337 21188
rect 95423 21148 95440 21188
rect 95480 21148 95489 21188
rect 95103 21125 95169 21148
rect 95255 21125 95337 21148
rect 95423 21125 95489 21148
rect 95103 21106 95489 21125
rect 99103 21211 99489 21230
rect 99103 21188 99169 21211
rect 99255 21188 99337 21211
rect 99423 21188 99489 21211
rect 99103 21148 99112 21188
rect 99152 21148 99169 21188
rect 99255 21148 99276 21188
rect 99316 21148 99337 21188
rect 99423 21148 99440 21188
rect 99480 21148 99489 21188
rect 99103 21125 99169 21148
rect 99255 21125 99337 21148
rect 99423 21125 99489 21148
rect 99103 21106 99489 21125
rect 4343 20455 4729 20474
rect 4343 20432 4409 20455
rect 4495 20432 4577 20455
rect 4663 20432 4729 20455
rect 4343 20392 4352 20432
rect 4392 20392 4409 20432
rect 4495 20392 4516 20432
rect 4556 20392 4577 20432
rect 4663 20392 4680 20432
rect 4720 20392 4729 20432
rect 4343 20369 4409 20392
rect 4495 20369 4577 20392
rect 4663 20369 4729 20392
rect 4343 20350 4729 20369
rect 8343 20455 8729 20474
rect 8343 20432 8409 20455
rect 8495 20432 8577 20455
rect 8663 20432 8729 20455
rect 8343 20392 8352 20432
rect 8392 20392 8409 20432
rect 8495 20392 8516 20432
rect 8556 20392 8577 20432
rect 8663 20392 8680 20432
rect 8720 20392 8729 20432
rect 8343 20369 8409 20392
rect 8495 20369 8577 20392
rect 8663 20369 8729 20392
rect 8343 20350 8729 20369
rect 12343 20455 12729 20474
rect 12343 20432 12409 20455
rect 12495 20432 12577 20455
rect 12663 20432 12729 20455
rect 12343 20392 12352 20432
rect 12392 20392 12409 20432
rect 12495 20392 12516 20432
rect 12556 20392 12577 20432
rect 12663 20392 12680 20432
rect 12720 20392 12729 20432
rect 12343 20369 12409 20392
rect 12495 20369 12577 20392
rect 12663 20369 12729 20392
rect 12343 20350 12729 20369
rect 16343 20455 16729 20474
rect 16343 20432 16409 20455
rect 16495 20432 16577 20455
rect 16663 20432 16729 20455
rect 16343 20392 16352 20432
rect 16392 20392 16409 20432
rect 16495 20392 16516 20432
rect 16556 20392 16577 20432
rect 16663 20392 16680 20432
rect 16720 20392 16729 20432
rect 16343 20369 16409 20392
rect 16495 20369 16577 20392
rect 16663 20369 16729 20392
rect 16343 20350 16729 20369
rect 20343 20455 20729 20474
rect 20343 20432 20409 20455
rect 20495 20432 20577 20455
rect 20663 20432 20729 20455
rect 20343 20392 20352 20432
rect 20392 20392 20409 20432
rect 20495 20392 20516 20432
rect 20556 20392 20577 20432
rect 20663 20392 20680 20432
rect 20720 20392 20729 20432
rect 20343 20369 20409 20392
rect 20495 20369 20577 20392
rect 20663 20369 20729 20392
rect 20343 20350 20729 20369
rect 24343 20455 24729 20474
rect 24343 20432 24409 20455
rect 24495 20432 24577 20455
rect 24663 20432 24729 20455
rect 24343 20392 24352 20432
rect 24392 20392 24409 20432
rect 24495 20392 24516 20432
rect 24556 20392 24577 20432
rect 24663 20392 24680 20432
rect 24720 20392 24729 20432
rect 24343 20369 24409 20392
rect 24495 20369 24577 20392
rect 24663 20369 24729 20392
rect 24343 20350 24729 20369
rect 28343 20455 28729 20474
rect 28343 20432 28409 20455
rect 28495 20432 28577 20455
rect 28663 20432 28729 20455
rect 28343 20392 28352 20432
rect 28392 20392 28409 20432
rect 28495 20392 28516 20432
rect 28556 20392 28577 20432
rect 28663 20392 28680 20432
rect 28720 20392 28729 20432
rect 28343 20369 28409 20392
rect 28495 20369 28577 20392
rect 28663 20369 28729 20392
rect 28343 20350 28729 20369
rect 32343 20455 32729 20474
rect 32343 20432 32409 20455
rect 32495 20432 32577 20455
rect 32663 20432 32729 20455
rect 32343 20392 32352 20432
rect 32392 20392 32409 20432
rect 32495 20392 32516 20432
rect 32556 20392 32577 20432
rect 32663 20392 32680 20432
rect 32720 20392 32729 20432
rect 32343 20369 32409 20392
rect 32495 20369 32577 20392
rect 32663 20369 32729 20392
rect 32343 20350 32729 20369
rect 36343 20455 36729 20474
rect 36343 20432 36409 20455
rect 36495 20432 36577 20455
rect 36663 20432 36729 20455
rect 36343 20392 36352 20432
rect 36392 20392 36409 20432
rect 36495 20392 36516 20432
rect 36556 20392 36577 20432
rect 36663 20392 36680 20432
rect 36720 20392 36729 20432
rect 36343 20369 36409 20392
rect 36495 20369 36577 20392
rect 36663 20369 36729 20392
rect 36343 20350 36729 20369
rect 40343 20455 40729 20474
rect 40343 20432 40409 20455
rect 40495 20432 40577 20455
rect 40663 20432 40729 20455
rect 40343 20392 40352 20432
rect 40392 20392 40409 20432
rect 40495 20392 40516 20432
rect 40556 20392 40577 20432
rect 40663 20392 40680 20432
rect 40720 20392 40729 20432
rect 40343 20369 40409 20392
rect 40495 20369 40577 20392
rect 40663 20369 40729 20392
rect 40343 20350 40729 20369
rect 44343 20455 44729 20474
rect 44343 20432 44409 20455
rect 44495 20432 44577 20455
rect 44663 20432 44729 20455
rect 44343 20392 44352 20432
rect 44392 20392 44409 20432
rect 44495 20392 44516 20432
rect 44556 20392 44577 20432
rect 44663 20392 44680 20432
rect 44720 20392 44729 20432
rect 44343 20369 44409 20392
rect 44495 20369 44577 20392
rect 44663 20369 44729 20392
rect 44343 20350 44729 20369
rect 48343 20455 48729 20474
rect 48343 20432 48409 20455
rect 48495 20432 48577 20455
rect 48663 20432 48729 20455
rect 48343 20392 48352 20432
rect 48392 20392 48409 20432
rect 48495 20392 48516 20432
rect 48556 20392 48577 20432
rect 48663 20392 48680 20432
rect 48720 20392 48729 20432
rect 48343 20369 48409 20392
rect 48495 20369 48577 20392
rect 48663 20369 48729 20392
rect 48343 20350 48729 20369
rect 52343 20455 52729 20474
rect 52343 20432 52409 20455
rect 52495 20432 52577 20455
rect 52663 20432 52729 20455
rect 52343 20392 52352 20432
rect 52392 20392 52409 20432
rect 52495 20392 52516 20432
rect 52556 20392 52577 20432
rect 52663 20392 52680 20432
rect 52720 20392 52729 20432
rect 52343 20369 52409 20392
rect 52495 20369 52577 20392
rect 52663 20369 52729 20392
rect 52343 20350 52729 20369
rect 56343 20455 56729 20474
rect 56343 20432 56409 20455
rect 56495 20432 56577 20455
rect 56663 20432 56729 20455
rect 56343 20392 56352 20432
rect 56392 20392 56409 20432
rect 56495 20392 56516 20432
rect 56556 20392 56577 20432
rect 56663 20392 56680 20432
rect 56720 20392 56729 20432
rect 56343 20369 56409 20392
rect 56495 20369 56577 20392
rect 56663 20369 56729 20392
rect 56343 20350 56729 20369
rect 60343 20455 60729 20474
rect 60343 20432 60409 20455
rect 60495 20432 60577 20455
rect 60663 20432 60729 20455
rect 60343 20392 60352 20432
rect 60392 20392 60409 20432
rect 60495 20392 60516 20432
rect 60556 20392 60577 20432
rect 60663 20392 60680 20432
rect 60720 20392 60729 20432
rect 60343 20369 60409 20392
rect 60495 20369 60577 20392
rect 60663 20369 60729 20392
rect 60343 20350 60729 20369
rect 64343 20455 64729 20474
rect 64343 20432 64409 20455
rect 64495 20432 64577 20455
rect 64663 20432 64729 20455
rect 64343 20392 64352 20432
rect 64392 20392 64409 20432
rect 64495 20392 64516 20432
rect 64556 20392 64577 20432
rect 64663 20392 64680 20432
rect 64720 20392 64729 20432
rect 64343 20369 64409 20392
rect 64495 20369 64577 20392
rect 64663 20369 64729 20392
rect 64343 20350 64729 20369
rect 68343 20455 68729 20474
rect 68343 20432 68409 20455
rect 68495 20432 68577 20455
rect 68663 20432 68729 20455
rect 68343 20392 68352 20432
rect 68392 20392 68409 20432
rect 68495 20392 68516 20432
rect 68556 20392 68577 20432
rect 68663 20392 68680 20432
rect 68720 20392 68729 20432
rect 68343 20369 68409 20392
rect 68495 20369 68577 20392
rect 68663 20369 68729 20392
rect 68343 20350 68729 20369
rect 72343 20455 72729 20474
rect 72343 20432 72409 20455
rect 72495 20432 72577 20455
rect 72663 20432 72729 20455
rect 72343 20392 72352 20432
rect 72392 20392 72409 20432
rect 72495 20392 72516 20432
rect 72556 20392 72577 20432
rect 72663 20392 72680 20432
rect 72720 20392 72729 20432
rect 72343 20369 72409 20392
rect 72495 20369 72577 20392
rect 72663 20369 72729 20392
rect 72343 20350 72729 20369
rect 76343 20455 76729 20474
rect 76343 20432 76409 20455
rect 76495 20432 76577 20455
rect 76663 20432 76729 20455
rect 76343 20392 76352 20432
rect 76392 20392 76409 20432
rect 76495 20392 76516 20432
rect 76556 20392 76577 20432
rect 76663 20392 76680 20432
rect 76720 20392 76729 20432
rect 76343 20369 76409 20392
rect 76495 20369 76577 20392
rect 76663 20369 76729 20392
rect 76343 20350 76729 20369
rect 80343 20455 80729 20474
rect 80343 20432 80409 20455
rect 80495 20432 80577 20455
rect 80663 20432 80729 20455
rect 80343 20392 80352 20432
rect 80392 20392 80409 20432
rect 80495 20392 80516 20432
rect 80556 20392 80577 20432
rect 80663 20392 80680 20432
rect 80720 20392 80729 20432
rect 80343 20369 80409 20392
rect 80495 20369 80577 20392
rect 80663 20369 80729 20392
rect 80343 20350 80729 20369
rect 84343 20455 84729 20474
rect 84343 20432 84409 20455
rect 84495 20432 84577 20455
rect 84663 20432 84729 20455
rect 84343 20392 84352 20432
rect 84392 20392 84409 20432
rect 84495 20392 84516 20432
rect 84556 20392 84577 20432
rect 84663 20392 84680 20432
rect 84720 20392 84729 20432
rect 84343 20369 84409 20392
rect 84495 20369 84577 20392
rect 84663 20369 84729 20392
rect 84343 20350 84729 20369
rect 88343 20455 88729 20474
rect 88343 20432 88409 20455
rect 88495 20432 88577 20455
rect 88663 20432 88729 20455
rect 88343 20392 88352 20432
rect 88392 20392 88409 20432
rect 88495 20392 88516 20432
rect 88556 20392 88577 20432
rect 88663 20392 88680 20432
rect 88720 20392 88729 20432
rect 88343 20369 88409 20392
rect 88495 20369 88577 20392
rect 88663 20369 88729 20392
rect 88343 20350 88729 20369
rect 92343 20455 92729 20474
rect 92343 20432 92409 20455
rect 92495 20432 92577 20455
rect 92663 20432 92729 20455
rect 92343 20392 92352 20432
rect 92392 20392 92409 20432
rect 92495 20392 92516 20432
rect 92556 20392 92577 20432
rect 92663 20392 92680 20432
rect 92720 20392 92729 20432
rect 92343 20369 92409 20392
rect 92495 20369 92577 20392
rect 92663 20369 92729 20392
rect 92343 20350 92729 20369
rect 96343 20455 96729 20474
rect 96343 20432 96409 20455
rect 96495 20432 96577 20455
rect 96663 20432 96729 20455
rect 96343 20392 96352 20432
rect 96392 20392 96409 20432
rect 96495 20392 96516 20432
rect 96556 20392 96577 20432
rect 96663 20392 96680 20432
rect 96720 20392 96729 20432
rect 96343 20369 96409 20392
rect 96495 20369 96577 20392
rect 96663 20369 96729 20392
rect 96343 20350 96729 20369
rect 3103 19699 3489 19718
rect 3103 19676 3169 19699
rect 3255 19676 3337 19699
rect 3423 19676 3489 19699
rect 3103 19636 3112 19676
rect 3152 19636 3169 19676
rect 3255 19636 3276 19676
rect 3316 19636 3337 19676
rect 3423 19636 3440 19676
rect 3480 19636 3489 19676
rect 3103 19613 3169 19636
rect 3255 19613 3337 19636
rect 3423 19613 3489 19636
rect 3103 19594 3489 19613
rect 7103 19699 7489 19718
rect 7103 19676 7169 19699
rect 7255 19676 7337 19699
rect 7423 19676 7489 19699
rect 7103 19636 7112 19676
rect 7152 19636 7169 19676
rect 7255 19636 7276 19676
rect 7316 19636 7337 19676
rect 7423 19636 7440 19676
rect 7480 19636 7489 19676
rect 7103 19613 7169 19636
rect 7255 19613 7337 19636
rect 7423 19613 7489 19636
rect 7103 19594 7489 19613
rect 11103 19699 11489 19718
rect 11103 19676 11169 19699
rect 11255 19676 11337 19699
rect 11423 19676 11489 19699
rect 11103 19636 11112 19676
rect 11152 19636 11169 19676
rect 11255 19636 11276 19676
rect 11316 19636 11337 19676
rect 11423 19636 11440 19676
rect 11480 19636 11489 19676
rect 11103 19613 11169 19636
rect 11255 19613 11337 19636
rect 11423 19613 11489 19636
rect 11103 19594 11489 19613
rect 15103 19699 15489 19718
rect 15103 19676 15169 19699
rect 15255 19676 15337 19699
rect 15423 19676 15489 19699
rect 15103 19636 15112 19676
rect 15152 19636 15169 19676
rect 15255 19636 15276 19676
rect 15316 19636 15337 19676
rect 15423 19636 15440 19676
rect 15480 19636 15489 19676
rect 15103 19613 15169 19636
rect 15255 19613 15337 19636
rect 15423 19613 15489 19636
rect 15103 19594 15489 19613
rect 19103 19699 19489 19718
rect 19103 19676 19169 19699
rect 19255 19676 19337 19699
rect 19423 19676 19489 19699
rect 19103 19636 19112 19676
rect 19152 19636 19169 19676
rect 19255 19636 19276 19676
rect 19316 19636 19337 19676
rect 19423 19636 19440 19676
rect 19480 19636 19489 19676
rect 19103 19613 19169 19636
rect 19255 19613 19337 19636
rect 19423 19613 19489 19636
rect 19103 19594 19489 19613
rect 23103 19699 23489 19718
rect 23103 19676 23169 19699
rect 23255 19676 23337 19699
rect 23423 19676 23489 19699
rect 23103 19636 23112 19676
rect 23152 19636 23169 19676
rect 23255 19636 23276 19676
rect 23316 19636 23337 19676
rect 23423 19636 23440 19676
rect 23480 19636 23489 19676
rect 23103 19613 23169 19636
rect 23255 19613 23337 19636
rect 23423 19613 23489 19636
rect 23103 19594 23489 19613
rect 27103 19699 27489 19718
rect 27103 19676 27169 19699
rect 27255 19676 27337 19699
rect 27423 19676 27489 19699
rect 27103 19636 27112 19676
rect 27152 19636 27169 19676
rect 27255 19636 27276 19676
rect 27316 19636 27337 19676
rect 27423 19636 27440 19676
rect 27480 19636 27489 19676
rect 27103 19613 27169 19636
rect 27255 19613 27337 19636
rect 27423 19613 27489 19636
rect 27103 19594 27489 19613
rect 31103 19699 31489 19718
rect 31103 19676 31169 19699
rect 31255 19676 31337 19699
rect 31423 19676 31489 19699
rect 31103 19636 31112 19676
rect 31152 19636 31169 19676
rect 31255 19636 31276 19676
rect 31316 19636 31337 19676
rect 31423 19636 31440 19676
rect 31480 19636 31489 19676
rect 31103 19613 31169 19636
rect 31255 19613 31337 19636
rect 31423 19613 31489 19636
rect 31103 19594 31489 19613
rect 35103 19699 35489 19718
rect 35103 19676 35169 19699
rect 35255 19676 35337 19699
rect 35423 19676 35489 19699
rect 35103 19636 35112 19676
rect 35152 19636 35169 19676
rect 35255 19636 35276 19676
rect 35316 19636 35337 19676
rect 35423 19636 35440 19676
rect 35480 19636 35489 19676
rect 35103 19613 35169 19636
rect 35255 19613 35337 19636
rect 35423 19613 35489 19636
rect 35103 19594 35489 19613
rect 39103 19699 39489 19718
rect 39103 19676 39169 19699
rect 39255 19676 39337 19699
rect 39423 19676 39489 19699
rect 39103 19636 39112 19676
rect 39152 19636 39169 19676
rect 39255 19636 39276 19676
rect 39316 19636 39337 19676
rect 39423 19636 39440 19676
rect 39480 19636 39489 19676
rect 39103 19613 39169 19636
rect 39255 19613 39337 19636
rect 39423 19613 39489 19636
rect 39103 19594 39489 19613
rect 43103 19699 43489 19718
rect 43103 19676 43169 19699
rect 43255 19676 43337 19699
rect 43423 19676 43489 19699
rect 43103 19636 43112 19676
rect 43152 19636 43169 19676
rect 43255 19636 43276 19676
rect 43316 19636 43337 19676
rect 43423 19636 43440 19676
rect 43480 19636 43489 19676
rect 43103 19613 43169 19636
rect 43255 19613 43337 19636
rect 43423 19613 43489 19636
rect 43103 19594 43489 19613
rect 47103 19699 47489 19718
rect 47103 19676 47169 19699
rect 47255 19676 47337 19699
rect 47423 19676 47489 19699
rect 47103 19636 47112 19676
rect 47152 19636 47169 19676
rect 47255 19636 47276 19676
rect 47316 19636 47337 19676
rect 47423 19636 47440 19676
rect 47480 19636 47489 19676
rect 47103 19613 47169 19636
rect 47255 19613 47337 19636
rect 47423 19613 47489 19636
rect 47103 19594 47489 19613
rect 51103 19699 51489 19718
rect 51103 19676 51169 19699
rect 51255 19676 51337 19699
rect 51423 19676 51489 19699
rect 51103 19636 51112 19676
rect 51152 19636 51169 19676
rect 51255 19636 51276 19676
rect 51316 19636 51337 19676
rect 51423 19636 51440 19676
rect 51480 19636 51489 19676
rect 51103 19613 51169 19636
rect 51255 19613 51337 19636
rect 51423 19613 51489 19636
rect 51103 19594 51489 19613
rect 55103 19699 55489 19718
rect 55103 19676 55169 19699
rect 55255 19676 55337 19699
rect 55423 19676 55489 19699
rect 55103 19636 55112 19676
rect 55152 19636 55169 19676
rect 55255 19636 55276 19676
rect 55316 19636 55337 19676
rect 55423 19636 55440 19676
rect 55480 19636 55489 19676
rect 55103 19613 55169 19636
rect 55255 19613 55337 19636
rect 55423 19613 55489 19636
rect 55103 19594 55489 19613
rect 59103 19699 59489 19718
rect 59103 19676 59169 19699
rect 59255 19676 59337 19699
rect 59423 19676 59489 19699
rect 59103 19636 59112 19676
rect 59152 19636 59169 19676
rect 59255 19636 59276 19676
rect 59316 19636 59337 19676
rect 59423 19636 59440 19676
rect 59480 19636 59489 19676
rect 59103 19613 59169 19636
rect 59255 19613 59337 19636
rect 59423 19613 59489 19636
rect 59103 19594 59489 19613
rect 63103 19699 63489 19718
rect 63103 19676 63169 19699
rect 63255 19676 63337 19699
rect 63423 19676 63489 19699
rect 63103 19636 63112 19676
rect 63152 19636 63169 19676
rect 63255 19636 63276 19676
rect 63316 19636 63337 19676
rect 63423 19636 63440 19676
rect 63480 19636 63489 19676
rect 63103 19613 63169 19636
rect 63255 19613 63337 19636
rect 63423 19613 63489 19636
rect 63103 19594 63489 19613
rect 67103 19699 67489 19718
rect 67103 19676 67169 19699
rect 67255 19676 67337 19699
rect 67423 19676 67489 19699
rect 67103 19636 67112 19676
rect 67152 19636 67169 19676
rect 67255 19636 67276 19676
rect 67316 19636 67337 19676
rect 67423 19636 67440 19676
rect 67480 19636 67489 19676
rect 67103 19613 67169 19636
rect 67255 19613 67337 19636
rect 67423 19613 67489 19636
rect 67103 19594 67489 19613
rect 71103 19699 71489 19718
rect 71103 19676 71169 19699
rect 71255 19676 71337 19699
rect 71423 19676 71489 19699
rect 71103 19636 71112 19676
rect 71152 19636 71169 19676
rect 71255 19636 71276 19676
rect 71316 19636 71337 19676
rect 71423 19636 71440 19676
rect 71480 19636 71489 19676
rect 71103 19613 71169 19636
rect 71255 19613 71337 19636
rect 71423 19613 71489 19636
rect 71103 19594 71489 19613
rect 75103 19699 75489 19718
rect 75103 19676 75169 19699
rect 75255 19676 75337 19699
rect 75423 19676 75489 19699
rect 75103 19636 75112 19676
rect 75152 19636 75169 19676
rect 75255 19636 75276 19676
rect 75316 19636 75337 19676
rect 75423 19636 75440 19676
rect 75480 19636 75489 19676
rect 75103 19613 75169 19636
rect 75255 19613 75337 19636
rect 75423 19613 75489 19636
rect 75103 19594 75489 19613
rect 79103 19699 79489 19718
rect 79103 19676 79169 19699
rect 79255 19676 79337 19699
rect 79423 19676 79489 19699
rect 79103 19636 79112 19676
rect 79152 19636 79169 19676
rect 79255 19636 79276 19676
rect 79316 19636 79337 19676
rect 79423 19636 79440 19676
rect 79480 19636 79489 19676
rect 79103 19613 79169 19636
rect 79255 19613 79337 19636
rect 79423 19613 79489 19636
rect 79103 19594 79489 19613
rect 83103 19699 83489 19718
rect 83103 19676 83169 19699
rect 83255 19676 83337 19699
rect 83423 19676 83489 19699
rect 83103 19636 83112 19676
rect 83152 19636 83169 19676
rect 83255 19636 83276 19676
rect 83316 19636 83337 19676
rect 83423 19636 83440 19676
rect 83480 19636 83489 19676
rect 83103 19613 83169 19636
rect 83255 19613 83337 19636
rect 83423 19613 83489 19636
rect 83103 19594 83489 19613
rect 87103 19699 87489 19718
rect 87103 19676 87169 19699
rect 87255 19676 87337 19699
rect 87423 19676 87489 19699
rect 87103 19636 87112 19676
rect 87152 19636 87169 19676
rect 87255 19636 87276 19676
rect 87316 19636 87337 19676
rect 87423 19636 87440 19676
rect 87480 19636 87489 19676
rect 87103 19613 87169 19636
rect 87255 19613 87337 19636
rect 87423 19613 87489 19636
rect 87103 19594 87489 19613
rect 91103 19699 91489 19718
rect 91103 19676 91169 19699
rect 91255 19676 91337 19699
rect 91423 19676 91489 19699
rect 91103 19636 91112 19676
rect 91152 19636 91169 19676
rect 91255 19636 91276 19676
rect 91316 19636 91337 19676
rect 91423 19636 91440 19676
rect 91480 19636 91489 19676
rect 91103 19613 91169 19636
rect 91255 19613 91337 19636
rect 91423 19613 91489 19636
rect 91103 19594 91489 19613
rect 95103 19699 95489 19718
rect 95103 19676 95169 19699
rect 95255 19676 95337 19699
rect 95423 19676 95489 19699
rect 95103 19636 95112 19676
rect 95152 19636 95169 19676
rect 95255 19636 95276 19676
rect 95316 19636 95337 19676
rect 95423 19636 95440 19676
rect 95480 19636 95489 19676
rect 95103 19613 95169 19636
rect 95255 19613 95337 19636
rect 95423 19613 95489 19636
rect 95103 19594 95489 19613
rect 99103 19699 99489 19718
rect 99103 19676 99169 19699
rect 99255 19676 99337 19699
rect 99423 19676 99489 19699
rect 99103 19636 99112 19676
rect 99152 19636 99169 19676
rect 99255 19636 99276 19676
rect 99316 19636 99337 19676
rect 99423 19636 99440 19676
rect 99480 19636 99489 19676
rect 99103 19613 99169 19636
rect 99255 19613 99337 19636
rect 99423 19613 99489 19636
rect 99103 19594 99489 19613
rect 4343 18943 4729 18962
rect 4343 18920 4409 18943
rect 4495 18920 4577 18943
rect 4663 18920 4729 18943
rect 4343 18880 4352 18920
rect 4392 18880 4409 18920
rect 4495 18880 4516 18920
rect 4556 18880 4577 18920
rect 4663 18880 4680 18920
rect 4720 18880 4729 18920
rect 4343 18857 4409 18880
rect 4495 18857 4577 18880
rect 4663 18857 4729 18880
rect 4343 18838 4729 18857
rect 8343 18943 8729 18962
rect 8343 18920 8409 18943
rect 8495 18920 8577 18943
rect 8663 18920 8729 18943
rect 8343 18880 8352 18920
rect 8392 18880 8409 18920
rect 8495 18880 8516 18920
rect 8556 18880 8577 18920
rect 8663 18880 8680 18920
rect 8720 18880 8729 18920
rect 8343 18857 8409 18880
rect 8495 18857 8577 18880
rect 8663 18857 8729 18880
rect 8343 18838 8729 18857
rect 12343 18943 12729 18962
rect 12343 18920 12409 18943
rect 12495 18920 12577 18943
rect 12663 18920 12729 18943
rect 12343 18880 12352 18920
rect 12392 18880 12409 18920
rect 12495 18880 12516 18920
rect 12556 18880 12577 18920
rect 12663 18880 12680 18920
rect 12720 18880 12729 18920
rect 12343 18857 12409 18880
rect 12495 18857 12577 18880
rect 12663 18857 12729 18880
rect 12343 18838 12729 18857
rect 16343 18943 16729 18962
rect 16343 18920 16409 18943
rect 16495 18920 16577 18943
rect 16663 18920 16729 18943
rect 16343 18880 16352 18920
rect 16392 18880 16409 18920
rect 16495 18880 16516 18920
rect 16556 18880 16577 18920
rect 16663 18880 16680 18920
rect 16720 18880 16729 18920
rect 16343 18857 16409 18880
rect 16495 18857 16577 18880
rect 16663 18857 16729 18880
rect 16343 18838 16729 18857
rect 20343 18943 20729 18962
rect 20343 18920 20409 18943
rect 20495 18920 20577 18943
rect 20663 18920 20729 18943
rect 20343 18880 20352 18920
rect 20392 18880 20409 18920
rect 20495 18880 20516 18920
rect 20556 18880 20577 18920
rect 20663 18880 20680 18920
rect 20720 18880 20729 18920
rect 20343 18857 20409 18880
rect 20495 18857 20577 18880
rect 20663 18857 20729 18880
rect 20343 18838 20729 18857
rect 24343 18943 24729 18962
rect 24343 18920 24409 18943
rect 24495 18920 24577 18943
rect 24663 18920 24729 18943
rect 24343 18880 24352 18920
rect 24392 18880 24409 18920
rect 24495 18880 24516 18920
rect 24556 18880 24577 18920
rect 24663 18880 24680 18920
rect 24720 18880 24729 18920
rect 24343 18857 24409 18880
rect 24495 18857 24577 18880
rect 24663 18857 24729 18880
rect 24343 18838 24729 18857
rect 28343 18943 28729 18962
rect 28343 18920 28409 18943
rect 28495 18920 28577 18943
rect 28663 18920 28729 18943
rect 28343 18880 28352 18920
rect 28392 18880 28409 18920
rect 28495 18880 28516 18920
rect 28556 18880 28577 18920
rect 28663 18880 28680 18920
rect 28720 18880 28729 18920
rect 28343 18857 28409 18880
rect 28495 18857 28577 18880
rect 28663 18857 28729 18880
rect 28343 18838 28729 18857
rect 32343 18943 32729 18962
rect 32343 18920 32409 18943
rect 32495 18920 32577 18943
rect 32663 18920 32729 18943
rect 32343 18880 32352 18920
rect 32392 18880 32409 18920
rect 32495 18880 32516 18920
rect 32556 18880 32577 18920
rect 32663 18880 32680 18920
rect 32720 18880 32729 18920
rect 32343 18857 32409 18880
rect 32495 18857 32577 18880
rect 32663 18857 32729 18880
rect 32343 18838 32729 18857
rect 36343 18943 36729 18962
rect 36343 18920 36409 18943
rect 36495 18920 36577 18943
rect 36663 18920 36729 18943
rect 36343 18880 36352 18920
rect 36392 18880 36409 18920
rect 36495 18880 36516 18920
rect 36556 18880 36577 18920
rect 36663 18880 36680 18920
rect 36720 18880 36729 18920
rect 36343 18857 36409 18880
rect 36495 18857 36577 18880
rect 36663 18857 36729 18880
rect 36343 18838 36729 18857
rect 40343 18943 40729 18962
rect 40343 18920 40409 18943
rect 40495 18920 40577 18943
rect 40663 18920 40729 18943
rect 40343 18880 40352 18920
rect 40392 18880 40409 18920
rect 40495 18880 40516 18920
rect 40556 18880 40577 18920
rect 40663 18880 40680 18920
rect 40720 18880 40729 18920
rect 40343 18857 40409 18880
rect 40495 18857 40577 18880
rect 40663 18857 40729 18880
rect 40343 18838 40729 18857
rect 44343 18943 44729 18962
rect 44343 18920 44409 18943
rect 44495 18920 44577 18943
rect 44663 18920 44729 18943
rect 44343 18880 44352 18920
rect 44392 18880 44409 18920
rect 44495 18880 44516 18920
rect 44556 18880 44577 18920
rect 44663 18880 44680 18920
rect 44720 18880 44729 18920
rect 44343 18857 44409 18880
rect 44495 18857 44577 18880
rect 44663 18857 44729 18880
rect 44343 18838 44729 18857
rect 48343 18943 48729 18962
rect 48343 18920 48409 18943
rect 48495 18920 48577 18943
rect 48663 18920 48729 18943
rect 48343 18880 48352 18920
rect 48392 18880 48409 18920
rect 48495 18880 48516 18920
rect 48556 18880 48577 18920
rect 48663 18880 48680 18920
rect 48720 18880 48729 18920
rect 48343 18857 48409 18880
rect 48495 18857 48577 18880
rect 48663 18857 48729 18880
rect 48343 18838 48729 18857
rect 52343 18943 52729 18962
rect 52343 18920 52409 18943
rect 52495 18920 52577 18943
rect 52663 18920 52729 18943
rect 52343 18880 52352 18920
rect 52392 18880 52409 18920
rect 52495 18880 52516 18920
rect 52556 18880 52577 18920
rect 52663 18880 52680 18920
rect 52720 18880 52729 18920
rect 52343 18857 52409 18880
rect 52495 18857 52577 18880
rect 52663 18857 52729 18880
rect 52343 18838 52729 18857
rect 56343 18943 56729 18962
rect 56343 18920 56409 18943
rect 56495 18920 56577 18943
rect 56663 18920 56729 18943
rect 56343 18880 56352 18920
rect 56392 18880 56409 18920
rect 56495 18880 56516 18920
rect 56556 18880 56577 18920
rect 56663 18880 56680 18920
rect 56720 18880 56729 18920
rect 56343 18857 56409 18880
rect 56495 18857 56577 18880
rect 56663 18857 56729 18880
rect 56343 18838 56729 18857
rect 60343 18943 60729 18962
rect 60343 18920 60409 18943
rect 60495 18920 60577 18943
rect 60663 18920 60729 18943
rect 60343 18880 60352 18920
rect 60392 18880 60409 18920
rect 60495 18880 60516 18920
rect 60556 18880 60577 18920
rect 60663 18880 60680 18920
rect 60720 18880 60729 18920
rect 60343 18857 60409 18880
rect 60495 18857 60577 18880
rect 60663 18857 60729 18880
rect 60343 18838 60729 18857
rect 64343 18943 64729 18962
rect 64343 18920 64409 18943
rect 64495 18920 64577 18943
rect 64663 18920 64729 18943
rect 64343 18880 64352 18920
rect 64392 18880 64409 18920
rect 64495 18880 64516 18920
rect 64556 18880 64577 18920
rect 64663 18880 64680 18920
rect 64720 18880 64729 18920
rect 64343 18857 64409 18880
rect 64495 18857 64577 18880
rect 64663 18857 64729 18880
rect 64343 18838 64729 18857
rect 68343 18943 68729 18962
rect 68343 18920 68409 18943
rect 68495 18920 68577 18943
rect 68663 18920 68729 18943
rect 68343 18880 68352 18920
rect 68392 18880 68409 18920
rect 68495 18880 68516 18920
rect 68556 18880 68577 18920
rect 68663 18880 68680 18920
rect 68720 18880 68729 18920
rect 68343 18857 68409 18880
rect 68495 18857 68577 18880
rect 68663 18857 68729 18880
rect 68343 18838 68729 18857
rect 72343 18943 72729 18962
rect 72343 18920 72409 18943
rect 72495 18920 72577 18943
rect 72663 18920 72729 18943
rect 72343 18880 72352 18920
rect 72392 18880 72409 18920
rect 72495 18880 72516 18920
rect 72556 18880 72577 18920
rect 72663 18880 72680 18920
rect 72720 18880 72729 18920
rect 72343 18857 72409 18880
rect 72495 18857 72577 18880
rect 72663 18857 72729 18880
rect 72343 18838 72729 18857
rect 76343 18943 76729 18962
rect 76343 18920 76409 18943
rect 76495 18920 76577 18943
rect 76663 18920 76729 18943
rect 76343 18880 76352 18920
rect 76392 18880 76409 18920
rect 76495 18880 76516 18920
rect 76556 18880 76577 18920
rect 76663 18880 76680 18920
rect 76720 18880 76729 18920
rect 76343 18857 76409 18880
rect 76495 18857 76577 18880
rect 76663 18857 76729 18880
rect 76343 18838 76729 18857
rect 80343 18943 80729 18962
rect 80343 18920 80409 18943
rect 80495 18920 80577 18943
rect 80663 18920 80729 18943
rect 80343 18880 80352 18920
rect 80392 18880 80409 18920
rect 80495 18880 80516 18920
rect 80556 18880 80577 18920
rect 80663 18880 80680 18920
rect 80720 18880 80729 18920
rect 80343 18857 80409 18880
rect 80495 18857 80577 18880
rect 80663 18857 80729 18880
rect 80343 18838 80729 18857
rect 84343 18943 84729 18962
rect 84343 18920 84409 18943
rect 84495 18920 84577 18943
rect 84663 18920 84729 18943
rect 84343 18880 84352 18920
rect 84392 18880 84409 18920
rect 84495 18880 84516 18920
rect 84556 18880 84577 18920
rect 84663 18880 84680 18920
rect 84720 18880 84729 18920
rect 84343 18857 84409 18880
rect 84495 18857 84577 18880
rect 84663 18857 84729 18880
rect 84343 18838 84729 18857
rect 88343 18943 88729 18962
rect 88343 18920 88409 18943
rect 88495 18920 88577 18943
rect 88663 18920 88729 18943
rect 88343 18880 88352 18920
rect 88392 18880 88409 18920
rect 88495 18880 88516 18920
rect 88556 18880 88577 18920
rect 88663 18880 88680 18920
rect 88720 18880 88729 18920
rect 88343 18857 88409 18880
rect 88495 18857 88577 18880
rect 88663 18857 88729 18880
rect 88343 18838 88729 18857
rect 92343 18943 92729 18962
rect 92343 18920 92409 18943
rect 92495 18920 92577 18943
rect 92663 18920 92729 18943
rect 92343 18880 92352 18920
rect 92392 18880 92409 18920
rect 92495 18880 92516 18920
rect 92556 18880 92577 18920
rect 92663 18880 92680 18920
rect 92720 18880 92729 18920
rect 92343 18857 92409 18880
rect 92495 18857 92577 18880
rect 92663 18857 92729 18880
rect 92343 18838 92729 18857
rect 96343 18943 96729 18962
rect 96343 18920 96409 18943
rect 96495 18920 96577 18943
rect 96663 18920 96729 18943
rect 96343 18880 96352 18920
rect 96392 18880 96409 18920
rect 96495 18880 96516 18920
rect 96556 18880 96577 18920
rect 96663 18880 96680 18920
rect 96720 18880 96729 18920
rect 96343 18857 96409 18880
rect 96495 18857 96577 18880
rect 96663 18857 96729 18880
rect 96343 18838 96729 18857
rect 3103 18187 3489 18206
rect 3103 18164 3169 18187
rect 3255 18164 3337 18187
rect 3423 18164 3489 18187
rect 3103 18124 3112 18164
rect 3152 18124 3169 18164
rect 3255 18124 3276 18164
rect 3316 18124 3337 18164
rect 3423 18124 3440 18164
rect 3480 18124 3489 18164
rect 3103 18101 3169 18124
rect 3255 18101 3337 18124
rect 3423 18101 3489 18124
rect 3103 18082 3489 18101
rect 7103 18187 7489 18206
rect 7103 18164 7169 18187
rect 7255 18164 7337 18187
rect 7423 18164 7489 18187
rect 7103 18124 7112 18164
rect 7152 18124 7169 18164
rect 7255 18124 7276 18164
rect 7316 18124 7337 18164
rect 7423 18124 7440 18164
rect 7480 18124 7489 18164
rect 7103 18101 7169 18124
rect 7255 18101 7337 18124
rect 7423 18101 7489 18124
rect 7103 18082 7489 18101
rect 11103 18187 11489 18206
rect 11103 18164 11169 18187
rect 11255 18164 11337 18187
rect 11423 18164 11489 18187
rect 11103 18124 11112 18164
rect 11152 18124 11169 18164
rect 11255 18124 11276 18164
rect 11316 18124 11337 18164
rect 11423 18124 11440 18164
rect 11480 18124 11489 18164
rect 11103 18101 11169 18124
rect 11255 18101 11337 18124
rect 11423 18101 11489 18124
rect 11103 18082 11489 18101
rect 15103 18187 15489 18206
rect 15103 18164 15169 18187
rect 15255 18164 15337 18187
rect 15423 18164 15489 18187
rect 15103 18124 15112 18164
rect 15152 18124 15169 18164
rect 15255 18124 15276 18164
rect 15316 18124 15337 18164
rect 15423 18124 15440 18164
rect 15480 18124 15489 18164
rect 15103 18101 15169 18124
rect 15255 18101 15337 18124
rect 15423 18101 15489 18124
rect 15103 18082 15489 18101
rect 19103 18187 19489 18206
rect 19103 18164 19169 18187
rect 19255 18164 19337 18187
rect 19423 18164 19489 18187
rect 19103 18124 19112 18164
rect 19152 18124 19169 18164
rect 19255 18124 19276 18164
rect 19316 18124 19337 18164
rect 19423 18124 19440 18164
rect 19480 18124 19489 18164
rect 19103 18101 19169 18124
rect 19255 18101 19337 18124
rect 19423 18101 19489 18124
rect 19103 18082 19489 18101
rect 23103 18187 23489 18206
rect 23103 18164 23169 18187
rect 23255 18164 23337 18187
rect 23423 18164 23489 18187
rect 23103 18124 23112 18164
rect 23152 18124 23169 18164
rect 23255 18124 23276 18164
rect 23316 18124 23337 18164
rect 23423 18124 23440 18164
rect 23480 18124 23489 18164
rect 23103 18101 23169 18124
rect 23255 18101 23337 18124
rect 23423 18101 23489 18124
rect 23103 18082 23489 18101
rect 27103 18187 27489 18206
rect 27103 18164 27169 18187
rect 27255 18164 27337 18187
rect 27423 18164 27489 18187
rect 27103 18124 27112 18164
rect 27152 18124 27169 18164
rect 27255 18124 27276 18164
rect 27316 18124 27337 18164
rect 27423 18124 27440 18164
rect 27480 18124 27489 18164
rect 27103 18101 27169 18124
rect 27255 18101 27337 18124
rect 27423 18101 27489 18124
rect 27103 18082 27489 18101
rect 31103 18187 31489 18206
rect 31103 18164 31169 18187
rect 31255 18164 31337 18187
rect 31423 18164 31489 18187
rect 31103 18124 31112 18164
rect 31152 18124 31169 18164
rect 31255 18124 31276 18164
rect 31316 18124 31337 18164
rect 31423 18124 31440 18164
rect 31480 18124 31489 18164
rect 31103 18101 31169 18124
rect 31255 18101 31337 18124
rect 31423 18101 31489 18124
rect 31103 18082 31489 18101
rect 35103 18187 35489 18206
rect 35103 18164 35169 18187
rect 35255 18164 35337 18187
rect 35423 18164 35489 18187
rect 35103 18124 35112 18164
rect 35152 18124 35169 18164
rect 35255 18124 35276 18164
rect 35316 18124 35337 18164
rect 35423 18124 35440 18164
rect 35480 18124 35489 18164
rect 35103 18101 35169 18124
rect 35255 18101 35337 18124
rect 35423 18101 35489 18124
rect 35103 18082 35489 18101
rect 39103 18187 39489 18206
rect 39103 18164 39169 18187
rect 39255 18164 39337 18187
rect 39423 18164 39489 18187
rect 39103 18124 39112 18164
rect 39152 18124 39169 18164
rect 39255 18124 39276 18164
rect 39316 18124 39337 18164
rect 39423 18124 39440 18164
rect 39480 18124 39489 18164
rect 39103 18101 39169 18124
rect 39255 18101 39337 18124
rect 39423 18101 39489 18124
rect 39103 18082 39489 18101
rect 43103 18187 43489 18206
rect 43103 18164 43169 18187
rect 43255 18164 43337 18187
rect 43423 18164 43489 18187
rect 43103 18124 43112 18164
rect 43152 18124 43169 18164
rect 43255 18124 43276 18164
rect 43316 18124 43337 18164
rect 43423 18124 43440 18164
rect 43480 18124 43489 18164
rect 43103 18101 43169 18124
rect 43255 18101 43337 18124
rect 43423 18101 43489 18124
rect 43103 18082 43489 18101
rect 47103 18187 47489 18206
rect 47103 18164 47169 18187
rect 47255 18164 47337 18187
rect 47423 18164 47489 18187
rect 47103 18124 47112 18164
rect 47152 18124 47169 18164
rect 47255 18124 47276 18164
rect 47316 18124 47337 18164
rect 47423 18124 47440 18164
rect 47480 18124 47489 18164
rect 47103 18101 47169 18124
rect 47255 18101 47337 18124
rect 47423 18101 47489 18124
rect 47103 18082 47489 18101
rect 51103 18187 51489 18206
rect 51103 18164 51169 18187
rect 51255 18164 51337 18187
rect 51423 18164 51489 18187
rect 51103 18124 51112 18164
rect 51152 18124 51169 18164
rect 51255 18124 51276 18164
rect 51316 18124 51337 18164
rect 51423 18124 51440 18164
rect 51480 18124 51489 18164
rect 51103 18101 51169 18124
rect 51255 18101 51337 18124
rect 51423 18101 51489 18124
rect 51103 18082 51489 18101
rect 55103 18187 55489 18206
rect 55103 18164 55169 18187
rect 55255 18164 55337 18187
rect 55423 18164 55489 18187
rect 55103 18124 55112 18164
rect 55152 18124 55169 18164
rect 55255 18124 55276 18164
rect 55316 18124 55337 18164
rect 55423 18124 55440 18164
rect 55480 18124 55489 18164
rect 55103 18101 55169 18124
rect 55255 18101 55337 18124
rect 55423 18101 55489 18124
rect 55103 18082 55489 18101
rect 59103 18187 59489 18206
rect 59103 18164 59169 18187
rect 59255 18164 59337 18187
rect 59423 18164 59489 18187
rect 59103 18124 59112 18164
rect 59152 18124 59169 18164
rect 59255 18124 59276 18164
rect 59316 18124 59337 18164
rect 59423 18124 59440 18164
rect 59480 18124 59489 18164
rect 59103 18101 59169 18124
rect 59255 18101 59337 18124
rect 59423 18101 59489 18124
rect 59103 18082 59489 18101
rect 63103 18187 63489 18206
rect 63103 18164 63169 18187
rect 63255 18164 63337 18187
rect 63423 18164 63489 18187
rect 63103 18124 63112 18164
rect 63152 18124 63169 18164
rect 63255 18124 63276 18164
rect 63316 18124 63337 18164
rect 63423 18124 63440 18164
rect 63480 18124 63489 18164
rect 63103 18101 63169 18124
rect 63255 18101 63337 18124
rect 63423 18101 63489 18124
rect 63103 18082 63489 18101
rect 67103 18187 67489 18206
rect 67103 18164 67169 18187
rect 67255 18164 67337 18187
rect 67423 18164 67489 18187
rect 67103 18124 67112 18164
rect 67152 18124 67169 18164
rect 67255 18124 67276 18164
rect 67316 18124 67337 18164
rect 67423 18124 67440 18164
rect 67480 18124 67489 18164
rect 67103 18101 67169 18124
rect 67255 18101 67337 18124
rect 67423 18101 67489 18124
rect 67103 18082 67489 18101
rect 71103 18187 71489 18206
rect 71103 18164 71169 18187
rect 71255 18164 71337 18187
rect 71423 18164 71489 18187
rect 71103 18124 71112 18164
rect 71152 18124 71169 18164
rect 71255 18124 71276 18164
rect 71316 18124 71337 18164
rect 71423 18124 71440 18164
rect 71480 18124 71489 18164
rect 71103 18101 71169 18124
rect 71255 18101 71337 18124
rect 71423 18101 71489 18124
rect 71103 18082 71489 18101
rect 75103 18187 75489 18206
rect 75103 18164 75169 18187
rect 75255 18164 75337 18187
rect 75423 18164 75489 18187
rect 75103 18124 75112 18164
rect 75152 18124 75169 18164
rect 75255 18124 75276 18164
rect 75316 18124 75337 18164
rect 75423 18124 75440 18164
rect 75480 18124 75489 18164
rect 75103 18101 75169 18124
rect 75255 18101 75337 18124
rect 75423 18101 75489 18124
rect 75103 18082 75489 18101
rect 79103 18187 79489 18206
rect 79103 18164 79169 18187
rect 79255 18164 79337 18187
rect 79423 18164 79489 18187
rect 79103 18124 79112 18164
rect 79152 18124 79169 18164
rect 79255 18124 79276 18164
rect 79316 18124 79337 18164
rect 79423 18124 79440 18164
rect 79480 18124 79489 18164
rect 79103 18101 79169 18124
rect 79255 18101 79337 18124
rect 79423 18101 79489 18124
rect 79103 18082 79489 18101
rect 83103 18187 83489 18206
rect 83103 18164 83169 18187
rect 83255 18164 83337 18187
rect 83423 18164 83489 18187
rect 83103 18124 83112 18164
rect 83152 18124 83169 18164
rect 83255 18124 83276 18164
rect 83316 18124 83337 18164
rect 83423 18124 83440 18164
rect 83480 18124 83489 18164
rect 83103 18101 83169 18124
rect 83255 18101 83337 18124
rect 83423 18101 83489 18124
rect 83103 18082 83489 18101
rect 87103 18187 87489 18206
rect 87103 18164 87169 18187
rect 87255 18164 87337 18187
rect 87423 18164 87489 18187
rect 87103 18124 87112 18164
rect 87152 18124 87169 18164
rect 87255 18124 87276 18164
rect 87316 18124 87337 18164
rect 87423 18124 87440 18164
rect 87480 18124 87489 18164
rect 87103 18101 87169 18124
rect 87255 18101 87337 18124
rect 87423 18101 87489 18124
rect 87103 18082 87489 18101
rect 91103 18187 91489 18206
rect 91103 18164 91169 18187
rect 91255 18164 91337 18187
rect 91423 18164 91489 18187
rect 91103 18124 91112 18164
rect 91152 18124 91169 18164
rect 91255 18124 91276 18164
rect 91316 18124 91337 18164
rect 91423 18124 91440 18164
rect 91480 18124 91489 18164
rect 91103 18101 91169 18124
rect 91255 18101 91337 18124
rect 91423 18101 91489 18124
rect 91103 18082 91489 18101
rect 95103 18187 95489 18206
rect 95103 18164 95169 18187
rect 95255 18164 95337 18187
rect 95423 18164 95489 18187
rect 95103 18124 95112 18164
rect 95152 18124 95169 18164
rect 95255 18124 95276 18164
rect 95316 18124 95337 18164
rect 95423 18124 95440 18164
rect 95480 18124 95489 18164
rect 95103 18101 95169 18124
rect 95255 18101 95337 18124
rect 95423 18101 95489 18124
rect 95103 18082 95489 18101
rect 99103 18187 99489 18206
rect 99103 18164 99169 18187
rect 99255 18164 99337 18187
rect 99423 18164 99489 18187
rect 99103 18124 99112 18164
rect 99152 18124 99169 18164
rect 99255 18124 99276 18164
rect 99316 18124 99337 18164
rect 99423 18124 99440 18164
rect 99480 18124 99489 18164
rect 99103 18101 99169 18124
rect 99255 18101 99337 18124
rect 99423 18101 99489 18124
rect 99103 18082 99489 18101
rect 4343 17431 4729 17450
rect 4343 17408 4409 17431
rect 4495 17408 4577 17431
rect 4663 17408 4729 17431
rect 4343 17368 4352 17408
rect 4392 17368 4409 17408
rect 4495 17368 4516 17408
rect 4556 17368 4577 17408
rect 4663 17368 4680 17408
rect 4720 17368 4729 17408
rect 4343 17345 4409 17368
rect 4495 17345 4577 17368
rect 4663 17345 4729 17368
rect 4343 17326 4729 17345
rect 8343 17431 8729 17450
rect 8343 17408 8409 17431
rect 8495 17408 8577 17431
rect 8663 17408 8729 17431
rect 8343 17368 8352 17408
rect 8392 17368 8409 17408
rect 8495 17368 8516 17408
rect 8556 17368 8577 17408
rect 8663 17368 8680 17408
rect 8720 17368 8729 17408
rect 8343 17345 8409 17368
rect 8495 17345 8577 17368
rect 8663 17345 8729 17368
rect 8343 17326 8729 17345
rect 12343 17431 12729 17450
rect 12343 17408 12409 17431
rect 12495 17408 12577 17431
rect 12663 17408 12729 17431
rect 12343 17368 12352 17408
rect 12392 17368 12409 17408
rect 12495 17368 12516 17408
rect 12556 17368 12577 17408
rect 12663 17368 12680 17408
rect 12720 17368 12729 17408
rect 12343 17345 12409 17368
rect 12495 17345 12577 17368
rect 12663 17345 12729 17368
rect 12343 17326 12729 17345
rect 16343 17431 16729 17450
rect 16343 17408 16409 17431
rect 16495 17408 16577 17431
rect 16663 17408 16729 17431
rect 16343 17368 16352 17408
rect 16392 17368 16409 17408
rect 16495 17368 16516 17408
rect 16556 17368 16577 17408
rect 16663 17368 16680 17408
rect 16720 17368 16729 17408
rect 16343 17345 16409 17368
rect 16495 17345 16577 17368
rect 16663 17345 16729 17368
rect 16343 17326 16729 17345
rect 20343 17431 20729 17450
rect 20343 17408 20409 17431
rect 20495 17408 20577 17431
rect 20663 17408 20729 17431
rect 20343 17368 20352 17408
rect 20392 17368 20409 17408
rect 20495 17368 20516 17408
rect 20556 17368 20577 17408
rect 20663 17368 20680 17408
rect 20720 17368 20729 17408
rect 20343 17345 20409 17368
rect 20495 17345 20577 17368
rect 20663 17345 20729 17368
rect 20343 17326 20729 17345
rect 24343 17431 24729 17450
rect 24343 17408 24409 17431
rect 24495 17408 24577 17431
rect 24663 17408 24729 17431
rect 24343 17368 24352 17408
rect 24392 17368 24409 17408
rect 24495 17368 24516 17408
rect 24556 17368 24577 17408
rect 24663 17368 24680 17408
rect 24720 17368 24729 17408
rect 24343 17345 24409 17368
rect 24495 17345 24577 17368
rect 24663 17345 24729 17368
rect 24343 17326 24729 17345
rect 28343 17431 28729 17450
rect 28343 17408 28409 17431
rect 28495 17408 28577 17431
rect 28663 17408 28729 17431
rect 28343 17368 28352 17408
rect 28392 17368 28409 17408
rect 28495 17368 28516 17408
rect 28556 17368 28577 17408
rect 28663 17368 28680 17408
rect 28720 17368 28729 17408
rect 28343 17345 28409 17368
rect 28495 17345 28577 17368
rect 28663 17345 28729 17368
rect 28343 17326 28729 17345
rect 32343 17431 32729 17450
rect 32343 17408 32409 17431
rect 32495 17408 32577 17431
rect 32663 17408 32729 17431
rect 32343 17368 32352 17408
rect 32392 17368 32409 17408
rect 32495 17368 32516 17408
rect 32556 17368 32577 17408
rect 32663 17368 32680 17408
rect 32720 17368 32729 17408
rect 32343 17345 32409 17368
rect 32495 17345 32577 17368
rect 32663 17345 32729 17368
rect 32343 17326 32729 17345
rect 36343 17431 36729 17450
rect 36343 17408 36409 17431
rect 36495 17408 36577 17431
rect 36663 17408 36729 17431
rect 36343 17368 36352 17408
rect 36392 17368 36409 17408
rect 36495 17368 36516 17408
rect 36556 17368 36577 17408
rect 36663 17368 36680 17408
rect 36720 17368 36729 17408
rect 36343 17345 36409 17368
rect 36495 17345 36577 17368
rect 36663 17345 36729 17368
rect 36343 17326 36729 17345
rect 40343 17431 40729 17450
rect 40343 17408 40409 17431
rect 40495 17408 40577 17431
rect 40663 17408 40729 17431
rect 40343 17368 40352 17408
rect 40392 17368 40409 17408
rect 40495 17368 40516 17408
rect 40556 17368 40577 17408
rect 40663 17368 40680 17408
rect 40720 17368 40729 17408
rect 40343 17345 40409 17368
rect 40495 17345 40577 17368
rect 40663 17345 40729 17368
rect 40343 17326 40729 17345
rect 44343 17431 44729 17450
rect 44343 17408 44409 17431
rect 44495 17408 44577 17431
rect 44663 17408 44729 17431
rect 44343 17368 44352 17408
rect 44392 17368 44409 17408
rect 44495 17368 44516 17408
rect 44556 17368 44577 17408
rect 44663 17368 44680 17408
rect 44720 17368 44729 17408
rect 44343 17345 44409 17368
rect 44495 17345 44577 17368
rect 44663 17345 44729 17368
rect 44343 17326 44729 17345
rect 48343 17431 48729 17450
rect 48343 17408 48409 17431
rect 48495 17408 48577 17431
rect 48663 17408 48729 17431
rect 48343 17368 48352 17408
rect 48392 17368 48409 17408
rect 48495 17368 48516 17408
rect 48556 17368 48577 17408
rect 48663 17368 48680 17408
rect 48720 17368 48729 17408
rect 48343 17345 48409 17368
rect 48495 17345 48577 17368
rect 48663 17345 48729 17368
rect 48343 17326 48729 17345
rect 52343 17431 52729 17450
rect 52343 17408 52409 17431
rect 52495 17408 52577 17431
rect 52663 17408 52729 17431
rect 52343 17368 52352 17408
rect 52392 17368 52409 17408
rect 52495 17368 52516 17408
rect 52556 17368 52577 17408
rect 52663 17368 52680 17408
rect 52720 17368 52729 17408
rect 52343 17345 52409 17368
rect 52495 17345 52577 17368
rect 52663 17345 52729 17368
rect 52343 17326 52729 17345
rect 56343 17431 56729 17450
rect 56343 17408 56409 17431
rect 56495 17408 56577 17431
rect 56663 17408 56729 17431
rect 56343 17368 56352 17408
rect 56392 17368 56409 17408
rect 56495 17368 56516 17408
rect 56556 17368 56577 17408
rect 56663 17368 56680 17408
rect 56720 17368 56729 17408
rect 56343 17345 56409 17368
rect 56495 17345 56577 17368
rect 56663 17345 56729 17368
rect 56343 17326 56729 17345
rect 60343 17431 60729 17450
rect 60343 17408 60409 17431
rect 60495 17408 60577 17431
rect 60663 17408 60729 17431
rect 60343 17368 60352 17408
rect 60392 17368 60409 17408
rect 60495 17368 60516 17408
rect 60556 17368 60577 17408
rect 60663 17368 60680 17408
rect 60720 17368 60729 17408
rect 60343 17345 60409 17368
rect 60495 17345 60577 17368
rect 60663 17345 60729 17368
rect 60343 17326 60729 17345
rect 64343 17431 64729 17450
rect 64343 17408 64409 17431
rect 64495 17408 64577 17431
rect 64663 17408 64729 17431
rect 64343 17368 64352 17408
rect 64392 17368 64409 17408
rect 64495 17368 64516 17408
rect 64556 17368 64577 17408
rect 64663 17368 64680 17408
rect 64720 17368 64729 17408
rect 64343 17345 64409 17368
rect 64495 17345 64577 17368
rect 64663 17345 64729 17368
rect 64343 17326 64729 17345
rect 68343 17431 68729 17450
rect 68343 17408 68409 17431
rect 68495 17408 68577 17431
rect 68663 17408 68729 17431
rect 68343 17368 68352 17408
rect 68392 17368 68409 17408
rect 68495 17368 68516 17408
rect 68556 17368 68577 17408
rect 68663 17368 68680 17408
rect 68720 17368 68729 17408
rect 68343 17345 68409 17368
rect 68495 17345 68577 17368
rect 68663 17345 68729 17368
rect 68343 17326 68729 17345
rect 72343 17431 72729 17450
rect 72343 17408 72409 17431
rect 72495 17408 72577 17431
rect 72663 17408 72729 17431
rect 72343 17368 72352 17408
rect 72392 17368 72409 17408
rect 72495 17368 72516 17408
rect 72556 17368 72577 17408
rect 72663 17368 72680 17408
rect 72720 17368 72729 17408
rect 72343 17345 72409 17368
rect 72495 17345 72577 17368
rect 72663 17345 72729 17368
rect 72343 17326 72729 17345
rect 76343 17431 76729 17450
rect 76343 17408 76409 17431
rect 76495 17408 76577 17431
rect 76663 17408 76729 17431
rect 76343 17368 76352 17408
rect 76392 17368 76409 17408
rect 76495 17368 76516 17408
rect 76556 17368 76577 17408
rect 76663 17368 76680 17408
rect 76720 17368 76729 17408
rect 76343 17345 76409 17368
rect 76495 17345 76577 17368
rect 76663 17345 76729 17368
rect 76343 17326 76729 17345
rect 80343 17431 80729 17450
rect 80343 17408 80409 17431
rect 80495 17408 80577 17431
rect 80663 17408 80729 17431
rect 80343 17368 80352 17408
rect 80392 17368 80409 17408
rect 80495 17368 80516 17408
rect 80556 17368 80577 17408
rect 80663 17368 80680 17408
rect 80720 17368 80729 17408
rect 80343 17345 80409 17368
rect 80495 17345 80577 17368
rect 80663 17345 80729 17368
rect 80343 17326 80729 17345
rect 84343 17431 84729 17450
rect 84343 17408 84409 17431
rect 84495 17408 84577 17431
rect 84663 17408 84729 17431
rect 84343 17368 84352 17408
rect 84392 17368 84409 17408
rect 84495 17368 84516 17408
rect 84556 17368 84577 17408
rect 84663 17368 84680 17408
rect 84720 17368 84729 17408
rect 84343 17345 84409 17368
rect 84495 17345 84577 17368
rect 84663 17345 84729 17368
rect 84343 17326 84729 17345
rect 88343 17431 88729 17450
rect 88343 17408 88409 17431
rect 88495 17408 88577 17431
rect 88663 17408 88729 17431
rect 88343 17368 88352 17408
rect 88392 17368 88409 17408
rect 88495 17368 88516 17408
rect 88556 17368 88577 17408
rect 88663 17368 88680 17408
rect 88720 17368 88729 17408
rect 88343 17345 88409 17368
rect 88495 17345 88577 17368
rect 88663 17345 88729 17368
rect 88343 17326 88729 17345
rect 92343 17431 92729 17450
rect 92343 17408 92409 17431
rect 92495 17408 92577 17431
rect 92663 17408 92729 17431
rect 92343 17368 92352 17408
rect 92392 17368 92409 17408
rect 92495 17368 92516 17408
rect 92556 17368 92577 17408
rect 92663 17368 92680 17408
rect 92720 17368 92729 17408
rect 92343 17345 92409 17368
rect 92495 17345 92577 17368
rect 92663 17345 92729 17368
rect 92343 17326 92729 17345
rect 96343 17431 96729 17450
rect 96343 17408 96409 17431
rect 96495 17408 96577 17431
rect 96663 17408 96729 17431
rect 96343 17368 96352 17408
rect 96392 17368 96409 17408
rect 96495 17368 96516 17408
rect 96556 17368 96577 17408
rect 96663 17368 96680 17408
rect 96720 17368 96729 17408
rect 96343 17345 96409 17368
rect 96495 17345 96577 17368
rect 96663 17345 96729 17368
rect 96343 17326 96729 17345
rect 3103 16675 3489 16694
rect 3103 16652 3169 16675
rect 3255 16652 3337 16675
rect 3423 16652 3489 16675
rect 3103 16612 3112 16652
rect 3152 16612 3169 16652
rect 3255 16612 3276 16652
rect 3316 16612 3337 16652
rect 3423 16612 3440 16652
rect 3480 16612 3489 16652
rect 3103 16589 3169 16612
rect 3255 16589 3337 16612
rect 3423 16589 3489 16612
rect 3103 16570 3489 16589
rect 7103 16675 7489 16694
rect 7103 16652 7169 16675
rect 7255 16652 7337 16675
rect 7423 16652 7489 16675
rect 7103 16612 7112 16652
rect 7152 16612 7169 16652
rect 7255 16612 7276 16652
rect 7316 16612 7337 16652
rect 7423 16612 7440 16652
rect 7480 16612 7489 16652
rect 7103 16589 7169 16612
rect 7255 16589 7337 16612
rect 7423 16589 7489 16612
rect 7103 16570 7489 16589
rect 11103 16675 11489 16694
rect 11103 16652 11169 16675
rect 11255 16652 11337 16675
rect 11423 16652 11489 16675
rect 11103 16612 11112 16652
rect 11152 16612 11169 16652
rect 11255 16612 11276 16652
rect 11316 16612 11337 16652
rect 11423 16612 11440 16652
rect 11480 16612 11489 16652
rect 11103 16589 11169 16612
rect 11255 16589 11337 16612
rect 11423 16589 11489 16612
rect 11103 16570 11489 16589
rect 15103 16675 15489 16694
rect 15103 16652 15169 16675
rect 15255 16652 15337 16675
rect 15423 16652 15489 16675
rect 15103 16612 15112 16652
rect 15152 16612 15169 16652
rect 15255 16612 15276 16652
rect 15316 16612 15337 16652
rect 15423 16612 15440 16652
rect 15480 16612 15489 16652
rect 15103 16589 15169 16612
rect 15255 16589 15337 16612
rect 15423 16589 15489 16612
rect 15103 16570 15489 16589
rect 19103 16675 19489 16694
rect 19103 16652 19169 16675
rect 19255 16652 19337 16675
rect 19423 16652 19489 16675
rect 19103 16612 19112 16652
rect 19152 16612 19169 16652
rect 19255 16612 19276 16652
rect 19316 16612 19337 16652
rect 19423 16612 19440 16652
rect 19480 16612 19489 16652
rect 19103 16589 19169 16612
rect 19255 16589 19337 16612
rect 19423 16589 19489 16612
rect 19103 16570 19489 16589
rect 23103 16675 23489 16694
rect 23103 16652 23169 16675
rect 23255 16652 23337 16675
rect 23423 16652 23489 16675
rect 23103 16612 23112 16652
rect 23152 16612 23169 16652
rect 23255 16612 23276 16652
rect 23316 16612 23337 16652
rect 23423 16612 23440 16652
rect 23480 16612 23489 16652
rect 23103 16589 23169 16612
rect 23255 16589 23337 16612
rect 23423 16589 23489 16612
rect 23103 16570 23489 16589
rect 27103 16675 27489 16694
rect 27103 16652 27169 16675
rect 27255 16652 27337 16675
rect 27423 16652 27489 16675
rect 27103 16612 27112 16652
rect 27152 16612 27169 16652
rect 27255 16612 27276 16652
rect 27316 16612 27337 16652
rect 27423 16612 27440 16652
rect 27480 16612 27489 16652
rect 27103 16589 27169 16612
rect 27255 16589 27337 16612
rect 27423 16589 27489 16612
rect 27103 16570 27489 16589
rect 31103 16675 31489 16694
rect 31103 16652 31169 16675
rect 31255 16652 31337 16675
rect 31423 16652 31489 16675
rect 31103 16612 31112 16652
rect 31152 16612 31169 16652
rect 31255 16612 31276 16652
rect 31316 16612 31337 16652
rect 31423 16612 31440 16652
rect 31480 16612 31489 16652
rect 31103 16589 31169 16612
rect 31255 16589 31337 16612
rect 31423 16589 31489 16612
rect 31103 16570 31489 16589
rect 35103 16675 35489 16694
rect 35103 16652 35169 16675
rect 35255 16652 35337 16675
rect 35423 16652 35489 16675
rect 35103 16612 35112 16652
rect 35152 16612 35169 16652
rect 35255 16612 35276 16652
rect 35316 16612 35337 16652
rect 35423 16612 35440 16652
rect 35480 16612 35489 16652
rect 35103 16589 35169 16612
rect 35255 16589 35337 16612
rect 35423 16589 35489 16612
rect 35103 16570 35489 16589
rect 39103 16675 39489 16694
rect 39103 16652 39169 16675
rect 39255 16652 39337 16675
rect 39423 16652 39489 16675
rect 39103 16612 39112 16652
rect 39152 16612 39169 16652
rect 39255 16612 39276 16652
rect 39316 16612 39337 16652
rect 39423 16612 39440 16652
rect 39480 16612 39489 16652
rect 39103 16589 39169 16612
rect 39255 16589 39337 16612
rect 39423 16589 39489 16612
rect 39103 16570 39489 16589
rect 43103 16675 43489 16694
rect 43103 16652 43169 16675
rect 43255 16652 43337 16675
rect 43423 16652 43489 16675
rect 43103 16612 43112 16652
rect 43152 16612 43169 16652
rect 43255 16612 43276 16652
rect 43316 16612 43337 16652
rect 43423 16612 43440 16652
rect 43480 16612 43489 16652
rect 43103 16589 43169 16612
rect 43255 16589 43337 16612
rect 43423 16589 43489 16612
rect 43103 16570 43489 16589
rect 47103 16675 47489 16694
rect 47103 16652 47169 16675
rect 47255 16652 47337 16675
rect 47423 16652 47489 16675
rect 47103 16612 47112 16652
rect 47152 16612 47169 16652
rect 47255 16612 47276 16652
rect 47316 16612 47337 16652
rect 47423 16612 47440 16652
rect 47480 16612 47489 16652
rect 47103 16589 47169 16612
rect 47255 16589 47337 16612
rect 47423 16589 47489 16612
rect 47103 16570 47489 16589
rect 51103 16675 51489 16694
rect 51103 16652 51169 16675
rect 51255 16652 51337 16675
rect 51423 16652 51489 16675
rect 51103 16612 51112 16652
rect 51152 16612 51169 16652
rect 51255 16612 51276 16652
rect 51316 16612 51337 16652
rect 51423 16612 51440 16652
rect 51480 16612 51489 16652
rect 51103 16589 51169 16612
rect 51255 16589 51337 16612
rect 51423 16589 51489 16612
rect 51103 16570 51489 16589
rect 55103 16675 55489 16694
rect 55103 16652 55169 16675
rect 55255 16652 55337 16675
rect 55423 16652 55489 16675
rect 55103 16612 55112 16652
rect 55152 16612 55169 16652
rect 55255 16612 55276 16652
rect 55316 16612 55337 16652
rect 55423 16612 55440 16652
rect 55480 16612 55489 16652
rect 55103 16589 55169 16612
rect 55255 16589 55337 16612
rect 55423 16589 55489 16612
rect 55103 16570 55489 16589
rect 59103 16675 59489 16694
rect 59103 16652 59169 16675
rect 59255 16652 59337 16675
rect 59423 16652 59489 16675
rect 59103 16612 59112 16652
rect 59152 16612 59169 16652
rect 59255 16612 59276 16652
rect 59316 16612 59337 16652
rect 59423 16612 59440 16652
rect 59480 16612 59489 16652
rect 59103 16589 59169 16612
rect 59255 16589 59337 16612
rect 59423 16589 59489 16612
rect 59103 16570 59489 16589
rect 63103 16675 63489 16694
rect 63103 16652 63169 16675
rect 63255 16652 63337 16675
rect 63423 16652 63489 16675
rect 63103 16612 63112 16652
rect 63152 16612 63169 16652
rect 63255 16612 63276 16652
rect 63316 16612 63337 16652
rect 63423 16612 63440 16652
rect 63480 16612 63489 16652
rect 63103 16589 63169 16612
rect 63255 16589 63337 16612
rect 63423 16589 63489 16612
rect 63103 16570 63489 16589
rect 67103 16675 67489 16694
rect 67103 16652 67169 16675
rect 67255 16652 67337 16675
rect 67423 16652 67489 16675
rect 67103 16612 67112 16652
rect 67152 16612 67169 16652
rect 67255 16612 67276 16652
rect 67316 16612 67337 16652
rect 67423 16612 67440 16652
rect 67480 16612 67489 16652
rect 67103 16589 67169 16612
rect 67255 16589 67337 16612
rect 67423 16589 67489 16612
rect 67103 16570 67489 16589
rect 71103 16675 71489 16694
rect 71103 16652 71169 16675
rect 71255 16652 71337 16675
rect 71423 16652 71489 16675
rect 71103 16612 71112 16652
rect 71152 16612 71169 16652
rect 71255 16612 71276 16652
rect 71316 16612 71337 16652
rect 71423 16612 71440 16652
rect 71480 16612 71489 16652
rect 71103 16589 71169 16612
rect 71255 16589 71337 16612
rect 71423 16589 71489 16612
rect 71103 16570 71489 16589
rect 75103 16675 75489 16694
rect 75103 16652 75169 16675
rect 75255 16652 75337 16675
rect 75423 16652 75489 16675
rect 75103 16612 75112 16652
rect 75152 16612 75169 16652
rect 75255 16612 75276 16652
rect 75316 16612 75337 16652
rect 75423 16612 75440 16652
rect 75480 16612 75489 16652
rect 75103 16589 75169 16612
rect 75255 16589 75337 16612
rect 75423 16589 75489 16612
rect 75103 16570 75489 16589
rect 79103 16675 79489 16694
rect 79103 16652 79169 16675
rect 79255 16652 79337 16675
rect 79423 16652 79489 16675
rect 79103 16612 79112 16652
rect 79152 16612 79169 16652
rect 79255 16612 79276 16652
rect 79316 16612 79337 16652
rect 79423 16612 79440 16652
rect 79480 16612 79489 16652
rect 79103 16589 79169 16612
rect 79255 16589 79337 16612
rect 79423 16589 79489 16612
rect 79103 16570 79489 16589
rect 83103 16675 83489 16694
rect 83103 16652 83169 16675
rect 83255 16652 83337 16675
rect 83423 16652 83489 16675
rect 83103 16612 83112 16652
rect 83152 16612 83169 16652
rect 83255 16612 83276 16652
rect 83316 16612 83337 16652
rect 83423 16612 83440 16652
rect 83480 16612 83489 16652
rect 83103 16589 83169 16612
rect 83255 16589 83337 16612
rect 83423 16589 83489 16612
rect 83103 16570 83489 16589
rect 87103 16675 87489 16694
rect 87103 16652 87169 16675
rect 87255 16652 87337 16675
rect 87423 16652 87489 16675
rect 87103 16612 87112 16652
rect 87152 16612 87169 16652
rect 87255 16612 87276 16652
rect 87316 16612 87337 16652
rect 87423 16612 87440 16652
rect 87480 16612 87489 16652
rect 87103 16589 87169 16612
rect 87255 16589 87337 16612
rect 87423 16589 87489 16612
rect 87103 16570 87489 16589
rect 91103 16675 91489 16694
rect 91103 16652 91169 16675
rect 91255 16652 91337 16675
rect 91423 16652 91489 16675
rect 91103 16612 91112 16652
rect 91152 16612 91169 16652
rect 91255 16612 91276 16652
rect 91316 16612 91337 16652
rect 91423 16612 91440 16652
rect 91480 16612 91489 16652
rect 91103 16589 91169 16612
rect 91255 16589 91337 16612
rect 91423 16589 91489 16612
rect 91103 16570 91489 16589
rect 95103 16675 95489 16694
rect 95103 16652 95169 16675
rect 95255 16652 95337 16675
rect 95423 16652 95489 16675
rect 95103 16612 95112 16652
rect 95152 16612 95169 16652
rect 95255 16612 95276 16652
rect 95316 16612 95337 16652
rect 95423 16612 95440 16652
rect 95480 16612 95489 16652
rect 95103 16589 95169 16612
rect 95255 16589 95337 16612
rect 95423 16589 95489 16612
rect 95103 16570 95489 16589
rect 99103 16675 99489 16694
rect 99103 16652 99169 16675
rect 99255 16652 99337 16675
rect 99423 16652 99489 16675
rect 99103 16612 99112 16652
rect 99152 16612 99169 16652
rect 99255 16612 99276 16652
rect 99316 16612 99337 16652
rect 99423 16612 99440 16652
rect 99480 16612 99489 16652
rect 99103 16589 99169 16612
rect 99255 16589 99337 16612
rect 99423 16589 99489 16612
rect 99103 16570 99489 16589
rect 86450 16423 86574 16442
rect 86450 16400 86469 16423
rect 86179 16360 86188 16400
rect 86228 16360 86469 16400
rect 86450 16337 86469 16360
rect 86555 16337 86574 16423
rect 86450 16318 86574 16337
rect 4343 15919 4729 15938
rect 4343 15896 4409 15919
rect 4495 15896 4577 15919
rect 4663 15896 4729 15919
rect 4343 15856 4352 15896
rect 4392 15856 4409 15896
rect 4495 15856 4516 15896
rect 4556 15856 4577 15896
rect 4663 15856 4680 15896
rect 4720 15856 4729 15896
rect 4343 15833 4409 15856
rect 4495 15833 4577 15856
rect 4663 15833 4729 15856
rect 4343 15814 4729 15833
rect 8343 15919 8729 15938
rect 8343 15896 8409 15919
rect 8495 15896 8577 15919
rect 8663 15896 8729 15919
rect 8343 15856 8352 15896
rect 8392 15856 8409 15896
rect 8495 15856 8516 15896
rect 8556 15856 8577 15896
rect 8663 15856 8680 15896
rect 8720 15856 8729 15896
rect 8343 15833 8409 15856
rect 8495 15833 8577 15856
rect 8663 15833 8729 15856
rect 8343 15814 8729 15833
rect 12343 15919 12729 15938
rect 12343 15896 12409 15919
rect 12495 15896 12577 15919
rect 12663 15896 12729 15919
rect 12343 15856 12352 15896
rect 12392 15856 12409 15896
rect 12495 15856 12516 15896
rect 12556 15856 12577 15896
rect 12663 15856 12680 15896
rect 12720 15856 12729 15896
rect 12343 15833 12409 15856
rect 12495 15833 12577 15856
rect 12663 15833 12729 15856
rect 12343 15814 12729 15833
rect 16343 15919 16729 15938
rect 16343 15896 16409 15919
rect 16495 15896 16577 15919
rect 16663 15896 16729 15919
rect 16343 15856 16352 15896
rect 16392 15856 16409 15896
rect 16495 15856 16516 15896
rect 16556 15856 16577 15896
rect 16663 15856 16680 15896
rect 16720 15856 16729 15896
rect 16343 15833 16409 15856
rect 16495 15833 16577 15856
rect 16663 15833 16729 15856
rect 16343 15814 16729 15833
rect 20343 15919 20729 15938
rect 20343 15896 20409 15919
rect 20495 15896 20577 15919
rect 20663 15896 20729 15919
rect 20343 15856 20352 15896
rect 20392 15856 20409 15896
rect 20495 15856 20516 15896
rect 20556 15856 20577 15896
rect 20663 15856 20680 15896
rect 20720 15856 20729 15896
rect 20343 15833 20409 15856
rect 20495 15833 20577 15856
rect 20663 15833 20729 15856
rect 20343 15814 20729 15833
rect 24343 15919 24729 15938
rect 24343 15896 24409 15919
rect 24495 15896 24577 15919
rect 24663 15896 24729 15919
rect 24343 15856 24352 15896
rect 24392 15856 24409 15896
rect 24495 15856 24516 15896
rect 24556 15856 24577 15896
rect 24663 15856 24680 15896
rect 24720 15856 24729 15896
rect 24343 15833 24409 15856
rect 24495 15833 24577 15856
rect 24663 15833 24729 15856
rect 24343 15814 24729 15833
rect 28343 15919 28729 15938
rect 28343 15896 28409 15919
rect 28495 15896 28577 15919
rect 28663 15896 28729 15919
rect 28343 15856 28352 15896
rect 28392 15856 28409 15896
rect 28495 15856 28516 15896
rect 28556 15856 28577 15896
rect 28663 15856 28680 15896
rect 28720 15856 28729 15896
rect 28343 15833 28409 15856
rect 28495 15833 28577 15856
rect 28663 15833 28729 15856
rect 28343 15814 28729 15833
rect 32343 15919 32729 15938
rect 32343 15896 32409 15919
rect 32495 15896 32577 15919
rect 32663 15896 32729 15919
rect 32343 15856 32352 15896
rect 32392 15856 32409 15896
rect 32495 15856 32516 15896
rect 32556 15856 32577 15896
rect 32663 15856 32680 15896
rect 32720 15856 32729 15896
rect 32343 15833 32409 15856
rect 32495 15833 32577 15856
rect 32663 15833 32729 15856
rect 32343 15814 32729 15833
rect 36343 15919 36729 15938
rect 36343 15896 36409 15919
rect 36495 15896 36577 15919
rect 36663 15896 36729 15919
rect 36343 15856 36352 15896
rect 36392 15856 36409 15896
rect 36495 15856 36516 15896
rect 36556 15856 36577 15896
rect 36663 15856 36680 15896
rect 36720 15856 36729 15896
rect 36343 15833 36409 15856
rect 36495 15833 36577 15856
rect 36663 15833 36729 15856
rect 36343 15814 36729 15833
rect 40343 15919 40729 15938
rect 40343 15896 40409 15919
rect 40495 15896 40577 15919
rect 40663 15896 40729 15919
rect 40343 15856 40352 15896
rect 40392 15856 40409 15896
rect 40495 15856 40516 15896
rect 40556 15856 40577 15896
rect 40663 15856 40680 15896
rect 40720 15856 40729 15896
rect 40343 15833 40409 15856
rect 40495 15833 40577 15856
rect 40663 15833 40729 15856
rect 40343 15814 40729 15833
rect 44343 15919 44729 15938
rect 44343 15896 44409 15919
rect 44495 15896 44577 15919
rect 44663 15896 44729 15919
rect 44343 15856 44352 15896
rect 44392 15856 44409 15896
rect 44495 15856 44516 15896
rect 44556 15856 44577 15896
rect 44663 15856 44680 15896
rect 44720 15856 44729 15896
rect 44343 15833 44409 15856
rect 44495 15833 44577 15856
rect 44663 15833 44729 15856
rect 44343 15814 44729 15833
rect 48343 15919 48729 15938
rect 48343 15896 48409 15919
rect 48495 15896 48577 15919
rect 48663 15896 48729 15919
rect 48343 15856 48352 15896
rect 48392 15856 48409 15896
rect 48495 15856 48516 15896
rect 48556 15856 48577 15896
rect 48663 15856 48680 15896
rect 48720 15856 48729 15896
rect 48343 15833 48409 15856
rect 48495 15833 48577 15856
rect 48663 15833 48729 15856
rect 48343 15814 48729 15833
rect 52343 15919 52729 15938
rect 52343 15896 52409 15919
rect 52495 15896 52577 15919
rect 52663 15896 52729 15919
rect 52343 15856 52352 15896
rect 52392 15856 52409 15896
rect 52495 15856 52516 15896
rect 52556 15856 52577 15896
rect 52663 15856 52680 15896
rect 52720 15856 52729 15896
rect 52343 15833 52409 15856
rect 52495 15833 52577 15856
rect 52663 15833 52729 15856
rect 52343 15814 52729 15833
rect 56343 15919 56729 15938
rect 56343 15896 56409 15919
rect 56495 15896 56577 15919
rect 56663 15896 56729 15919
rect 56343 15856 56352 15896
rect 56392 15856 56409 15896
rect 56495 15856 56516 15896
rect 56556 15856 56577 15896
rect 56663 15856 56680 15896
rect 56720 15856 56729 15896
rect 56343 15833 56409 15856
rect 56495 15833 56577 15856
rect 56663 15833 56729 15856
rect 56343 15814 56729 15833
rect 60343 15919 60729 15938
rect 60343 15896 60409 15919
rect 60495 15896 60577 15919
rect 60663 15896 60729 15919
rect 60343 15856 60352 15896
rect 60392 15856 60409 15896
rect 60495 15856 60516 15896
rect 60556 15856 60577 15896
rect 60663 15856 60680 15896
rect 60720 15856 60729 15896
rect 60343 15833 60409 15856
rect 60495 15833 60577 15856
rect 60663 15833 60729 15856
rect 60343 15814 60729 15833
rect 64343 15919 64729 15938
rect 64343 15896 64409 15919
rect 64495 15896 64577 15919
rect 64663 15896 64729 15919
rect 64343 15856 64352 15896
rect 64392 15856 64409 15896
rect 64495 15856 64516 15896
rect 64556 15856 64577 15896
rect 64663 15856 64680 15896
rect 64720 15856 64729 15896
rect 64343 15833 64409 15856
rect 64495 15833 64577 15856
rect 64663 15833 64729 15856
rect 64343 15814 64729 15833
rect 68343 15919 68729 15938
rect 68343 15896 68409 15919
rect 68495 15896 68577 15919
rect 68663 15896 68729 15919
rect 68343 15856 68352 15896
rect 68392 15856 68409 15896
rect 68495 15856 68516 15896
rect 68556 15856 68577 15896
rect 68663 15856 68680 15896
rect 68720 15856 68729 15896
rect 68343 15833 68409 15856
rect 68495 15833 68577 15856
rect 68663 15833 68729 15856
rect 68343 15814 68729 15833
rect 72343 15919 72729 15938
rect 72343 15896 72409 15919
rect 72495 15896 72577 15919
rect 72663 15896 72729 15919
rect 72343 15856 72352 15896
rect 72392 15856 72409 15896
rect 72495 15856 72516 15896
rect 72556 15856 72577 15896
rect 72663 15856 72680 15896
rect 72720 15856 72729 15896
rect 72343 15833 72409 15856
rect 72495 15833 72577 15856
rect 72663 15833 72729 15856
rect 72343 15814 72729 15833
rect 76343 15919 76729 15938
rect 76343 15896 76409 15919
rect 76495 15896 76577 15919
rect 76663 15896 76729 15919
rect 76343 15856 76352 15896
rect 76392 15856 76409 15896
rect 76495 15856 76516 15896
rect 76556 15856 76577 15896
rect 76663 15856 76680 15896
rect 76720 15856 76729 15896
rect 76343 15833 76409 15856
rect 76495 15833 76577 15856
rect 76663 15833 76729 15856
rect 76343 15814 76729 15833
rect 80343 15919 80729 15938
rect 80343 15896 80409 15919
rect 80495 15896 80577 15919
rect 80663 15896 80729 15919
rect 80343 15856 80352 15896
rect 80392 15856 80409 15896
rect 80495 15856 80516 15896
rect 80556 15856 80577 15896
rect 80663 15856 80680 15896
rect 80720 15856 80729 15896
rect 80343 15833 80409 15856
rect 80495 15833 80577 15856
rect 80663 15833 80729 15856
rect 80343 15814 80729 15833
rect 84343 15919 84729 15938
rect 84343 15896 84409 15919
rect 84495 15896 84577 15919
rect 84663 15896 84729 15919
rect 84343 15856 84352 15896
rect 84392 15856 84409 15896
rect 84495 15856 84516 15896
rect 84556 15856 84577 15896
rect 84663 15856 84680 15896
rect 84720 15856 84729 15896
rect 84343 15833 84409 15856
rect 84495 15833 84577 15856
rect 84663 15833 84729 15856
rect 84343 15814 84729 15833
rect 88343 15919 88729 15938
rect 88343 15896 88409 15919
rect 88495 15896 88577 15919
rect 88663 15896 88729 15919
rect 88343 15856 88352 15896
rect 88392 15856 88409 15896
rect 88495 15856 88516 15896
rect 88556 15856 88577 15896
rect 88663 15856 88680 15896
rect 88720 15856 88729 15896
rect 88343 15833 88409 15856
rect 88495 15833 88577 15856
rect 88663 15833 88729 15856
rect 88343 15814 88729 15833
rect 92343 15919 92729 15938
rect 92343 15896 92409 15919
rect 92495 15896 92577 15919
rect 92663 15896 92729 15919
rect 92343 15856 92352 15896
rect 92392 15856 92409 15896
rect 92495 15856 92516 15896
rect 92556 15856 92577 15896
rect 92663 15856 92680 15896
rect 92720 15856 92729 15896
rect 92343 15833 92409 15856
rect 92495 15833 92577 15856
rect 92663 15833 92729 15856
rect 92343 15814 92729 15833
rect 96343 15919 96729 15938
rect 96343 15896 96409 15919
rect 96495 15896 96577 15919
rect 96663 15896 96729 15919
rect 96343 15856 96352 15896
rect 96392 15856 96409 15896
rect 96495 15856 96516 15896
rect 96556 15856 96577 15896
rect 96663 15856 96680 15896
rect 96720 15856 96729 15896
rect 96343 15833 96409 15856
rect 96495 15833 96577 15856
rect 96663 15833 96729 15856
rect 96343 15814 96729 15833
rect 3103 15163 3489 15182
rect 3103 15140 3169 15163
rect 3255 15140 3337 15163
rect 3423 15140 3489 15163
rect 3103 15100 3112 15140
rect 3152 15100 3169 15140
rect 3255 15100 3276 15140
rect 3316 15100 3337 15140
rect 3423 15100 3440 15140
rect 3480 15100 3489 15140
rect 3103 15077 3169 15100
rect 3255 15077 3337 15100
rect 3423 15077 3489 15100
rect 3103 15058 3489 15077
rect 7103 15163 7489 15182
rect 7103 15140 7169 15163
rect 7255 15140 7337 15163
rect 7423 15140 7489 15163
rect 7103 15100 7112 15140
rect 7152 15100 7169 15140
rect 7255 15100 7276 15140
rect 7316 15100 7337 15140
rect 7423 15100 7440 15140
rect 7480 15100 7489 15140
rect 7103 15077 7169 15100
rect 7255 15077 7337 15100
rect 7423 15077 7489 15100
rect 7103 15058 7489 15077
rect 11103 15163 11489 15182
rect 11103 15140 11169 15163
rect 11255 15140 11337 15163
rect 11423 15140 11489 15163
rect 11103 15100 11112 15140
rect 11152 15100 11169 15140
rect 11255 15100 11276 15140
rect 11316 15100 11337 15140
rect 11423 15100 11440 15140
rect 11480 15100 11489 15140
rect 11103 15077 11169 15100
rect 11255 15077 11337 15100
rect 11423 15077 11489 15100
rect 11103 15058 11489 15077
rect 15103 15163 15489 15182
rect 15103 15140 15169 15163
rect 15255 15140 15337 15163
rect 15423 15140 15489 15163
rect 15103 15100 15112 15140
rect 15152 15100 15169 15140
rect 15255 15100 15276 15140
rect 15316 15100 15337 15140
rect 15423 15100 15440 15140
rect 15480 15100 15489 15140
rect 15103 15077 15169 15100
rect 15255 15077 15337 15100
rect 15423 15077 15489 15100
rect 15103 15058 15489 15077
rect 19103 15163 19489 15182
rect 19103 15140 19169 15163
rect 19255 15140 19337 15163
rect 19423 15140 19489 15163
rect 19103 15100 19112 15140
rect 19152 15100 19169 15140
rect 19255 15100 19276 15140
rect 19316 15100 19337 15140
rect 19423 15100 19440 15140
rect 19480 15100 19489 15140
rect 19103 15077 19169 15100
rect 19255 15077 19337 15100
rect 19423 15077 19489 15100
rect 19103 15058 19489 15077
rect 23103 15163 23489 15182
rect 23103 15140 23169 15163
rect 23255 15140 23337 15163
rect 23423 15140 23489 15163
rect 23103 15100 23112 15140
rect 23152 15100 23169 15140
rect 23255 15100 23276 15140
rect 23316 15100 23337 15140
rect 23423 15100 23440 15140
rect 23480 15100 23489 15140
rect 23103 15077 23169 15100
rect 23255 15077 23337 15100
rect 23423 15077 23489 15100
rect 23103 15058 23489 15077
rect 27103 15163 27489 15182
rect 27103 15140 27169 15163
rect 27255 15140 27337 15163
rect 27423 15140 27489 15163
rect 27103 15100 27112 15140
rect 27152 15100 27169 15140
rect 27255 15100 27276 15140
rect 27316 15100 27337 15140
rect 27423 15100 27440 15140
rect 27480 15100 27489 15140
rect 27103 15077 27169 15100
rect 27255 15077 27337 15100
rect 27423 15077 27489 15100
rect 27103 15058 27489 15077
rect 31103 15163 31489 15182
rect 31103 15140 31169 15163
rect 31255 15140 31337 15163
rect 31423 15140 31489 15163
rect 31103 15100 31112 15140
rect 31152 15100 31169 15140
rect 31255 15100 31276 15140
rect 31316 15100 31337 15140
rect 31423 15100 31440 15140
rect 31480 15100 31489 15140
rect 31103 15077 31169 15100
rect 31255 15077 31337 15100
rect 31423 15077 31489 15100
rect 31103 15058 31489 15077
rect 35103 15163 35489 15182
rect 35103 15140 35169 15163
rect 35255 15140 35337 15163
rect 35423 15140 35489 15163
rect 35103 15100 35112 15140
rect 35152 15100 35169 15140
rect 35255 15100 35276 15140
rect 35316 15100 35337 15140
rect 35423 15100 35440 15140
rect 35480 15100 35489 15140
rect 35103 15077 35169 15100
rect 35255 15077 35337 15100
rect 35423 15077 35489 15100
rect 35103 15058 35489 15077
rect 39103 15163 39489 15182
rect 39103 15140 39169 15163
rect 39255 15140 39337 15163
rect 39423 15140 39489 15163
rect 39103 15100 39112 15140
rect 39152 15100 39169 15140
rect 39255 15100 39276 15140
rect 39316 15100 39337 15140
rect 39423 15100 39440 15140
rect 39480 15100 39489 15140
rect 39103 15077 39169 15100
rect 39255 15077 39337 15100
rect 39423 15077 39489 15100
rect 39103 15058 39489 15077
rect 43103 15163 43489 15182
rect 43103 15140 43169 15163
rect 43255 15140 43337 15163
rect 43423 15140 43489 15163
rect 43103 15100 43112 15140
rect 43152 15100 43169 15140
rect 43255 15100 43276 15140
rect 43316 15100 43337 15140
rect 43423 15100 43440 15140
rect 43480 15100 43489 15140
rect 43103 15077 43169 15100
rect 43255 15077 43337 15100
rect 43423 15077 43489 15100
rect 43103 15058 43489 15077
rect 47103 15163 47489 15182
rect 47103 15140 47169 15163
rect 47255 15140 47337 15163
rect 47423 15140 47489 15163
rect 47103 15100 47112 15140
rect 47152 15100 47169 15140
rect 47255 15100 47276 15140
rect 47316 15100 47337 15140
rect 47423 15100 47440 15140
rect 47480 15100 47489 15140
rect 47103 15077 47169 15100
rect 47255 15077 47337 15100
rect 47423 15077 47489 15100
rect 47103 15058 47489 15077
rect 51103 15163 51489 15182
rect 51103 15140 51169 15163
rect 51255 15140 51337 15163
rect 51423 15140 51489 15163
rect 51103 15100 51112 15140
rect 51152 15100 51169 15140
rect 51255 15100 51276 15140
rect 51316 15100 51337 15140
rect 51423 15100 51440 15140
rect 51480 15100 51489 15140
rect 51103 15077 51169 15100
rect 51255 15077 51337 15100
rect 51423 15077 51489 15100
rect 51103 15058 51489 15077
rect 55103 15163 55489 15182
rect 55103 15140 55169 15163
rect 55255 15140 55337 15163
rect 55423 15140 55489 15163
rect 55103 15100 55112 15140
rect 55152 15100 55169 15140
rect 55255 15100 55276 15140
rect 55316 15100 55337 15140
rect 55423 15100 55440 15140
rect 55480 15100 55489 15140
rect 55103 15077 55169 15100
rect 55255 15077 55337 15100
rect 55423 15077 55489 15100
rect 55103 15058 55489 15077
rect 59103 15163 59489 15182
rect 59103 15140 59169 15163
rect 59255 15140 59337 15163
rect 59423 15140 59489 15163
rect 59103 15100 59112 15140
rect 59152 15100 59169 15140
rect 59255 15100 59276 15140
rect 59316 15100 59337 15140
rect 59423 15100 59440 15140
rect 59480 15100 59489 15140
rect 59103 15077 59169 15100
rect 59255 15077 59337 15100
rect 59423 15077 59489 15100
rect 59103 15058 59489 15077
rect 63103 15163 63489 15182
rect 63103 15140 63169 15163
rect 63255 15140 63337 15163
rect 63423 15140 63489 15163
rect 63103 15100 63112 15140
rect 63152 15100 63169 15140
rect 63255 15100 63276 15140
rect 63316 15100 63337 15140
rect 63423 15100 63440 15140
rect 63480 15100 63489 15140
rect 63103 15077 63169 15100
rect 63255 15077 63337 15100
rect 63423 15077 63489 15100
rect 63103 15058 63489 15077
rect 67103 15163 67489 15182
rect 67103 15140 67169 15163
rect 67255 15140 67337 15163
rect 67423 15140 67489 15163
rect 67103 15100 67112 15140
rect 67152 15100 67169 15140
rect 67255 15100 67276 15140
rect 67316 15100 67337 15140
rect 67423 15100 67440 15140
rect 67480 15100 67489 15140
rect 67103 15077 67169 15100
rect 67255 15077 67337 15100
rect 67423 15077 67489 15100
rect 67103 15058 67489 15077
rect 4343 14407 4729 14426
rect 4343 14384 4409 14407
rect 4495 14384 4577 14407
rect 4663 14384 4729 14407
rect 4343 14344 4352 14384
rect 4392 14344 4409 14384
rect 4495 14344 4516 14384
rect 4556 14344 4577 14384
rect 4663 14344 4680 14384
rect 4720 14344 4729 14384
rect 4343 14321 4409 14344
rect 4495 14321 4577 14344
rect 4663 14321 4729 14344
rect 4343 14302 4729 14321
rect 8343 14407 8729 14426
rect 8343 14384 8409 14407
rect 8495 14384 8577 14407
rect 8663 14384 8729 14407
rect 8343 14344 8352 14384
rect 8392 14344 8409 14384
rect 8495 14344 8516 14384
rect 8556 14344 8577 14384
rect 8663 14344 8680 14384
rect 8720 14344 8729 14384
rect 8343 14321 8409 14344
rect 8495 14321 8577 14344
rect 8663 14321 8729 14344
rect 8343 14302 8729 14321
rect 12343 14407 12729 14426
rect 12343 14384 12409 14407
rect 12495 14384 12577 14407
rect 12663 14384 12729 14407
rect 12343 14344 12352 14384
rect 12392 14344 12409 14384
rect 12495 14344 12516 14384
rect 12556 14344 12577 14384
rect 12663 14344 12680 14384
rect 12720 14344 12729 14384
rect 12343 14321 12409 14344
rect 12495 14321 12577 14344
rect 12663 14321 12729 14344
rect 12343 14302 12729 14321
rect 16343 14407 16729 14426
rect 16343 14384 16409 14407
rect 16495 14384 16577 14407
rect 16663 14384 16729 14407
rect 16343 14344 16352 14384
rect 16392 14344 16409 14384
rect 16495 14344 16516 14384
rect 16556 14344 16577 14384
rect 16663 14344 16680 14384
rect 16720 14344 16729 14384
rect 16343 14321 16409 14344
rect 16495 14321 16577 14344
rect 16663 14321 16729 14344
rect 16343 14302 16729 14321
rect 20343 14407 20729 14426
rect 20343 14384 20409 14407
rect 20495 14384 20577 14407
rect 20663 14384 20729 14407
rect 20343 14344 20352 14384
rect 20392 14344 20409 14384
rect 20495 14344 20516 14384
rect 20556 14344 20577 14384
rect 20663 14344 20680 14384
rect 20720 14344 20729 14384
rect 20343 14321 20409 14344
rect 20495 14321 20577 14344
rect 20663 14321 20729 14344
rect 20343 14302 20729 14321
rect 24343 14407 24729 14426
rect 24343 14384 24409 14407
rect 24495 14384 24577 14407
rect 24663 14384 24729 14407
rect 24343 14344 24352 14384
rect 24392 14344 24409 14384
rect 24495 14344 24516 14384
rect 24556 14344 24577 14384
rect 24663 14344 24680 14384
rect 24720 14344 24729 14384
rect 24343 14321 24409 14344
rect 24495 14321 24577 14344
rect 24663 14321 24729 14344
rect 24343 14302 24729 14321
rect 28343 14407 28729 14426
rect 28343 14384 28409 14407
rect 28495 14384 28577 14407
rect 28663 14384 28729 14407
rect 28343 14344 28352 14384
rect 28392 14344 28409 14384
rect 28495 14344 28516 14384
rect 28556 14344 28577 14384
rect 28663 14344 28680 14384
rect 28720 14344 28729 14384
rect 28343 14321 28409 14344
rect 28495 14321 28577 14344
rect 28663 14321 28729 14344
rect 28343 14302 28729 14321
rect 32343 14407 32729 14426
rect 32343 14384 32409 14407
rect 32495 14384 32577 14407
rect 32663 14384 32729 14407
rect 32343 14344 32352 14384
rect 32392 14344 32409 14384
rect 32495 14344 32516 14384
rect 32556 14344 32577 14384
rect 32663 14344 32680 14384
rect 32720 14344 32729 14384
rect 32343 14321 32409 14344
rect 32495 14321 32577 14344
rect 32663 14321 32729 14344
rect 32343 14302 32729 14321
rect 36343 14407 36729 14426
rect 36343 14384 36409 14407
rect 36495 14384 36577 14407
rect 36663 14384 36729 14407
rect 36343 14344 36352 14384
rect 36392 14344 36409 14384
rect 36495 14344 36516 14384
rect 36556 14344 36577 14384
rect 36663 14344 36680 14384
rect 36720 14344 36729 14384
rect 36343 14321 36409 14344
rect 36495 14321 36577 14344
rect 36663 14321 36729 14344
rect 36343 14302 36729 14321
rect 40343 14407 40729 14426
rect 40343 14384 40409 14407
rect 40495 14384 40577 14407
rect 40663 14384 40729 14407
rect 40343 14344 40352 14384
rect 40392 14344 40409 14384
rect 40495 14344 40516 14384
rect 40556 14344 40577 14384
rect 40663 14344 40680 14384
rect 40720 14344 40729 14384
rect 40343 14321 40409 14344
rect 40495 14321 40577 14344
rect 40663 14321 40729 14344
rect 40343 14302 40729 14321
rect 44343 14407 44729 14426
rect 44343 14384 44409 14407
rect 44495 14384 44577 14407
rect 44663 14384 44729 14407
rect 44343 14344 44352 14384
rect 44392 14344 44409 14384
rect 44495 14344 44516 14384
rect 44556 14344 44577 14384
rect 44663 14344 44680 14384
rect 44720 14344 44729 14384
rect 44343 14321 44409 14344
rect 44495 14321 44577 14344
rect 44663 14321 44729 14344
rect 44343 14302 44729 14321
rect 48343 14407 48729 14426
rect 48343 14384 48409 14407
rect 48495 14384 48577 14407
rect 48663 14384 48729 14407
rect 48343 14344 48352 14384
rect 48392 14344 48409 14384
rect 48495 14344 48516 14384
rect 48556 14344 48577 14384
rect 48663 14344 48680 14384
rect 48720 14344 48729 14384
rect 48343 14321 48409 14344
rect 48495 14321 48577 14344
rect 48663 14321 48729 14344
rect 48343 14302 48729 14321
rect 52343 14407 52729 14426
rect 52343 14384 52409 14407
rect 52495 14384 52577 14407
rect 52663 14384 52729 14407
rect 52343 14344 52352 14384
rect 52392 14344 52409 14384
rect 52495 14344 52516 14384
rect 52556 14344 52577 14384
rect 52663 14344 52680 14384
rect 52720 14344 52729 14384
rect 52343 14321 52409 14344
rect 52495 14321 52577 14344
rect 52663 14321 52729 14344
rect 52343 14302 52729 14321
rect 56343 14407 56729 14426
rect 56343 14384 56409 14407
rect 56495 14384 56577 14407
rect 56663 14384 56729 14407
rect 56343 14344 56352 14384
rect 56392 14344 56409 14384
rect 56495 14344 56516 14384
rect 56556 14344 56577 14384
rect 56663 14344 56680 14384
rect 56720 14344 56729 14384
rect 56343 14321 56409 14344
rect 56495 14321 56577 14344
rect 56663 14321 56729 14344
rect 56343 14302 56729 14321
rect 60343 14407 60729 14426
rect 60343 14384 60409 14407
rect 60495 14384 60577 14407
rect 60663 14384 60729 14407
rect 60343 14344 60352 14384
rect 60392 14344 60409 14384
rect 60495 14344 60516 14384
rect 60556 14344 60577 14384
rect 60663 14344 60680 14384
rect 60720 14344 60729 14384
rect 60343 14321 60409 14344
rect 60495 14321 60577 14344
rect 60663 14321 60729 14344
rect 60343 14302 60729 14321
rect 64343 14407 64729 14426
rect 64343 14384 64409 14407
rect 64495 14384 64577 14407
rect 64663 14384 64729 14407
rect 64343 14344 64352 14384
rect 64392 14344 64409 14384
rect 64495 14344 64516 14384
rect 64556 14344 64577 14384
rect 64663 14344 64680 14384
rect 64720 14344 64729 14384
rect 64343 14321 64409 14344
rect 64495 14321 64577 14344
rect 64663 14321 64729 14344
rect 64343 14302 64729 14321
rect 68343 14407 68729 14426
rect 68343 14384 68409 14407
rect 68495 14384 68577 14407
rect 68663 14384 68729 14407
rect 68343 14344 68352 14384
rect 68392 14344 68409 14384
rect 68495 14344 68516 14384
rect 68556 14344 68577 14384
rect 68663 14344 68680 14384
rect 68720 14344 68729 14384
rect 68343 14321 68409 14344
rect 68495 14321 68577 14344
rect 68663 14321 68729 14344
rect 68343 14302 68729 14321
rect 3103 13651 3489 13670
rect 3103 13628 3169 13651
rect 3255 13628 3337 13651
rect 3423 13628 3489 13651
rect 3103 13588 3112 13628
rect 3152 13588 3169 13628
rect 3255 13588 3276 13628
rect 3316 13588 3337 13628
rect 3423 13588 3440 13628
rect 3480 13588 3489 13628
rect 3103 13565 3169 13588
rect 3255 13565 3337 13588
rect 3423 13565 3489 13588
rect 3103 13546 3489 13565
rect 7103 13651 7489 13670
rect 7103 13628 7169 13651
rect 7255 13628 7337 13651
rect 7423 13628 7489 13651
rect 7103 13588 7112 13628
rect 7152 13588 7169 13628
rect 7255 13588 7276 13628
rect 7316 13588 7337 13628
rect 7423 13588 7440 13628
rect 7480 13588 7489 13628
rect 7103 13565 7169 13588
rect 7255 13565 7337 13588
rect 7423 13565 7489 13588
rect 7103 13546 7489 13565
rect 11103 13651 11489 13670
rect 11103 13628 11169 13651
rect 11255 13628 11337 13651
rect 11423 13628 11489 13651
rect 11103 13588 11112 13628
rect 11152 13588 11169 13628
rect 11255 13588 11276 13628
rect 11316 13588 11337 13628
rect 11423 13588 11440 13628
rect 11480 13588 11489 13628
rect 11103 13565 11169 13588
rect 11255 13565 11337 13588
rect 11423 13565 11489 13588
rect 11103 13546 11489 13565
rect 15103 13651 15489 13670
rect 15103 13628 15169 13651
rect 15255 13628 15337 13651
rect 15423 13628 15489 13651
rect 15103 13588 15112 13628
rect 15152 13588 15169 13628
rect 15255 13588 15276 13628
rect 15316 13588 15337 13628
rect 15423 13588 15440 13628
rect 15480 13588 15489 13628
rect 15103 13565 15169 13588
rect 15255 13565 15337 13588
rect 15423 13565 15489 13588
rect 15103 13546 15489 13565
rect 19103 13651 19489 13670
rect 19103 13628 19169 13651
rect 19255 13628 19337 13651
rect 19423 13628 19489 13651
rect 19103 13588 19112 13628
rect 19152 13588 19169 13628
rect 19255 13588 19276 13628
rect 19316 13588 19337 13628
rect 19423 13588 19440 13628
rect 19480 13588 19489 13628
rect 19103 13565 19169 13588
rect 19255 13565 19337 13588
rect 19423 13565 19489 13588
rect 19103 13546 19489 13565
rect 23103 13651 23489 13670
rect 23103 13628 23169 13651
rect 23255 13628 23337 13651
rect 23423 13628 23489 13651
rect 23103 13588 23112 13628
rect 23152 13588 23169 13628
rect 23255 13588 23276 13628
rect 23316 13588 23337 13628
rect 23423 13588 23440 13628
rect 23480 13588 23489 13628
rect 23103 13565 23169 13588
rect 23255 13565 23337 13588
rect 23423 13565 23489 13588
rect 23103 13546 23489 13565
rect 27103 13651 27489 13670
rect 27103 13628 27169 13651
rect 27255 13628 27337 13651
rect 27423 13628 27489 13651
rect 27103 13588 27112 13628
rect 27152 13588 27169 13628
rect 27255 13588 27276 13628
rect 27316 13588 27337 13628
rect 27423 13588 27440 13628
rect 27480 13588 27489 13628
rect 27103 13565 27169 13588
rect 27255 13565 27337 13588
rect 27423 13565 27489 13588
rect 27103 13546 27489 13565
rect 31103 13651 31489 13670
rect 31103 13628 31169 13651
rect 31255 13628 31337 13651
rect 31423 13628 31489 13651
rect 31103 13588 31112 13628
rect 31152 13588 31169 13628
rect 31255 13588 31276 13628
rect 31316 13588 31337 13628
rect 31423 13588 31440 13628
rect 31480 13588 31489 13628
rect 31103 13565 31169 13588
rect 31255 13565 31337 13588
rect 31423 13565 31489 13588
rect 31103 13546 31489 13565
rect 35103 13651 35489 13670
rect 35103 13628 35169 13651
rect 35255 13628 35337 13651
rect 35423 13628 35489 13651
rect 35103 13588 35112 13628
rect 35152 13588 35169 13628
rect 35255 13588 35276 13628
rect 35316 13588 35337 13628
rect 35423 13588 35440 13628
rect 35480 13588 35489 13628
rect 35103 13565 35169 13588
rect 35255 13565 35337 13588
rect 35423 13565 35489 13588
rect 35103 13546 35489 13565
rect 39103 13651 39489 13670
rect 39103 13628 39169 13651
rect 39255 13628 39337 13651
rect 39423 13628 39489 13651
rect 39103 13588 39112 13628
rect 39152 13588 39169 13628
rect 39255 13588 39276 13628
rect 39316 13588 39337 13628
rect 39423 13588 39440 13628
rect 39480 13588 39489 13628
rect 39103 13565 39169 13588
rect 39255 13565 39337 13588
rect 39423 13565 39489 13588
rect 39103 13546 39489 13565
rect 43103 13651 43489 13670
rect 43103 13628 43169 13651
rect 43255 13628 43337 13651
rect 43423 13628 43489 13651
rect 43103 13588 43112 13628
rect 43152 13588 43169 13628
rect 43255 13588 43276 13628
rect 43316 13588 43337 13628
rect 43423 13588 43440 13628
rect 43480 13588 43489 13628
rect 43103 13565 43169 13588
rect 43255 13565 43337 13588
rect 43423 13565 43489 13588
rect 43103 13546 43489 13565
rect 47103 13651 47489 13670
rect 47103 13628 47169 13651
rect 47255 13628 47337 13651
rect 47423 13628 47489 13651
rect 47103 13588 47112 13628
rect 47152 13588 47169 13628
rect 47255 13588 47276 13628
rect 47316 13588 47337 13628
rect 47423 13588 47440 13628
rect 47480 13588 47489 13628
rect 47103 13565 47169 13588
rect 47255 13565 47337 13588
rect 47423 13565 47489 13588
rect 47103 13546 47489 13565
rect 51103 13651 51489 13670
rect 51103 13628 51169 13651
rect 51255 13628 51337 13651
rect 51423 13628 51489 13651
rect 51103 13588 51112 13628
rect 51152 13588 51169 13628
rect 51255 13588 51276 13628
rect 51316 13588 51337 13628
rect 51423 13588 51440 13628
rect 51480 13588 51489 13628
rect 51103 13565 51169 13588
rect 51255 13565 51337 13588
rect 51423 13565 51489 13588
rect 51103 13546 51489 13565
rect 55103 13651 55489 13670
rect 55103 13628 55169 13651
rect 55255 13628 55337 13651
rect 55423 13628 55489 13651
rect 55103 13588 55112 13628
rect 55152 13588 55169 13628
rect 55255 13588 55276 13628
rect 55316 13588 55337 13628
rect 55423 13588 55440 13628
rect 55480 13588 55489 13628
rect 55103 13565 55169 13588
rect 55255 13565 55337 13588
rect 55423 13565 55489 13588
rect 55103 13546 55489 13565
rect 59103 13651 59489 13670
rect 59103 13628 59169 13651
rect 59255 13628 59337 13651
rect 59423 13628 59489 13651
rect 59103 13588 59112 13628
rect 59152 13588 59169 13628
rect 59255 13588 59276 13628
rect 59316 13588 59337 13628
rect 59423 13588 59440 13628
rect 59480 13588 59489 13628
rect 59103 13565 59169 13588
rect 59255 13565 59337 13588
rect 59423 13565 59489 13588
rect 59103 13546 59489 13565
rect 63103 13651 63489 13670
rect 63103 13628 63169 13651
rect 63255 13628 63337 13651
rect 63423 13628 63489 13651
rect 63103 13588 63112 13628
rect 63152 13588 63169 13628
rect 63255 13588 63276 13628
rect 63316 13588 63337 13628
rect 63423 13588 63440 13628
rect 63480 13588 63489 13628
rect 63103 13565 63169 13588
rect 63255 13565 63337 13588
rect 63423 13565 63489 13588
rect 63103 13546 63489 13565
rect 67103 13651 67489 13670
rect 67103 13628 67169 13651
rect 67255 13628 67337 13651
rect 67423 13628 67489 13651
rect 67103 13588 67112 13628
rect 67152 13588 67169 13628
rect 67255 13588 67276 13628
rect 67316 13588 67337 13628
rect 67423 13588 67440 13628
rect 67480 13588 67489 13628
rect 67103 13565 67169 13588
rect 67255 13565 67337 13588
rect 67423 13565 67489 13588
rect 67103 13546 67489 13565
rect 72316 13122 72756 13252
rect 72316 13036 72409 13122
rect 72495 13036 72577 13122
rect 72663 13036 72756 13122
rect 72316 12954 72756 13036
rect 4343 12895 4729 12914
rect 4343 12872 4409 12895
rect 4495 12872 4577 12895
rect 4663 12872 4729 12895
rect 4343 12832 4352 12872
rect 4392 12832 4409 12872
rect 4495 12832 4516 12872
rect 4556 12832 4577 12872
rect 4663 12832 4680 12872
rect 4720 12832 4729 12872
rect 4343 12809 4409 12832
rect 4495 12809 4577 12832
rect 4663 12809 4729 12832
rect 4343 12790 4729 12809
rect 8343 12895 8729 12914
rect 8343 12872 8409 12895
rect 8495 12872 8577 12895
rect 8663 12872 8729 12895
rect 8343 12832 8352 12872
rect 8392 12832 8409 12872
rect 8495 12832 8516 12872
rect 8556 12832 8577 12872
rect 8663 12832 8680 12872
rect 8720 12832 8729 12872
rect 8343 12809 8409 12832
rect 8495 12809 8577 12832
rect 8663 12809 8729 12832
rect 8343 12790 8729 12809
rect 12343 12895 12729 12914
rect 12343 12872 12409 12895
rect 12495 12872 12577 12895
rect 12663 12872 12729 12895
rect 12343 12832 12352 12872
rect 12392 12832 12409 12872
rect 12495 12832 12516 12872
rect 12556 12832 12577 12872
rect 12663 12832 12680 12872
rect 12720 12832 12729 12872
rect 12343 12809 12409 12832
rect 12495 12809 12577 12832
rect 12663 12809 12729 12832
rect 12343 12790 12729 12809
rect 16343 12895 16729 12914
rect 16343 12872 16409 12895
rect 16495 12872 16577 12895
rect 16663 12872 16729 12895
rect 16343 12832 16352 12872
rect 16392 12832 16409 12872
rect 16495 12832 16516 12872
rect 16556 12832 16577 12872
rect 16663 12832 16680 12872
rect 16720 12832 16729 12872
rect 16343 12809 16409 12832
rect 16495 12809 16577 12832
rect 16663 12809 16729 12832
rect 16343 12790 16729 12809
rect 20343 12895 20729 12914
rect 20343 12872 20409 12895
rect 20495 12872 20577 12895
rect 20663 12872 20729 12895
rect 20343 12832 20352 12872
rect 20392 12832 20409 12872
rect 20495 12832 20516 12872
rect 20556 12832 20577 12872
rect 20663 12832 20680 12872
rect 20720 12832 20729 12872
rect 20343 12809 20409 12832
rect 20495 12809 20577 12832
rect 20663 12809 20729 12832
rect 20343 12790 20729 12809
rect 24343 12895 24729 12914
rect 24343 12872 24409 12895
rect 24495 12872 24577 12895
rect 24663 12872 24729 12895
rect 24343 12832 24352 12872
rect 24392 12832 24409 12872
rect 24495 12832 24516 12872
rect 24556 12832 24577 12872
rect 24663 12832 24680 12872
rect 24720 12832 24729 12872
rect 24343 12809 24409 12832
rect 24495 12809 24577 12832
rect 24663 12809 24729 12832
rect 24343 12790 24729 12809
rect 28343 12895 28729 12914
rect 28343 12872 28409 12895
rect 28495 12872 28577 12895
rect 28663 12872 28729 12895
rect 28343 12832 28352 12872
rect 28392 12832 28409 12872
rect 28495 12832 28516 12872
rect 28556 12832 28577 12872
rect 28663 12832 28680 12872
rect 28720 12832 28729 12872
rect 28343 12809 28409 12832
rect 28495 12809 28577 12832
rect 28663 12809 28729 12832
rect 28343 12790 28729 12809
rect 32343 12895 32729 12914
rect 32343 12872 32409 12895
rect 32495 12872 32577 12895
rect 32663 12872 32729 12895
rect 32343 12832 32352 12872
rect 32392 12832 32409 12872
rect 32495 12832 32516 12872
rect 32556 12832 32577 12872
rect 32663 12832 32680 12872
rect 32720 12832 32729 12872
rect 32343 12809 32409 12832
rect 32495 12809 32577 12832
rect 32663 12809 32729 12832
rect 32343 12790 32729 12809
rect 36343 12895 36729 12914
rect 36343 12872 36409 12895
rect 36495 12872 36577 12895
rect 36663 12872 36729 12895
rect 36343 12832 36352 12872
rect 36392 12832 36409 12872
rect 36495 12832 36516 12872
rect 36556 12832 36577 12872
rect 36663 12832 36680 12872
rect 36720 12832 36729 12872
rect 36343 12809 36409 12832
rect 36495 12809 36577 12832
rect 36663 12809 36729 12832
rect 36343 12790 36729 12809
rect 40343 12895 40729 12914
rect 40343 12872 40409 12895
rect 40495 12872 40577 12895
rect 40663 12872 40729 12895
rect 40343 12832 40352 12872
rect 40392 12832 40409 12872
rect 40495 12832 40516 12872
rect 40556 12832 40577 12872
rect 40663 12832 40680 12872
rect 40720 12832 40729 12872
rect 40343 12809 40409 12832
rect 40495 12809 40577 12832
rect 40663 12809 40729 12832
rect 40343 12790 40729 12809
rect 44343 12895 44729 12914
rect 44343 12872 44409 12895
rect 44495 12872 44577 12895
rect 44663 12872 44729 12895
rect 44343 12832 44352 12872
rect 44392 12832 44409 12872
rect 44495 12832 44516 12872
rect 44556 12832 44577 12872
rect 44663 12832 44680 12872
rect 44720 12832 44729 12872
rect 44343 12809 44409 12832
rect 44495 12809 44577 12832
rect 44663 12809 44729 12832
rect 44343 12790 44729 12809
rect 48343 12895 48729 12914
rect 48343 12872 48409 12895
rect 48495 12872 48577 12895
rect 48663 12872 48729 12895
rect 48343 12832 48352 12872
rect 48392 12832 48409 12872
rect 48495 12832 48516 12872
rect 48556 12832 48577 12872
rect 48663 12832 48680 12872
rect 48720 12832 48729 12872
rect 48343 12809 48409 12832
rect 48495 12809 48577 12832
rect 48663 12809 48729 12832
rect 48343 12790 48729 12809
rect 52343 12895 52729 12914
rect 52343 12872 52409 12895
rect 52495 12872 52577 12895
rect 52663 12872 52729 12895
rect 52343 12832 52352 12872
rect 52392 12832 52409 12872
rect 52495 12832 52516 12872
rect 52556 12832 52577 12872
rect 52663 12832 52680 12872
rect 52720 12832 52729 12872
rect 52343 12809 52409 12832
rect 52495 12809 52577 12832
rect 52663 12809 52729 12832
rect 52343 12790 52729 12809
rect 56343 12895 56729 12914
rect 56343 12872 56409 12895
rect 56495 12872 56577 12895
rect 56663 12872 56729 12895
rect 56343 12832 56352 12872
rect 56392 12832 56409 12872
rect 56495 12832 56516 12872
rect 56556 12832 56577 12872
rect 56663 12832 56680 12872
rect 56720 12832 56729 12872
rect 56343 12809 56409 12832
rect 56495 12809 56577 12832
rect 56663 12809 56729 12832
rect 56343 12790 56729 12809
rect 60343 12895 60729 12914
rect 60343 12872 60409 12895
rect 60495 12872 60577 12895
rect 60663 12872 60729 12895
rect 60343 12832 60352 12872
rect 60392 12832 60409 12872
rect 60495 12832 60516 12872
rect 60556 12832 60577 12872
rect 60663 12832 60680 12872
rect 60720 12832 60729 12872
rect 60343 12809 60409 12832
rect 60495 12809 60577 12832
rect 60663 12809 60729 12832
rect 60343 12790 60729 12809
rect 64343 12895 64729 12914
rect 64343 12872 64409 12895
rect 64495 12872 64577 12895
rect 64663 12872 64729 12895
rect 64343 12832 64352 12872
rect 64392 12832 64409 12872
rect 64495 12832 64516 12872
rect 64556 12832 64577 12872
rect 64663 12832 64680 12872
rect 64720 12832 64729 12872
rect 64343 12809 64409 12832
rect 64495 12809 64577 12832
rect 64663 12809 64729 12832
rect 64343 12790 64729 12809
rect 68343 12895 68729 12914
rect 68343 12872 68409 12895
rect 68495 12872 68577 12895
rect 68663 12872 68729 12895
rect 68343 12832 68352 12872
rect 68392 12832 68409 12872
rect 68495 12832 68516 12872
rect 68556 12832 68577 12872
rect 68663 12832 68680 12872
rect 68720 12832 68729 12872
rect 68343 12809 68409 12832
rect 68495 12809 68577 12832
rect 68663 12809 68729 12832
rect 68343 12790 68729 12809
rect 72316 12868 72409 12954
rect 72495 12868 72577 12954
rect 72663 12868 72756 12954
rect 72316 12786 72756 12868
rect 72316 12700 72409 12786
rect 72495 12700 72577 12786
rect 72663 12700 72756 12786
rect 72316 12618 72756 12700
rect 72316 12532 72409 12618
rect 72495 12532 72577 12618
rect 72663 12532 72756 12618
rect 72316 12450 72756 12532
rect 72316 12364 72409 12450
rect 72495 12364 72577 12450
rect 72663 12364 72756 12450
rect 72316 12282 72756 12364
rect 72316 12196 72409 12282
rect 72495 12196 72577 12282
rect 72663 12196 72756 12282
rect 3103 12139 3489 12158
rect 3103 12116 3169 12139
rect 3255 12116 3337 12139
rect 3423 12116 3489 12139
rect 3103 12076 3112 12116
rect 3152 12076 3169 12116
rect 3255 12076 3276 12116
rect 3316 12076 3337 12116
rect 3423 12076 3440 12116
rect 3480 12076 3489 12116
rect 3103 12053 3169 12076
rect 3255 12053 3337 12076
rect 3423 12053 3489 12076
rect 3103 12034 3489 12053
rect 7103 12139 7489 12158
rect 7103 12116 7169 12139
rect 7255 12116 7337 12139
rect 7423 12116 7489 12139
rect 7103 12076 7112 12116
rect 7152 12076 7169 12116
rect 7255 12076 7276 12116
rect 7316 12076 7337 12116
rect 7423 12076 7440 12116
rect 7480 12076 7489 12116
rect 7103 12053 7169 12076
rect 7255 12053 7337 12076
rect 7423 12053 7489 12076
rect 7103 12034 7489 12053
rect 11103 12139 11489 12158
rect 11103 12116 11169 12139
rect 11255 12116 11337 12139
rect 11423 12116 11489 12139
rect 11103 12076 11112 12116
rect 11152 12076 11169 12116
rect 11255 12076 11276 12116
rect 11316 12076 11337 12116
rect 11423 12076 11440 12116
rect 11480 12076 11489 12116
rect 11103 12053 11169 12076
rect 11255 12053 11337 12076
rect 11423 12053 11489 12076
rect 11103 12034 11489 12053
rect 15103 12139 15489 12158
rect 15103 12116 15169 12139
rect 15255 12116 15337 12139
rect 15423 12116 15489 12139
rect 15103 12076 15112 12116
rect 15152 12076 15169 12116
rect 15255 12076 15276 12116
rect 15316 12076 15337 12116
rect 15423 12076 15440 12116
rect 15480 12076 15489 12116
rect 15103 12053 15169 12076
rect 15255 12053 15337 12076
rect 15423 12053 15489 12076
rect 15103 12034 15489 12053
rect 19103 12139 19489 12158
rect 19103 12116 19169 12139
rect 19255 12116 19337 12139
rect 19423 12116 19489 12139
rect 19103 12076 19112 12116
rect 19152 12076 19169 12116
rect 19255 12076 19276 12116
rect 19316 12076 19337 12116
rect 19423 12076 19440 12116
rect 19480 12076 19489 12116
rect 19103 12053 19169 12076
rect 19255 12053 19337 12076
rect 19423 12053 19489 12076
rect 19103 12034 19489 12053
rect 23103 12139 23489 12158
rect 23103 12116 23169 12139
rect 23255 12116 23337 12139
rect 23423 12116 23489 12139
rect 23103 12076 23112 12116
rect 23152 12076 23169 12116
rect 23255 12076 23276 12116
rect 23316 12076 23337 12116
rect 23423 12076 23440 12116
rect 23480 12076 23489 12116
rect 23103 12053 23169 12076
rect 23255 12053 23337 12076
rect 23423 12053 23489 12076
rect 23103 12034 23489 12053
rect 27103 12139 27489 12158
rect 27103 12116 27169 12139
rect 27255 12116 27337 12139
rect 27423 12116 27489 12139
rect 27103 12076 27112 12116
rect 27152 12076 27169 12116
rect 27255 12076 27276 12116
rect 27316 12076 27337 12116
rect 27423 12076 27440 12116
rect 27480 12076 27489 12116
rect 27103 12053 27169 12076
rect 27255 12053 27337 12076
rect 27423 12053 27489 12076
rect 27103 12034 27489 12053
rect 31103 12139 31489 12158
rect 31103 12116 31169 12139
rect 31255 12116 31337 12139
rect 31423 12116 31489 12139
rect 31103 12076 31112 12116
rect 31152 12076 31169 12116
rect 31255 12076 31276 12116
rect 31316 12076 31337 12116
rect 31423 12076 31440 12116
rect 31480 12076 31489 12116
rect 31103 12053 31169 12076
rect 31255 12053 31337 12076
rect 31423 12053 31489 12076
rect 31103 12034 31489 12053
rect 35103 12139 35489 12158
rect 35103 12116 35169 12139
rect 35255 12116 35337 12139
rect 35423 12116 35489 12139
rect 35103 12076 35112 12116
rect 35152 12076 35169 12116
rect 35255 12076 35276 12116
rect 35316 12076 35337 12116
rect 35423 12076 35440 12116
rect 35480 12076 35489 12116
rect 35103 12053 35169 12076
rect 35255 12053 35337 12076
rect 35423 12053 35489 12076
rect 35103 12034 35489 12053
rect 39103 12139 39489 12158
rect 39103 12116 39169 12139
rect 39255 12116 39337 12139
rect 39423 12116 39489 12139
rect 39103 12076 39112 12116
rect 39152 12076 39169 12116
rect 39255 12076 39276 12116
rect 39316 12076 39337 12116
rect 39423 12076 39440 12116
rect 39480 12076 39489 12116
rect 39103 12053 39169 12076
rect 39255 12053 39337 12076
rect 39423 12053 39489 12076
rect 39103 12034 39489 12053
rect 43103 12139 43489 12158
rect 43103 12116 43169 12139
rect 43255 12116 43337 12139
rect 43423 12116 43489 12139
rect 43103 12076 43112 12116
rect 43152 12076 43169 12116
rect 43255 12076 43276 12116
rect 43316 12076 43337 12116
rect 43423 12076 43440 12116
rect 43480 12076 43489 12116
rect 43103 12053 43169 12076
rect 43255 12053 43337 12076
rect 43423 12053 43489 12076
rect 43103 12034 43489 12053
rect 47103 12139 47489 12158
rect 47103 12116 47169 12139
rect 47255 12116 47337 12139
rect 47423 12116 47489 12139
rect 47103 12076 47112 12116
rect 47152 12076 47169 12116
rect 47255 12076 47276 12116
rect 47316 12076 47337 12116
rect 47423 12076 47440 12116
rect 47480 12076 47489 12116
rect 47103 12053 47169 12076
rect 47255 12053 47337 12076
rect 47423 12053 47489 12076
rect 47103 12034 47489 12053
rect 51103 12139 51489 12158
rect 51103 12116 51169 12139
rect 51255 12116 51337 12139
rect 51423 12116 51489 12139
rect 51103 12076 51112 12116
rect 51152 12076 51169 12116
rect 51255 12076 51276 12116
rect 51316 12076 51337 12116
rect 51423 12076 51440 12116
rect 51480 12076 51489 12116
rect 51103 12053 51169 12076
rect 51255 12053 51337 12076
rect 51423 12053 51489 12076
rect 51103 12034 51489 12053
rect 55103 12139 55489 12158
rect 55103 12116 55169 12139
rect 55255 12116 55337 12139
rect 55423 12116 55489 12139
rect 55103 12076 55112 12116
rect 55152 12076 55169 12116
rect 55255 12076 55276 12116
rect 55316 12076 55337 12116
rect 55423 12076 55440 12116
rect 55480 12076 55489 12116
rect 55103 12053 55169 12076
rect 55255 12053 55337 12076
rect 55423 12053 55489 12076
rect 55103 12034 55489 12053
rect 59103 12139 59489 12158
rect 59103 12116 59169 12139
rect 59255 12116 59337 12139
rect 59423 12116 59489 12139
rect 59103 12076 59112 12116
rect 59152 12076 59169 12116
rect 59255 12076 59276 12116
rect 59316 12076 59337 12116
rect 59423 12076 59440 12116
rect 59480 12076 59489 12116
rect 59103 12053 59169 12076
rect 59255 12053 59337 12076
rect 59423 12053 59489 12076
rect 59103 12034 59489 12053
rect 63103 12139 63489 12158
rect 63103 12116 63169 12139
rect 63255 12116 63337 12139
rect 63423 12116 63489 12139
rect 63103 12076 63112 12116
rect 63152 12076 63169 12116
rect 63255 12076 63276 12116
rect 63316 12076 63337 12116
rect 63423 12076 63440 12116
rect 63480 12076 63489 12116
rect 63103 12053 63169 12076
rect 63255 12053 63337 12076
rect 63423 12053 63489 12076
rect 63103 12034 63489 12053
rect 67103 12139 67489 12158
rect 67103 12116 67169 12139
rect 67255 12116 67337 12139
rect 67423 12116 67489 12139
rect 67103 12076 67112 12116
rect 67152 12076 67169 12116
rect 67255 12076 67276 12116
rect 67316 12076 67337 12116
rect 67423 12076 67440 12116
rect 67480 12076 67489 12116
rect 67103 12053 67169 12076
rect 67255 12053 67337 12076
rect 67423 12053 67489 12076
rect 67103 12034 67489 12053
rect 72316 12114 72756 12196
rect 72316 12028 72409 12114
rect 72495 12028 72577 12114
rect 72663 12028 72756 12114
rect 72316 11946 72756 12028
rect 72316 11860 72409 11946
rect 72495 11860 72577 11946
rect 72663 11860 72756 11946
rect 72316 11778 72756 11860
rect 72316 11692 72409 11778
rect 72495 11692 72577 11778
rect 72663 11692 72756 11778
rect 72316 11610 72756 11692
rect 72316 11524 72409 11610
rect 72495 11524 72577 11610
rect 72663 11524 72756 11610
rect 72316 11442 72756 11524
rect 4343 11383 4729 11402
rect 4343 11360 4409 11383
rect 4495 11360 4577 11383
rect 4663 11360 4729 11383
rect 4343 11320 4352 11360
rect 4392 11320 4409 11360
rect 4495 11320 4516 11360
rect 4556 11320 4577 11360
rect 4663 11320 4680 11360
rect 4720 11320 4729 11360
rect 4343 11297 4409 11320
rect 4495 11297 4577 11320
rect 4663 11297 4729 11320
rect 4343 11278 4729 11297
rect 8343 11383 8729 11402
rect 8343 11360 8409 11383
rect 8495 11360 8577 11383
rect 8663 11360 8729 11383
rect 8343 11320 8352 11360
rect 8392 11320 8409 11360
rect 8495 11320 8516 11360
rect 8556 11320 8577 11360
rect 8663 11320 8680 11360
rect 8720 11320 8729 11360
rect 8343 11297 8409 11320
rect 8495 11297 8577 11320
rect 8663 11297 8729 11320
rect 8343 11278 8729 11297
rect 12343 11383 12729 11402
rect 12343 11360 12409 11383
rect 12495 11360 12577 11383
rect 12663 11360 12729 11383
rect 12343 11320 12352 11360
rect 12392 11320 12409 11360
rect 12495 11320 12516 11360
rect 12556 11320 12577 11360
rect 12663 11320 12680 11360
rect 12720 11320 12729 11360
rect 12343 11297 12409 11320
rect 12495 11297 12577 11320
rect 12663 11297 12729 11320
rect 12343 11278 12729 11297
rect 16343 11383 16729 11402
rect 16343 11360 16409 11383
rect 16495 11360 16577 11383
rect 16663 11360 16729 11383
rect 16343 11320 16352 11360
rect 16392 11320 16409 11360
rect 16495 11320 16516 11360
rect 16556 11320 16577 11360
rect 16663 11320 16680 11360
rect 16720 11320 16729 11360
rect 16343 11297 16409 11320
rect 16495 11297 16577 11320
rect 16663 11297 16729 11320
rect 16343 11278 16729 11297
rect 20343 11383 20729 11402
rect 20343 11360 20409 11383
rect 20495 11360 20577 11383
rect 20663 11360 20729 11383
rect 20343 11320 20352 11360
rect 20392 11320 20409 11360
rect 20495 11320 20516 11360
rect 20556 11320 20577 11360
rect 20663 11320 20680 11360
rect 20720 11320 20729 11360
rect 20343 11297 20409 11320
rect 20495 11297 20577 11320
rect 20663 11297 20729 11320
rect 20343 11278 20729 11297
rect 24343 11383 24729 11402
rect 24343 11360 24409 11383
rect 24495 11360 24577 11383
rect 24663 11360 24729 11383
rect 24343 11320 24352 11360
rect 24392 11320 24409 11360
rect 24495 11320 24516 11360
rect 24556 11320 24577 11360
rect 24663 11320 24680 11360
rect 24720 11320 24729 11360
rect 24343 11297 24409 11320
rect 24495 11297 24577 11320
rect 24663 11297 24729 11320
rect 24343 11278 24729 11297
rect 28343 11383 28729 11402
rect 28343 11360 28409 11383
rect 28495 11360 28577 11383
rect 28663 11360 28729 11383
rect 28343 11320 28352 11360
rect 28392 11320 28409 11360
rect 28495 11320 28516 11360
rect 28556 11320 28577 11360
rect 28663 11320 28680 11360
rect 28720 11320 28729 11360
rect 28343 11297 28409 11320
rect 28495 11297 28577 11320
rect 28663 11297 28729 11320
rect 28343 11278 28729 11297
rect 32343 11383 32729 11402
rect 32343 11360 32409 11383
rect 32495 11360 32577 11383
rect 32663 11360 32729 11383
rect 32343 11320 32352 11360
rect 32392 11320 32409 11360
rect 32495 11320 32516 11360
rect 32556 11320 32577 11360
rect 32663 11320 32680 11360
rect 32720 11320 32729 11360
rect 32343 11297 32409 11320
rect 32495 11297 32577 11320
rect 32663 11297 32729 11320
rect 32343 11278 32729 11297
rect 36343 11383 36729 11402
rect 36343 11360 36409 11383
rect 36495 11360 36577 11383
rect 36663 11360 36729 11383
rect 36343 11320 36352 11360
rect 36392 11320 36409 11360
rect 36495 11320 36516 11360
rect 36556 11320 36577 11360
rect 36663 11320 36680 11360
rect 36720 11320 36729 11360
rect 36343 11297 36409 11320
rect 36495 11297 36577 11320
rect 36663 11297 36729 11320
rect 36343 11278 36729 11297
rect 40343 11383 40729 11402
rect 40343 11360 40409 11383
rect 40495 11360 40577 11383
rect 40663 11360 40729 11383
rect 40343 11320 40352 11360
rect 40392 11320 40409 11360
rect 40495 11320 40516 11360
rect 40556 11320 40577 11360
rect 40663 11320 40680 11360
rect 40720 11320 40729 11360
rect 40343 11297 40409 11320
rect 40495 11297 40577 11320
rect 40663 11297 40729 11320
rect 40343 11278 40729 11297
rect 44343 11383 44729 11402
rect 44343 11360 44409 11383
rect 44495 11360 44577 11383
rect 44663 11360 44729 11383
rect 44343 11320 44352 11360
rect 44392 11320 44409 11360
rect 44495 11320 44516 11360
rect 44556 11320 44577 11360
rect 44663 11320 44680 11360
rect 44720 11320 44729 11360
rect 44343 11297 44409 11320
rect 44495 11297 44577 11320
rect 44663 11297 44729 11320
rect 44343 11278 44729 11297
rect 48343 11383 48729 11402
rect 48343 11360 48409 11383
rect 48495 11360 48577 11383
rect 48663 11360 48729 11383
rect 48343 11320 48352 11360
rect 48392 11320 48409 11360
rect 48495 11320 48516 11360
rect 48556 11320 48577 11360
rect 48663 11320 48680 11360
rect 48720 11320 48729 11360
rect 48343 11297 48409 11320
rect 48495 11297 48577 11320
rect 48663 11297 48729 11320
rect 48343 11278 48729 11297
rect 52343 11383 52729 11402
rect 52343 11360 52409 11383
rect 52495 11360 52577 11383
rect 52663 11360 52729 11383
rect 52343 11320 52352 11360
rect 52392 11320 52409 11360
rect 52495 11320 52516 11360
rect 52556 11320 52577 11360
rect 52663 11320 52680 11360
rect 52720 11320 52729 11360
rect 52343 11297 52409 11320
rect 52495 11297 52577 11320
rect 52663 11297 52729 11320
rect 52343 11278 52729 11297
rect 56343 11383 56729 11402
rect 56343 11360 56409 11383
rect 56495 11360 56577 11383
rect 56663 11360 56729 11383
rect 56343 11320 56352 11360
rect 56392 11320 56409 11360
rect 56495 11320 56516 11360
rect 56556 11320 56577 11360
rect 56663 11320 56680 11360
rect 56720 11320 56729 11360
rect 56343 11297 56409 11320
rect 56495 11297 56577 11320
rect 56663 11297 56729 11320
rect 56343 11278 56729 11297
rect 60343 11383 60729 11402
rect 60343 11360 60409 11383
rect 60495 11360 60577 11383
rect 60663 11360 60729 11383
rect 60343 11320 60352 11360
rect 60392 11320 60409 11360
rect 60495 11320 60516 11360
rect 60556 11320 60577 11360
rect 60663 11320 60680 11360
rect 60720 11320 60729 11360
rect 60343 11297 60409 11320
rect 60495 11297 60577 11320
rect 60663 11297 60729 11320
rect 60343 11278 60729 11297
rect 64343 11383 64729 11402
rect 64343 11360 64409 11383
rect 64495 11360 64577 11383
rect 64663 11360 64729 11383
rect 64343 11320 64352 11360
rect 64392 11320 64409 11360
rect 64495 11320 64516 11360
rect 64556 11320 64577 11360
rect 64663 11320 64680 11360
rect 64720 11320 64729 11360
rect 64343 11297 64409 11320
rect 64495 11297 64577 11320
rect 64663 11297 64729 11320
rect 64343 11278 64729 11297
rect 68343 11383 68729 11402
rect 68343 11360 68409 11383
rect 68495 11360 68577 11383
rect 68663 11360 68729 11383
rect 68343 11320 68352 11360
rect 68392 11320 68409 11360
rect 68495 11320 68516 11360
rect 68556 11320 68577 11360
rect 68663 11320 68680 11360
rect 68720 11320 68729 11360
rect 68343 11297 68409 11320
rect 68495 11297 68577 11320
rect 68663 11297 68729 11320
rect 68343 11278 68729 11297
rect 72316 11356 72409 11442
rect 72495 11356 72577 11442
rect 72663 11356 72756 11442
rect 72316 11274 72756 11356
rect 72316 11188 72409 11274
rect 72495 11188 72577 11274
rect 72663 11188 72756 11274
rect 72316 11106 72756 11188
rect 72316 11020 72409 11106
rect 72495 11020 72577 11106
rect 72663 11020 72756 11106
rect 72316 10890 72756 11020
rect 76316 13122 76756 13252
rect 76316 13036 76409 13122
rect 76495 13036 76577 13122
rect 76663 13036 76756 13122
rect 76316 12954 76756 13036
rect 76316 12868 76409 12954
rect 76495 12868 76577 12954
rect 76663 12868 76756 12954
rect 76316 12786 76756 12868
rect 76316 12700 76409 12786
rect 76495 12700 76577 12786
rect 76663 12700 76756 12786
rect 76316 12618 76756 12700
rect 76316 12532 76409 12618
rect 76495 12532 76577 12618
rect 76663 12532 76756 12618
rect 76316 12450 76756 12532
rect 76316 12364 76409 12450
rect 76495 12364 76577 12450
rect 76663 12364 76756 12450
rect 76316 12282 76756 12364
rect 76316 12196 76409 12282
rect 76495 12196 76577 12282
rect 76663 12196 76756 12282
rect 76316 12114 76756 12196
rect 76316 12028 76409 12114
rect 76495 12028 76577 12114
rect 76663 12028 76756 12114
rect 76316 11946 76756 12028
rect 76316 11860 76409 11946
rect 76495 11860 76577 11946
rect 76663 11860 76756 11946
rect 76316 11778 76756 11860
rect 76316 11692 76409 11778
rect 76495 11692 76577 11778
rect 76663 11692 76756 11778
rect 76316 11610 76756 11692
rect 76316 11524 76409 11610
rect 76495 11524 76577 11610
rect 76663 11524 76756 11610
rect 76316 11442 76756 11524
rect 76316 11356 76409 11442
rect 76495 11356 76577 11442
rect 76663 11356 76756 11442
rect 76316 11274 76756 11356
rect 76316 11188 76409 11274
rect 76495 11188 76577 11274
rect 76663 11188 76756 11274
rect 76316 11106 76756 11188
rect 76316 11020 76409 11106
rect 76495 11020 76577 11106
rect 76663 11020 76756 11106
rect 76316 10890 76756 11020
rect 80316 13122 80756 13252
rect 80316 13036 80409 13122
rect 80495 13036 80577 13122
rect 80663 13036 80756 13122
rect 80316 12954 80756 13036
rect 80316 12868 80409 12954
rect 80495 12868 80577 12954
rect 80663 12868 80756 12954
rect 80316 12786 80756 12868
rect 80316 12700 80409 12786
rect 80495 12700 80577 12786
rect 80663 12700 80756 12786
rect 80316 12618 80756 12700
rect 80316 12532 80409 12618
rect 80495 12532 80577 12618
rect 80663 12532 80756 12618
rect 80316 12450 80756 12532
rect 80316 12364 80409 12450
rect 80495 12364 80577 12450
rect 80663 12364 80756 12450
rect 80316 12282 80756 12364
rect 80316 12196 80409 12282
rect 80495 12196 80577 12282
rect 80663 12196 80756 12282
rect 80316 12114 80756 12196
rect 80316 12028 80409 12114
rect 80495 12028 80577 12114
rect 80663 12028 80756 12114
rect 80316 11946 80756 12028
rect 80316 11860 80409 11946
rect 80495 11860 80577 11946
rect 80663 11860 80756 11946
rect 80316 11778 80756 11860
rect 80316 11692 80409 11778
rect 80495 11692 80577 11778
rect 80663 11692 80756 11778
rect 80316 11610 80756 11692
rect 80316 11524 80409 11610
rect 80495 11524 80577 11610
rect 80663 11524 80756 11610
rect 80316 11442 80756 11524
rect 80316 11356 80409 11442
rect 80495 11356 80577 11442
rect 80663 11356 80756 11442
rect 80316 11274 80756 11356
rect 80316 11188 80409 11274
rect 80495 11188 80577 11274
rect 80663 11188 80756 11274
rect 80316 11106 80756 11188
rect 80316 11020 80409 11106
rect 80495 11020 80577 11106
rect 80663 11020 80756 11106
rect 80316 10890 80756 11020
rect 84316 13122 84756 13252
rect 84316 13036 84409 13122
rect 84495 13036 84577 13122
rect 84663 13036 84756 13122
rect 84316 12954 84756 13036
rect 84316 12868 84409 12954
rect 84495 12868 84577 12954
rect 84663 12868 84756 12954
rect 84316 12786 84756 12868
rect 84316 12700 84409 12786
rect 84495 12700 84577 12786
rect 84663 12700 84756 12786
rect 84316 12618 84756 12700
rect 84316 12532 84409 12618
rect 84495 12532 84577 12618
rect 84663 12532 84756 12618
rect 84316 12450 84756 12532
rect 84316 12364 84409 12450
rect 84495 12364 84577 12450
rect 84663 12364 84756 12450
rect 84316 12282 84756 12364
rect 84316 12196 84409 12282
rect 84495 12196 84577 12282
rect 84663 12196 84756 12282
rect 84316 12114 84756 12196
rect 84316 12028 84409 12114
rect 84495 12028 84577 12114
rect 84663 12028 84756 12114
rect 84316 11946 84756 12028
rect 84316 11860 84409 11946
rect 84495 11860 84577 11946
rect 84663 11860 84756 11946
rect 84316 11778 84756 11860
rect 84316 11692 84409 11778
rect 84495 11692 84577 11778
rect 84663 11692 84756 11778
rect 84316 11610 84756 11692
rect 84316 11524 84409 11610
rect 84495 11524 84577 11610
rect 84663 11524 84756 11610
rect 84316 11442 84756 11524
rect 84316 11356 84409 11442
rect 84495 11356 84577 11442
rect 84663 11356 84756 11442
rect 84316 11274 84756 11356
rect 84316 11188 84409 11274
rect 84495 11188 84577 11274
rect 84663 11188 84756 11274
rect 84316 11106 84756 11188
rect 84316 11020 84409 11106
rect 84495 11020 84577 11106
rect 84663 11020 84756 11106
rect 84316 10890 84756 11020
rect 88316 13122 88756 13252
rect 88316 13036 88409 13122
rect 88495 13036 88577 13122
rect 88663 13036 88756 13122
rect 88316 12954 88756 13036
rect 88316 12868 88409 12954
rect 88495 12868 88577 12954
rect 88663 12868 88756 12954
rect 88316 12786 88756 12868
rect 88316 12700 88409 12786
rect 88495 12700 88577 12786
rect 88663 12700 88756 12786
rect 88316 12618 88756 12700
rect 88316 12532 88409 12618
rect 88495 12532 88577 12618
rect 88663 12532 88756 12618
rect 88316 12450 88756 12532
rect 88316 12364 88409 12450
rect 88495 12364 88577 12450
rect 88663 12364 88756 12450
rect 88316 12282 88756 12364
rect 88316 12196 88409 12282
rect 88495 12196 88577 12282
rect 88663 12196 88756 12282
rect 88316 12114 88756 12196
rect 88316 12028 88409 12114
rect 88495 12028 88577 12114
rect 88663 12028 88756 12114
rect 88316 11946 88756 12028
rect 88316 11860 88409 11946
rect 88495 11860 88577 11946
rect 88663 11860 88756 11946
rect 88316 11778 88756 11860
rect 88316 11692 88409 11778
rect 88495 11692 88577 11778
rect 88663 11692 88756 11778
rect 88316 11610 88756 11692
rect 88316 11524 88409 11610
rect 88495 11524 88577 11610
rect 88663 11524 88756 11610
rect 88316 11442 88756 11524
rect 88316 11356 88409 11442
rect 88495 11356 88577 11442
rect 88663 11356 88756 11442
rect 88316 11274 88756 11356
rect 88316 11188 88409 11274
rect 88495 11188 88577 11274
rect 88663 11188 88756 11274
rect 88316 11106 88756 11188
rect 88316 11020 88409 11106
rect 88495 11020 88577 11106
rect 88663 11020 88756 11106
rect 88316 10890 88756 11020
rect 92316 13122 92756 13252
rect 92316 13036 92409 13122
rect 92495 13036 92577 13122
rect 92663 13036 92756 13122
rect 92316 12954 92756 13036
rect 92316 12868 92409 12954
rect 92495 12868 92577 12954
rect 92663 12868 92756 12954
rect 92316 12786 92756 12868
rect 92316 12700 92409 12786
rect 92495 12700 92577 12786
rect 92663 12700 92756 12786
rect 92316 12618 92756 12700
rect 92316 12532 92409 12618
rect 92495 12532 92577 12618
rect 92663 12532 92756 12618
rect 92316 12450 92756 12532
rect 92316 12364 92409 12450
rect 92495 12364 92577 12450
rect 92663 12364 92756 12450
rect 92316 12282 92756 12364
rect 92316 12196 92409 12282
rect 92495 12196 92577 12282
rect 92663 12196 92756 12282
rect 92316 12114 92756 12196
rect 92316 12028 92409 12114
rect 92495 12028 92577 12114
rect 92663 12028 92756 12114
rect 92316 11946 92756 12028
rect 92316 11860 92409 11946
rect 92495 11860 92577 11946
rect 92663 11860 92756 11946
rect 92316 11778 92756 11860
rect 92316 11692 92409 11778
rect 92495 11692 92577 11778
rect 92663 11692 92756 11778
rect 92316 11610 92756 11692
rect 92316 11524 92409 11610
rect 92495 11524 92577 11610
rect 92663 11524 92756 11610
rect 92316 11442 92756 11524
rect 92316 11356 92409 11442
rect 92495 11356 92577 11442
rect 92663 11356 92756 11442
rect 92316 11274 92756 11356
rect 92316 11188 92409 11274
rect 92495 11188 92577 11274
rect 92663 11188 92756 11274
rect 92316 11106 92756 11188
rect 92316 11020 92409 11106
rect 92495 11020 92577 11106
rect 92663 11020 92756 11106
rect 92316 10890 92756 11020
rect 96316 13122 96756 13252
rect 96316 13036 96409 13122
rect 96495 13036 96577 13122
rect 96663 13036 96756 13122
rect 96316 12954 96756 13036
rect 96316 12868 96409 12954
rect 96495 12868 96577 12954
rect 96663 12868 96756 12954
rect 96316 12786 96756 12868
rect 96316 12700 96409 12786
rect 96495 12700 96577 12786
rect 96663 12700 96756 12786
rect 96316 12618 96756 12700
rect 96316 12532 96409 12618
rect 96495 12532 96577 12618
rect 96663 12532 96756 12618
rect 96316 12450 96756 12532
rect 96316 12364 96409 12450
rect 96495 12364 96577 12450
rect 96663 12364 96756 12450
rect 96316 12282 96756 12364
rect 96316 12196 96409 12282
rect 96495 12196 96577 12282
rect 96663 12196 96756 12282
rect 96316 12114 96756 12196
rect 96316 12028 96409 12114
rect 96495 12028 96577 12114
rect 96663 12028 96756 12114
rect 96316 11946 96756 12028
rect 96316 11860 96409 11946
rect 96495 11860 96577 11946
rect 96663 11860 96756 11946
rect 96316 11778 96756 11860
rect 96316 11692 96409 11778
rect 96495 11692 96577 11778
rect 96663 11692 96756 11778
rect 96316 11610 96756 11692
rect 96316 11524 96409 11610
rect 96495 11524 96577 11610
rect 96663 11524 96756 11610
rect 96316 11442 96756 11524
rect 96316 11356 96409 11442
rect 96495 11356 96577 11442
rect 96663 11356 96756 11442
rect 96316 11274 96756 11356
rect 96316 11188 96409 11274
rect 96495 11188 96577 11274
rect 96663 11188 96756 11274
rect 96316 11106 96756 11188
rect 96316 11020 96409 11106
rect 96495 11020 96577 11106
rect 96663 11020 96756 11106
rect 96316 10890 96756 11020
rect 3103 10627 3489 10646
rect 3103 10604 3169 10627
rect 3255 10604 3337 10627
rect 3423 10604 3489 10627
rect 3103 10564 3112 10604
rect 3152 10564 3169 10604
rect 3255 10564 3276 10604
rect 3316 10564 3337 10604
rect 3423 10564 3440 10604
rect 3480 10564 3489 10604
rect 3103 10541 3169 10564
rect 3255 10541 3337 10564
rect 3423 10541 3489 10564
rect 3103 10522 3489 10541
rect 7103 10627 7489 10646
rect 7103 10604 7169 10627
rect 7255 10604 7337 10627
rect 7423 10604 7489 10627
rect 7103 10564 7112 10604
rect 7152 10564 7169 10604
rect 7255 10564 7276 10604
rect 7316 10564 7337 10604
rect 7423 10564 7440 10604
rect 7480 10564 7489 10604
rect 7103 10541 7169 10564
rect 7255 10541 7337 10564
rect 7423 10541 7489 10564
rect 7103 10522 7489 10541
rect 11103 10627 11489 10646
rect 11103 10604 11169 10627
rect 11255 10604 11337 10627
rect 11423 10604 11489 10627
rect 11103 10564 11112 10604
rect 11152 10564 11169 10604
rect 11255 10564 11276 10604
rect 11316 10564 11337 10604
rect 11423 10564 11440 10604
rect 11480 10564 11489 10604
rect 11103 10541 11169 10564
rect 11255 10541 11337 10564
rect 11423 10541 11489 10564
rect 11103 10522 11489 10541
rect 15103 10627 15489 10646
rect 15103 10604 15169 10627
rect 15255 10604 15337 10627
rect 15423 10604 15489 10627
rect 15103 10564 15112 10604
rect 15152 10564 15169 10604
rect 15255 10564 15276 10604
rect 15316 10564 15337 10604
rect 15423 10564 15440 10604
rect 15480 10564 15489 10604
rect 15103 10541 15169 10564
rect 15255 10541 15337 10564
rect 15423 10541 15489 10564
rect 15103 10522 15489 10541
rect 19103 10627 19489 10646
rect 19103 10604 19169 10627
rect 19255 10604 19337 10627
rect 19423 10604 19489 10627
rect 19103 10564 19112 10604
rect 19152 10564 19169 10604
rect 19255 10564 19276 10604
rect 19316 10564 19337 10604
rect 19423 10564 19440 10604
rect 19480 10564 19489 10604
rect 19103 10541 19169 10564
rect 19255 10541 19337 10564
rect 19423 10541 19489 10564
rect 19103 10522 19489 10541
rect 23103 10627 23489 10646
rect 23103 10604 23169 10627
rect 23255 10604 23337 10627
rect 23423 10604 23489 10627
rect 23103 10564 23112 10604
rect 23152 10564 23169 10604
rect 23255 10564 23276 10604
rect 23316 10564 23337 10604
rect 23423 10564 23440 10604
rect 23480 10564 23489 10604
rect 23103 10541 23169 10564
rect 23255 10541 23337 10564
rect 23423 10541 23489 10564
rect 23103 10522 23489 10541
rect 27103 10627 27489 10646
rect 27103 10604 27169 10627
rect 27255 10604 27337 10627
rect 27423 10604 27489 10627
rect 27103 10564 27112 10604
rect 27152 10564 27169 10604
rect 27255 10564 27276 10604
rect 27316 10564 27337 10604
rect 27423 10564 27440 10604
rect 27480 10564 27489 10604
rect 27103 10541 27169 10564
rect 27255 10541 27337 10564
rect 27423 10541 27489 10564
rect 27103 10522 27489 10541
rect 31103 10627 31489 10646
rect 31103 10604 31169 10627
rect 31255 10604 31337 10627
rect 31423 10604 31489 10627
rect 31103 10564 31112 10604
rect 31152 10564 31169 10604
rect 31255 10564 31276 10604
rect 31316 10564 31337 10604
rect 31423 10564 31440 10604
rect 31480 10564 31489 10604
rect 31103 10541 31169 10564
rect 31255 10541 31337 10564
rect 31423 10541 31489 10564
rect 31103 10522 31489 10541
rect 35103 10627 35489 10646
rect 35103 10604 35169 10627
rect 35255 10604 35337 10627
rect 35423 10604 35489 10627
rect 35103 10564 35112 10604
rect 35152 10564 35169 10604
rect 35255 10564 35276 10604
rect 35316 10564 35337 10604
rect 35423 10564 35440 10604
rect 35480 10564 35489 10604
rect 35103 10541 35169 10564
rect 35255 10541 35337 10564
rect 35423 10541 35489 10564
rect 35103 10522 35489 10541
rect 39103 10627 39489 10646
rect 39103 10604 39169 10627
rect 39255 10604 39337 10627
rect 39423 10604 39489 10627
rect 39103 10564 39112 10604
rect 39152 10564 39169 10604
rect 39255 10564 39276 10604
rect 39316 10564 39337 10604
rect 39423 10564 39440 10604
rect 39480 10564 39489 10604
rect 39103 10541 39169 10564
rect 39255 10541 39337 10564
rect 39423 10541 39489 10564
rect 39103 10522 39489 10541
rect 43103 10627 43489 10646
rect 43103 10604 43169 10627
rect 43255 10604 43337 10627
rect 43423 10604 43489 10627
rect 43103 10564 43112 10604
rect 43152 10564 43169 10604
rect 43255 10564 43276 10604
rect 43316 10564 43337 10604
rect 43423 10564 43440 10604
rect 43480 10564 43489 10604
rect 43103 10541 43169 10564
rect 43255 10541 43337 10564
rect 43423 10541 43489 10564
rect 43103 10522 43489 10541
rect 47103 10627 47489 10646
rect 47103 10604 47169 10627
rect 47255 10604 47337 10627
rect 47423 10604 47489 10627
rect 47103 10564 47112 10604
rect 47152 10564 47169 10604
rect 47255 10564 47276 10604
rect 47316 10564 47337 10604
rect 47423 10564 47440 10604
rect 47480 10564 47489 10604
rect 47103 10541 47169 10564
rect 47255 10541 47337 10564
rect 47423 10541 47489 10564
rect 47103 10522 47489 10541
rect 51103 10627 51489 10646
rect 51103 10604 51169 10627
rect 51255 10604 51337 10627
rect 51423 10604 51489 10627
rect 51103 10564 51112 10604
rect 51152 10564 51169 10604
rect 51255 10564 51276 10604
rect 51316 10564 51337 10604
rect 51423 10564 51440 10604
rect 51480 10564 51489 10604
rect 51103 10541 51169 10564
rect 51255 10541 51337 10564
rect 51423 10541 51489 10564
rect 51103 10522 51489 10541
rect 55103 10627 55489 10646
rect 55103 10604 55169 10627
rect 55255 10604 55337 10627
rect 55423 10604 55489 10627
rect 55103 10564 55112 10604
rect 55152 10564 55169 10604
rect 55255 10564 55276 10604
rect 55316 10564 55337 10604
rect 55423 10564 55440 10604
rect 55480 10564 55489 10604
rect 55103 10541 55169 10564
rect 55255 10541 55337 10564
rect 55423 10541 55489 10564
rect 55103 10522 55489 10541
rect 59103 10627 59489 10646
rect 59103 10604 59169 10627
rect 59255 10604 59337 10627
rect 59423 10604 59489 10627
rect 59103 10564 59112 10604
rect 59152 10564 59169 10604
rect 59255 10564 59276 10604
rect 59316 10564 59337 10604
rect 59423 10564 59440 10604
rect 59480 10564 59489 10604
rect 59103 10541 59169 10564
rect 59255 10541 59337 10564
rect 59423 10541 59489 10564
rect 59103 10522 59489 10541
rect 63103 10627 63489 10646
rect 63103 10604 63169 10627
rect 63255 10604 63337 10627
rect 63423 10604 63489 10627
rect 63103 10564 63112 10604
rect 63152 10564 63169 10604
rect 63255 10564 63276 10604
rect 63316 10564 63337 10604
rect 63423 10564 63440 10604
rect 63480 10564 63489 10604
rect 63103 10541 63169 10564
rect 63255 10541 63337 10564
rect 63423 10541 63489 10564
rect 63103 10522 63489 10541
rect 67103 10627 67489 10646
rect 67103 10604 67169 10627
rect 67255 10604 67337 10627
rect 67423 10604 67489 10627
rect 67103 10564 67112 10604
rect 67152 10564 67169 10604
rect 67255 10564 67276 10604
rect 67316 10564 67337 10604
rect 67423 10564 67440 10604
rect 67480 10564 67489 10604
rect 67103 10541 67169 10564
rect 67255 10541 67337 10564
rect 67423 10541 67489 10564
rect 67103 10522 67489 10541
rect 75076 10246 75516 10376
rect 75076 10160 75169 10246
rect 75255 10160 75337 10246
rect 75423 10160 75516 10246
rect 75076 10078 75516 10160
rect 75076 9992 75169 10078
rect 75255 9992 75337 10078
rect 75423 9992 75516 10078
rect 75076 9910 75516 9992
rect 4343 9871 4729 9890
rect 4343 9848 4409 9871
rect 4495 9848 4577 9871
rect 4663 9848 4729 9871
rect 4343 9808 4352 9848
rect 4392 9808 4409 9848
rect 4495 9808 4516 9848
rect 4556 9808 4577 9848
rect 4663 9808 4680 9848
rect 4720 9808 4729 9848
rect 4343 9785 4409 9808
rect 4495 9785 4577 9808
rect 4663 9785 4729 9808
rect 4343 9766 4729 9785
rect 8343 9871 8729 9890
rect 8343 9848 8409 9871
rect 8495 9848 8577 9871
rect 8663 9848 8729 9871
rect 8343 9808 8352 9848
rect 8392 9808 8409 9848
rect 8495 9808 8516 9848
rect 8556 9808 8577 9848
rect 8663 9808 8680 9848
rect 8720 9808 8729 9848
rect 8343 9785 8409 9808
rect 8495 9785 8577 9808
rect 8663 9785 8729 9808
rect 8343 9766 8729 9785
rect 12343 9871 12729 9890
rect 12343 9848 12409 9871
rect 12495 9848 12577 9871
rect 12663 9848 12729 9871
rect 12343 9808 12352 9848
rect 12392 9808 12409 9848
rect 12495 9808 12516 9848
rect 12556 9808 12577 9848
rect 12663 9808 12680 9848
rect 12720 9808 12729 9848
rect 12343 9785 12409 9808
rect 12495 9785 12577 9808
rect 12663 9785 12729 9808
rect 12343 9766 12729 9785
rect 16343 9871 16729 9890
rect 16343 9848 16409 9871
rect 16495 9848 16577 9871
rect 16663 9848 16729 9871
rect 16343 9808 16352 9848
rect 16392 9808 16409 9848
rect 16495 9808 16516 9848
rect 16556 9808 16577 9848
rect 16663 9808 16680 9848
rect 16720 9808 16729 9848
rect 16343 9785 16409 9808
rect 16495 9785 16577 9808
rect 16663 9785 16729 9808
rect 16343 9766 16729 9785
rect 20343 9871 20729 9890
rect 20343 9848 20409 9871
rect 20495 9848 20577 9871
rect 20663 9848 20729 9871
rect 20343 9808 20352 9848
rect 20392 9808 20409 9848
rect 20495 9808 20516 9848
rect 20556 9808 20577 9848
rect 20663 9808 20680 9848
rect 20720 9808 20729 9848
rect 20343 9785 20409 9808
rect 20495 9785 20577 9808
rect 20663 9785 20729 9808
rect 20343 9766 20729 9785
rect 24343 9871 24729 9890
rect 24343 9848 24409 9871
rect 24495 9848 24577 9871
rect 24663 9848 24729 9871
rect 24343 9808 24352 9848
rect 24392 9808 24409 9848
rect 24495 9808 24516 9848
rect 24556 9808 24577 9848
rect 24663 9808 24680 9848
rect 24720 9808 24729 9848
rect 24343 9785 24409 9808
rect 24495 9785 24577 9808
rect 24663 9785 24729 9808
rect 24343 9766 24729 9785
rect 28343 9871 28729 9890
rect 28343 9848 28409 9871
rect 28495 9848 28577 9871
rect 28663 9848 28729 9871
rect 28343 9808 28352 9848
rect 28392 9808 28409 9848
rect 28495 9808 28516 9848
rect 28556 9808 28577 9848
rect 28663 9808 28680 9848
rect 28720 9808 28729 9848
rect 28343 9785 28409 9808
rect 28495 9785 28577 9808
rect 28663 9785 28729 9808
rect 28343 9766 28729 9785
rect 32343 9871 32729 9890
rect 32343 9848 32409 9871
rect 32495 9848 32577 9871
rect 32663 9848 32729 9871
rect 32343 9808 32352 9848
rect 32392 9808 32409 9848
rect 32495 9808 32516 9848
rect 32556 9808 32577 9848
rect 32663 9808 32680 9848
rect 32720 9808 32729 9848
rect 32343 9785 32409 9808
rect 32495 9785 32577 9808
rect 32663 9785 32729 9808
rect 32343 9766 32729 9785
rect 36343 9871 36729 9890
rect 36343 9848 36409 9871
rect 36495 9848 36577 9871
rect 36663 9848 36729 9871
rect 36343 9808 36352 9848
rect 36392 9808 36409 9848
rect 36495 9808 36516 9848
rect 36556 9808 36577 9848
rect 36663 9808 36680 9848
rect 36720 9808 36729 9848
rect 36343 9785 36409 9808
rect 36495 9785 36577 9808
rect 36663 9785 36729 9808
rect 36343 9766 36729 9785
rect 40343 9871 40729 9890
rect 40343 9848 40409 9871
rect 40495 9848 40577 9871
rect 40663 9848 40729 9871
rect 40343 9808 40352 9848
rect 40392 9808 40409 9848
rect 40495 9808 40516 9848
rect 40556 9808 40577 9848
rect 40663 9808 40680 9848
rect 40720 9808 40729 9848
rect 40343 9785 40409 9808
rect 40495 9785 40577 9808
rect 40663 9785 40729 9808
rect 40343 9766 40729 9785
rect 44343 9871 44729 9890
rect 44343 9848 44409 9871
rect 44495 9848 44577 9871
rect 44663 9848 44729 9871
rect 44343 9808 44352 9848
rect 44392 9808 44409 9848
rect 44495 9808 44516 9848
rect 44556 9808 44577 9848
rect 44663 9808 44680 9848
rect 44720 9808 44729 9848
rect 44343 9785 44409 9808
rect 44495 9785 44577 9808
rect 44663 9785 44729 9808
rect 44343 9766 44729 9785
rect 48343 9871 48729 9890
rect 48343 9848 48409 9871
rect 48495 9848 48577 9871
rect 48663 9848 48729 9871
rect 48343 9808 48352 9848
rect 48392 9808 48409 9848
rect 48495 9808 48516 9848
rect 48556 9808 48577 9848
rect 48663 9808 48680 9848
rect 48720 9808 48729 9848
rect 48343 9785 48409 9808
rect 48495 9785 48577 9808
rect 48663 9785 48729 9808
rect 48343 9766 48729 9785
rect 52343 9871 52729 9890
rect 52343 9848 52409 9871
rect 52495 9848 52577 9871
rect 52663 9848 52729 9871
rect 52343 9808 52352 9848
rect 52392 9808 52409 9848
rect 52495 9808 52516 9848
rect 52556 9808 52577 9848
rect 52663 9808 52680 9848
rect 52720 9808 52729 9848
rect 52343 9785 52409 9808
rect 52495 9785 52577 9808
rect 52663 9785 52729 9808
rect 52343 9766 52729 9785
rect 56343 9871 56729 9890
rect 56343 9848 56409 9871
rect 56495 9848 56577 9871
rect 56663 9848 56729 9871
rect 56343 9808 56352 9848
rect 56392 9808 56409 9848
rect 56495 9808 56516 9848
rect 56556 9808 56577 9848
rect 56663 9808 56680 9848
rect 56720 9808 56729 9848
rect 56343 9785 56409 9808
rect 56495 9785 56577 9808
rect 56663 9785 56729 9808
rect 56343 9766 56729 9785
rect 60343 9871 60729 9890
rect 60343 9848 60409 9871
rect 60495 9848 60577 9871
rect 60663 9848 60729 9871
rect 60343 9808 60352 9848
rect 60392 9808 60409 9848
rect 60495 9808 60516 9848
rect 60556 9808 60577 9848
rect 60663 9808 60680 9848
rect 60720 9808 60729 9848
rect 60343 9785 60409 9808
rect 60495 9785 60577 9808
rect 60663 9785 60729 9808
rect 60343 9766 60729 9785
rect 64343 9871 64729 9890
rect 64343 9848 64409 9871
rect 64495 9848 64577 9871
rect 64663 9848 64729 9871
rect 64343 9808 64352 9848
rect 64392 9808 64409 9848
rect 64495 9808 64516 9848
rect 64556 9808 64577 9848
rect 64663 9808 64680 9848
rect 64720 9808 64729 9848
rect 64343 9785 64409 9808
rect 64495 9785 64577 9808
rect 64663 9785 64729 9808
rect 64343 9766 64729 9785
rect 68343 9871 68729 9890
rect 68343 9848 68409 9871
rect 68495 9848 68577 9871
rect 68663 9848 68729 9871
rect 68343 9808 68352 9848
rect 68392 9808 68409 9848
rect 68495 9808 68516 9848
rect 68556 9808 68577 9848
rect 68663 9808 68680 9848
rect 68720 9808 68729 9848
rect 68343 9785 68409 9808
rect 68495 9785 68577 9808
rect 68663 9785 68729 9808
rect 68343 9766 68729 9785
rect 75076 9824 75169 9910
rect 75255 9824 75337 9910
rect 75423 9824 75516 9910
rect 75076 9742 75516 9824
rect 75076 9656 75169 9742
rect 75255 9656 75337 9742
rect 75423 9656 75516 9742
rect 75076 9574 75516 9656
rect 75076 9488 75169 9574
rect 75255 9488 75337 9574
rect 75423 9488 75516 9574
rect 75076 9406 75516 9488
rect 75076 9320 75169 9406
rect 75255 9320 75337 9406
rect 75423 9320 75516 9406
rect 75076 9238 75516 9320
rect 75076 9152 75169 9238
rect 75255 9152 75337 9238
rect 75423 9152 75516 9238
rect 3103 9115 3489 9134
rect 3103 9092 3169 9115
rect 3255 9092 3337 9115
rect 3423 9092 3489 9115
rect 3103 9052 3112 9092
rect 3152 9052 3169 9092
rect 3255 9052 3276 9092
rect 3316 9052 3337 9092
rect 3423 9052 3440 9092
rect 3480 9052 3489 9092
rect 3103 9029 3169 9052
rect 3255 9029 3337 9052
rect 3423 9029 3489 9052
rect 3103 9010 3489 9029
rect 7103 9115 7489 9134
rect 7103 9092 7169 9115
rect 7255 9092 7337 9115
rect 7423 9092 7489 9115
rect 7103 9052 7112 9092
rect 7152 9052 7169 9092
rect 7255 9052 7276 9092
rect 7316 9052 7337 9092
rect 7423 9052 7440 9092
rect 7480 9052 7489 9092
rect 7103 9029 7169 9052
rect 7255 9029 7337 9052
rect 7423 9029 7489 9052
rect 7103 9010 7489 9029
rect 11103 9115 11489 9134
rect 11103 9092 11169 9115
rect 11255 9092 11337 9115
rect 11423 9092 11489 9115
rect 11103 9052 11112 9092
rect 11152 9052 11169 9092
rect 11255 9052 11276 9092
rect 11316 9052 11337 9092
rect 11423 9052 11440 9092
rect 11480 9052 11489 9092
rect 11103 9029 11169 9052
rect 11255 9029 11337 9052
rect 11423 9029 11489 9052
rect 11103 9010 11489 9029
rect 15103 9115 15489 9134
rect 15103 9092 15169 9115
rect 15255 9092 15337 9115
rect 15423 9092 15489 9115
rect 15103 9052 15112 9092
rect 15152 9052 15169 9092
rect 15255 9052 15276 9092
rect 15316 9052 15337 9092
rect 15423 9052 15440 9092
rect 15480 9052 15489 9092
rect 15103 9029 15169 9052
rect 15255 9029 15337 9052
rect 15423 9029 15489 9052
rect 15103 9010 15489 9029
rect 19103 9115 19489 9134
rect 19103 9092 19169 9115
rect 19255 9092 19337 9115
rect 19423 9092 19489 9115
rect 19103 9052 19112 9092
rect 19152 9052 19169 9092
rect 19255 9052 19276 9092
rect 19316 9052 19337 9092
rect 19423 9052 19440 9092
rect 19480 9052 19489 9092
rect 19103 9029 19169 9052
rect 19255 9029 19337 9052
rect 19423 9029 19489 9052
rect 19103 9010 19489 9029
rect 23103 9115 23489 9134
rect 23103 9092 23169 9115
rect 23255 9092 23337 9115
rect 23423 9092 23489 9115
rect 23103 9052 23112 9092
rect 23152 9052 23169 9092
rect 23255 9052 23276 9092
rect 23316 9052 23337 9092
rect 23423 9052 23440 9092
rect 23480 9052 23489 9092
rect 23103 9029 23169 9052
rect 23255 9029 23337 9052
rect 23423 9029 23489 9052
rect 23103 9010 23489 9029
rect 27103 9115 27489 9134
rect 27103 9092 27169 9115
rect 27255 9092 27337 9115
rect 27423 9092 27489 9115
rect 27103 9052 27112 9092
rect 27152 9052 27169 9092
rect 27255 9052 27276 9092
rect 27316 9052 27337 9092
rect 27423 9052 27440 9092
rect 27480 9052 27489 9092
rect 27103 9029 27169 9052
rect 27255 9029 27337 9052
rect 27423 9029 27489 9052
rect 27103 9010 27489 9029
rect 31103 9115 31489 9134
rect 31103 9092 31169 9115
rect 31255 9092 31337 9115
rect 31423 9092 31489 9115
rect 31103 9052 31112 9092
rect 31152 9052 31169 9092
rect 31255 9052 31276 9092
rect 31316 9052 31337 9092
rect 31423 9052 31440 9092
rect 31480 9052 31489 9092
rect 31103 9029 31169 9052
rect 31255 9029 31337 9052
rect 31423 9029 31489 9052
rect 31103 9010 31489 9029
rect 35103 9115 35489 9134
rect 35103 9092 35169 9115
rect 35255 9092 35337 9115
rect 35423 9092 35489 9115
rect 35103 9052 35112 9092
rect 35152 9052 35169 9092
rect 35255 9052 35276 9092
rect 35316 9052 35337 9092
rect 35423 9052 35440 9092
rect 35480 9052 35489 9092
rect 35103 9029 35169 9052
rect 35255 9029 35337 9052
rect 35423 9029 35489 9052
rect 35103 9010 35489 9029
rect 39103 9115 39489 9134
rect 39103 9092 39169 9115
rect 39255 9092 39337 9115
rect 39423 9092 39489 9115
rect 39103 9052 39112 9092
rect 39152 9052 39169 9092
rect 39255 9052 39276 9092
rect 39316 9052 39337 9092
rect 39423 9052 39440 9092
rect 39480 9052 39489 9092
rect 39103 9029 39169 9052
rect 39255 9029 39337 9052
rect 39423 9029 39489 9052
rect 39103 9010 39489 9029
rect 43103 9115 43489 9134
rect 43103 9092 43169 9115
rect 43255 9092 43337 9115
rect 43423 9092 43489 9115
rect 43103 9052 43112 9092
rect 43152 9052 43169 9092
rect 43255 9052 43276 9092
rect 43316 9052 43337 9092
rect 43423 9052 43440 9092
rect 43480 9052 43489 9092
rect 43103 9029 43169 9052
rect 43255 9029 43337 9052
rect 43423 9029 43489 9052
rect 43103 9010 43489 9029
rect 47103 9115 47489 9134
rect 47103 9092 47169 9115
rect 47255 9092 47337 9115
rect 47423 9092 47489 9115
rect 47103 9052 47112 9092
rect 47152 9052 47169 9092
rect 47255 9052 47276 9092
rect 47316 9052 47337 9092
rect 47423 9052 47440 9092
rect 47480 9052 47489 9092
rect 47103 9029 47169 9052
rect 47255 9029 47337 9052
rect 47423 9029 47489 9052
rect 47103 9010 47489 9029
rect 51103 9115 51489 9134
rect 51103 9092 51169 9115
rect 51255 9092 51337 9115
rect 51423 9092 51489 9115
rect 51103 9052 51112 9092
rect 51152 9052 51169 9092
rect 51255 9052 51276 9092
rect 51316 9052 51337 9092
rect 51423 9052 51440 9092
rect 51480 9052 51489 9092
rect 51103 9029 51169 9052
rect 51255 9029 51337 9052
rect 51423 9029 51489 9052
rect 51103 9010 51489 9029
rect 55103 9115 55489 9134
rect 55103 9092 55169 9115
rect 55255 9092 55337 9115
rect 55423 9092 55489 9115
rect 55103 9052 55112 9092
rect 55152 9052 55169 9092
rect 55255 9052 55276 9092
rect 55316 9052 55337 9092
rect 55423 9052 55440 9092
rect 55480 9052 55489 9092
rect 55103 9029 55169 9052
rect 55255 9029 55337 9052
rect 55423 9029 55489 9052
rect 55103 9010 55489 9029
rect 59103 9115 59489 9134
rect 59103 9092 59169 9115
rect 59255 9092 59337 9115
rect 59423 9092 59489 9115
rect 59103 9052 59112 9092
rect 59152 9052 59169 9092
rect 59255 9052 59276 9092
rect 59316 9052 59337 9092
rect 59423 9052 59440 9092
rect 59480 9052 59489 9092
rect 59103 9029 59169 9052
rect 59255 9029 59337 9052
rect 59423 9029 59489 9052
rect 59103 9010 59489 9029
rect 63103 9115 63489 9134
rect 63103 9092 63169 9115
rect 63255 9092 63337 9115
rect 63423 9092 63489 9115
rect 63103 9052 63112 9092
rect 63152 9052 63169 9092
rect 63255 9052 63276 9092
rect 63316 9052 63337 9092
rect 63423 9052 63440 9092
rect 63480 9052 63489 9092
rect 63103 9029 63169 9052
rect 63255 9029 63337 9052
rect 63423 9029 63489 9052
rect 63103 9010 63489 9029
rect 67103 9115 67489 9134
rect 67103 9092 67169 9115
rect 67255 9092 67337 9115
rect 67423 9092 67489 9115
rect 67103 9052 67112 9092
rect 67152 9052 67169 9092
rect 67255 9052 67276 9092
rect 67316 9052 67337 9092
rect 67423 9052 67440 9092
rect 67480 9052 67489 9092
rect 67103 9029 67169 9052
rect 67255 9029 67337 9052
rect 67423 9029 67489 9052
rect 67103 9010 67489 9029
rect 75076 9070 75516 9152
rect 75076 8984 75169 9070
rect 75255 8984 75337 9070
rect 75423 8984 75516 9070
rect 75076 8902 75516 8984
rect 75076 8816 75169 8902
rect 75255 8816 75337 8902
rect 75423 8816 75516 8902
rect 75076 8734 75516 8816
rect 75076 8648 75169 8734
rect 75255 8648 75337 8734
rect 75423 8648 75516 8734
rect 75076 8566 75516 8648
rect 75076 8480 75169 8566
rect 75255 8480 75337 8566
rect 75423 8480 75516 8566
rect 75076 8398 75516 8480
rect 4343 8359 4729 8378
rect 4343 8336 4409 8359
rect 4495 8336 4577 8359
rect 4663 8336 4729 8359
rect 4343 8296 4352 8336
rect 4392 8296 4409 8336
rect 4495 8296 4516 8336
rect 4556 8296 4577 8336
rect 4663 8296 4680 8336
rect 4720 8296 4729 8336
rect 4343 8273 4409 8296
rect 4495 8273 4577 8296
rect 4663 8273 4729 8296
rect 4343 8254 4729 8273
rect 8343 8359 8729 8378
rect 8343 8336 8409 8359
rect 8495 8336 8577 8359
rect 8663 8336 8729 8359
rect 8343 8296 8352 8336
rect 8392 8296 8409 8336
rect 8495 8296 8516 8336
rect 8556 8296 8577 8336
rect 8663 8296 8680 8336
rect 8720 8296 8729 8336
rect 8343 8273 8409 8296
rect 8495 8273 8577 8296
rect 8663 8273 8729 8296
rect 8343 8254 8729 8273
rect 12343 8359 12729 8378
rect 12343 8336 12409 8359
rect 12495 8336 12577 8359
rect 12663 8336 12729 8359
rect 12343 8296 12352 8336
rect 12392 8296 12409 8336
rect 12495 8296 12516 8336
rect 12556 8296 12577 8336
rect 12663 8296 12680 8336
rect 12720 8296 12729 8336
rect 12343 8273 12409 8296
rect 12495 8273 12577 8296
rect 12663 8273 12729 8296
rect 12343 8254 12729 8273
rect 16343 8359 16729 8378
rect 16343 8336 16409 8359
rect 16495 8336 16577 8359
rect 16663 8336 16729 8359
rect 16343 8296 16352 8336
rect 16392 8296 16409 8336
rect 16495 8296 16516 8336
rect 16556 8296 16577 8336
rect 16663 8296 16680 8336
rect 16720 8296 16729 8336
rect 16343 8273 16409 8296
rect 16495 8273 16577 8296
rect 16663 8273 16729 8296
rect 16343 8254 16729 8273
rect 20343 8359 20729 8378
rect 20343 8336 20409 8359
rect 20495 8336 20577 8359
rect 20663 8336 20729 8359
rect 20343 8296 20352 8336
rect 20392 8296 20409 8336
rect 20495 8296 20516 8336
rect 20556 8296 20577 8336
rect 20663 8296 20680 8336
rect 20720 8296 20729 8336
rect 20343 8273 20409 8296
rect 20495 8273 20577 8296
rect 20663 8273 20729 8296
rect 20343 8254 20729 8273
rect 24343 8359 24729 8378
rect 24343 8336 24409 8359
rect 24495 8336 24577 8359
rect 24663 8336 24729 8359
rect 24343 8296 24352 8336
rect 24392 8296 24409 8336
rect 24495 8296 24516 8336
rect 24556 8296 24577 8336
rect 24663 8296 24680 8336
rect 24720 8296 24729 8336
rect 24343 8273 24409 8296
rect 24495 8273 24577 8296
rect 24663 8273 24729 8296
rect 24343 8254 24729 8273
rect 28343 8359 28729 8378
rect 28343 8336 28409 8359
rect 28495 8336 28577 8359
rect 28663 8336 28729 8359
rect 28343 8296 28352 8336
rect 28392 8296 28409 8336
rect 28495 8296 28516 8336
rect 28556 8296 28577 8336
rect 28663 8296 28680 8336
rect 28720 8296 28729 8336
rect 28343 8273 28409 8296
rect 28495 8273 28577 8296
rect 28663 8273 28729 8296
rect 28343 8254 28729 8273
rect 32343 8359 32729 8378
rect 32343 8336 32409 8359
rect 32495 8336 32577 8359
rect 32663 8336 32729 8359
rect 32343 8296 32352 8336
rect 32392 8296 32409 8336
rect 32495 8296 32516 8336
rect 32556 8296 32577 8336
rect 32663 8296 32680 8336
rect 32720 8296 32729 8336
rect 32343 8273 32409 8296
rect 32495 8273 32577 8296
rect 32663 8273 32729 8296
rect 32343 8254 32729 8273
rect 36343 8359 36729 8378
rect 36343 8336 36409 8359
rect 36495 8336 36577 8359
rect 36663 8336 36729 8359
rect 36343 8296 36352 8336
rect 36392 8296 36409 8336
rect 36495 8296 36516 8336
rect 36556 8296 36577 8336
rect 36663 8296 36680 8336
rect 36720 8296 36729 8336
rect 36343 8273 36409 8296
rect 36495 8273 36577 8296
rect 36663 8273 36729 8296
rect 36343 8254 36729 8273
rect 40343 8359 40729 8378
rect 40343 8336 40409 8359
rect 40495 8336 40577 8359
rect 40663 8336 40729 8359
rect 40343 8296 40352 8336
rect 40392 8296 40409 8336
rect 40495 8296 40516 8336
rect 40556 8296 40577 8336
rect 40663 8296 40680 8336
rect 40720 8296 40729 8336
rect 40343 8273 40409 8296
rect 40495 8273 40577 8296
rect 40663 8273 40729 8296
rect 40343 8254 40729 8273
rect 44343 8359 44729 8378
rect 44343 8336 44409 8359
rect 44495 8336 44577 8359
rect 44663 8336 44729 8359
rect 44343 8296 44352 8336
rect 44392 8296 44409 8336
rect 44495 8296 44516 8336
rect 44556 8296 44577 8336
rect 44663 8296 44680 8336
rect 44720 8296 44729 8336
rect 44343 8273 44409 8296
rect 44495 8273 44577 8296
rect 44663 8273 44729 8296
rect 44343 8254 44729 8273
rect 48343 8359 48729 8378
rect 48343 8336 48409 8359
rect 48495 8336 48577 8359
rect 48663 8336 48729 8359
rect 48343 8296 48352 8336
rect 48392 8296 48409 8336
rect 48495 8296 48516 8336
rect 48556 8296 48577 8336
rect 48663 8296 48680 8336
rect 48720 8296 48729 8336
rect 48343 8273 48409 8296
rect 48495 8273 48577 8296
rect 48663 8273 48729 8296
rect 48343 8254 48729 8273
rect 52343 8359 52729 8378
rect 52343 8336 52409 8359
rect 52495 8336 52577 8359
rect 52663 8336 52729 8359
rect 52343 8296 52352 8336
rect 52392 8296 52409 8336
rect 52495 8296 52516 8336
rect 52556 8296 52577 8336
rect 52663 8296 52680 8336
rect 52720 8296 52729 8336
rect 52343 8273 52409 8296
rect 52495 8273 52577 8296
rect 52663 8273 52729 8296
rect 52343 8254 52729 8273
rect 56343 8359 56729 8378
rect 56343 8336 56409 8359
rect 56495 8336 56577 8359
rect 56663 8336 56729 8359
rect 56343 8296 56352 8336
rect 56392 8296 56409 8336
rect 56495 8296 56516 8336
rect 56556 8296 56577 8336
rect 56663 8296 56680 8336
rect 56720 8296 56729 8336
rect 56343 8273 56409 8296
rect 56495 8273 56577 8296
rect 56663 8273 56729 8296
rect 56343 8254 56729 8273
rect 60343 8359 60729 8378
rect 60343 8336 60409 8359
rect 60495 8336 60577 8359
rect 60663 8336 60729 8359
rect 60343 8296 60352 8336
rect 60392 8296 60409 8336
rect 60495 8296 60516 8336
rect 60556 8296 60577 8336
rect 60663 8296 60680 8336
rect 60720 8296 60729 8336
rect 60343 8273 60409 8296
rect 60495 8273 60577 8296
rect 60663 8273 60729 8296
rect 60343 8254 60729 8273
rect 64343 8359 64729 8378
rect 64343 8336 64409 8359
rect 64495 8336 64577 8359
rect 64663 8336 64729 8359
rect 64343 8296 64352 8336
rect 64392 8296 64409 8336
rect 64495 8296 64516 8336
rect 64556 8296 64577 8336
rect 64663 8296 64680 8336
rect 64720 8296 64729 8336
rect 64343 8273 64409 8296
rect 64495 8273 64577 8296
rect 64663 8273 64729 8296
rect 64343 8254 64729 8273
rect 68343 8359 68729 8378
rect 68343 8336 68409 8359
rect 68495 8336 68577 8359
rect 68663 8336 68729 8359
rect 68343 8296 68352 8336
rect 68392 8296 68409 8336
rect 68495 8296 68516 8336
rect 68556 8296 68577 8336
rect 68663 8296 68680 8336
rect 68720 8296 68729 8336
rect 68343 8273 68409 8296
rect 68495 8273 68577 8296
rect 68663 8273 68729 8296
rect 68343 8254 68729 8273
rect 75076 8312 75169 8398
rect 75255 8312 75337 8398
rect 75423 8312 75516 8398
rect 75076 8230 75516 8312
rect 75076 8144 75169 8230
rect 75255 8144 75337 8230
rect 75423 8144 75516 8230
rect 75076 8014 75516 8144
rect 79076 10246 79516 10376
rect 79076 10160 79169 10246
rect 79255 10160 79337 10246
rect 79423 10160 79516 10246
rect 79076 10078 79516 10160
rect 79076 9992 79169 10078
rect 79255 9992 79337 10078
rect 79423 9992 79516 10078
rect 79076 9910 79516 9992
rect 79076 9824 79169 9910
rect 79255 9824 79337 9910
rect 79423 9824 79516 9910
rect 79076 9742 79516 9824
rect 79076 9656 79169 9742
rect 79255 9656 79337 9742
rect 79423 9656 79516 9742
rect 79076 9574 79516 9656
rect 79076 9488 79169 9574
rect 79255 9488 79337 9574
rect 79423 9488 79516 9574
rect 79076 9406 79516 9488
rect 79076 9320 79169 9406
rect 79255 9320 79337 9406
rect 79423 9320 79516 9406
rect 79076 9238 79516 9320
rect 79076 9152 79169 9238
rect 79255 9152 79337 9238
rect 79423 9152 79516 9238
rect 79076 9070 79516 9152
rect 79076 8984 79169 9070
rect 79255 8984 79337 9070
rect 79423 8984 79516 9070
rect 79076 8902 79516 8984
rect 79076 8816 79169 8902
rect 79255 8816 79337 8902
rect 79423 8816 79516 8902
rect 79076 8734 79516 8816
rect 79076 8648 79169 8734
rect 79255 8648 79337 8734
rect 79423 8648 79516 8734
rect 79076 8566 79516 8648
rect 79076 8480 79169 8566
rect 79255 8480 79337 8566
rect 79423 8480 79516 8566
rect 79076 8398 79516 8480
rect 79076 8312 79169 8398
rect 79255 8312 79337 8398
rect 79423 8312 79516 8398
rect 79076 8230 79516 8312
rect 79076 8144 79169 8230
rect 79255 8144 79337 8230
rect 79423 8144 79516 8230
rect 79076 8014 79516 8144
rect 83076 10246 83516 10376
rect 83076 10160 83169 10246
rect 83255 10160 83337 10246
rect 83423 10160 83516 10246
rect 83076 10078 83516 10160
rect 83076 9992 83169 10078
rect 83255 9992 83337 10078
rect 83423 9992 83516 10078
rect 83076 9910 83516 9992
rect 83076 9824 83169 9910
rect 83255 9824 83337 9910
rect 83423 9824 83516 9910
rect 83076 9742 83516 9824
rect 83076 9656 83169 9742
rect 83255 9656 83337 9742
rect 83423 9656 83516 9742
rect 83076 9574 83516 9656
rect 83076 9488 83169 9574
rect 83255 9488 83337 9574
rect 83423 9488 83516 9574
rect 83076 9406 83516 9488
rect 83076 9320 83169 9406
rect 83255 9320 83337 9406
rect 83423 9320 83516 9406
rect 83076 9238 83516 9320
rect 83076 9152 83169 9238
rect 83255 9152 83337 9238
rect 83423 9152 83516 9238
rect 83076 9070 83516 9152
rect 83076 8984 83169 9070
rect 83255 8984 83337 9070
rect 83423 8984 83516 9070
rect 83076 8902 83516 8984
rect 83076 8816 83169 8902
rect 83255 8816 83337 8902
rect 83423 8816 83516 8902
rect 83076 8734 83516 8816
rect 83076 8648 83169 8734
rect 83255 8648 83337 8734
rect 83423 8648 83516 8734
rect 83076 8566 83516 8648
rect 83076 8480 83169 8566
rect 83255 8480 83337 8566
rect 83423 8480 83516 8566
rect 83076 8398 83516 8480
rect 83076 8312 83169 8398
rect 83255 8312 83337 8398
rect 83423 8312 83516 8398
rect 83076 8230 83516 8312
rect 83076 8144 83169 8230
rect 83255 8144 83337 8230
rect 83423 8144 83516 8230
rect 83076 8014 83516 8144
rect 87076 10246 87516 10376
rect 87076 10160 87169 10246
rect 87255 10160 87337 10246
rect 87423 10160 87516 10246
rect 87076 10078 87516 10160
rect 87076 9992 87169 10078
rect 87255 9992 87337 10078
rect 87423 9992 87516 10078
rect 87076 9910 87516 9992
rect 87076 9824 87169 9910
rect 87255 9824 87337 9910
rect 87423 9824 87516 9910
rect 87076 9742 87516 9824
rect 87076 9656 87169 9742
rect 87255 9656 87337 9742
rect 87423 9656 87516 9742
rect 87076 9574 87516 9656
rect 87076 9488 87169 9574
rect 87255 9488 87337 9574
rect 87423 9488 87516 9574
rect 87076 9406 87516 9488
rect 87076 9320 87169 9406
rect 87255 9320 87337 9406
rect 87423 9320 87516 9406
rect 87076 9238 87516 9320
rect 87076 9152 87169 9238
rect 87255 9152 87337 9238
rect 87423 9152 87516 9238
rect 87076 9070 87516 9152
rect 87076 8984 87169 9070
rect 87255 8984 87337 9070
rect 87423 8984 87516 9070
rect 87076 8902 87516 8984
rect 87076 8816 87169 8902
rect 87255 8816 87337 8902
rect 87423 8816 87516 8902
rect 87076 8734 87516 8816
rect 87076 8648 87169 8734
rect 87255 8648 87337 8734
rect 87423 8648 87516 8734
rect 87076 8566 87516 8648
rect 87076 8480 87169 8566
rect 87255 8480 87337 8566
rect 87423 8480 87516 8566
rect 87076 8398 87516 8480
rect 87076 8312 87169 8398
rect 87255 8312 87337 8398
rect 87423 8312 87516 8398
rect 87076 8230 87516 8312
rect 87076 8144 87169 8230
rect 87255 8144 87337 8230
rect 87423 8144 87516 8230
rect 87076 8014 87516 8144
rect 91076 10246 91516 10376
rect 91076 10160 91169 10246
rect 91255 10160 91337 10246
rect 91423 10160 91516 10246
rect 91076 10078 91516 10160
rect 91076 9992 91169 10078
rect 91255 9992 91337 10078
rect 91423 9992 91516 10078
rect 91076 9910 91516 9992
rect 91076 9824 91169 9910
rect 91255 9824 91337 9910
rect 91423 9824 91516 9910
rect 91076 9742 91516 9824
rect 91076 9656 91169 9742
rect 91255 9656 91337 9742
rect 91423 9656 91516 9742
rect 91076 9574 91516 9656
rect 91076 9488 91169 9574
rect 91255 9488 91337 9574
rect 91423 9488 91516 9574
rect 91076 9406 91516 9488
rect 91076 9320 91169 9406
rect 91255 9320 91337 9406
rect 91423 9320 91516 9406
rect 91076 9238 91516 9320
rect 91076 9152 91169 9238
rect 91255 9152 91337 9238
rect 91423 9152 91516 9238
rect 91076 9070 91516 9152
rect 91076 8984 91169 9070
rect 91255 8984 91337 9070
rect 91423 8984 91516 9070
rect 91076 8902 91516 8984
rect 91076 8816 91169 8902
rect 91255 8816 91337 8902
rect 91423 8816 91516 8902
rect 91076 8734 91516 8816
rect 91076 8648 91169 8734
rect 91255 8648 91337 8734
rect 91423 8648 91516 8734
rect 91076 8566 91516 8648
rect 91076 8480 91169 8566
rect 91255 8480 91337 8566
rect 91423 8480 91516 8566
rect 91076 8398 91516 8480
rect 91076 8312 91169 8398
rect 91255 8312 91337 8398
rect 91423 8312 91516 8398
rect 91076 8230 91516 8312
rect 91076 8144 91169 8230
rect 91255 8144 91337 8230
rect 91423 8144 91516 8230
rect 91076 8014 91516 8144
rect 95076 10246 95516 10376
rect 95076 10160 95169 10246
rect 95255 10160 95337 10246
rect 95423 10160 95516 10246
rect 95076 10078 95516 10160
rect 95076 9992 95169 10078
rect 95255 9992 95337 10078
rect 95423 9992 95516 10078
rect 95076 9910 95516 9992
rect 95076 9824 95169 9910
rect 95255 9824 95337 9910
rect 95423 9824 95516 9910
rect 95076 9742 95516 9824
rect 95076 9656 95169 9742
rect 95255 9656 95337 9742
rect 95423 9656 95516 9742
rect 95076 9574 95516 9656
rect 95076 9488 95169 9574
rect 95255 9488 95337 9574
rect 95423 9488 95516 9574
rect 95076 9406 95516 9488
rect 95076 9320 95169 9406
rect 95255 9320 95337 9406
rect 95423 9320 95516 9406
rect 95076 9238 95516 9320
rect 95076 9152 95169 9238
rect 95255 9152 95337 9238
rect 95423 9152 95516 9238
rect 95076 9070 95516 9152
rect 95076 8984 95169 9070
rect 95255 8984 95337 9070
rect 95423 8984 95516 9070
rect 95076 8902 95516 8984
rect 95076 8816 95169 8902
rect 95255 8816 95337 8902
rect 95423 8816 95516 8902
rect 95076 8734 95516 8816
rect 95076 8648 95169 8734
rect 95255 8648 95337 8734
rect 95423 8648 95516 8734
rect 95076 8566 95516 8648
rect 95076 8480 95169 8566
rect 95255 8480 95337 8566
rect 95423 8480 95516 8566
rect 95076 8398 95516 8480
rect 95076 8312 95169 8398
rect 95255 8312 95337 8398
rect 95423 8312 95516 8398
rect 95076 8230 95516 8312
rect 95076 8144 95169 8230
rect 95255 8144 95337 8230
rect 95423 8144 95516 8230
rect 95076 8014 95516 8144
rect 3103 7603 3489 7622
rect 3103 7580 3169 7603
rect 3255 7580 3337 7603
rect 3423 7580 3489 7603
rect 3103 7540 3112 7580
rect 3152 7540 3169 7580
rect 3255 7540 3276 7580
rect 3316 7540 3337 7580
rect 3423 7540 3440 7580
rect 3480 7540 3489 7580
rect 3103 7517 3169 7540
rect 3255 7517 3337 7540
rect 3423 7517 3489 7540
rect 3103 7498 3489 7517
rect 7103 7603 7489 7622
rect 7103 7580 7169 7603
rect 7255 7580 7337 7603
rect 7423 7580 7489 7603
rect 7103 7540 7112 7580
rect 7152 7540 7169 7580
rect 7255 7540 7276 7580
rect 7316 7540 7337 7580
rect 7423 7540 7440 7580
rect 7480 7540 7489 7580
rect 7103 7517 7169 7540
rect 7255 7517 7337 7540
rect 7423 7517 7489 7540
rect 7103 7498 7489 7517
rect 11103 7603 11489 7622
rect 11103 7580 11169 7603
rect 11255 7580 11337 7603
rect 11423 7580 11489 7603
rect 11103 7540 11112 7580
rect 11152 7540 11169 7580
rect 11255 7540 11276 7580
rect 11316 7540 11337 7580
rect 11423 7540 11440 7580
rect 11480 7540 11489 7580
rect 11103 7517 11169 7540
rect 11255 7517 11337 7540
rect 11423 7517 11489 7540
rect 11103 7498 11489 7517
rect 15103 7603 15489 7622
rect 15103 7580 15169 7603
rect 15255 7580 15337 7603
rect 15423 7580 15489 7603
rect 15103 7540 15112 7580
rect 15152 7540 15169 7580
rect 15255 7540 15276 7580
rect 15316 7540 15337 7580
rect 15423 7540 15440 7580
rect 15480 7540 15489 7580
rect 15103 7517 15169 7540
rect 15255 7517 15337 7540
rect 15423 7517 15489 7540
rect 15103 7498 15489 7517
rect 19103 7603 19489 7622
rect 19103 7580 19169 7603
rect 19255 7580 19337 7603
rect 19423 7580 19489 7603
rect 19103 7540 19112 7580
rect 19152 7540 19169 7580
rect 19255 7540 19276 7580
rect 19316 7540 19337 7580
rect 19423 7540 19440 7580
rect 19480 7540 19489 7580
rect 19103 7517 19169 7540
rect 19255 7517 19337 7540
rect 19423 7517 19489 7540
rect 19103 7498 19489 7517
rect 23103 7603 23489 7622
rect 23103 7580 23169 7603
rect 23255 7580 23337 7603
rect 23423 7580 23489 7603
rect 23103 7540 23112 7580
rect 23152 7540 23169 7580
rect 23255 7540 23276 7580
rect 23316 7540 23337 7580
rect 23423 7540 23440 7580
rect 23480 7540 23489 7580
rect 23103 7517 23169 7540
rect 23255 7517 23337 7540
rect 23423 7517 23489 7540
rect 23103 7498 23489 7517
rect 27103 7603 27489 7622
rect 27103 7580 27169 7603
rect 27255 7580 27337 7603
rect 27423 7580 27489 7603
rect 27103 7540 27112 7580
rect 27152 7540 27169 7580
rect 27255 7540 27276 7580
rect 27316 7540 27337 7580
rect 27423 7540 27440 7580
rect 27480 7540 27489 7580
rect 27103 7517 27169 7540
rect 27255 7517 27337 7540
rect 27423 7517 27489 7540
rect 27103 7498 27489 7517
rect 31103 7603 31489 7622
rect 31103 7580 31169 7603
rect 31255 7580 31337 7603
rect 31423 7580 31489 7603
rect 31103 7540 31112 7580
rect 31152 7540 31169 7580
rect 31255 7540 31276 7580
rect 31316 7540 31337 7580
rect 31423 7540 31440 7580
rect 31480 7540 31489 7580
rect 31103 7517 31169 7540
rect 31255 7517 31337 7540
rect 31423 7517 31489 7540
rect 31103 7498 31489 7517
rect 35103 7603 35489 7622
rect 35103 7580 35169 7603
rect 35255 7580 35337 7603
rect 35423 7580 35489 7603
rect 35103 7540 35112 7580
rect 35152 7540 35169 7580
rect 35255 7540 35276 7580
rect 35316 7540 35337 7580
rect 35423 7540 35440 7580
rect 35480 7540 35489 7580
rect 35103 7517 35169 7540
rect 35255 7517 35337 7540
rect 35423 7517 35489 7540
rect 35103 7498 35489 7517
rect 39103 7603 39489 7622
rect 39103 7580 39169 7603
rect 39255 7580 39337 7603
rect 39423 7580 39489 7603
rect 39103 7540 39112 7580
rect 39152 7540 39169 7580
rect 39255 7540 39276 7580
rect 39316 7540 39337 7580
rect 39423 7540 39440 7580
rect 39480 7540 39489 7580
rect 39103 7517 39169 7540
rect 39255 7517 39337 7540
rect 39423 7517 39489 7540
rect 39103 7498 39489 7517
rect 43103 7603 43489 7622
rect 43103 7580 43169 7603
rect 43255 7580 43337 7603
rect 43423 7580 43489 7603
rect 43103 7540 43112 7580
rect 43152 7540 43169 7580
rect 43255 7540 43276 7580
rect 43316 7540 43337 7580
rect 43423 7540 43440 7580
rect 43480 7540 43489 7580
rect 43103 7517 43169 7540
rect 43255 7517 43337 7540
rect 43423 7517 43489 7540
rect 43103 7498 43489 7517
rect 47103 7603 47489 7622
rect 47103 7580 47169 7603
rect 47255 7580 47337 7603
rect 47423 7580 47489 7603
rect 47103 7540 47112 7580
rect 47152 7540 47169 7580
rect 47255 7540 47276 7580
rect 47316 7540 47337 7580
rect 47423 7540 47440 7580
rect 47480 7540 47489 7580
rect 47103 7517 47169 7540
rect 47255 7517 47337 7540
rect 47423 7517 47489 7540
rect 47103 7498 47489 7517
rect 51103 7603 51489 7622
rect 51103 7580 51169 7603
rect 51255 7580 51337 7603
rect 51423 7580 51489 7603
rect 51103 7540 51112 7580
rect 51152 7540 51169 7580
rect 51255 7540 51276 7580
rect 51316 7540 51337 7580
rect 51423 7540 51440 7580
rect 51480 7540 51489 7580
rect 51103 7517 51169 7540
rect 51255 7517 51337 7540
rect 51423 7517 51489 7540
rect 51103 7498 51489 7517
rect 55103 7603 55489 7622
rect 55103 7580 55169 7603
rect 55255 7580 55337 7603
rect 55423 7580 55489 7603
rect 55103 7540 55112 7580
rect 55152 7540 55169 7580
rect 55255 7540 55276 7580
rect 55316 7540 55337 7580
rect 55423 7540 55440 7580
rect 55480 7540 55489 7580
rect 55103 7517 55169 7540
rect 55255 7517 55337 7540
rect 55423 7517 55489 7540
rect 55103 7498 55489 7517
rect 59103 7603 59489 7622
rect 59103 7580 59169 7603
rect 59255 7580 59337 7603
rect 59423 7580 59489 7603
rect 59103 7540 59112 7580
rect 59152 7540 59169 7580
rect 59255 7540 59276 7580
rect 59316 7540 59337 7580
rect 59423 7540 59440 7580
rect 59480 7540 59489 7580
rect 59103 7517 59169 7540
rect 59255 7517 59337 7540
rect 59423 7517 59489 7540
rect 59103 7498 59489 7517
rect 63103 7603 63489 7622
rect 63103 7580 63169 7603
rect 63255 7580 63337 7603
rect 63423 7580 63489 7603
rect 63103 7540 63112 7580
rect 63152 7540 63169 7580
rect 63255 7540 63276 7580
rect 63316 7540 63337 7580
rect 63423 7540 63440 7580
rect 63480 7540 63489 7580
rect 63103 7517 63169 7540
rect 63255 7517 63337 7540
rect 63423 7517 63489 7540
rect 63103 7498 63489 7517
rect 67103 7603 67489 7622
rect 67103 7580 67169 7603
rect 67255 7580 67337 7603
rect 67423 7580 67489 7603
rect 67103 7540 67112 7580
rect 67152 7540 67169 7580
rect 67255 7540 67276 7580
rect 67316 7540 67337 7580
rect 67423 7540 67440 7580
rect 67480 7540 67489 7580
rect 67103 7517 67169 7540
rect 67255 7517 67337 7540
rect 67423 7517 67489 7540
rect 67103 7498 67489 7517
rect 86450 7519 86574 7538
rect 86450 7433 86469 7519
rect 86555 7496 86574 7519
rect 86555 7456 86668 7496
rect 86708 7456 86717 7496
rect 86555 7433 86574 7456
rect 86450 7414 86574 7433
rect 4343 6847 4729 6866
rect 4343 6824 4409 6847
rect 4495 6824 4577 6847
rect 4663 6824 4729 6847
rect 4343 6784 4352 6824
rect 4392 6784 4409 6824
rect 4495 6784 4516 6824
rect 4556 6784 4577 6824
rect 4663 6784 4680 6824
rect 4720 6784 4729 6824
rect 4343 6761 4409 6784
rect 4495 6761 4577 6784
rect 4663 6761 4729 6784
rect 4343 6742 4729 6761
rect 8343 6847 8729 6866
rect 8343 6824 8409 6847
rect 8495 6824 8577 6847
rect 8663 6824 8729 6847
rect 8343 6784 8352 6824
rect 8392 6784 8409 6824
rect 8495 6784 8516 6824
rect 8556 6784 8577 6824
rect 8663 6784 8680 6824
rect 8720 6784 8729 6824
rect 8343 6761 8409 6784
rect 8495 6761 8577 6784
rect 8663 6761 8729 6784
rect 8343 6742 8729 6761
rect 12343 6847 12729 6866
rect 12343 6824 12409 6847
rect 12495 6824 12577 6847
rect 12663 6824 12729 6847
rect 12343 6784 12352 6824
rect 12392 6784 12409 6824
rect 12495 6784 12516 6824
rect 12556 6784 12577 6824
rect 12663 6784 12680 6824
rect 12720 6784 12729 6824
rect 12343 6761 12409 6784
rect 12495 6761 12577 6784
rect 12663 6761 12729 6784
rect 12343 6742 12729 6761
rect 16343 6847 16729 6866
rect 16343 6824 16409 6847
rect 16495 6824 16577 6847
rect 16663 6824 16729 6847
rect 16343 6784 16352 6824
rect 16392 6784 16409 6824
rect 16495 6784 16516 6824
rect 16556 6784 16577 6824
rect 16663 6784 16680 6824
rect 16720 6784 16729 6824
rect 16343 6761 16409 6784
rect 16495 6761 16577 6784
rect 16663 6761 16729 6784
rect 16343 6742 16729 6761
rect 20343 6847 20729 6866
rect 20343 6824 20409 6847
rect 20495 6824 20577 6847
rect 20663 6824 20729 6847
rect 20343 6784 20352 6824
rect 20392 6784 20409 6824
rect 20495 6784 20516 6824
rect 20556 6784 20577 6824
rect 20663 6784 20680 6824
rect 20720 6784 20729 6824
rect 20343 6761 20409 6784
rect 20495 6761 20577 6784
rect 20663 6761 20729 6784
rect 20343 6742 20729 6761
rect 24343 6847 24729 6866
rect 24343 6824 24409 6847
rect 24495 6824 24577 6847
rect 24663 6824 24729 6847
rect 24343 6784 24352 6824
rect 24392 6784 24409 6824
rect 24495 6784 24516 6824
rect 24556 6784 24577 6824
rect 24663 6784 24680 6824
rect 24720 6784 24729 6824
rect 24343 6761 24409 6784
rect 24495 6761 24577 6784
rect 24663 6761 24729 6784
rect 24343 6742 24729 6761
rect 28343 6847 28729 6866
rect 28343 6824 28409 6847
rect 28495 6824 28577 6847
rect 28663 6824 28729 6847
rect 28343 6784 28352 6824
rect 28392 6784 28409 6824
rect 28495 6784 28516 6824
rect 28556 6784 28577 6824
rect 28663 6784 28680 6824
rect 28720 6784 28729 6824
rect 28343 6761 28409 6784
rect 28495 6761 28577 6784
rect 28663 6761 28729 6784
rect 28343 6742 28729 6761
rect 32343 6847 32729 6866
rect 32343 6824 32409 6847
rect 32495 6824 32577 6847
rect 32663 6824 32729 6847
rect 32343 6784 32352 6824
rect 32392 6784 32409 6824
rect 32495 6784 32516 6824
rect 32556 6784 32577 6824
rect 32663 6784 32680 6824
rect 32720 6784 32729 6824
rect 32343 6761 32409 6784
rect 32495 6761 32577 6784
rect 32663 6761 32729 6784
rect 32343 6742 32729 6761
rect 36343 6847 36729 6866
rect 36343 6824 36409 6847
rect 36495 6824 36577 6847
rect 36663 6824 36729 6847
rect 36343 6784 36352 6824
rect 36392 6784 36409 6824
rect 36495 6784 36516 6824
rect 36556 6784 36577 6824
rect 36663 6784 36680 6824
rect 36720 6784 36729 6824
rect 36343 6761 36409 6784
rect 36495 6761 36577 6784
rect 36663 6761 36729 6784
rect 36343 6742 36729 6761
rect 40343 6847 40729 6866
rect 40343 6824 40409 6847
rect 40495 6824 40577 6847
rect 40663 6824 40729 6847
rect 40343 6784 40352 6824
rect 40392 6784 40409 6824
rect 40495 6784 40516 6824
rect 40556 6784 40577 6824
rect 40663 6784 40680 6824
rect 40720 6784 40729 6824
rect 40343 6761 40409 6784
rect 40495 6761 40577 6784
rect 40663 6761 40729 6784
rect 40343 6742 40729 6761
rect 44343 6847 44729 6866
rect 44343 6824 44409 6847
rect 44495 6824 44577 6847
rect 44663 6824 44729 6847
rect 44343 6784 44352 6824
rect 44392 6784 44409 6824
rect 44495 6784 44516 6824
rect 44556 6784 44577 6824
rect 44663 6784 44680 6824
rect 44720 6784 44729 6824
rect 44343 6761 44409 6784
rect 44495 6761 44577 6784
rect 44663 6761 44729 6784
rect 44343 6742 44729 6761
rect 48343 6847 48729 6866
rect 48343 6824 48409 6847
rect 48495 6824 48577 6847
rect 48663 6824 48729 6847
rect 48343 6784 48352 6824
rect 48392 6784 48409 6824
rect 48495 6784 48516 6824
rect 48556 6784 48577 6824
rect 48663 6784 48680 6824
rect 48720 6784 48729 6824
rect 48343 6761 48409 6784
rect 48495 6761 48577 6784
rect 48663 6761 48729 6784
rect 48343 6742 48729 6761
rect 52343 6847 52729 6866
rect 52343 6824 52409 6847
rect 52495 6824 52577 6847
rect 52663 6824 52729 6847
rect 52343 6784 52352 6824
rect 52392 6784 52409 6824
rect 52495 6784 52516 6824
rect 52556 6784 52577 6824
rect 52663 6784 52680 6824
rect 52720 6784 52729 6824
rect 52343 6761 52409 6784
rect 52495 6761 52577 6784
rect 52663 6761 52729 6784
rect 52343 6742 52729 6761
rect 56343 6847 56729 6866
rect 56343 6824 56409 6847
rect 56495 6824 56577 6847
rect 56663 6824 56729 6847
rect 56343 6784 56352 6824
rect 56392 6784 56409 6824
rect 56495 6784 56516 6824
rect 56556 6784 56577 6824
rect 56663 6784 56680 6824
rect 56720 6784 56729 6824
rect 56343 6761 56409 6784
rect 56495 6761 56577 6784
rect 56663 6761 56729 6784
rect 56343 6742 56729 6761
rect 60343 6847 60729 6866
rect 60343 6824 60409 6847
rect 60495 6824 60577 6847
rect 60663 6824 60729 6847
rect 60343 6784 60352 6824
rect 60392 6784 60409 6824
rect 60495 6784 60516 6824
rect 60556 6784 60577 6824
rect 60663 6784 60680 6824
rect 60720 6784 60729 6824
rect 60343 6761 60409 6784
rect 60495 6761 60577 6784
rect 60663 6761 60729 6784
rect 60343 6742 60729 6761
rect 64343 6847 64729 6866
rect 64343 6824 64409 6847
rect 64495 6824 64577 6847
rect 64663 6824 64729 6847
rect 64343 6784 64352 6824
rect 64392 6784 64409 6824
rect 64495 6784 64516 6824
rect 64556 6784 64577 6824
rect 64663 6784 64680 6824
rect 64720 6784 64729 6824
rect 64343 6761 64409 6784
rect 64495 6761 64577 6784
rect 64663 6761 64729 6784
rect 64343 6742 64729 6761
rect 68343 6847 68729 6866
rect 68343 6824 68409 6847
rect 68495 6824 68577 6847
rect 68663 6824 68729 6847
rect 68343 6784 68352 6824
rect 68392 6784 68409 6824
rect 68495 6784 68516 6824
rect 68556 6784 68577 6824
rect 68663 6784 68680 6824
rect 68720 6784 68729 6824
rect 68343 6761 68409 6784
rect 68495 6761 68577 6784
rect 68663 6761 68729 6784
rect 68343 6742 68729 6761
rect 3103 6091 3489 6110
rect 3103 6068 3169 6091
rect 3255 6068 3337 6091
rect 3423 6068 3489 6091
rect 3103 6028 3112 6068
rect 3152 6028 3169 6068
rect 3255 6028 3276 6068
rect 3316 6028 3337 6068
rect 3423 6028 3440 6068
rect 3480 6028 3489 6068
rect 3103 6005 3169 6028
rect 3255 6005 3337 6028
rect 3423 6005 3489 6028
rect 3103 5986 3489 6005
rect 7103 6091 7489 6110
rect 7103 6068 7169 6091
rect 7255 6068 7337 6091
rect 7423 6068 7489 6091
rect 7103 6028 7112 6068
rect 7152 6028 7169 6068
rect 7255 6028 7276 6068
rect 7316 6028 7337 6068
rect 7423 6028 7440 6068
rect 7480 6028 7489 6068
rect 7103 6005 7169 6028
rect 7255 6005 7337 6028
rect 7423 6005 7489 6028
rect 7103 5986 7489 6005
rect 11103 6091 11489 6110
rect 11103 6068 11169 6091
rect 11255 6068 11337 6091
rect 11423 6068 11489 6091
rect 11103 6028 11112 6068
rect 11152 6028 11169 6068
rect 11255 6028 11276 6068
rect 11316 6028 11337 6068
rect 11423 6028 11440 6068
rect 11480 6028 11489 6068
rect 11103 6005 11169 6028
rect 11255 6005 11337 6028
rect 11423 6005 11489 6028
rect 11103 5986 11489 6005
rect 15103 6091 15489 6110
rect 15103 6068 15169 6091
rect 15255 6068 15337 6091
rect 15423 6068 15489 6091
rect 15103 6028 15112 6068
rect 15152 6028 15169 6068
rect 15255 6028 15276 6068
rect 15316 6028 15337 6068
rect 15423 6028 15440 6068
rect 15480 6028 15489 6068
rect 15103 6005 15169 6028
rect 15255 6005 15337 6028
rect 15423 6005 15489 6028
rect 15103 5986 15489 6005
rect 19103 6091 19489 6110
rect 19103 6068 19169 6091
rect 19255 6068 19337 6091
rect 19423 6068 19489 6091
rect 19103 6028 19112 6068
rect 19152 6028 19169 6068
rect 19255 6028 19276 6068
rect 19316 6028 19337 6068
rect 19423 6028 19440 6068
rect 19480 6028 19489 6068
rect 19103 6005 19169 6028
rect 19255 6005 19337 6028
rect 19423 6005 19489 6028
rect 19103 5986 19489 6005
rect 23103 6091 23489 6110
rect 23103 6068 23169 6091
rect 23255 6068 23337 6091
rect 23423 6068 23489 6091
rect 23103 6028 23112 6068
rect 23152 6028 23169 6068
rect 23255 6028 23276 6068
rect 23316 6028 23337 6068
rect 23423 6028 23440 6068
rect 23480 6028 23489 6068
rect 23103 6005 23169 6028
rect 23255 6005 23337 6028
rect 23423 6005 23489 6028
rect 23103 5986 23489 6005
rect 27103 6091 27489 6110
rect 27103 6068 27169 6091
rect 27255 6068 27337 6091
rect 27423 6068 27489 6091
rect 27103 6028 27112 6068
rect 27152 6028 27169 6068
rect 27255 6028 27276 6068
rect 27316 6028 27337 6068
rect 27423 6028 27440 6068
rect 27480 6028 27489 6068
rect 27103 6005 27169 6028
rect 27255 6005 27337 6028
rect 27423 6005 27489 6028
rect 27103 5986 27489 6005
rect 31103 6091 31489 6110
rect 31103 6068 31169 6091
rect 31255 6068 31337 6091
rect 31423 6068 31489 6091
rect 31103 6028 31112 6068
rect 31152 6028 31169 6068
rect 31255 6028 31276 6068
rect 31316 6028 31337 6068
rect 31423 6028 31440 6068
rect 31480 6028 31489 6068
rect 31103 6005 31169 6028
rect 31255 6005 31337 6028
rect 31423 6005 31489 6028
rect 31103 5986 31489 6005
rect 35103 6091 35489 6110
rect 35103 6068 35169 6091
rect 35255 6068 35337 6091
rect 35423 6068 35489 6091
rect 35103 6028 35112 6068
rect 35152 6028 35169 6068
rect 35255 6028 35276 6068
rect 35316 6028 35337 6068
rect 35423 6028 35440 6068
rect 35480 6028 35489 6068
rect 35103 6005 35169 6028
rect 35255 6005 35337 6028
rect 35423 6005 35489 6028
rect 35103 5986 35489 6005
rect 39103 6091 39489 6110
rect 39103 6068 39169 6091
rect 39255 6068 39337 6091
rect 39423 6068 39489 6091
rect 39103 6028 39112 6068
rect 39152 6028 39169 6068
rect 39255 6028 39276 6068
rect 39316 6028 39337 6068
rect 39423 6028 39440 6068
rect 39480 6028 39489 6068
rect 39103 6005 39169 6028
rect 39255 6005 39337 6028
rect 39423 6005 39489 6028
rect 39103 5986 39489 6005
rect 43103 6091 43489 6110
rect 43103 6068 43169 6091
rect 43255 6068 43337 6091
rect 43423 6068 43489 6091
rect 43103 6028 43112 6068
rect 43152 6028 43169 6068
rect 43255 6028 43276 6068
rect 43316 6028 43337 6068
rect 43423 6028 43440 6068
rect 43480 6028 43489 6068
rect 43103 6005 43169 6028
rect 43255 6005 43337 6028
rect 43423 6005 43489 6028
rect 43103 5986 43489 6005
rect 47103 6091 47489 6110
rect 47103 6068 47169 6091
rect 47255 6068 47337 6091
rect 47423 6068 47489 6091
rect 47103 6028 47112 6068
rect 47152 6028 47169 6068
rect 47255 6028 47276 6068
rect 47316 6028 47337 6068
rect 47423 6028 47440 6068
rect 47480 6028 47489 6068
rect 47103 6005 47169 6028
rect 47255 6005 47337 6028
rect 47423 6005 47489 6028
rect 47103 5986 47489 6005
rect 51103 6091 51489 6110
rect 51103 6068 51169 6091
rect 51255 6068 51337 6091
rect 51423 6068 51489 6091
rect 51103 6028 51112 6068
rect 51152 6028 51169 6068
rect 51255 6028 51276 6068
rect 51316 6028 51337 6068
rect 51423 6028 51440 6068
rect 51480 6028 51489 6068
rect 51103 6005 51169 6028
rect 51255 6005 51337 6028
rect 51423 6005 51489 6028
rect 51103 5986 51489 6005
rect 55103 6091 55489 6110
rect 55103 6068 55169 6091
rect 55255 6068 55337 6091
rect 55423 6068 55489 6091
rect 55103 6028 55112 6068
rect 55152 6028 55169 6068
rect 55255 6028 55276 6068
rect 55316 6028 55337 6068
rect 55423 6028 55440 6068
rect 55480 6028 55489 6068
rect 55103 6005 55169 6028
rect 55255 6005 55337 6028
rect 55423 6005 55489 6028
rect 55103 5986 55489 6005
rect 59103 6091 59489 6110
rect 59103 6068 59169 6091
rect 59255 6068 59337 6091
rect 59423 6068 59489 6091
rect 59103 6028 59112 6068
rect 59152 6028 59169 6068
rect 59255 6028 59276 6068
rect 59316 6028 59337 6068
rect 59423 6028 59440 6068
rect 59480 6028 59489 6068
rect 59103 6005 59169 6028
rect 59255 6005 59337 6028
rect 59423 6005 59489 6028
rect 59103 5986 59489 6005
rect 63103 6091 63489 6110
rect 63103 6068 63169 6091
rect 63255 6068 63337 6091
rect 63423 6068 63489 6091
rect 63103 6028 63112 6068
rect 63152 6028 63169 6068
rect 63255 6028 63276 6068
rect 63316 6028 63337 6068
rect 63423 6028 63440 6068
rect 63480 6028 63489 6068
rect 63103 6005 63169 6028
rect 63255 6005 63337 6028
rect 63423 6005 63489 6028
rect 63103 5986 63489 6005
rect 67103 6091 67489 6110
rect 67103 6068 67169 6091
rect 67255 6068 67337 6091
rect 67423 6068 67489 6091
rect 67103 6028 67112 6068
rect 67152 6028 67169 6068
rect 67255 6028 67276 6068
rect 67316 6028 67337 6068
rect 67423 6028 67440 6068
rect 67480 6028 67489 6068
rect 67103 6005 67169 6028
rect 67255 6005 67337 6028
rect 67423 6005 67489 6028
rect 67103 5986 67489 6005
rect 4343 5335 4729 5354
rect 4343 5312 4409 5335
rect 4495 5312 4577 5335
rect 4663 5312 4729 5335
rect 4343 5272 4352 5312
rect 4392 5272 4409 5312
rect 4495 5272 4516 5312
rect 4556 5272 4577 5312
rect 4663 5272 4680 5312
rect 4720 5272 4729 5312
rect 4343 5249 4409 5272
rect 4495 5249 4577 5272
rect 4663 5249 4729 5272
rect 4343 5230 4729 5249
rect 8343 5335 8729 5354
rect 8343 5312 8409 5335
rect 8495 5312 8577 5335
rect 8663 5312 8729 5335
rect 8343 5272 8352 5312
rect 8392 5272 8409 5312
rect 8495 5272 8516 5312
rect 8556 5272 8577 5312
rect 8663 5272 8680 5312
rect 8720 5272 8729 5312
rect 8343 5249 8409 5272
rect 8495 5249 8577 5272
rect 8663 5249 8729 5272
rect 8343 5230 8729 5249
rect 12343 5335 12729 5354
rect 12343 5312 12409 5335
rect 12495 5312 12577 5335
rect 12663 5312 12729 5335
rect 12343 5272 12352 5312
rect 12392 5272 12409 5312
rect 12495 5272 12516 5312
rect 12556 5272 12577 5312
rect 12663 5272 12680 5312
rect 12720 5272 12729 5312
rect 12343 5249 12409 5272
rect 12495 5249 12577 5272
rect 12663 5249 12729 5272
rect 12343 5230 12729 5249
rect 16343 5335 16729 5354
rect 16343 5312 16409 5335
rect 16495 5312 16577 5335
rect 16663 5312 16729 5335
rect 16343 5272 16352 5312
rect 16392 5272 16409 5312
rect 16495 5272 16516 5312
rect 16556 5272 16577 5312
rect 16663 5272 16680 5312
rect 16720 5272 16729 5312
rect 16343 5249 16409 5272
rect 16495 5249 16577 5272
rect 16663 5249 16729 5272
rect 16343 5230 16729 5249
rect 20343 5335 20729 5354
rect 20343 5312 20409 5335
rect 20495 5312 20577 5335
rect 20663 5312 20729 5335
rect 20343 5272 20352 5312
rect 20392 5272 20409 5312
rect 20495 5272 20516 5312
rect 20556 5272 20577 5312
rect 20663 5272 20680 5312
rect 20720 5272 20729 5312
rect 20343 5249 20409 5272
rect 20495 5249 20577 5272
rect 20663 5249 20729 5272
rect 20343 5230 20729 5249
rect 24343 5335 24729 5354
rect 24343 5312 24409 5335
rect 24495 5312 24577 5335
rect 24663 5312 24729 5335
rect 24343 5272 24352 5312
rect 24392 5272 24409 5312
rect 24495 5272 24516 5312
rect 24556 5272 24577 5312
rect 24663 5272 24680 5312
rect 24720 5272 24729 5312
rect 24343 5249 24409 5272
rect 24495 5249 24577 5272
rect 24663 5249 24729 5272
rect 24343 5230 24729 5249
rect 28343 5335 28729 5354
rect 28343 5312 28409 5335
rect 28495 5312 28577 5335
rect 28663 5312 28729 5335
rect 28343 5272 28352 5312
rect 28392 5272 28409 5312
rect 28495 5272 28516 5312
rect 28556 5272 28577 5312
rect 28663 5272 28680 5312
rect 28720 5272 28729 5312
rect 28343 5249 28409 5272
rect 28495 5249 28577 5272
rect 28663 5249 28729 5272
rect 28343 5230 28729 5249
rect 32343 5335 32729 5354
rect 32343 5312 32409 5335
rect 32495 5312 32577 5335
rect 32663 5312 32729 5335
rect 32343 5272 32352 5312
rect 32392 5272 32409 5312
rect 32495 5272 32516 5312
rect 32556 5272 32577 5312
rect 32663 5272 32680 5312
rect 32720 5272 32729 5312
rect 32343 5249 32409 5272
rect 32495 5249 32577 5272
rect 32663 5249 32729 5272
rect 32343 5230 32729 5249
rect 36343 5335 36729 5354
rect 36343 5312 36409 5335
rect 36495 5312 36577 5335
rect 36663 5312 36729 5335
rect 36343 5272 36352 5312
rect 36392 5272 36409 5312
rect 36495 5272 36516 5312
rect 36556 5272 36577 5312
rect 36663 5272 36680 5312
rect 36720 5272 36729 5312
rect 36343 5249 36409 5272
rect 36495 5249 36577 5272
rect 36663 5249 36729 5272
rect 36343 5230 36729 5249
rect 40343 5335 40729 5354
rect 40343 5312 40409 5335
rect 40495 5312 40577 5335
rect 40663 5312 40729 5335
rect 40343 5272 40352 5312
rect 40392 5272 40409 5312
rect 40495 5272 40516 5312
rect 40556 5272 40577 5312
rect 40663 5272 40680 5312
rect 40720 5272 40729 5312
rect 40343 5249 40409 5272
rect 40495 5249 40577 5272
rect 40663 5249 40729 5272
rect 40343 5230 40729 5249
rect 44343 5335 44729 5354
rect 44343 5312 44409 5335
rect 44495 5312 44577 5335
rect 44663 5312 44729 5335
rect 44343 5272 44352 5312
rect 44392 5272 44409 5312
rect 44495 5272 44516 5312
rect 44556 5272 44577 5312
rect 44663 5272 44680 5312
rect 44720 5272 44729 5312
rect 44343 5249 44409 5272
rect 44495 5249 44577 5272
rect 44663 5249 44729 5272
rect 44343 5230 44729 5249
rect 48343 5335 48729 5354
rect 48343 5312 48409 5335
rect 48495 5312 48577 5335
rect 48663 5312 48729 5335
rect 48343 5272 48352 5312
rect 48392 5272 48409 5312
rect 48495 5272 48516 5312
rect 48556 5272 48577 5312
rect 48663 5272 48680 5312
rect 48720 5272 48729 5312
rect 48343 5249 48409 5272
rect 48495 5249 48577 5272
rect 48663 5249 48729 5272
rect 48343 5230 48729 5249
rect 52343 5335 52729 5354
rect 52343 5312 52409 5335
rect 52495 5312 52577 5335
rect 52663 5312 52729 5335
rect 52343 5272 52352 5312
rect 52392 5272 52409 5312
rect 52495 5272 52516 5312
rect 52556 5272 52577 5312
rect 52663 5272 52680 5312
rect 52720 5272 52729 5312
rect 52343 5249 52409 5272
rect 52495 5249 52577 5272
rect 52663 5249 52729 5272
rect 52343 5230 52729 5249
rect 56343 5335 56729 5354
rect 56343 5312 56409 5335
rect 56495 5312 56577 5335
rect 56663 5312 56729 5335
rect 56343 5272 56352 5312
rect 56392 5272 56409 5312
rect 56495 5272 56516 5312
rect 56556 5272 56577 5312
rect 56663 5272 56680 5312
rect 56720 5272 56729 5312
rect 56343 5249 56409 5272
rect 56495 5249 56577 5272
rect 56663 5249 56729 5272
rect 56343 5230 56729 5249
rect 60343 5335 60729 5354
rect 60343 5312 60409 5335
rect 60495 5312 60577 5335
rect 60663 5312 60729 5335
rect 60343 5272 60352 5312
rect 60392 5272 60409 5312
rect 60495 5272 60516 5312
rect 60556 5272 60577 5312
rect 60663 5272 60680 5312
rect 60720 5272 60729 5312
rect 60343 5249 60409 5272
rect 60495 5249 60577 5272
rect 60663 5249 60729 5272
rect 60343 5230 60729 5249
rect 64343 5335 64729 5354
rect 64343 5312 64409 5335
rect 64495 5312 64577 5335
rect 64663 5312 64729 5335
rect 64343 5272 64352 5312
rect 64392 5272 64409 5312
rect 64495 5272 64516 5312
rect 64556 5272 64577 5312
rect 64663 5272 64680 5312
rect 64720 5272 64729 5312
rect 64343 5249 64409 5272
rect 64495 5249 64577 5272
rect 64663 5249 64729 5272
rect 64343 5230 64729 5249
rect 68343 5335 68729 5354
rect 68343 5312 68409 5335
rect 68495 5312 68577 5335
rect 68663 5312 68729 5335
rect 68343 5272 68352 5312
rect 68392 5272 68409 5312
rect 68495 5272 68516 5312
rect 68556 5272 68577 5312
rect 68663 5272 68680 5312
rect 68720 5272 68729 5312
rect 68343 5249 68409 5272
rect 68495 5249 68577 5272
rect 68663 5249 68729 5272
rect 68343 5230 68729 5249
rect 72343 5335 72729 5354
rect 72343 5312 72409 5335
rect 72495 5312 72577 5335
rect 72663 5312 72729 5335
rect 72343 5272 72352 5312
rect 72392 5272 72409 5312
rect 72495 5272 72516 5312
rect 72556 5272 72577 5312
rect 72663 5272 72680 5312
rect 72720 5272 72729 5312
rect 72343 5249 72409 5272
rect 72495 5249 72577 5272
rect 72663 5249 72729 5272
rect 72343 5230 72729 5249
rect 76343 5335 76729 5354
rect 76343 5312 76409 5335
rect 76495 5312 76577 5335
rect 76663 5312 76729 5335
rect 76343 5272 76352 5312
rect 76392 5272 76409 5312
rect 76495 5272 76516 5312
rect 76556 5272 76577 5312
rect 76663 5272 76680 5312
rect 76720 5272 76729 5312
rect 76343 5249 76409 5272
rect 76495 5249 76577 5272
rect 76663 5249 76729 5272
rect 76343 5230 76729 5249
rect 80343 5335 80729 5354
rect 80343 5312 80409 5335
rect 80495 5312 80577 5335
rect 80663 5312 80729 5335
rect 80343 5272 80352 5312
rect 80392 5272 80409 5312
rect 80495 5272 80516 5312
rect 80556 5272 80577 5312
rect 80663 5272 80680 5312
rect 80720 5272 80729 5312
rect 80343 5249 80409 5272
rect 80495 5249 80577 5272
rect 80663 5249 80729 5272
rect 80343 5230 80729 5249
rect 84343 5335 84729 5354
rect 84343 5312 84409 5335
rect 84495 5312 84577 5335
rect 84663 5312 84729 5335
rect 84343 5272 84352 5312
rect 84392 5272 84409 5312
rect 84495 5272 84516 5312
rect 84556 5272 84577 5312
rect 84663 5272 84680 5312
rect 84720 5272 84729 5312
rect 84343 5249 84409 5272
rect 84495 5249 84577 5272
rect 84663 5249 84729 5272
rect 84343 5230 84729 5249
rect 88343 5335 88729 5354
rect 88343 5312 88409 5335
rect 88495 5312 88577 5335
rect 88663 5312 88729 5335
rect 88343 5272 88352 5312
rect 88392 5272 88409 5312
rect 88495 5272 88516 5312
rect 88556 5272 88577 5312
rect 88663 5272 88680 5312
rect 88720 5272 88729 5312
rect 88343 5249 88409 5272
rect 88495 5249 88577 5272
rect 88663 5249 88729 5272
rect 88343 5230 88729 5249
rect 92343 5335 92729 5354
rect 92343 5312 92409 5335
rect 92495 5312 92577 5335
rect 92663 5312 92729 5335
rect 92343 5272 92352 5312
rect 92392 5272 92409 5312
rect 92495 5272 92516 5312
rect 92556 5272 92577 5312
rect 92663 5272 92680 5312
rect 92720 5272 92729 5312
rect 92343 5249 92409 5272
rect 92495 5249 92577 5272
rect 92663 5249 92729 5272
rect 92343 5230 92729 5249
rect 96343 5335 96729 5354
rect 96343 5312 96409 5335
rect 96495 5312 96577 5335
rect 96663 5312 96729 5335
rect 96343 5272 96352 5312
rect 96392 5272 96409 5312
rect 96495 5272 96516 5312
rect 96556 5272 96577 5312
rect 96663 5272 96680 5312
rect 96720 5272 96729 5312
rect 96343 5249 96409 5272
rect 96495 5249 96577 5272
rect 96663 5249 96729 5272
rect 96343 5230 96729 5249
rect 3103 4579 3489 4598
rect 3103 4556 3169 4579
rect 3255 4556 3337 4579
rect 3423 4556 3489 4579
rect 3103 4516 3112 4556
rect 3152 4516 3169 4556
rect 3255 4516 3276 4556
rect 3316 4516 3337 4556
rect 3423 4516 3440 4556
rect 3480 4516 3489 4556
rect 3103 4493 3169 4516
rect 3255 4493 3337 4516
rect 3423 4493 3489 4516
rect 3103 4474 3489 4493
rect 7103 4579 7489 4598
rect 7103 4556 7169 4579
rect 7255 4556 7337 4579
rect 7423 4556 7489 4579
rect 7103 4516 7112 4556
rect 7152 4516 7169 4556
rect 7255 4516 7276 4556
rect 7316 4516 7337 4556
rect 7423 4516 7440 4556
rect 7480 4516 7489 4556
rect 7103 4493 7169 4516
rect 7255 4493 7337 4516
rect 7423 4493 7489 4516
rect 7103 4474 7489 4493
rect 11103 4579 11489 4598
rect 11103 4556 11169 4579
rect 11255 4556 11337 4579
rect 11423 4556 11489 4579
rect 11103 4516 11112 4556
rect 11152 4516 11169 4556
rect 11255 4516 11276 4556
rect 11316 4516 11337 4556
rect 11423 4516 11440 4556
rect 11480 4516 11489 4556
rect 11103 4493 11169 4516
rect 11255 4493 11337 4516
rect 11423 4493 11489 4516
rect 11103 4474 11489 4493
rect 15103 4579 15489 4598
rect 15103 4556 15169 4579
rect 15255 4556 15337 4579
rect 15423 4556 15489 4579
rect 15103 4516 15112 4556
rect 15152 4516 15169 4556
rect 15255 4516 15276 4556
rect 15316 4516 15337 4556
rect 15423 4516 15440 4556
rect 15480 4516 15489 4556
rect 15103 4493 15169 4516
rect 15255 4493 15337 4516
rect 15423 4493 15489 4516
rect 15103 4474 15489 4493
rect 19103 4579 19489 4598
rect 19103 4556 19169 4579
rect 19255 4556 19337 4579
rect 19423 4556 19489 4579
rect 19103 4516 19112 4556
rect 19152 4516 19169 4556
rect 19255 4516 19276 4556
rect 19316 4516 19337 4556
rect 19423 4516 19440 4556
rect 19480 4516 19489 4556
rect 19103 4493 19169 4516
rect 19255 4493 19337 4516
rect 19423 4493 19489 4516
rect 19103 4474 19489 4493
rect 23103 4579 23489 4598
rect 23103 4556 23169 4579
rect 23255 4556 23337 4579
rect 23423 4556 23489 4579
rect 23103 4516 23112 4556
rect 23152 4516 23169 4556
rect 23255 4516 23276 4556
rect 23316 4516 23337 4556
rect 23423 4516 23440 4556
rect 23480 4516 23489 4556
rect 23103 4493 23169 4516
rect 23255 4493 23337 4516
rect 23423 4493 23489 4516
rect 23103 4474 23489 4493
rect 27103 4579 27489 4598
rect 27103 4556 27169 4579
rect 27255 4556 27337 4579
rect 27423 4556 27489 4579
rect 27103 4516 27112 4556
rect 27152 4516 27169 4556
rect 27255 4516 27276 4556
rect 27316 4516 27337 4556
rect 27423 4516 27440 4556
rect 27480 4516 27489 4556
rect 27103 4493 27169 4516
rect 27255 4493 27337 4516
rect 27423 4493 27489 4516
rect 27103 4474 27489 4493
rect 31103 4579 31489 4598
rect 31103 4556 31169 4579
rect 31255 4556 31337 4579
rect 31423 4556 31489 4579
rect 31103 4516 31112 4556
rect 31152 4516 31169 4556
rect 31255 4516 31276 4556
rect 31316 4516 31337 4556
rect 31423 4516 31440 4556
rect 31480 4516 31489 4556
rect 31103 4493 31169 4516
rect 31255 4493 31337 4516
rect 31423 4493 31489 4516
rect 31103 4474 31489 4493
rect 35103 4579 35489 4598
rect 35103 4556 35169 4579
rect 35255 4556 35337 4579
rect 35423 4556 35489 4579
rect 35103 4516 35112 4556
rect 35152 4516 35169 4556
rect 35255 4516 35276 4556
rect 35316 4516 35337 4556
rect 35423 4516 35440 4556
rect 35480 4516 35489 4556
rect 35103 4493 35169 4516
rect 35255 4493 35337 4516
rect 35423 4493 35489 4516
rect 35103 4474 35489 4493
rect 39103 4579 39489 4598
rect 39103 4556 39169 4579
rect 39255 4556 39337 4579
rect 39423 4556 39489 4579
rect 39103 4516 39112 4556
rect 39152 4516 39169 4556
rect 39255 4516 39276 4556
rect 39316 4516 39337 4556
rect 39423 4516 39440 4556
rect 39480 4516 39489 4556
rect 39103 4493 39169 4516
rect 39255 4493 39337 4516
rect 39423 4493 39489 4516
rect 39103 4474 39489 4493
rect 43103 4579 43489 4598
rect 43103 4556 43169 4579
rect 43255 4556 43337 4579
rect 43423 4556 43489 4579
rect 43103 4516 43112 4556
rect 43152 4516 43169 4556
rect 43255 4516 43276 4556
rect 43316 4516 43337 4556
rect 43423 4516 43440 4556
rect 43480 4516 43489 4556
rect 43103 4493 43169 4516
rect 43255 4493 43337 4516
rect 43423 4493 43489 4516
rect 43103 4474 43489 4493
rect 47103 4579 47489 4598
rect 47103 4556 47169 4579
rect 47255 4556 47337 4579
rect 47423 4556 47489 4579
rect 47103 4516 47112 4556
rect 47152 4516 47169 4556
rect 47255 4516 47276 4556
rect 47316 4516 47337 4556
rect 47423 4516 47440 4556
rect 47480 4516 47489 4556
rect 47103 4493 47169 4516
rect 47255 4493 47337 4516
rect 47423 4493 47489 4516
rect 47103 4474 47489 4493
rect 51103 4579 51489 4598
rect 51103 4556 51169 4579
rect 51255 4556 51337 4579
rect 51423 4556 51489 4579
rect 51103 4516 51112 4556
rect 51152 4516 51169 4556
rect 51255 4516 51276 4556
rect 51316 4516 51337 4556
rect 51423 4516 51440 4556
rect 51480 4516 51489 4556
rect 51103 4493 51169 4516
rect 51255 4493 51337 4516
rect 51423 4493 51489 4516
rect 51103 4474 51489 4493
rect 55103 4579 55489 4598
rect 55103 4556 55169 4579
rect 55255 4556 55337 4579
rect 55423 4556 55489 4579
rect 55103 4516 55112 4556
rect 55152 4516 55169 4556
rect 55255 4516 55276 4556
rect 55316 4516 55337 4556
rect 55423 4516 55440 4556
rect 55480 4516 55489 4556
rect 55103 4493 55169 4516
rect 55255 4493 55337 4516
rect 55423 4493 55489 4516
rect 55103 4474 55489 4493
rect 59103 4579 59489 4598
rect 59103 4556 59169 4579
rect 59255 4556 59337 4579
rect 59423 4556 59489 4579
rect 59103 4516 59112 4556
rect 59152 4516 59169 4556
rect 59255 4516 59276 4556
rect 59316 4516 59337 4556
rect 59423 4516 59440 4556
rect 59480 4516 59489 4556
rect 59103 4493 59169 4516
rect 59255 4493 59337 4516
rect 59423 4493 59489 4516
rect 59103 4474 59489 4493
rect 63103 4579 63489 4598
rect 63103 4556 63169 4579
rect 63255 4556 63337 4579
rect 63423 4556 63489 4579
rect 63103 4516 63112 4556
rect 63152 4516 63169 4556
rect 63255 4516 63276 4556
rect 63316 4516 63337 4556
rect 63423 4516 63440 4556
rect 63480 4516 63489 4556
rect 63103 4493 63169 4516
rect 63255 4493 63337 4516
rect 63423 4493 63489 4516
rect 63103 4474 63489 4493
rect 67103 4579 67489 4598
rect 67103 4556 67169 4579
rect 67255 4556 67337 4579
rect 67423 4556 67489 4579
rect 67103 4516 67112 4556
rect 67152 4516 67169 4556
rect 67255 4516 67276 4556
rect 67316 4516 67337 4556
rect 67423 4516 67440 4556
rect 67480 4516 67489 4556
rect 67103 4493 67169 4516
rect 67255 4493 67337 4516
rect 67423 4493 67489 4516
rect 67103 4474 67489 4493
rect 71103 4579 71489 4598
rect 71103 4556 71169 4579
rect 71255 4556 71337 4579
rect 71423 4556 71489 4579
rect 71103 4516 71112 4556
rect 71152 4516 71169 4556
rect 71255 4516 71276 4556
rect 71316 4516 71337 4556
rect 71423 4516 71440 4556
rect 71480 4516 71489 4556
rect 71103 4493 71169 4516
rect 71255 4493 71337 4516
rect 71423 4493 71489 4516
rect 71103 4474 71489 4493
rect 75103 4579 75489 4598
rect 75103 4556 75169 4579
rect 75255 4556 75337 4579
rect 75423 4556 75489 4579
rect 75103 4516 75112 4556
rect 75152 4516 75169 4556
rect 75255 4516 75276 4556
rect 75316 4516 75337 4556
rect 75423 4516 75440 4556
rect 75480 4516 75489 4556
rect 75103 4493 75169 4516
rect 75255 4493 75337 4516
rect 75423 4493 75489 4516
rect 75103 4474 75489 4493
rect 79103 4579 79489 4598
rect 79103 4556 79169 4579
rect 79255 4556 79337 4579
rect 79423 4556 79489 4579
rect 79103 4516 79112 4556
rect 79152 4516 79169 4556
rect 79255 4516 79276 4556
rect 79316 4516 79337 4556
rect 79423 4516 79440 4556
rect 79480 4516 79489 4556
rect 79103 4493 79169 4516
rect 79255 4493 79337 4516
rect 79423 4493 79489 4516
rect 79103 4474 79489 4493
rect 83103 4579 83489 4598
rect 83103 4556 83169 4579
rect 83255 4556 83337 4579
rect 83423 4556 83489 4579
rect 83103 4516 83112 4556
rect 83152 4516 83169 4556
rect 83255 4516 83276 4556
rect 83316 4516 83337 4556
rect 83423 4516 83440 4556
rect 83480 4516 83489 4556
rect 83103 4493 83169 4516
rect 83255 4493 83337 4516
rect 83423 4493 83489 4516
rect 83103 4474 83489 4493
rect 87103 4579 87489 4598
rect 87103 4556 87169 4579
rect 87255 4556 87337 4579
rect 87423 4556 87489 4579
rect 87103 4516 87112 4556
rect 87152 4516 87169 4556
rect 87255 4516 87276 4556
rect 87316 4516 87337 4556
rect 87423 4516 87440 4556
rect 87480 4516 87489 4556
rect 87103 4493 87169 4516
rect 87255 4493 87337 4516
rect 87423 4493 87489 4516
rect 87103 4474 87489 4493
rect 91103 4579 91489 4598
rect 91103 4556 91169 4579
rect 91255 4556 91337 4579
rect 91423 4556 91489 4579
rect 91103 4516 91112 4556
rect 91152 4516 91169 4556
rect 91255 4516 91276 4556
rect 91316 4516 91337 4556
rect 91423 4516 91440 4556
rect 91480 4516 91489 4556
rect 91103 4493 91169 4516
rect 91255 4493 91337 4516
rect 91423 4493 91489 4516
rect 91103 4474 91489 4493
rect 95103 4579 95489 4598
rect 95103 4556 95169 4579
rect 95255 4556 95337 4579
rect 95423 4556 95489 4579
rect 95103 4516 95112 4556
rect 95152 4516 95169 4556
rect 95255 4516 95276 4556
rect 95316 4516 95337 4556
rect 95423 4516 95440 4556
rect 95480 4516 95489 4556
rect 95103 4493 95169 4516
rect 95255 4493 95337 4516
rect 95423 4493 95489 4516
rect 95103 4474 95489 4493
rect 99103 4579 99489 4598
rect 99103 4556 99169 4579
rect 99255 4556 99337 4579
rect 99423 4556 99489 4579
rect 99103 4516 99112 4556
rect 99152 4516 99169 4556
rect 99255 4516 99276 4556
rect 99316 4516 99337 4556
rect 99423 4516 99440 4556
rect 99480 4516 99489 4556
rect 99103 4493 99169 4516
rect 99255 4493 99337 4516
rect 99423 4493 99489 4516
rect 99103 4474 99489 4493
rect 4343 3823 4729 3842
rect 4343 3800 4409 3823
rect 4495 3800 4577 3823
rect 4663 3800 4729 3823
rect 4343 3760 4352 3800
rect 4392 3760 4409 3800
rect 4495 3760 4516 3800
rect 4556 3760 4577 3800
rect 4663 3760 4680 3800
rect 4720 3760 4729 3800
rect 4343 3737 4409 3760
rect 4495 3737 4577 3760
rect 4663 3737 4729 3760
rect 4343 3718 4729 3737
rect 8343 3823 8729 3842
rect 8343 3800 8409 3823
rect 8495 3800 8577 3823
rect 8663 3800 8729 3823
rect 8343 3760 8352 3800
rect 8392 3760 8409 3800
rect 8495 3760 8516 3800
rect 8556 3760 8577 3800
rect 8663 3760 8680 3800
rect 8720 3760 8729 3800
rect 8343 3737 8409 3760
rect 8495 3737 8577 3760
rect 8663 3737 8729 3760
rect 8343 3718 8729 3737
rect 12343 3823 12729 3842
rect 12343 3800 12409 3823
rect 12495 3800 12577 3823
rect 12663 3800 12729 3823
rect 12343 3760 12352 3800
rect 12392 3760 12409 3800
rect 12495 3760 12516 3800
rect 12556 3760 12577 3800
rect 12663 3760 12680 3800
rect 12720 3760 12729 3800
rect 12343 3737 12409 3760
rect 12495 3737 12577 3760
rect 12663 3737 12729 3760
rect 12343 3718 12729 3737
rect 16343 3823 16729 3842
rect 16343 3800 16409 3823
rect 16495 3800 16577 3823
rect 16663 3800 16729 3823
rect 16343 3760 16352 3800
rect 16392 3760 16409 3800
rect 16495 3760 16516 3800
rect 16556 3760 16577 3800
rect 16663 3760 16680 3800
rect 16720 3760 16729 3800
rect 16343 3737 16409 3760
rect 16495 3737 16577 3760
rect 16663 3737 16729 3760
rect 16343 3718 16729 3737
rect 20343 3823 20729 3842
rect 20343 3800 20409 3823
rect 20495 3800 20577 3823
rect 20663 3800 20729 3823
rect 20343 3760 20352 3800
rect 20392 3760 20409 3800
rect 20495 3760 20516 3800
rect 20556 3760 20577 3800
rect 20663 3760 20680 3800
rect 20720 3760 20729 3800
rect 20343 3737 20409 3760
rect 20495 3737 20577 3760
rect 20663 3737 20729 3760
rect 20343 3718 20729 3737
rect 24343 3823 24729 3842
rect 24343 3800 24409 3823
rect 24495 3800 24577 3823
rect 24663 3800 24729 3823
rect 24343 3760 24352 3800
rect 24392 3760 24409 3800
rect 24495 3760 24516 3800
rect 24556 3760 24577 3800
rect 24663 3760 24680 3800
rect 24720 3760 24729 3800
rect 24343 3737 24409 3760
rect 24495 3737 24577 3760
rect 24663 3737 24729 3760
rect 24343 3718 24729 3737
rect 28343 3823 28729 3842
rect 28343 3800 28409 3823
rect 28495 3800 28577 3823
rect 28663 3800 28729 3823
rect 28343 3760 28352 3800
rect 28392 3760 28409 3800
rect 28495 3760 28516 3800
rect 28556 3760 28577 3800
rect 28663 3760 28680 3800
rect 28720 3760 28729 3800
rect 28343 3737 28409 3760
rect 28495 3737 28577 3760
rect 28663 3737 28729 3760
rect 28343 3718 28729 3737
rect 32343 3823 32729 3842
rect 32343 3800 32409 3823
rect 32495 3800 32577 3823
rect 32663 3800 32729 3823
rect 32343 3760 32352 3800
rect 32392 3760 32409 3800
rect 32495 3760 32516 3800
rect 32556 3760 32577 3800
rect 32663 3760 32680 3800
rect 32720 3760 32729 3800
rect 32343 3737 32409 3760
rect 32495 3737 32577 3760
rect 32663 3737 32729 3760
rect 32343 3718 32729 3737
rect 36343 3823 36729 3842
rect 36343 3800 36409 3823
rect 36495 3800 36577 3823
rect 36663 3800 36729 3823
rect 36343 3760 36352 3800
rect 36392 3760 36409 3800
rect 36495 3760 36516 3800
rect 36556 3760 36577 3800
rect 36663 3760 36680 3800
rect 36720 3760 36729 3800
rect 36343 3737 36409 3760
rect 36495 3737 36577 3760
rect 36663 3737 36729 3760
rect 36343 3718 36729 3737
rect 40343 3823 40729 3842
rect 40343 3800 40409 3823
rect 40495 3800 40577 3823
rect 40663 3800 40729 3823
rect 40343 3760 40352 3800
rect 40392 3760 40409 3800
rect 40495 3760 40516 3800
rect 40556 3760 40577 3800
rect 40663 3760 40680 3800
rect 40720 3760 40729 3800
rect 40343 3737 40409 3760
rect 40495 3737 40577 3760
rect 40663 3737 40729 3760
rect 40343 3718 40729 3737
rect 44343 3823 44729 3842
rect 44343 3800 44409 3823
rect 44495 3800 44577 3823
rect 44663 3800 44729 3823
rect 44343 3760 44352 3800
rect 44392 3760 44409 3800
rect 44495 3760 44516 3800
rect 44556 3760 44577 3800
rect 44663 3760 44680 3800
rect 44720 3760 44729 3800
rect 44343 3737 44409 3760
rect 44495 3737 44577 3760
rect 44663 3737 44729 3760
rect 44343 3718 44729 3737
rect 48343 3823 48729 3842
rect 48343 3800 48409 3823
rect 48495 3800 48577 3823
rect 48663 3800 48729 3823
rect 48343 3760 48352 3800
rect 48392 3760 48409 3800
rect 48495 3760 48516 3800
rect 48556 3760 48577 3800
rect 48663 3760 48680 3800
rect 48720 3760 48729 3800
rect 48343 3737 48409 3760
rect 48495 3737 48577 3760
rect 48663 3737 48729 3760
rect 48343 3718 48729 3737
rect 52343 3823 52729 3842
rect 52343 3800 52409 3823
rect 52495 3800 52577 3823
rect 52663 3800 52729 3823
rect 52343 3760 52352 3800
rect 52392 3760 52409 3800
rect 52495 3760 52516 3800
rect 52556 3760 52577 3800
rect 52663 3760 52680 3800
rect 52720 3760 52729 3800
rect 52343 3737 52409 3760
rect 52495 3737 52577 3760
rect 52663 3737 52729 3760
rect 52343 3718 52729 3737
rect 56343 3823 56729 3842
rect 56343 3800 56409 3823
rect 56495 3800 56577 3823
rect 56663 3800 56729 3823
rect 56343 3760 56352 3800
rect 56392 3760 56409 3800
rect 56495 3760 56516 3800
rect 56556 3760 56577 3800
rect 56663 3760 56680 3800
rect 56720 3760 56729 3800
rect 56343 3737 56409 3760
rect 56495 3737 56577 3760
rect 56663 3737 56729 3760
rect 56343 3718 56729 3737
rect 60343 3823 60729 3842
rect 60343 3800 60409 3823
rect 60495 3800 60577 3823
rect 60663 3800 60729 3823
rect 60343 3760 60352 3800
rect 60392 3760 60409 3800
rect 60495 3760 60516 3800
rect 60556 3760 60577 3800
rect 60663 3760 60680 3800
rect 60720 3760 60729 3800
rect 60343 3737 60409 3760
rect 60495 3737 60577 3760
rect 60663 3737 60729 3760
rect 60343 3718 60729 3737
rect 64343 3823 64729 3842
rect 64343 3800 64409 3823
rect 64495 3800 64577 3823
rect 64663 3800 64729 3823
rect 64343 3760 64352 3800
rect 64392 3760 64409 3800
rect 64495 3760 64516 3800
rect 64556 3760 64577 3800
rect 64663 3760 64680 3800
rect 64720 3760 64729 3800
rect 64343 3737 64409 3760
rect 64495 3737 64577 3760
rect 64663 3737 64729 3760
rect 64343 3718 64729 3737
rect 68343 3823 68729 3842
rect 68343 3800 68409 3823
rect 68495 3800 68577 3823
rect 68663 3800 68729 3823
rect 68343 3760 68352 3800
rect 68392 3760 68409 3800
rect 68495 3760 68516 3800
rect 68556 3760 68577 3800
rect 68663 3760 68680 3800
rect 68720 3760 68729 3800
rect 68343 3737 68409 3760
rect 68495 3737 68577 3760
rect 68663 3737 68729 3760
rect 68343 3718 68729 3737
rect 72343 3823 72729 3842
rect 72343 3800 72409 3823
rect 72495 3800 72577 3823
rect 72663 3800 72729 3823
rect 72343 3760 72352 3800
rect 72392 3760 72409 3800
rect 72495 3760 72516 3800
rect 72556 3760 72577 3800
rect 72663 3760 72680 3800
rect 72720 3760 72729 3800
rect 72343 3737 72409 3760
rect 72495 3737 72577 3760
rect 72663 3737 72729 3760
rect 72343 3718 72729 3737
rect 76343 3823 76729 3842
rect 76343 3800 76409 3823
rect 76495 3800 76577 3823
rect 76663 3800 76729 3823
rect 76343 3760 76352 3800
rect 76392 3760 76409 3800
rect 76495 3760 76516 3800
rect 76556 3760 76577 3800
rect 76663 3760 76680 3800
rect 76720 3760 76729 3800
rect 76343 3737 76409 3760
rect 76495 3737 76577 3760
rect 76663 3737 76729 3760
rect 76343 3718 76729 3737
rect 80343 3823 80729 3842
rect 80343 3800 80409 3823
rect 80495 3800 80577 3823
rect 80663 3800 80729 3823
rect 80343 3760 80352 3800
rect 80392 3760 80409 3800
rect 80495 3760 80516 3800
rect 80556 3760 80577 3800
rect 80663 3760 80680 3800
rect 80720 3760 80729 3800
rect 80343 3737 80409 3760
rect 80495 3737 80577 3760
rect 80663 3737 80729 3760
rect 80343 3718 80729 3737
rect 84343 3823 84729 3842
rect 84343 3800 84409 3823
rect 84495 3800 84577 3823
rect 84663 3800 84729 3823
rect 84343 3760 84352 3800
rect 84392 3760 84409 3800
rect 84495 3760 84516 3800
rect 84556 3760 84577 3800
rect 84663 3760 84680 3800
rect 84720 3760 84729 3800
rect 84343 3737 84409 3760
rect 84495 3737 84577 3760
rect 84663 3737 84729 3760
rect 84343 3718 84729 3737
rect 88343 3823 88729 3842
rect 88343 3800 88409 3823
rect 88495 3800 88577 3823
rect 88663 3800 88729 3823
rect 88343 3760 88352 3800
rect 88392 3760 88409 3800
rect 88495 3760 88516 3800
rect 88556 3760 88577 3800
rect 88663 3760 88680 3800
rect 88720 3760 88729 3800
rect 88343 3737 88409 3760
rect 88495 3737 88577 3760
rect 88663 3737 88729 3760
rect 88343 3718 88729 3737
rect 92343 3823 92729 3842
rect 92343 3800 92409 3823
rect 92495 3800 92577 3823
rect 92663 3800 92729 3823
rect 92343 3760 92352 3800
rect 92392 3760 92409 3800
rect 92495 3760 92516 3800
rect 92556 3760 92577 3800
rect 92663 3760 92680 3800
rect 92720 3760 92729 3800
rect 92343 3737 92409 3760
rect 92495 3737 92577 3760
rect 92663 3737 92729 3760
rect 92343 3718 92729 3737
rect 96343 3823 96729 3842
rect 96343 3800 96409 3823
rect 96495 3800 96577 3823
rect 96663 3800 96729 3823
rect 96343 3760 96352 3800
rect 96392 3760 96409 3800
rect 96495 3760 96516 3800
rect 96556 3760 96577 3800
rect 96663 3760 96680 3800
rect 96720 3760 96729 3800
rect 96343 3737 96409 3760
rect 96495 3737 96577 3760
rect 96663 3737 96729 3760
rect 96343 3718 96729 3737
rect 3103 3067 3489 3086
rect 3103 3044 3169 3067
rect 3255 3044 3337 3067
rect 3423 3044 3489 3067
rect 3103 3004 3112 3044
rect 3152 3004 3169 3044
rect 3255 3004 3276 3044
rect 3316 3004 3337 3044
rect 3423 3004 3440 3044
rect 3480 3004 3489 3044
rect 3103 2981 3169 3004
rect 3255 2981 3337 3004
rect 3423 2981 3489 3004
rect 3103 2962 3489 2981
rect 7103 3067 7489 3086
rect 7103 3044 7169 3067
rect 7255 3044 7337 3067
rect 7423 3044 7489 3067
rect 7103 3004 7112 3044
rect 7152 3004 7169 3044
rect 7255 3004 7276 3044
rect 7316 3004 7337 3044
rect 7423 3004 7440 3044
rect 7480 3004 7489 3044
rect 7103 2981 7169 3004
rect 7255 2981 7337 3004
rect 7423 2981 7489 3004
rect 7103 2962 7489 2981
rect 11103 3067 11489 3086
rect 11103 3044 11169 3067
rect 11255 3044 11337 3067
rect 11423 3044 11489 3067
rect 11103 3004 11112 3044
rect 11152 3004 11169 3044
rect 11255 3004 11276 3044
rect 11316 3004 11337 3044
rect 11423 3004 11440 3044
rect 11480 3004 11489 3044
rect 11103 2981 11169 3004
rect 11255 2981 11337 3004
rect 11423 2981 11489 3004
rect 11103 2962 11489 2981
rect 15103 3067 15489 3086
rect 15103 3044 15169 3067
rect 15255 3044 15337 3067
rect 15423 3044 15489 3067
rect 15103 3004 15112 3044
rect 15152 3004 15169 3044
rect 15255 3004 15276 3044
rect 15316 3004 15337 3044
rect 15423 3004 15440 3044
rect 15480 3004 15489 3044
rect 15103 2981 15169 3004
rect 15255 2981 15337 3004
rect 15423 2981 15489 3004
rect 15103 2962 15489 2981
rect 19103 3067 19489 3086
rect 19103 3044 19169 3067
rect 19255 3044 19337 3067
rect 19423 3044 19489 3067
rect 19103 3004 19112 3044
rect 19152 3004 19169 3044
rect 19255 3004 19276 3044
rect 19316 3004 19337 3044
rect 19423 3004 19440 3044
rect 19480 3004 19489 3044
rect 19103 2981 19169 3004
rect 19255 2981 19337 3004
rect 19423 2981 19489 3004
rect 19103 2962 19489 2981
rect 23103 3067 23489 3086
rect 23103 3044 23169 3067
rect 23255 3044 23337 3067
rect 23423 3044 23489 3067
rect 23103 3004 23112 3044
rect 23152 3004 23169 3044
rect 23255 3004 23276 3044
rect 23316 3004 23337 3044
rect 23423 3004 23440 3044
rect 23480 3004 23489 3044
rect 23103 2981 23169 3004
rect 23255 2981 23337 3004
rect 23423 2981 23489 3004
rect 23103 2962 23489 2981
rect 27103 3067 27489 3086
rect 27103 3044 27169 3067
rect 27255 3044 27337 3067
rect 27423 3044 27489 3067
rect 27103 3004 27112 3044
rect 27152 3004 27169 3044
rect 27255 3004 27276 3044
rect 27316 3004 27337 3044
rect 27423 3004 27440 3044
rect 27480 3004 27489 3044
rect 27103 2981 27169 3004
rect 27255 2981 27337 3004
rect 27423 2981 27489 3004
rect 27103 2962 27489 2981
rect 31103 3067 31489 3086
rect 31103 3044 31169 3067
rect 31255 3044 31337 3067
rect 31423 3044 31489 3067
rect 31103 3004 31112 3044
rect 31152 3004 31169 3044
rect 31255 3004 31276 3044
rect 31316 3004 31337 3044
rect 31423 3004 31440 3044
rect 31480 3004 31489 3044
rect 31103 2981 31169 3004
rect 31255 2981 31337 3004
rect 31423 2981 31489 3004
rect 31103 2962 31489 2981
rect 35103 3067 35489 3086
rect 35103 3044 35169 3067
rect 35255 3044 35337 3067
rect 35423 3044 35489 3067
rect 35103 3004 35112 3044
rect 35152 3004 35169 3044
rect 35255 3004 35276 3044
rect 35316 3004 35337 3044
rect 35423 3004 35440 3044
rect 35480 3004 35489 3044
rect 35103 2981 35169 3004
rect 35255 2981 35337 3004
rect 35423 2981 35489 3004
rect 35103 2962 35489 2981
rect 39103 3067 39489 3086
rect 39103 3044 39169 3067
rect 39255 3044 39337 3067
rect 39423 3044 39489 3067
rect 39103 3004 39112 3044
rect 39152 3004 39169 3044
rect 39255 3004 39276 3044
rect 39316 3004 39337 3044
rect 39423 3004 39440 3044
rect 39480 3004 39489 3044
rect 39103 2981 39169 3004
rect 39255 2981 39337 3004
rect 39423 2981 39489 3004
rect 39103 2962 39489 2981
rect 43103 3067 43489 3086
rect 43103 3044 43169 3067
rect 43255 3044 43337 3067
rect 43423 3044 43489 3067
rect 43103 3004 43112 3044
rect 43152 3004 43169 3044
rect 43255 3004 43276 3044
rect 43316 3004 43337 3044
rect 43423 3004 43440 3044
rect 43480 3004 43489 3044
rect 43103 2981 43169 3004
rect 43255 2981 43337 3004
rect 43423 2981 43489 3004
rect 43103 2962 43489 2981
rect 47103 3067 47489 3086
rect 47103 3044 47169 3067
rect 47255 3044 47337 3067
rect 47423 3044 47489 3067
rect 47103 3004 47112 3044
rect 47152 3004 47169 3044
rect 47255 3004 47276 3044
rect 47316 3004 47337 3044
rect 47423 3004 47440 3044
rect 47480 3004 47489 3044
rect 47103 2981 47169 3004
rect 47255 2981 47337 3004
rect 47423 2981 47489 3004
rect 47103 2962 47489 2981
rect 51103 3067 51489 3086
rect 51103 3044 51169 3067
rect 51255 3044 51337 3067
rect 51423 3044 51489 3067
rect 51103 3004 51112 3044
rect 51152 3004 51169 3044
rect 51255 3004 51276 3044
rect 51316 3004 51337 3044
rect 51423 3004 51440 3044
rect 51480 3004 51489 3044
rect 51103 2981 51169 3004
rect 51255 2981 51337 3004
rect 51423 2981 51489 3004
rect 51103 2962 51489 2981
rect 55103 3067 55489 3086
rect 55103 3044 55169 3067
rect 55255 3044 55337 3067
rect 55423 3044 55489 3067
rect 55103 3004 55112 3044
rect 55152 3004 55169 3044
rect 55255 3004 55276 3044
rect 55316 3004 55337 3044
rect 55423 3004 55440 3044
rect 55480 3004 55489 3044
rect 55103 2981 55169 3004
rect 55255 2981 55337 3004
rect 55423 2981 55489 3004
rect 55103 2962 55489 2981
rect 59103 3067 59489 3086
rect 59103 3044 59169 3067
rect 59255 3044 59337 3067
rect 59423 3044 59489 3067
rect 59103 3004 59112 3044
rect 59152 3004 59169 3044
rect 59255 3004 59276 3044
rect 59316 3004 59337 3044
rect 59423 3004 59440 3044
rect 59480 3004 59489 3044
rect 59103 2981 59169 3004
rect 59255 2981 59337 3004
rect 59423 2981 59489 3004
rect 59103 2962 59489 2981
rect 63103 3067 63489 3086
rect 63103 3044 63169 3067
rect 63255 3044 63337 3067
rect 63423 3044 63489 3067
rect 63103 3004 63112 3044
rect 63152 3004 63169 3044
rect 63255 3004 63276 3044
rect 63316 3004 63337 3044
rect 63423 3004 63440 3044
rect 63480 3004 63489 3044
rect 63103 2981 63169 3004
rect 63255 2981 63337 3004
rect 63423 2981 63489 3004
rect 63103 2962 63489 2981
rect 67103 3067 67489 3086
rect 67103 3044 67169 3067
rect 67255 3044 67337 3067
rect 67423 3044 67489 3067
rect 67103 3004 67112 3044
rect 67152 3004 67169 3044
rect 67255 3004 67276 3044
rect 67316 3004 67337 3044
rect 67423 3004 67440 3044
rect 67480 3004 67489 3044
rect 67103 2981 67169 3004
rect 67255 2981 67337 3004
rect 67423 2981 67489 3004
rect 67103 2962 67489 2981
rect 71103 3067 71489 3086
rect 71103 3044 71169 3067
rect 71255 3044 71337 3067
rect 71423 3044 71489 3067
rect 71103 3004 71112 3044
rect 71152 3004 71169 3044
rect 71255 3004 71276 3044
rect 71316 3004 71337 3044
rect 71423 3004 71440 3044
rect 71480 3004 71489 3044
rect 71103 2981 71169 3004
rect 71255 2981 71337 3004
rect 71423 2981 71489 3004
rect 71103 2962 71489 2981
rect 75103 3067 75489 3086
rect 75103 3044 75169 3067
rect 75255 3044 75337 3067
rect 75423 3044 75489 3067
rect 75103 3004 75112 3044
rect 75152 3004 75169 3044
rect 75255 3004 75276 3044
rect 75316 3004 75337 3044
rect 75423 3004 75440 3044
rect 75480 3004 75489 3044
rect 75103 2981 75169 3004
rect 75255 2981 75337 3004
rect 75423 2981 75489 3004
rect 75103 2962 75489 2981
rect 79103 3067 79489 3086
rect 79103 3044 79169 3067
rect 79255 3044 79337 3067
rect 79423 3044 79489 3067
rect 79103 3004 79112 3044
rect 79152 3004 79169 3044
rect 79255 3004 79276 3044
rect 79316 3004 79337 3044
rect 79423 3004 79440 3044
rect 79480 3004 79489 3044
rect 79103 2981 79169 3004
rect 79255 2981 79337 3004
rect 79423 2981 79489 3004
rect 79103 2962 79489 2981
rect 83103 3067 83489 3086
rect 83103 3044 83169 3067
rect 83255 3044 83337 3067
rect 83423 3044 83489 3067
rect 83103 3004 83112 3044
rect 83152 3004 83169 3044
rect 83255 3004 83276 3044
rect 83316 3004 83337 3044
rect 83423 3004 83440 3044
rect 83480 3004 83489 3044
rect 83103 2981 83169 3004
rect 83255 2981 83337 3004
rect 83423 2981 83489 3004
rect 83103 2962 83489 2981
rect 87103 3067 87489 3086
rect 87103 3044 87169 3067
rect 87255 3044 87337 3067
rect 87423 3044 87489 3067
rect 87103 3004 87112 3044
rect 87152 3004 87169 3044
rect 87255 3004 87276 3044
rect 87316 3004 87337 3044
rect 87423 3004 87440 3044
rect 87480 3004 87489 3044
rect 87103 2981 87169 3004
rect 87255 2981 87337 3004
rect 87423 2981 87489 3004
rect 87103 2962 87489 2981
rect 91103 3067 91489 3086
rect 91103 3044 91169 3067
rect 91255 3044 91337 3067
rect 91423 3044 91489 3067
rect 91103 3004 91112 3044
rect 91152 3004 91169 3044
rect 91255 3004 91276 3044
rect 91316 3004 91337 3044
rect 91423 3004 91440 3044
rect 91480 3004 91489 3044
rect 91103 2981 91169 3004
rect 91255 2981 91337 3004
rect 91423 2981 91489 3004
rect 91103 2962 91489 2981
rect 95103 3067 95489 3086
rect 95103 3044 95169 3067
rect 95255 3044 95337 3067
rect 95423 3044 95489 3067
rect 95103 3004 95112 3044
rect 95152 3004 95169 3044
rect 95255 3004 95276 3044
rect 95316 3004 95337 3044
rect 95423 3004 95440 3044
rect 95480 3004 95489 3044
rect 95103 2981 95169 3004
rect 95255 2981 95337 3004
rect 95423 2981 95489 3004
rect 95103 2962 95489 2981
rect 99103 3067 99489 3086
rect 99103 3044 99169 3067
rect 99255 3044 99337 3067
rect 99423 3044 99489 3067
rect 99103 3004 99112 3044
rect 99152 3004 99169 3044
rect 99255 3004 99276 3044
rect 99316 3004 99337 3044
rect 99423 3004 99440 3044
rect 99480 3004 99489 3044
rect 99103 2981 99169 3004
rect 99255 2981 99337 3004
rect 99423 2981 99489 3004
rect 99103 2962 99489 2981
rect 4343 2311 4729 2330
rect 4343 2288 4409 2311
rect 4495 2288 4577 2311
rect 4663 2288 4729 2311
rect 4343 2248 4352 2288
rect 4392 2248 4409 2288
rect 4495 2248 4516 2288
rect 4556 2248 4577 2288
rect 4663 2248 4680 2288
rect 4720 2248 4729 2288
rect 4343 2225 4409 2248
rect 4495 2225 4577 2248
rect 4663 2225 4729 2248
rect 4343 2206 4729 2225
rect 8343 2311 8729 2330
rect 8343 2288 8409 2311
rect 8495 2288 8577 2311
rect 8663 2288 8729 2311
rect 8343 2248 8352 2288
rect 8392 2248 8409 2288
rect 8495 2248 8516 2288
rect 8556 2248 8577 2288
rect 8663 2248 8680 2288
rect 8720 2248 8729 2288
rect 8343 2225 8409 2248
rect 8495 2225 8577 2248
rect 8663 2225 8729 2248
rect 8343 2206 8729 2225
rect 12343 2311 12729 2330
rect 12343 2288 12409 2311
rect 12495 2288 12577 2311
rect 12663 2288 12729 2311
rect 12343 2248 12352 2288
rect 12392 2248 12409 2288
rect 12495 2248 12516 2288
rect 12556 2248 12577 2288
rect 12663 2248 12680 2288
rect 12720 2248 12729 2288
rect 12343 2225 12409 2248
rect 12495 2225 12577 2248
rect 12663 2225 12729 2248
rect 12343 2206 12729 2225
rect 16343 2311 16729 2330
rect 16343 2288 16409 2311
rect 16495 2288 16577 2311
rect 16663 2288 16729 2311
rect 16343 2248 16352 2288
rect 16392 2248 16409 2288
rect 16495 2248 16516 2288
rect 16556 2248 16577 2288
rect 16663 2248 16680 2288
rect 16720 2248 16729 2288
rect 16343 2225 16409 2248
rect 16495 2225 16577 2248
rect 16663 2225 16729 2248
rect 16343 2206 16729 2225
rect 20343 2311 20729 2330
rect 20343 2288 20409 2311
rect 20495 2288 20577 2311
rect 20663 2288 20729 2311
rect 20343 2248 20352 2288
rect 20392 2248 20409 2288
rect 20495 2248 20516 2288
rect 20556 2248 20577 2288
rect 20663 2248 20680 2288
rect 20720 2248 20729 2288
rect 20343 2225 20409 2248
rect 20495 2225 20577 2248
rect 20663 2225 20729 2248
rect 20343 2206 20729 2225
rect 24343 2311 24729 2330
rect 24343 2288 24409 2311
rect 24495 2288 24577 2311
rect 24663 2288 24729 2311
rect 24343 2248 24352 2288
rect 24392 2248 24409 2288
rect 24495 2248 24516 2288
rect 24556 2248 24577 2288
rect 24663 2248 24680 2288
rect 24720 2248 24729 2288
rect 24343 2225 24409 2248
rect 24495 2225 24577 2248
rect 24663 2225 24729 2248
rect 24343 2206 24729 2225
rect 28343 2311 28729 2330
rect 28343 2288 28409 2311
rect 28495 2288 28577 2311
rect 28663 2288 28729 2311
rect 28343 2248 28352 2288
rect 28392 2248 28409 2288
rect 28495 2248 28516 2288
rect 28556 2248 28577 2288
rect 28663 2248 28680 2288
rect 28720 2248 28729 2288
rect 28343 2225 28409 2248
rect 28495 2225 28577 2248
rect 28663 2225 28729 2248
rect 28343 2206 28729 2225
rect 32343 2311 32729 2330
rect 32343 2288 32409 2311
rect 32495 2288 32577 2311
rect 32663 2288 32729 2311
rect 32343 2248 32352 2288
rect 32392 2248 32409 2288
rect 32495 2248 32516 2288
rect 32556 2248 32577 2288
rect 32663 2248 32680 2288
rect 32720 2248 32729 2288
rect 32343 2225 32409 2248
rect 32495 2225 32577 2248
rect 32663 2225 32729 2248
rect 32343 2206 32729 2225
rect 36343 2311 36729 2330
rect 36343 2288 36409 2311
rect 36495 2288 36577 2311
rect 36663 2288 36729 2311
rect 36343 2248 36352 2288
rect 36392 2248 36409 2288
rect 36495 2248 36516 2288
rect 36556 2248 36577 2288
rect 36663 2248 36680 2288
rect 36720 2248 36729 2288
rect 36343 2225 36409 2248
rect 36495 2225 36577 2248
rect 36663 2225 36729 2248
rect 36343 2206 36729 2225
rect 40343 2311 40729 2330
rect 40343 2288 40409 2311
rect 40495 2288 40577 2311
rect 40663 2288 40729 2311
rect 40343 2248 40352 2288
rect 40392 2248 40409 2288
rect 40495 2248 40516 2288
rect 40556 2248 40577 2288
rect 40663 2248 40680 2288
rect 40720 2248 40729 2288
rect 40343 2225 40409 2248
rect 40495 2225 40577 2248
rect 40663 2225 40729 2248
rect 40343 2206 40729 2225
rect 44343 2311 44729 2330
rect 44343 2288 44409 2311
rect 44495 2288 44577 2311
rect 44663 2288 44729 2311
rect 44343 2248 44352 2288
rect 44392 2248 44409 2288
rect 44495 2248 44516 2288
rect 44556 2248 44577 2288
rect 44663 2248 44680 2288
rect 44720 2248 44729 2288
rect 44343 2225 44409 2248
rect 44495 2225 44577 2248
rect 44663 2225 44729 2248
rect 44343 2206 44729 2225
rect 48343 2311 48729 2330
rect 48343 2288 48409 2311
rect 48495 2288 48577 2311
rect 48663 2288 48729 2311
rect 48343 2248 48352 2288
rect 48392 2248 48409 2288
rect 48495 2248 48516 2288
rect 48556 2248 48577 2288
rect 48663 2248 48680 2288
rect 48720 2248 48729 2288
rect 48343 2225 48409 2248
rect 48495 2225 48577 2248
rect 48663 2225 48729 2248
rect 48343 2206 48729 2225
rect 52343 2311 52729 2330
rect 52343 2288 52409 2311
rect 52495 2288 52577 2311
rect 52663 2288 52729 2311
rect 52343 2248 52352 2288
rect 52392 2248 52409 2288
rect 52495 2248 52516 2288
rect 52556 2248 52577 2288
rect 52663 2248 52680 2288
rect 52720 2248 52729 2288
rect 52343 2225 52409 2248
rect 52495 2225 52577 2248
rect 52663 2225 52729 2248
rect 52343 2206 52729 2225
rect 56343 2311 56729 2330
rect 56343 2288 56409 2311
rect 56495 2288 56577 2311
rect 56663 2288 56729 2311
rect 56343 2248 56352 2288
rect 56392 2248 56409 2288
rect 56495 2248 56516 2288
rect 56556 2248 56577 2288
rect 56663 2248 56680 2288
rect 56720 2248 56729 2288
rect 56343 2225 56409 2248
rect 56495 2225 56577 2248
rect 56663 2225 56729 2248
rect 56343 2206 56729 2225
rect 60343 2311 60729 2330
rect 60343 2288 60409 2311
rect 60495 2288 60577 2311
rect 60663 2288 60729 2311
rect 60343 2248 60352 2288
rect 60392 2248 60409 2288
rect 60495 2248 60516 2288
rect 60556 2248 60577 2288
rect 60663 2248 60680 2288
rect 60720 2248 60729 2288
rect 60343 2225 60409 2248
rect 60495 2225 60577 2248
rect 60663 2225 60729 2248
rect 60343 2206 60729 2225
rect 64343 2311 64729 2330
rect 64343 2288 64409 2311
rect 64495 2288 64577 2311
rect 64663 2288 64729 2311
rect 64343 2248 64352 2288
rect 64392 2248 64409 2288
rect 64495 2248 64516 2288
rect 64556 2248 64577 2288
rect 64663 2248 64680 2288
rect 64720 2248 64729 2288
rect 64343 2225 64409 2248
rect 64495 2225 64577 2248
rect 64663 2225 64729 2248
rect 64343 2206 64729 2225
rect 68343 2311 68729 2330
rect 68343 2288 68409 2311
rect 68495 2288 68577 2311
rect 68663 2288 68729 2311
rect 68343 2248 68352 2288
rect 68392 2248 68409 2288
rect 68495 2248 68516 2288
rect 68556 2248 68577 2288
rect 68663 2248 68680 2288
rect 68720 2248 68729 2288
rect 68343 2225 68409 2248
rect 68495 2225 68577 2248
rect 68663 2225 68729 2248
rect 68343 2206 68729 2225
rect 72343 2311 72729 2330
rect 72343 2288 72409 2311
rect 72495 2288 72577 2311
rect 72663 2288 72729 2311
rect 72343 2248 72352 2288
rect 72392 2248 72409 2288
rect 72495 2248 72516 2288
rect 72556 2248 72577 2288
rect 72663 2248 72680 2288
rect 72720 2248 72729 2288
rect 72343 2225 72409 2248
rect 72495 2225 72577 2248
rect 72663 2225 72729 2248
rect 72343 2206 72729 2225
rect 76343 2311 76729 2330
rect 76343 2288 76409 2311
rect 76495 2288 76577 2311
rect 76663 2288 76729 2311
rect 76343 2248 76352 2288
rect 76392 2248 76409 2288
rect 76495 2248 76516 2288
rect 76556 2248 76577 2288
rect 76663 2248 76680 2288
rect 76720 2248 76729 2288
rect 76343 2225 76409 2248
rect 76495 2225 76577 2248
rect 76663 2225 76729 2248
rect 76343 2206 76729 2225
rect 80343 2311 80729 2330
rect 80343 2288 80409 2311
rect 80495 2288 80577 2311
rect 80663 2288 80729 2311
rect 80343 2248 80352 2288
rect 80392 2248 80409 2288
rect 80495 2248 80516 2288
rect 80556 2248 80577 2288
rect 80663 2248 80680 2288
rect 80720 2248 80729 2288
rect 80343 2225 80409 2248
rect 80495 2225 80577 2248
rect 80663 2225 80729 2248
rect 80343 2206 80729 2225
rect 84343 2311 84729 2330
rect 84343 2288 84409 2311
rect 84495 2288 84577 2311
rect 84663 2288 84729 2311
rect 84343 2248 84352 2288
rect 84392 2248 84409 2288
rect 84495 2248 84516 2288
rect 84556 2248 84577 2288
rect 84663 2248 84680 2288
rect 84720 2248 84729 2288
rect 84343 2225 84409 2248
rect 84495 2225 84577 2248
rect 84663 2225 84729 2248
rect 84343 2206 84729 2225
rect 88343 2311 88729 2330
rect 88343 2288 88409 2311
rect 88495 2288 88577 2311
rect 88663 2288 88729 2311
rect 88343 2248 88352 2288
rect 88392 2248 88409 2288
rect 88495 2248 88516 2288
rect 88556 2248 88577 2288
rect 88663 2248 88680 2288
rect 88720 2248 88729 2288
rect 88343 2225 88409 2248
rect 88495 2225 88577 2248
rect 88663 2225 88729 2248
rect 88343 2206 88729 2225
rect 92343 2311 92729 2330
rect 92343 2288 92409 2311
rect 92495 2288 92577 2311
rect 92663 2288 92729 2311
rect 92343 2248 92352 2288
rect 92392 2248 92409 2288
rect 92495 2248 92516 2288
rect 92556 2248 92577 2288
rect 92663 2248 92680 2288
rect 92720 2248 92729 2288
rect 92343 2225 92409 2248
rect 92495 2225 92577 2248
rect 92663 2225 92729 2248
rect 92343 2206 92729 2225
rect 96343 2311 96729 2330
rect 96343 2288 96409 2311
rect 96495 2288 96577 2311
rect 96663 2288 96729 2311
rect 96343 2248 96352 2288
rect 96392 2248 96409 2288
rect 96495 2248 96516 2288
rect 96556 2248 96577 2288
rect 96663 2248 96680 2288
rect 96720 2248 96729 2288
rect 96343 2225 96409 2248
rect 96495 2225 96577 2248
rect 96663 2225 96729 2248
rect 96343 2206 96729 2225
rect 3103 1555 3489 1574
rect 3103 1532 3169 1555
rect 3255 1532 3337 1555
rect 3423 1532 3489 1555
rect 3103 1492 3112 1532
rect 3152 1492 3169 1532
rect 3255 1492 3276 1532
rect 3316 1492 3337 1532
rect 3423 1492 3440 1532
rect 3480 1492 3489 1532
rect 3103 1469 3169 1492
rect 3255 1469 3337 1492
rect 3423 1469 3489 1492
rect 3103 1450 3489 1469
rect 7103 1555 7489 1574
rect 7103 1532 7169 1555
rect 7255 1532 7337 1555
rect 7423 1532 7489 1555
rect 7103 1492 7112 1532
rect 7152 1492 7169 1532
rect 7255 1492 7276 1532
rect 7316 1492 7337 1532
rect 7423 1492 7440 1532
rect 7480 1492 7489 1532
rect 7103 1469 7169 1492
rect 7255 1469 7337 1492
rect 7423 1469 7489 1492
rect 7103 1450 7489 1469
rect 11103 1555 11489 1574
rect 11103 1532 11169 1555
rect 11255 1532 11337 1555
rect 11423 1532 11489 1555
rect 11103 1492 11112 1532
rect 11152 1492 11169 1532
rect 11255 1492 11276 1532
rect 11316 1492 11337 1532
rect 11423 1492 11440 1532
rect 11480 1492 11489 1532
rect 11103 1469 11169 1492
rect 11255 1469 11337 1492
rect 11423 1469 11489 1492
rect 11103 1450 11489 1469
rect 15103 1555 15489 1574
rect 15103 1532 15169 1555
rect 15255 1532 15337 1555
rect 15423 1532 15489 1555
rect 15103 1492 15112 1532
rect 15152 1492 15169 1532
rect 15255 1492 15276 1532
rect 15316 1492 15337 1532
rect 15423 1492 15440 1532
rect 15480 1492 15489 1532
rect 15103 1469 15169 1492
rect 15255 1469 15337 1492
rect 15423 1469 15489 1492
rect 15103 1450 15489 1469
rect 19103 1555 19489 1574
rect 19103 1532 19169 1555
rect 19255 1532 19337 1555
rect 19423 1532 19489 1555
rect 19103 1492 19112 1532
rect 19152 1492 19169 1532
rect 19255 1492 19276 1532
rect 19316 1492 19337 1532
rect 19423 1492 19440 1532
rect 19480 1492 19489 1532
rect 19103 1469 19169 1492
rect 19255 1469 19337 1492
rect 19423 1469 19489 1492
rect 19103 1450 19489 1469
rect 23103 1555 23489 1574
rect 23103 1532 23169 1555
rect 23255 1532 23337 1555
rect 23423 1532 23489 1555
rect 23103 1492 23112 1532
rect 23152 1492 23169 1532
rect 23255 1492 23276 1532
rect 23316 1492 23337 1532
rect 23423 1492 23440 1532
rect 23480 1492 23489 1532
rect 23103 1469 23169 1492
rect 23255 1469 23337 1492
rect 23423 1469 23489 1492
rect 23103 1450 23489 1469
rect 27103 1555 27489 1574
rect 27103 1532 27169 1555
rect 27255 1532 27337 1555
rect 27423 1532 27489 1555
rect 27103 1492 27112 1532
rect 27152 1492 27169 1532
rect 27255 1492 27276 1532
rect 27316 1492 27337 1532
rect 27423 1492 27440 1532
rect 27480 1492 27489 1532
rect 27103 1469 27169 1492
rect 27255 1469 27337 1492
rect 27423 1469 27489 1492
rect 27103 1450 27489 1469
rect 31103 1555 31489 1574
rect 31103 1532 31169 1555
rect 31255 1532 31337 1555
rect 31423 1532 31489 1555
rect 31103 1492 31112 1532
rect 31152 1492 31169 1532
rect 31255 1492 31276 1532
rect 31316 1492 31337 1532
rect 31423 1492 31440 1532
rect 31480 1492 31489 1532
rect 31103 1469 31169 1492
rect 31255 1469 31337 1492
rect 31423 1469 31489 1492
rect 31103 1450 31489 1469
rect 35103 1555 35489 1574
rect 35103 1532 35169 1555
rect 35255 1532 35337 1555
rect 35423 1532 35489 1555
rect 35103 1492 35112 1532
rect 35152 1492 35169 1532
rect 35255 1492 35276 1532
rect 35316 1492 35337 1532
rect 35423 1492 35440 1532
rect 35480 1492 35489 1532
rect 35103 1469 35169 1492
rect 35255 1469 35337 1492
rect 35423 1469 35489 1492
rect 35103 1450 35489 1469
rect 39103 1555 39489 1574
rect 39103 1532 39169 1555
rect 39255 1532 39337 1555
rect 39423 1532 39489 1555
rect 39103 1492 39112 1532
rect 39152 1492 39169 1532
rect 39255 1492 39276 1532
rect 39316 1492 39337 1532
rect 39423 1492 39440 1532
rect 39480 1492 39489 1532
rect 39103 1469 39169 1492
rect 39255 1469 39337 1492
rect 39423 1469 39489 1492
rect 39103 1450 39489 1469
rect 43103 1555 43489 1574
rect 43103 1532 43169 1555
rect 43255 1532 43337 1555
rect 43423 1532 43489 1555
rect 43103 1492 43112 1532
rect 43152 1492 43169 1532
rect 43255 1492 43276 1532
rect 43316 1492 43337 1532
rect 43423 1492 43440 1532
rect 43480 1492 43489 1532
rect 43103 1469 43169 1492
rect 43255 1469 43337 1492
rect 43423 1469 43489 1492
rect 43103 1450 43489 1469
rect 47103 1555 47489 1574
rect 47103 1532 47169 1555
rect 47255 1532 47337 1555
rect 47423 1532 47489 1555
rect 47103 1492 47112 1532
rect 47152 1492 47169 1532
rect 47255 1492 47276 1532
rect 47316 1492 47337 1532
rect 47423 1492 47440 1532
rect 47480 1492 47489 1532
rect 47103 1469 47169 1492
rect 47255 1469 47337 1492
rect 47423 1469 47489 1492
rect 47103 1450 47489 1469
rect 51103 1555 51489 1574
rect 51103 1532 51169 1555
rect 51255 1532 51337 1555
rect 51423 1532 51489 1555
rect 51103 1492 51112 1532
rect 51152 1492 51169 1532
rect 51255 1492 51276 1532
rect 51316 1492 51337 1532
rect 51423 1492 51440 1532
rect 51480 1492 51489 1532
rect 51103 1469 51169 1492
rect 51255 1469 51337 1492
rect 51423 1469 51489 1492
rect 51103 1450 51489 1469
rect 55103 1555 55489 1574
rect 55103 1532 55169 1555
rect 55255 1532 55337 1555
rect 55423 1532 55489 1555
rect 55103 1492 55112 1532
rect 55152 1492 55169 1532
rect 55255 1492 55276 1532
rect 55316 1492 55337 1532
rect 55423 1492 55440 1532
rect 55480 1492 55489 1532
rect 55103 1469 55169 1492
rect 55255 1469 55337 1492
rect 55423 1469 55489 1492
rect 55103 1450 55489 1469
rect 59103 1555 59489 1574
rect 59103 1532 59169 1555
rect 59255 1532 59337 1555
rect 59423 1532 59489 1555
rect 59103 1492 59112 1532
rect 59152 1492 59169 1532
rect 59255 1492 59276 1532
rect 59316 1492 59337 1532
rect 59423 1492 59440 1532
rect 59480 1492 59489 1532
rect 59103 1469 59169 1492
rect 59255 1469 59337 1492
rect 59423 1469 59489 1492
rect 59103 1450 59489 1469
rect 63103 1555 63489 1574
rect 63103 1532 63169 1555
rect 63255 1532 63337 1555
rect 63423 1532 63489 1555
rect 63103 1492 63112 1532
rect 63152 1492 63169 1532
rect 63255 1492 63276 1532
rect 63316 1492 63337 1532
rect 63423 1492 63440 1532
rect 63480 1492 63489 1532
rect 63103 1469 63169 1492
rect 63255 1469 63337 1492
rect 63423 1469 63489 1492
rect 63103 1450 63489 1469
rect 67103 1555 67489 1574
rect 67103 1532 67169 1555
rect 67255 1532 67337 1555
rect 67423 1532 67489 1555
rect 67103 1492 67112 1532
rect 67152 1492 67169 1532
rect 67255 1492 67276 1532
rect 67316 1492 67337 1532
rect 67423 1492 67440 1532
rect 67480 1492 67489 1532
rect 67103 1469 67169 1492
rect 67255 1469 67337 1492
rect 67423 1469 67489 1492
rect 67103 1450 67489 1469
rect 71103 1555 71489 1574
rect 71103 1532 71169 1555
rect 71255 1532 71337 1555
rect 71423 1532 71489 1555
rect 71103 1492 71112 1532
rect 71152 1492 71169 1532
rect 71255 1492 71276 1532
rect 71316 1492 71337 1532
rect 71423 1492 71440 1532
rect 71480 1492 71489 1532
rect 71103 1469 71169 1492
rect 71255 1469 71337 1492
rect 71423 1469 71489 1492
rect 71103 1450 71489 1469
rect 75103 1555 75489 1574
rect 75103 1532 75169 1555
rect 75255 1532 75337 1555
rect 75423 1532 75489 1555
rect 75103 1492 75112 1532
rect 75152 1492 75169 1532
rect 75255 1492 75276 1532
rect 75316 1492 75337 1532
rect 75423 1492 75440 1532
rect 75480 1492 75489 1532
rect 75103 1469 75169 1492
rect 75255 1469 75337 1492
rect 75423 1469 75489 1492
rect 75103 1450 75489 1469
rect 79103 1555 79489 1574
rect 79103 1532 79169 1555
rect 79255 1532 79337 1555
rect 79423 1532 79489 1555
rect 79103 1492 79112 1532
rect 79152 1492 79169 1532
rect 79255 1492 79276 1532
rect 79316 1492 79337 1532
rect 79423 1492 79440 1532
rect 79480 1492 79489 1532
rect 79103 1469 79169 1492
rect 79255 1469 79337 1492
rect 79423 1469 79489 1492
rect 79103 1450 79489 1469
rect 83103 1555 83489 1574
rect 83103 1532 83169 1555
rect 83255 1532 83337 1555
rect 83423 1532 83489 1555
rect 83103 1492 83112 1532
rect 83152 1492 83169 1532
rect 83255 1492 83276 1532
rect 83316 1492 83337 1532
rect 83423 1492 83440 1532
rect 83480 1492 83489 1532
rect 83103 1469 83169 1492
rect 83255 1469 83337 1492
rect 83423 1469 83489 1492
rect 83103 1450 83489 1469
rect 87103 1555 87489 1574
rect 87103 1532 87169 1555
rect 87255 1532 87337 1555
rect 87423 1532 87489 1555
rect 87103 1492 87112 1532
rect 87152 1492 87169 1532
rect 87255 1492 87276 1532
rect 87316 1492 87337 1532
rect 87423 1492 87440 1532
rect 87480 1492 87489 1532
rect 87103 1469 87169 1492
rect 87255 1469 87337 1492
rect 87423 1469 87489 1492
rect 87103 1450 87489 1469
rect 91103 1555 91489 1574
rect 91103 1532 91169 1555
rect 91255 1532 91337 1555
rect 91423 1532 91489 1555
rect 91103 1492 91112 1532
rect 91152 1492 91169 1532
rect 91255 1492 91276 1532
rect 91316 1492 91337 1532
rect 91423 1492 91440 1532
rect 91480 1492 91489 1532
rect 91103 1469 91169 1492
rect 91255 1469 91337 1492
rect 91423 1469 91489 1492
rect 91103 1450 91489 1469
rect 95103 1555 95489 1574
rect 95103 1532 95169 1555
rect 95255 1532 95337 1555
rect 95423 1532 95489 1555
rect 95103 1492 95112 1532
rect 95152 1492 95169 1532
rect 95255 1492 95276 1532
rect 95316 1492 95337 1532
rect 95423 1492 95440 1532
rect 95480 1492 95489 1532
rect 95103 1469 95169 1492
rect 95255 1469 95337 1492
rect 95423 1469 95489 1492
rect 95103 1450 95489 1469
rect 99103 1555 99489 1574
rect 99103 1532 99169 1555
rect 99255 1532 99337 1555
rect 99423 1532 99489 1555
rect 99103 1492 99112 1532
rect 99152 1492 99169 1532
rect 99255 1492 99276 1532
rect 99316 1492 99337 1532
rect 99423 1492 99440 1532
rect 99480 1492 99489 1532
rect 99103 1469 99169 1492
rect 99255 1469 99337 1492
rect 99423 1469 99489 1492
rect 99103 1450 99489 1469
rect 4343 799 4729 818
rect 4343 776 4409 799
rect 4495 776 4577 799
rect 4663 776 4729 799
rect 4343 736 4352 776
rect 4392 736 4409 776
rect 4495 736 4516 776
rect 4556 736 4577 776
rect 4663 736 4680 776
rect 4720 736 4729 776
rect 4343 713 4409 736
rect 4495 713 4577 736
rect 4663 713 4729 736
rect 4343 694 4729 713
rect 8343 799 8729 818
rect 8343 776 8409 799
rect 8495 776 8577 799
rect 8663 776 8729 799
rect 8343 736 8352 776
rect 8392 736 8409 776
rect 8495 736 8516 776
rect 8556 736 8577 776
rect 8663 736 8680 776
rect 8720 736 8729 776
rect 8343 713 8409 736
rect 8495 713 8577 736
rect 8663 713 8729 736
rect 8343 694 8729 713
rect 12343 799 12729 818
rect 12343 776 12409 799
rect 12495 776 12577 799
rect 12663 776 12729 799
rect 12343 736 12352 776
rect 12392 736 12409 776
rect 12495 736 12516 776
rect 12556 736 12577 776
rect 12663 736 12680 776
rect 12720 736 12729 776
rect 12343 713 12409 736
rect 12495 713 12577 736
rect 12663 713 12729 736
rect 12343 694 12729 713
rect 16343 799 16729 818
rect 16343 776 16409 799
rect 16495 776 16577 799
rect 16663 776 16729 799
rect 16343 736 16352 776
rect 16392 736 16409 776
rect 16495 736 16516 776
rect 16556 736 16577 776
rect 16663 736 16680 776
rect 16720 736 16729 776
rect 16343 713 16409 736
rect 16495 713 16577 736
rect 16663 713 16729 736
rect 16343 694 16729 713
rect 20343 799 20729 818
rect 20343 776 20409 799
rect 20495 776 20577 799
rect 20663 776 20729 799
rect 20343 736 20352 776
rect 20392 736 20409 776
rect 20495 736 20516 776
rect 20556 736 20577 776
rect 20663 736 20680 776
rect 20720 736 20729 776
rect 20343 713 20409 736
rect 20495 713 20577 736
rect 20663 713 20729 736
rect 20343 694 20729 713
rect 24343 799 24729 818
rect 24343 776 24409 799
rect 24495 776 24577 799
rect 24663 776 24729 799
rect 24343 736 24352 776
rect 24392 736 24409 776
rect 24495 736 24516 776
rect 24556 736 24577 776
rect 24663 736 24680 776
rect 24720 736 24729 776
rect 24343 713 24409 736
rect 24495 713 24577 736
rect 24663 713 24729 736
rect 24343 694 24729 713
rect 28343 799 28729 818
rect 28343 776 28409 799
rect 28495 776 28577 799
rect 28663 776 28729 799
rect 28343 736 28352 776
rect 28392 736 28409 776
rect 28495 736 28516 776
rect 28556 736 28577 776
rect 28663 736 28680 776
rect 28720 736 28729 776
rect 28343 713 28409 736
rect 28495 713 28577 736
rect 28663 713 28729 736
rect 28343 694 28729 713
rect 32343 799 32729 818
rect 32343 776 32409 799
rect 32495 776 32577 799
rect 32663 776 32729 799
rect 32343 736 32352 776
rect 32392 736 32409 776
rect 32495 736 32516 776
rect 32556 736 32577 776
rect 32663 736 32680 776
rect 32720 736 32729 776
rect 32343 713 32409 736
rect 32495 713 32577 736
rect 32663 713 32729 736
rect 32343 694 32729 713
rect 36343 799 36729 818
rect 36343 776 36409 799
rect 36495 776 36577 799
rect 36663 776 36729 799
rect 36343 736 36352 776
rect 36392 736 36409 776
rect 36495 736 36516 776
rect 36556 736 36577 776
rect 36663 736 36680 776
rect 36720 736 36729 776
rect 36343 713 36409 736
rect 36495 713 36577 736
rect 36663 713 36729 736
rect 36343 694 36729 713
rect 40343 799 40729 818
rect 40343 776 40409 799
rect 40495 776 40577 799
rect 40663 776 40729 799
rect 40343 736 40352 776
rect 40392 736 40409 776
rect 40495 736 40516 776
rect 40556 736 40577 776
rect 40663 736 40680 776
rect 40720 736 40729 776
rect 40343 713 40409 736
rect 40495 713 40577 736
rect 40663 713 40729 736
rect 40343 694 40729 713
rect 44343 799 44729 818
rect 44343 776 44409 799
rect 44495 776 44577 799
rect 44663 776 44729 799
rect 44343 736 44352 776
rect 44392 736 44409 776
rect 44495 736 44516 776
rect 44556 736 44577 776
rect 44663 736 44680 776
rect 44720 736 44729 776
rect 44343 713 44409 736
rect 44495 713 44577 736
rect 44663 713 44729 736
rect 44343 694 44729 713
rect 48343 799 48729 818
rect 48343 776 48409 799
rect 48495 776 48577 799
rect 48663 776 48729 799
rect 48343 736 48352 776
rect 48392 736 48409 776
rect 48495 736 48516 776
rect 48556 736 48577 776
rect 48663 736 48680 776
rect 48720 736 48729 776
rect 48343 713 48409 736
rect 48495 713 48577 736
rect 48663 713 48729 736
rect 48343 694 48729 713
rect 52343 799 52729 818
rect 52343 776 52409 799
rect 52495 776 52577 799
rect 52663 776 52729 799
rect 52343 736 52352 776
rect 52392 736 52409 776
rect 52495 736 52516 776
rect 52556 736 52577 776
rect 52663 736 52680 776
rect 52720 736 52729 776
rect 52343 713 52409 736
rect 52495 713 52577 736
rect 52663 713 52729 736
rect 52343 694 52729 713
rect 56343 799 56729 818
rect 56343 776 56409 799
rect 56495 776 56577 799
rect 56663 776 56729 799
rect 56343 736 56352 776
rect 56392 736 56409 776
rect 56495 736 56516 776
rect 56556 736 56577 776
rect 56663 736 56680 776
rect 56720 736 56729 776
rect 56343 713 56409 736
rect 56495 713 56577 736
rect 56663 713 56729 736
rect 56343 694 56729 713
rect 60343 799 60729 818
rect 60343 776 60409 799
rect 60495 776 60577 799
rect 60663 776 60729 799
rect 60343 736 60352 776
rect 60392 736 60409 776
rect 60495 736 60516 776
rect 60556 736 60577 776
rect 60663 736 60680 776
rect 60720 736 60729 776
rect 60343 713 60409 736
rect 60495 713 60577 736
rect 60663 713 60729 736
rect 60343 694 60729 713
rect 64343 799 64729 818
rect 64343 776 64409 799
rect 64495 776 64577 799
rect 64663 776 64729 799
rect 64343 736 64352 776
rect 64392 736 64409 776
rect 64495 736 64516 776
rect 64556 736 64577 776
rect 64663 736 64680 776
rect 64720 736 64729 776
rect 64343 713 64409 736
rect 64495 713 64577 736
rect 64663 713 64729 736
rect 64343 694 64729 713
rect 68343 799 68729 818
rect 68343 776 68409 799
rect 68495 776 68577 799
rect 68663 776 68729 799
rect 68343 736 68352 776
rect 68392 736 68409 776
rect 68495 736 68516 776
rect 68556 736 68577 776
rect 68663 736 68680 776
rect 68720 736 68729 776
rect 68343 713 68409 736
rect 68495 713 68577 736
rect 68663 713 68729 736
rect 68343 694 68729 713
rect 72343 799 72729 818
rect 72343 776 72409 799
rect 72495 776 72577 799
rect 72663 776 72729 799
rect 72343 736 72352 776
rect 72392 736 72409 776
rect 72495 736 72516 776
rect 72556 736 72577 776
rect 72663 736 72680 776
rect 72720 736 72729 776
rect 72343 713 72409 736
rect 72495 713 72577 736
rect 72663 713 72729 736
rect 72343 694 72729 713
rect 76343 799 76729 818
rect 76343 776 76409 799
rect 76495 776 76577 799
rect 76663 776 76729 799
rect 76343 736 76352 776
rect 76392 736 76409 776
rect 76495 736 76516 776
rect 76556 736 76577 776
rect 76663 736 76680 776
rect 76720 736 76729 776
rect 76343 713 76409 736
rect 76495 713 76577 736
rect 76663 713 76729 736
rect 76343 694 76729 713
rect 80343 799 80729 818
rect 80343 776 80409 799
rect 80495 776 80577 799
rect 80663 776 80729 799
rect 80343 736 80352 776
rect 80392 736 80409 776
rect 80495 736 80516 776
rect 80556 736 80577 776
rect 80663 736 80680 776
rect 80720 736 80729 776
rect 80343 713 80409 736
rect 80495 713 80577 736
rect 80663 713 80729 736
rect 80343 694 80729 713
rect 84343 799 84729 818
rect 84343 776 84409 799
rect 84495 776 84577 799
rect 84663 776 84729 799
rect 84343 736 84352 776
rect 84392 736 84409 776
rect 84495 736 84516 776
rect 84556 736 84577 776
rect 84663 736 84680 776
rect 84720 736 84729 776
rect 84343 713 84409 736
rect 84495 713 84577 736
rect 84663 713 84729 736
rect 84343 694 84729 713
rect 88343 799 88729 818
rect 88343 776 88409 799
rect 88495 776 88577 799
rect 88663 776 88729 799
rect 88343 736 88352 776
rect 88392 736 88409 776
rect 88495 736 88516 776
rect 88556 736 88577 776
rect 88663 736 88680 776
rect 88720 736 88729 776
rect 88343 713 88409 736
rect 88495 713 88577 736
rect 88663 713 88729 736
rect 88343 694 88729 713
rect 92343 799 92729 818
rect 92343 776 92409 799
rect 92495 776 92577 799
rect 92663 776 92729 799
rect 92343 736 92352 776
rect 92392 736 92409 776
rect 92495 736 92516 776
rect 92556 736 92577 776
rect 92663 736 92680 776
rect 92720 736 92729 776
rect 92343 713 92409 736
rect 92495 713 92577 736
rect 92663 713 92729 736
rect 92343 694 92729 713
rect 96343 799 96729 818
rect 96343 776 96409 799
rect 96495 776 96577 799
rect 96663 776 96729 799
rect 96343 736 96352 776
rect 96392 736 96409 776
rect 96495 736 96516 776
rect 96556 736 96577 776
rect 96663 736 96680 776
rect 96720 736 96729 776
rect 96343 713 96409 736
rect 96495 713 96577 736
rect 96663 713 96729 736
rect 96343 694 96729 713
<< via5 >>
rect 4409 38576 4495 38599
rect 4577 38576 4663 38599
rect 4409 38536 4434 38576
rect 4434 38536 4474 38576
rect 4474 38536 4495 38576
rect 4577 38536 4598 38576
rect 4598 38536 4638 38576
rect 4638 38536 4663 38576
rect 4409 38513 4495 38536
rect 4577 38513 4663 38536
rect 8409 38576 8495 38599
rect 8577 38576 8663 38599
rect 8409 38536 8434 38576
rect 8434 38536 8474 38576
rect 8474 38536 8495 38576
rect 8577 38536 8598 38576
rect 8598 38536 8638 38576
rect 8638 38536 8663 38576
rect 8409 38513 8495 38536
rect 8577 38513 8663 38536
rect 12409 38576 12495 38599
rect 12577 38576 12663 38599
rect 12409 38536 12434 38576
rect 12434 38536 12474 38576
rect 12474 38536 12495 38576
rect 12577 38536 12598 38576
rect 12598 38536 12638 38576
rect 12638 38536 12663 38576
rect 12409 38513 12495 38536
rect 12577 38513 12663 38536
rect 16409 38576 16495 38599
rect 16577 38576 16663 38599
rect 16409 38536 16434 38576
rect 16434 38536 16474 38576
rect 16474 38536 16495 38576
rect 16577 38536 16598 38576
rect 16598 38536 16638 38576
rect 16638 38536 16663 38576
rect 16409 38513 16495 38536
rect 16577 38513 16663 38536
rect 20409 38576 20495 38599
rect 20577 38576 20663 38599
rect 20409 38536 20434 38576
rect 20434 38536 20474 38576
rect 20474 38536 20495 38576
rect 20577 38536 20598 38576
rect 20598 38536 20638 38576
rect 20638 38536 20663 38576
rect 20409 38513 20495 38536
rect 20577 38513 20663 38536
rect 24409 38576 24495 38599
rect 24577 38576 24663 38599
rect 24409 38536 24434 38576
rect 24434 38536 24474 38576
rect 24474 38536 24495 38576
rect 24577 38536 24598 38576
rect 24598 38536 24638 38576
rect 24638 38536 24663 38576
rect 24409 38513 24495 38536
rect 24577 38513 24663 38536
rect 28409 38576 28495 38599
rect 28577 38576 28663 38599
rect 28409 38536 28434 38576
rect 28434 38536 28474 38576
rect 28474 38536 28495 38576
rect 28577 38536 28598 38576
rect 28598 38536 28638 38576
rect 28638 38536 28663 38576
rect 28409 38513 28495 38536
rect 28577 38513 28663 38536
rect 32409 38576 32495 38599
rect 32577 38576 32663 38599
rect 32409 38536 32434 38576
rect 32434 38536 32474 38576
rect 32474 38536 32495 38576
rect 32577 38536 32598 38576
rect 32598 38536 32638 38576
rect 32638 38536 32663 38576
rect 32409 38513 32495 38536
rect 32577 38513 32663 38536
rect 36409 38576 36495 38599
rect 36577 38576 36663 38599
rect 36409 38536 36434 38576
rect 36434 38536 36474 38576
rect 36474 38536 36495 38576
rect 36577 38536 36598 38576
rect 36598 38536 36638 38576
rect 36638 38536 36663 38576
rect 36409 38513 36495 38536
rect 36577 38513 36663 38536
rect 40409 38576 40495 38599
rect 40577 38576 40663 38599
rect 40409 38536 40434 38576
rect 40434 38536 40474 38576
rect 40474 38536 40495 38576
rect 40577 38536 40598 38576
rect 40598 38536 40638 38576
rect 40638 38536 40663 38576
rect 40409 38513 40495 38536
rect 40577 38513 40663 38536
rect 44409 38576 44495 38599
rect 44577 38576 44663 38599
rect 44409 38536 44434 38576
rect 44434 38536 44474 38576
rect 44474 38536 44495 38576
rect 44577 38536 44598 38576
rect 44598 38536 44638 38576
rect 44638 38536 44663 38576
rect 44409 38513 44495 38536
rect 44577 38513 44663 38536
rect 48409 38576 48495 38599
rect 48577 38576 48663 38599
rect 48409 38536 48434 38576
rect 48434 38536 48474 38576
rect 48474 38536 48495 38576
rect 48577 38536 48598 38576
rect 48598 38536 48638 38576
rect 48638 38536 48663 38576
rect 48409 38513 48495 38536
rect 48577 38513 48663 38536
rect 52409 38576 52495 38599
rect 52577 38576 52663 38599
rect 52409 38536 52434 38576
rect 52434 38536 52474 38576
rect 52474 38536 52495 38576
rect 52577 38536 52598 38576
rect 52598 38536 52638 38576
rect 52638 38536 52663 38576
rect 52409 38513 52495 38536
rect 52577 38513 52663 38536
rect 56409 38576 56495 38599
rect 56577 38576 56663 38599
rect 56409 38536 56434 38576
rect 56434 38536 56474 38576
rect 56474 38536 56495 38576
rect 56577 38536 56598 38576
rect 56598 38536 56638 38576
rect 56638 38536 56663 38576
rect 56409 38513 56495 38536
rect 56577 38513 56663 38536
rect 60409 38576 60495 38599
rect 60577 38576 60663 38599
rect 60409 38536 60434 38576
rect 60434 38536 60474 38576
rect 60474 38536 60495 38576
rect 60577 38536 60598 38576
rect 60598 38536 60638 38576
rect 60638 38536 60663 38576
rect 60409 38513 60495 38536
rect 60577 38513 60663 38536
rect 64409 38576 64495 38599
rect 64577 38576 64663 38599
rect 64409 38536 64434 38576
rect 64434 38536 64474 38576
rect 64474 38536 64495 38576
rect 64577 38536 64598 38576
rect 64598 38536 64638 38576
rect 64638 38536 64663 38576
rect 64409 38513 64495 38536
rect 64577 38513 64663 38536
rect 68409 38576 68495 38599
rect 68577 38576 68663 38599
rect 68409 38536 68434 38576
rect 68434 38536 68474 38576
rect 68474 38536 68495 38576
rect 68577 38536 68598 38576
rect 68598 38536 68638 38576
rect 68638 38536 68663 38576
rect 68409 38513 68495 38536
rect 68577 38513 68663 38536
rect 72409 38576 72495 38599
rect 72577 38576 72663 38599
rect 72409 38536 72434 38576
rect 72434 38536 72474 38576
rect 72474 38536 72495 38576
rect 72577 38536 72598 38576
rect 72598 38536 72638 38576
rect 72638 38536 72663 38576
rect 72409 38513 72495 38536
rect 72577 38513 72663 38536
rect 76409 38576 76495 38599
rect 76577 38576 76663 38599
rect 76409 38536 76434 38576
rect 76434 38536 76474 38576
rect 76474 38536 76495 38576
rect 76577 38536 76598 38576
rect 76598 38536 76638 38576
rect 76638 38536 76663 38576
rect 76409 38513 76495 38536
rect 76577 38513 76663 38536
rect 80409 38576 80495 38599
rect 80577 38576 80663 38599
rect 80409 38536 80434 38576
rect 80434 38536 80474 38576
rect 80474 38536 80495 38576
rect 80577 38536 80598 38576
rect 80598 38536 80638 38576
rect 80638 38536 80663 38576
rect 80409 38513 80495 38536
rect 80577 38513 80663 38536
rect 84409 38576 84495 38599
rect 84577 38576 84663 38599
rect 84409 38536 84434 38576
rect 84434 38536 84474 38576
rect 84474 38536 84495 38576
rect 84577 38536 84598 38576
rect 84598 38536 84638 38576
rect 84638 38536 84663 38576
rect 84409 38513 84495 38536
rect 84577 38513 84663 38536
rect 88409 38576 88495 38599
rect 88577 38576 88663 38599
rect 88409 38536 88434 38576
rect 88434 38536 88474 38576
rect 88474 38536 88495 38576
rect 88577 38536 88598 38576
rect 88598 38536 88638 38576
rect 88638 38536 88663 38576
rect 88409 38513 88495 38536
rect 88577 38513 88663 38536
rect 92409 38576 92495 38599
rect 92577 38576 92663 38599
rect 92409 38536 92434 38576
rect 92434 38536 92474 38576
rect 92474 38536 92495 38576
rect 92577 38536 92598 38576
rect 92598 38536 92638 38576
rect 92638 38536 92663 38576
rect 92409 38513 92495 38536
rect 92577 38513 92663 38536
rect 96409 38576 96495 38599
rect 96577 38576 96663 38599
rect 96409 38536 96434 38576
rect 96434 38536 96474 38576
rect 96474 38536 96495 38576
rect 96577 38536 96598 38576
rect 96598 38536 96638 38576
rect 96638 38536 96663 38576
rect 96409 38513 96495 38536
rect 96577 38513 96663 38536
rect 3169 37820 3255 37843
rect 3337 37820 3423 37843
rect 3169 37780 3194 37820
rect 3194 37780 3234 37820
rect 3234 37780 3255 37820
rect 3337 37780 3358 37820
rect 3358 37780 3398 37820
rect 3398 37780 3423 37820
rect 3169 37757 3255 37780
rect 3337 37757 3423 37780
rect 7169 37820 7255 37843
rect 7337 37820 7423 37843
rect 7169 37780 7194 37820
rect 7194 37780 7234 37820
rect 7234 37780 7255 37820
rect 7337 37780 7358 37820
rect 7358 37780 7398 37820
rect 7398 37780 7423 37820
rect 7169 37757 7255 37780
rect 7337 37757 7423 37780
rect 11169 37820 11255 37843
rect 11337 37820 11423 37843
rect 11169 37780 11194 37820
rect 11194 37780 11234 37820
rect 11234 37780 11255 37820
rect 11337 37780 11358 37820
rect 11358 37780 11398 37820
rect 11398 37780 11423 37820
rect 11169 37757 11255 37780
rect 11337 37757 11423 37780
rect 15169 37820 15255 37843
rect 15337 37820 15423 37843
rect 15169 37780 15194 37820
rect 15194 37780 15234 37820
rect 15234 37780 15255 37820
rect 15337 37780 15358 37820
rect 15358 37780 15398 37820
rect 15398 37780 15423 37820
rect 15169 37757 15255 37780
rect 15337 37757 15423 37780
rect 19169 37820 19255 37843
rect 19337 37820 19423 37843
rect 19169 37780 19194 37820
rect 19194 37780 19234 37820
rect 19234 37780 19255 37820
rect 19337 37780 19358 37820
rect 19358 37780 19398 37820
rect 19398 37780 19423 37820
rect 19169 37757 19255 37780
rect 19337 37757 19423 37780
rect 23169 37820 23255 37843
rect 23337 37820 23423 37843
rect 23169 37780 23194 37820
rect 23194 37780 23234 37820
rect 23234 37780 23255 37820
rect 23337 37780 23358 37820
rect 23358 37780 23398 37820
rect 23398 37780 23423 37820
rect 23169 37757 23255 37780
rect 23337 37757 23423 37780
rect 27169 37820 27255 37843
rect 27337 37820 27423 37843
rect 27169 37780 27194 37820
rect 27194 37780 27234 37820
rect 27234 37780 27255 37820
rect 27337 37780 27358 37820
rect 27358 37780 27398 37820
rect 27398 37780 27423 37820
rect 27169 37757 27255 37780
rect 27337 37757 27423 37780
rect 31169 37820 31255 37843
rect 31337 37820 31423 37843
rect 31169 37780 31194 37820
rect 31194 37780 31234 37820
rect 31234 37780 31255 37820
rect 31337 37780 31358 37820
rect 31358 37780 31398 37820
rect 31398 37780 31423 37820
rect 31169 37757 31255 37780
rect 31337 37757 31423 37780
rect 35169 37820 35255 37843
rect 35337 37820 35423 37843
rect 35169 37780 35194 37820
rect 35194 37780 35234 37820
rect 35234 37780 35255 37820
rect 35337 37780 35358 37820
rect 35358 37780 35398 37820
rect 35398 37780 35423 37820
rect 35169 37757 35255 37780
rect 35337 37757 35423 37780
rect 39169 37820 39255 37843
rect 39337 37820 39423 37843
rect 39169 37780 39194 37820
rect 39194 37780 39234 37820
rect 39234 37780 39255 37820
rect 39337 37780 39358 37820
rect 39358 37780 39398 37820
rect 39398 37780 39423 37820
rect 39169 37757 39255 37780
rect 39337 37757 39423 37780
rect 43169 37820 43255 37843
rect 43337 37820 43423 37843
rect 43169 37780 43194 37820
rect 43194 37780 43234 37820
rect 43234 37780 43255 37820
rect 43337 37780 43358 37820
rect 43358 37780 43398 37820
rect 43398 37780 43423 37820
rect 43169 37757 43255 37780
rect 43337 37757 43423 37780
rect 47169 37820 47255 37843
rect 47337 37820 47423 37843
rect 47169 37780 47194 37820
rect 47194 37780 47234 37820
rect 47234 37780 47255 37820
rect 47337 37780 47358 37820
rect 47358 37780 47398 37820
rect 47398 37780 47423 37820
rect 47169 37757 47255 37780
rect 47337 37757 47423 37780
rect 51169 37820 51255 37843
rect 51337 37820 51423 37843
rect 51169 37780 51194 37820
rect 51194 37780 51234 37820
rect 51234 37780 51255 37820
rect 51337 37780 51358 37820
rect 51358 37780 51398 37820
rect 51398 37780 51423 37820
rect 51169 37757 51255 37780
rect 51337 37757 51423 37780
rect 55169 37820 55255 37843
rect 55337 37820 55423 37843
rect 55169 37780 55194 37820
rect 55194 37780 55234 37820
rect 55234 37780 55255 37820
rect 55337 37780 55358 37820
rect 55358 37780 55398 37820
rect 55398 37780 55423 37820
rect 55169 37757 55255 37780
rect 55337 37757 55423 37780
rect 59169 37820 59255 37843
rect 59337 37820 59423 37843
rect 59169 37780 59194 37820
rect 59194 37780 59234 37820
rect 59234 37780 59255 37820
rect 59337 37780 59358 37820
rect 59358 37780 59398 37820
rect 59398 37780 59423 37820
rect 59169 37757 59255 37780
rect 59337 37757 59423 37780
rect 63169 37820 63255 37843
rect 63337 37820 63423 37843
rect 63169 37780 63194 37820
rect 63194 37780 63234 37820
rect 63234 37780 63255 37820
rect 63337 37780 63358 37820
rect 63358 37780 63398 37820
rect 63398 37780 63423 37820
rect 63169 37757 63255 37780
rect 63337 37757 63423 37780
rect 67169 37820 67255 37843
rect 67337 37820 67423 37843
rect 67169 37780 67194 37820
rect 67194 37780 67234 37820
rect 67234 37780 67255 37820
rect 67337 37780 67358 37820
rect 67358 37780 67398 37820
rect 67398 37780 67423 37820
rect 67169 37757 67255 37780
rect 67337 37757 67423 37780
rect 71169 37820 71255 37843
rect 71337 37820 71423 37843
rect 71169 37780 71194 37820
rect 71194 37780 71234 37820
rect 71234 37780 71255 37820
rect 71337 37780 71358 37820
rect 71358 37780 71398 37820
rect 71398 37780 71423 37820
rect 71169 37757 71255 37780
rect 71337 37757 71423 37780
rect 75169 37820 75255 37843
rect 75337 37820 75423 37843
rect 75169 37780 75194 37820
rect 75194 37780 75234 37820
rect 75234 37780 75255 37820
rect 75337 37780 75358 37820
rect 75358 37780 75398 37820
rect 75398 37780 75423 37820
rect 75169 37757 75255 37780
rect 75337 37757 75423 37780
rect 79169 37820 79255 37843
rect 79337 37820 79423 37843
rect 79169 37780 79194 37820
rect 79194 37780 79234 37820
rect 79234 37780 79255 37820
rect 79337 37780 79358 37820
rect 79358 37780 79398 37820
rect 79398 37780 79423 37820
rect 79169 37757 79255 37780
rect 79337 37757 79423 37780
rect 83169 37820 83255 37843
rect 83337 37820 83423 37843
rect 83169 37780 83194 37820
rect 83194 37780 83234 37820
rect 83234 37780 83255 37820
rect 83337 37780 83358 37820
rect 83358 37780 83398 37820
rect 83398 37780 83423 37820
rect 83169 37757 83255 37780
rect 83337 37757 83423 37780
rect 87169 37820 87255 37843
rect 87337 37820 87423 37843
rect 87169 37780 87194 37820
rect 87194 37780 87234 37820
rect 87234 37780 87255 37820
rect 87337 37780 87358 37820
rect 87358 37780 87398 37820
rect 87398 37780 87423 37820
rect 87169 37757 87255 37780
rect 87337 37757 87423 37780
rect 91169 37820 91255 37843
rect 91337 37820 91423 37843
rect 91169 37780 91194 37820
rect 91194 37780 91234 37820
rect 91234 37780 91255 37820
rect 91337 37780 91358 37820
rect 91358 37780 91398 37820
rect 91398 37780 91423 37820
rect 91169 37757 91255 37780
rect 91337 37757 91423 37780
rect 95169 37820 95255 37843
rect 95337 37820 95423 37843
rect 95169 37780 95194 37820
rect 95194 37780 95234 37820
rect 95234 37780 95255 37820
rect 95337 37780 95358 37820
rect 95358 37780 95398 37820
rect 95398 37780 95423 37820
rect 95169 37757 95255 37780
rect 95337 37757 95423 37780
rect 99169 37820 99255 37843
rect 99337 37820 99423 37843
rect 99169 37780 99194 37820
rect 99194 37780 99234 37820
rect 99234 37780 99255 37820
rect 99337 37780 99358 37820
rect 99358 37780 99398 37820
rect 99398 37780 99423 37820
rect 99169 37757 99255 37780
rect 99337 37757 99423 37780
rect 4409 37064 4495 37087
rect 4577 37064 4663 37087
rect 4409 37024 4434 37064
rect 4434 37024 4474 37064
rect 4474 37024 4495 37064
rect 4577 37024 4598 37064
rect 4598 37024 4638 37064
rect 4638 37024 4663 37064
rect 4409 37001 4495 37024
rect 4577 37001 4663 37024
rect 8409 37064 8495 37087
rect 8577 37064 8663 37087
rect 8409 37024 8434 37064
rect 8434 37024 8474 37064
rect 8474 37024 8495 37064
rect 8577 37024 8598 37064
rect 8598 37024 8638 37064
rect 8638 37024 8663 37064
rect 8409 37001 8495 37024
rect 8577 37001 8663 37024
rect 12409 37064 12495 37087
rect 12577 37064 12663 37087
rect 12409 37024 12434 37064
rect 12434 37024 12474 37064
rect 12474 37024 12495 37064
rect 12577 37024 12598 37064
rect 12598 37024 12638 37064
rect 12638 37024 12663 37064
rect 12409 37001 12495 37024
rect 12577 37001 12663 37024
rect 16409 37064 16495 37087
rect 16577 37064 16663 37087
rect 16409 37024 16434 37064
rect 16434 37024 16474 37064
rect 16474 37024 16495 37064
rect 16577 37024 16598 37064
rect 16598 37024 16638 37064
rect 16638 37024 16663 37064
rect 16409 37001 16495 37024
rect 16577 37001 16663 37024
rect 20409 37064 20495 37087
rect 20577 37064 20663 37087
rect 20409 37024 20434 37064
rect 20434 37024 20474 37064
rect 20474 37024 20495 37064
rect 20577 37024 20598 37064
rect 20598 37024 20638 37064
rect 20638 37024 20663 37064
rect 20409 37001 20495 37024
rect 20577 37001 20663 37024
rect 24409 37064 24495 37087
rect 24577 37064 24663 37087
rect 24409 37024 24434 37064
rect 24434 37024 24474 37064
rect 24474 37024 24495 37064
rect 24577 37024 24598 37064
rect 24598 37024 24638 37064
rect 24638 37024 24663 37064
rect 24409 37001 24495 37024
rect 24577 37001 24663 37024
rect 28409 37064 28495 37087
rect 28577 37064 28663 37087
rect 28409 37024 28434 37064
rect 28434 37024 28474 37064
rect 28474 37024 28495 37064
rect 28577 37024 28598 37064
rect 28598 37024 28638 37064
rect 28638 37024 28663 37064
rect 28409 37001 28495 37024
rect 28577 37001 28663 37024
rect 32409 37064 32495 37087
rect 32577 37064 32663 37087
rect 32409 37024 32434 37064
rect 32434 37024 32474 37064
rect 32474 37024 32495 37064
rect 32577 37024 32598 37064
rect 32598 37024 32638 37064
rect 32638 37024 32663 37064
rect 32409 37001 32495 37024
rect 32577 37001 32663 37024
rect 36409 37064 36495 37087
rect 36577 37064 36663 37087
rect 36409 37024 36434 37064
rect 36434 37024 36474 37064
rect 36474 37024 36495 37064
rect 36577 37024 36598 37064
rect 36598 37024 36638 37064
rect 36638 37024 36663 37064
rect 36409 37001 36495 37024
rect 36577 37001 36663 37024
rect 40409 37064 40495 37087
rect 40577 37064 40663 37087
rect 40409 37024 40434 37064
rect 40434 37024 40474 37064
rect 40474 37024 40495 37064
rect 40577 37024 40598 37064
rect 40598 37024 40638 37064
rect 40638 37024 40663 37064
rect 40409 37001 40495 37024
rect 40577 37001 40663 37024
rect 44409 37064 44495 37087
rect 44577 37064 44663 37087
rect 44409 37024 44434 37064
rect 44434 37024 44474 37064
rect 44474 37024 44495 37064
rect 44577 37024 44598 37064
rect 44598 37024 44638 37064
rect 44638 37024 44663 37064
rect 44409 37001 44495 37024
rect 44577 37001 44663 37024
rect 48409 37064 48495 37087
rect 48577 37064 48663 37087
rect 48409 37024 48434 37064
rect 48434 37024 48474 37064
rect 48474 37024 48495 37064
rect 48577 37024 48598 37064
rect 48598 37024 48638 37064
rect 48638 37024 48663 37064
rect 48409 37001 48495 37024
rect 48577 37001 48663 37024
rect 52409 37064 52495 37087
rect 52577 37064 52663 37087
rect 52409 37024 52434 37064
rect 52434 37024 52474 37064
rect 52474 37024 52495 37064
rect 52577 37024 52598 37064
rect 52598 37024 52638 37064
rect 52638 37024 52663 37064
rect 52409 37001 52495 37024
rect 52577 37001 52663 37024
rect 56409 37064 56495 37087
rect 56577 37064 56663 37087
rect 56409 37024 56434 37064
rect 56434 37024 56474 37064
rect 56474 37024 56495 37064
rect 56577 37024 56598 37064
rect 56598 37024 56638 37064
rect 56638 37024 56663 37064
rect 56409 37001 56495 37024
rect 56577 37001 56663 37024
rect 60409 37064 60495 37087
rect 60577 37064 60663 37087
rect 60409 37024 60434 37064
rect 60434 37024 60474 37064
rect 60474 37024 60495 37064
rect 60577 37024 60598 37064
rect 60598 37024 60638 37064
rect 60638 37024 60663 37064
rect 60409 37001 60495 37024
rect 60577 37001 60663 37024
rect 64409 37064 64495 37087
rect 64577 37064 64663 37087
rect 64409 37024 64434 37064
rect 64434 37024 64474 37064
rect 64474 37024 64495 37064
rect 64577 37024 64598 37064
rect 64598 37024 64638 37064
rect 64638 37024 64663 37064
rect 64409 37001 64495 37024
rect 64577 37001 64663 37024
rect 68409 37064 68495 37087
rect 68577 37064 68663 37087
rect 68409 37024 68434 37064
rect 68434 37024 68474 37064
rect 68474 37024 68495 37064
rect 68577 37024 68598 37064
rect 68598 37024 68638 37064
rect 68638 37024 68663 37064
rect 68409 37001 68495 37024
rect 68577 37001 68663 37024
rect 72409 37064 72495 37087
rect 72577 37064 72663 37087
rect 72409 37024 72434 37064
rect 72434 37024 72474 37064
rect 72474 37024 72495 37064
rect 72577 37024 72598 37064
rect 72598 37024 72638 37064
rect 72638 37024 72663 37064
rect 72409 37001 72495 37024
rect 72577 37001 72663 37024
rect 76409 37064 76495 37087
rect 76577 37064 76663 37087
rect 76409 37024 76434 37064
rect 76434 37024 76474 37064
rect 76474 37024 76495 37064
rect 76577 37024 76598 37064
rect 76598 37024 76638 37064
rect 76638 37024 76663 37064
rect 76409 37001 76495 37024
rect 76577 37001 76663 37024
rect 80409 37064 80495 37087
rect 80577 37064 80663 37087
rect 80409 37024 80434 37064
rect 80434 37024 80474 37064
rect 80474 37024 80495 37064
rect 80577 37024 80598 37064
rect 80598 37024 80638 37064
rect 80638 37024 80663 37064
rect 80409 37001 80495 37024
rect 80577 37001 80663 37024
rect 84409 37064 84495 37087
rect 84577 37064 84663 37087
rect 84409 37024 84434 37064
rect 84434 37024 84474 37064
rect 84474 37024 84495 37064
rect 84577 37024 84598 37064
rect 84598 37024 84638 37064
rect 84638 37024 84663 37064
rect 84409 37001 84495 37024
rect 84577 37001 84663 37024
rect 88409 37064 88495 37087
rect 88577 37064 88663 37087
rect 88409 37024 88434 37064
rect 88434 37024 88474 37064
rect 88474 37024 88495 37064
rect 88577 37024 88598 37064
rect 88598 37024 88638 37064
rect 88638 37024 88663 37064
rect 88409 37001 88495 37024
rect 88577 37001 88663 37024
rect 92409 37064 92495 37087
rect 92577 37064 92663 37087
rect 92409 37024 92434 37064
rect 92434 37024 92474 37064
rect 92474 37024 92495 37064
rect 92577 37024 92598 37064
rect 92598 37024 92638 37064
rect 92638 37024 92663 37064
rect 92409 37001 92495 37024
rect 92577 37001 92663 37024
rect 96409 37064 96495 37087
rect 96577 37064 96663 37087
rect 96409 37024 96434 37064
rect 96434 37024 96474 37064
rect 96474 37024 96495 37064
rect 96577 37024 96598 37064
rect 96598 37024 96638 37064
rect 96638 37024 96663 37064
rect 96409 37001 96495 37024
rect 96577 37001 96663 37024
rect 3169 36308 3255 36331
rect 3337 36308 3423 36331
rect 3169 36268 3194 36308
rect 3194 36268 3234 36308
rect 3234 36268 3255 36308
rect 3337 36268 3358 36308
rect 3358 36268 3398 36308
rect 3398 36268 3423 36308
rect 3169 36245 3255 36268
rect 3337 36245 3423 36268
rect 7169 36308 7255 36331
rect 7337 36308 7423 36331
rect 7169 36268 7194 36308
rect 7194 36268 7234 36308
rect 7234 36268 7255 36308
rect 7337 36268 7358 36308
rect 7358 36268 7398 36308
rect 7398 36268 7423 36308
rect 7169 36245 7255 36268
rect 7337 36245 7423 36268
rect 11169 36308 11255 36331
rect 11337 36308 11423 36331
rect 11169 36268 11194 36308
rect 11194 36268 11234 36308
rect 11234 36268 11255 36308
rect 11337 36268 11358 36308
rect 11358 36268 11398 36308
rect 11398 36268 11423 36308
rect 11169 36245 11255 36268
rect 11337 36245 11423 36268
rect 15169 36308 15255 36331
rect 15337 36308 15423 36331
rect 15169 36268 15194 36308
rect 15194 36268 15234 36308
rect 15234 36268 15255 36308
rect 15337 36268 15358 36308
rect 15358 36268 15398 36308
rect 15398 36268 15423 36308
rect 15169 36245 15255 36268
rect 15337 36245 15423 36268
rect 19169 36308 19255 36331
rect 19337 36308 19423 36331
rect 19169 36268 19194 36308
rect 19194 36268 19234 36308
rect 19234 36268 19255 36308
rect 19337 36268 19358 36308
rect 19358 36268 19398 36308
rect 19398 36268 19423 36308
rect 19169 36245 19255 36268
rect 19337 36245 19423 36268
rect 23169 36308 23255 36331
rect 23337 36308 23423 36331
rect 23169 36268 23194 36308
rect 23194 36268 23234 36308
rect 23234 36268 23255 36308
rect 23337 36268 23358 36308
rect 23358 36268 23398 36308
rect 23398 36268 23423 36308
rect 23169 36245 23255 36268
rect 23337 36245 23423 36268
rect 27169 36308 27255 36331
rect 27337 36308 27423 36331
rect 27169 36268 27194 36308
rect 27194 36268 27234 36308
rect 27234 36268 27255 36308
rect 27337 36268 27358 36308
rect 27358 36268 27398 36308
rect 27398 36268 27423 36308
rect 27169 36245 27255 36268
rect 27337 36245 27423 36268
rect 31169 36308 31255 36331
rect 31337 36308 31423 36331
rect 31169 36268 31194 36308
rect 31194 36268 31234 36308
rect 31234 36268 31255 36308
rect 31337 36268 31358 36308
rect 31358 36268 31398 36308
rect 31398 36268 31423 36308
rect 31169 36245 31255 36268
rect 31337 36245 31423 36268
rect 35169 36308 35255 36331
rect 35337 36308 35423 36331
rect 35169 36268 35194 36308
rect 35194 36268 35234 36308
rect 35234 36268 35255 36308
rect 35337 36268 35358 36308
rect 35358 36268 35398 36308
rect 35398 36268 35423 36308
rect 35169 36245 35255 36268
rect 35337 36245 35423 36268
rect 39169 36308 39255 36331
rect 39337 36308 39423 36331
rect 39169 36268 39194 36308
rect 39194 36268 39234 36308
rect 39234 36268 39255 36308
rect 39337 36268 39358 36308
rect 39358 36268 39398 36308
rect 39398 36268 39423 36308
rect 39169 36245 39255 36268
rect 39337 36245 39423 36268
rect 43169 36308 43255 36331
rect 43337 36308 43423 36331
rect 43169 36268 43194 36308
rect 43194 36268 43234 36308
rect 43234 36268 43255 36308
rect 43337 36268 43358 36308
rect 43358 36268 43398 36308
rect 43398 36268 43423 36308
rect 43169 36245 43255 36268
rect 43337 36245 43423 36268
rect 47169 36308 47255 36331
rect 47337 36308 47423 36331
rect 47169 36268 47194 36308
rect 47194 36268 47234 36308
rect 47234 36268 47255 36308
rect 47337 36268 47358 36308
rect 47358 36268 47398 36308
rect 47398 36268 47423 36308
rect 47169 36245 47255 36268
rect 47337 36245 47423 36268
rect 51169 36308 51255 36331
rect 51337 36308 51423 36331
rect 51169 36268 51194 36308
rect 51194 36268 51234 36308
rect 51234 36268 51255 36308
rect 51337 36268 51358 36308
rect 51358 36268 51398 36308
rect 51398 36268 51423 36308
rect 51169 36245 51255 36268
rect 51337 36245 51423 36268
rect 55169 36308 55255 36331
rect 55337 36308 55423 36331
rect 55169 36268 55194 36308
rect 55194 36268 55234 36308
rect 55234 36268 55255 36308
rect 55337 36268 55358 36308
rect 55358 36268 55398 36308
rect 55398 36268 55423 36308
rect 55169 36245 55255 36268
rect 55337 36245 55423 36268
rect 59169 36308 59255 36331
rect 59337 36308 59423 36331
rect 59169 36268 59194 36308
rect 59194 36268 59234 36308
rect 59234 36268 59255 36308
rect 59337 36268 59358 36308
rect 59358 36268 59398 36308
rect 59398 36268 59423 36308
rect 59169 36245 59255 36268
rect 59337 36245 59423 36268
rect 63169 36308 63255 36331
rect 63337 36308 63423 36331
rect 63169 36268 63194 36308
rect 63194 36268 63234 36308
rect 63234 36268 63255 36308
rect 63337 36268 63358 36308
rect 63358 36268 63398 36308
rect 63398 36268 63423 36308
rect 63169 36245 63255 36268
rect 63337 36245 63423 36268
rect 67169 36308 67255 36331
rect 67337 36308 67423 36331
rect 67169 36268 67194 36308
rect 67194 36268 67234 36308
rect 67234 36268 67255 36308
rect 67337 36268 67358 36308
rect 67358 36268 67398 36308
rect 67398 36268 67423 36308
rect 67169 36245 67255 36268
rect 67337 36245 67423 36268
rect 71169 36308 71255 36331
rect 71337 36308 71423 36331
rect 71169 36268 71194 36308
rect 71194 36268 71234 36308
rect 71234 36268 71255 36308
rect 71337 36268 71358 36308
rect 71358 36268 71398 36308
rect 71398 36268 71423 36308
rect 71169 36245 71255 36268
rect 71337 36245 71423 36268
rect 75169 36308 75255 36331
rect 75337 36308 75423 36331
rect 75169 36268 75194 36308
rect 75194 36268 75234 36308
rect 75234 36268 75255 36308
rect 75337 36268 75358 36308
rect 75358 36268 75398 36308
rect 75398 36268 75423 36308
rect 75169 36245 75255 36268
rect 75337 36245 75423 36268
rect 79169 36308 79255 36331
rect 79337 36308 79423 36331
rect 79169 36268 79194 36308
rect 79194 36268 79234 36308
rect 79234 36268 79255 36308
rect 79337 36268 79358 36308
rect 79358 36268 79398 36308
rect 79398 36268 79423 36308
rect 79169 36245 79255 36268
rect 79337 36245 79423 36268
rect 83169 36308 83255 36331
rect 83337 36308 83423 36331
rect 83169 36268 83194 36308
rect 83194 36268 83234 36308
rect 83234 36268 83255 36308
rect 83337 36268 83358 36308
rect 83358 36268 83398 36308
rect 83398 36268 83423 36308
rect 83169 36245 83255 36268
rect 83337 36245 83423 36268
rect 87169 36308 87255 36331
rect 87337 36308 87423 36331
rect 87169 36268 87194 36308
rect 87194 36268 87234 36308
rect 87234 36268 87255 36308
rect 87337 36268 87358 36308
rect 87358 36268 87398 36308
rect 87398 36268 87423 36308
rect 87169 36245 87255 36268
rect 87337 36245 87423 36268
rect 91169 36308 91255 36331
rect 91337 36308 91423 36331
rect 91169 36268 91194 36308
rect 91194 36268 91234 36308
rect 91234 36268 91255 36308
rect 91337 36268 91358 36308
rect 91358 36268 91398 36308
rect 91398 36268 91423 36308
rect 91169 36245 91255 36268
rect 91337 36245 91423 36268
rect 95169 36308 95255 36331
rect 95337 36308 95423 36331
rect 95169 36268 95194 36308
rect 95194 36268 95234 36308
rect 95234 36268 95255 36308
rect 95337 36268 95358 36308
rect 95358 36268 95398 36308
rect 95398 36268 95423 36308
rect 95169 36245 95255 36268
rect 95337 36245 95423 36268
rect 99169 36308 99255 36331
rect 99337 36308 99423 36331
rect 99169 36268 99194 36308
rect 99194 36268 99234 36308
rect 99234 36268 99255 36308
rect 99337 36268 99358 36308
rect 99358 36268 99398 36308
rect 99398 36268 99423 36308
rect 99169 36245 99255 36268
rect 99337 36245 99423 36268
rect 4409 35552 4495 35575
rect 4577 35552 4663 35575
rect 4409 35512 4434 35552
rect 4434 35512 4474 35552
rect 4474 35512 4495 35552
rect 4577 35512 4598 35552
rect 4598 35512 4638 35552
rect 4638 35512 4663 35552
rect 4409 35489 4495 35512
rect 4577 35489 4663 35512
rect 8409 35552 8495 35575
rect 8577 35552 8663 35575
rect 8409 35512 8434 35552
rect 8434 35512 8474 35552
rect 8474 35512 8495 35552
rect 8577 35512 8598 35552
rect 8598 35512 8638 35552
rect 8638 35512 8663 35552
rect 8409 35489 8495 35512
rect 8577 35489 8663 35512
rect 12409 35552 12495 35575
rect 12577 35552 12663 35575
rect 12409 35512 12434 35552
rect 12434 35512 12474 35552
rect 12474 35512 12495 35552
rect 12577 35512 12598 35552
rect 12598 35512 12638 35552
rect 12638 35512 12663 35552
rect 12409 35489 12495 35512
rect 12577 35489 12663 35512
rect 16409 35552 16495 35575
rect 16577 35552 16663 35575
rect 16409 35512 16434 35552
rect 16434 35512 16474 35552
rect 16474 35512 16495 35552
rect 16577 35512 16598 35552
rect 16598 35512 16638 35552
rect 16638 35512 16663 35552
rect 16409 35489 16495 35512
rect 16577 35489 16663 35512
rect 20409 35552 20495 35575
rect 20577 35552 20663 35575
rect 20409 35512 20434 35552
rect 20434 35512 20474 35552
rect 20474 35512 20495 35552
rect 20577 35512 20598 35552
rect 20598 35512 20638 35552
rect 20638 35512 20663 35552
rect 20409 35489 20495 35512
rect 20577 35489 20663 35512
rect 24409 35552 24495 35575
rect 24577 35552 24663 35575
rect 24409 35512 24434 35552
rect 24434 35512 24474 35552
rect 24474 35512 24495 35552
rect 24577 35512 24598 35552
rect 24598 35512 24638 35552
rect 24638 35512 24663 35552
rect 24409 35489 24495 35512
rect 24577 35489 24663 35512
rect 28409 35552 28495 35575
rect 28577 35552 28663 35575
rect 28409 35512 28434 35552
rect 28434 35512 28474 35552
rect 28474 35512 28495 35552
rect 28577 35512 28598 35552
rect 28598 35512 28638 35552
rect 28638 35512 28663 35552
rect 28409 35489 28495 35512
rect 28577 35489 28663 35512
rect 32409 35552 32495 35575
rect 32577 35552 32663 35575
rect 32409 35512 32434 35552
rect 32434 35512 32474 35552
rect 32474 35512 32495 35552
rect 32577 35512 32598 35552
rect 32598 35512 32638 35552
rect 32638 35512 32663 35552
rect 32409 35489 32495 35512
rect 32577 35489 32663 35512
rect 36409 35552 36495 35575
rect 36577 35552 36663 35575
rect 36409 35512 36434 35552
rect 36434 35512 36474 35552
rect 36474 35512 36495 35552
rect 36577 35512 36598 35552
rect 36598 35512 36638 35552
rect 36638 35512 36663 35552
rect 36409 35489 36495 35512
rect 36577 35489 36663 35512
rect 40409 35552 40495 35575
rect 40577 35552 40663 35575
rect 40409 35512 40434 35552
rect 40434 35512 40474 35552
rect 40474 35512 40495 35552
rect 40577 35512 40598 35552
rect 40598 35512 40638 35552
rect 40638 35512 40663 35552
rect 40409 35489 40495 35512
rect 40577 35489 40663 35512
rect 44409 35552 44495 35575
rect 44577 35552 44663 35575
rect 44409 35512 44434 35552
rect 44434 35512 44474 35552
rect 44474 35512 44495 35552
rect 44577 35512 44598 35552
rect 44598 35512 44638 35552
rect 44638 35512 44663 35552
rect 44409 35489 44495 35512
rect 44577 35489 44663 35512
rect 48409 35552 48495 35575
rect 48577 35552 48663 35575
rect 48409 35512 48434 35552
rect 48434 35512 48474 35552
rect 48474 35512 48495 35552
rect 48577 35512 48598 35552
rect 48598 35512 48638 35552
rect 48638 35512 48663 35552
rect 48409 35489 48495 35512
rect 48577 35489 48663 35512
rect 52409 35552 52495 35575
rect 52577 35552 52663 35575
rect 52409 35512 52434 35552
rect 52434 35512 52474 35552
rect 52474 35512 52495 35552
rect 52577 35512 52598 35552
rect 52598 35512 52638 35552
rect 52638 35512 52663 35552
rect 52409 35489 52495 35512
rect 52577 35489 52663 35512
rect 56409 35552 56495 35575
rect 56577 35552 56663 35575
rect 56409 35512 56434 35552
rect 56434 35512 56474 35552
rect 56474 35512 56495 35552
rect 56577 35512 56598 35552
rect 56598 35512 56638 35552
rect 56638 35512 56663 35552
rect 56409 35489 56495 35512
rect 56577 35489 56663 35512
rect 60409 35552 60495 35575
rect 60577 35552 60663 35575
rect 60409 35512 60434 35552
rect 60434 35512 60474 35552
rect 60474 35512 60495 35552
rect 60577 35512 60598 35552
rect 60598 35512 60638 35552
rect 60638 35512 60663 35552
rect 60409 35489 60495 35512
rect 60577 35489 60663 35512
rect 64409 35552 64495 35575
rect 64577 35552 64663 35575
rect 64409 35512 64434 35552
rect 64434 35512 64474 35552
rect 64474 35512 64495 35552
rect 64577 35512 64598 35552
rect 64598 35512 64638 35552
rect 64638 35512 64663 35552
rect 64409 35489 64495 35512
rect 64577 35489 64663 35512
rect 68409 35552 68495 35575
rect 68577 35552 68663 35575
rect 68409 35512 68434 35552
rect 68434 35512 68474 35552
rect 68474 35512 68495 35552
rect 68577 35512 68598 35552
rect 68598 35512 68638 35552
rect 68638 35512 68663 35552
rect 68409 35489 68495 35512
rect 68577 35489 68663 35512
rect 72409 35552 72495 35575
rect 72577 35552 72663 35575
rect 72409 35512 72434 35552
rect 72434 35512 72474 35552
rect 72474 35512 72495 35552
rect 72577 35512 72598 35552
rect 72598 35512 72638 35552
rect 72638 35512 72663 35552
rect 72409 35489 72495 35512
rect 72577 35489 72663 35512
rect 76409 35552 76495 35575
rect 76577 35552 76663 35575
rect 76409 35512 76434 35552
rect 76434 35512 76474 35552
rect 76474 35512 76495 35552
rect 76577 35512 76598 35552
rect 76598 35512 76638 35552
rect 76638 35512 76663 35552
rect 76409 35489 76495 35512
rect 76577 35489 76663 35512
rect 80409 35552 80495 35575
rect 80577 35552 80663 35575
rect 80409 35512 80434 35552
rect 80434 35512 80474 35552
rect 80474 35512 80495 35552
rect 80577 35512 80598 35552
rect 80598 35512 80638 35552
rect 80638 35512 80663 35552
rect 80409 35489 80495 35512
rect 80577 35489 80663 35512
rect 84409 35552 84495 35575
rect 84577 35552 84663 35575
rect 84409 35512 84434 35552
rect 84434 35512 84474 35552
rect 84474 35512 84495 35552
rect 84577 35512 84598 35552
rect 84598 35512 84638 35552
rect 84638 35512 84663 35552
rect 84409 35489 84495 35512
rect 84577 35489 84663 35512
rect 88409 35552 88495 35575
rect 88577 35552 88663 35575
rect 88409 35512 88434 35552
rect 88434 35512 88474 35552
rect 88474 35512 88495 35552
rect 88577 35512 88598 35552
rect 88598 35512 88638 35552
rect 88638 35512 88663 35552
rect 88409 35489 88495 35512
rect 88577 35489 88663 35512
rect 92409 35552 92495 35575
rect 92577 35552 92663 35575
rect 92409 35512 92434 35552
rect 92434 35512 92474 35552
rect 92474 35512 92495 35552
rect 92577 35512 92598 35552
rect 92598 35512 92638 35552
rect 92638 35512 92663 35552
rect 92409 35489 92495 35512
rect 92577 35489 92663 35512
rect 96409 35552 96495 35575
rect 96577 35552 96663 35575
rect 96409 35512 96434 35552
rect 96434 35512 96474 35552
rect 96474 35512 96495 35552
rect 96577 35512 96598 35552
rect 96598 35512 96638 35552
rect 96638 35512 96663 35552
rect 96409 35489 96495 35512
rect 96577 35489 96663 35512
rect 3169 34796 3255 34819
rect 3337 34796 3423 34819
rect 3169 34756 3194 34796
rect 3194 34756 3234 34796
rect 3234 34756 3255 34796
rect 3337 34756 3358 34796
rect 3358 34756 3398 34796
rect 3398 34756 3423 34796
rect 3169 34733 3255 34756
rect 3337 34733 3423 34756
rect 7169 34796 7255 34819
rect 7337 34796 7423 34819
rect 7169 34756 7194 34796
rect 7194 34756 7234 34796
rect 7234 34756 7255 34796
rect 7337 34756 7358 34796
rect 7358 34756 7398 34796
rect 7398 34756 7423 34796
rect 7169 34733 7255 34756
rect 7337 34733 7423 34756
rect 11169 34796 11255 34819
rect 11337 34796 11423 34819
rect 11169 34756 11194 34796
rect 11194 34756 11234 34796
rect 11234 34756 11255 34796
rect 11337 34756 11358 34796
rect 11358 34756 11398 34796
rect 11398 34756 11423 34796
rect 11169 34733 11255 34756
rect 11337 34733 11423 34756
rect 15169 34796 15255 34819
rect 15337 34796 15423 34819
rect 15169 34756 15194 34796
rect 15194 34756 15234 34796
rect 15234 34756 15255 34796
rect 15337 34756 15358 34796
rect 15358 34756 15398 34796
rect 15398 34756 15423 34796
rect 15169 34733 15255 34756
rect 15337 34733 15423 34756
rect 19169 34796 19255 34819
rect 19337 34796 19423 34819
rect 19169 34756 19194 34796
rect 19194 34756 19234 34796
rect 19234 34756 19255 34796
rect 19337 34756 19358 34796
rect 19358 34756 19398 34796
rect 19398 34756 19423 34796
rect 19169 34733 19255 34756
rect 19337 34733 19423 34756
rect 23169 34796 23255 34819
rect 23337 34796 23423 34819
rect 23169 34756 23194 34796
rect 23194 34756 23234 34796
rect 23234 34756 23255 34796
rect 23337 34756 23358 34796
rect 23358 34756 23398 34796
rect 23398 34756 23423 34796
rect 23169 34733 23255 34756
rect 23337 34733 23423 34756
rect 27169 34796 27255 34819
rect 27337 34796 27423 34819
rect 27169 34756 27194 34796
rect 27194 34756 27234 34796
rect 27234 34756 27255 34796
rect 27337 34756 27358 34796
rect 27358 34756 27398 34796
rect 27398 34756 27423 34796
rect 27169 34733 27255 34756
rect 27337 34733 27423 34756
rect 31169 34796 31255 34819
rect 31337 34796 31423 34819
rect 31169 34756 31194 34796
rect 31194 34756 31234 34796
rect 31234 34756 31255 34796
rect 31337 34756 31358 34796
rect 31358 34756 31398 34796
rect 31398 34756 31423 34796
rect 31169 34733 31255 34756
rect 31337 34733 31423 34756
rect 35169 34796 35255 34819
rect 35337 34796 35423 34819
rect 35169 34756 35194 34796
rect 35194 34756 35234 34796
rect 35234 34756 35255 34796
rect 35337 34756 35358 34796
rect 35358 34756 35398 34796
rect 35398 34756 35423 34796
rect 35169 34733 35255 34756
rect 35337 34733 35423 34756
rect 39169 34796 39255 34819
rect 39337 34796 39423 34819
rect 39169 34756 39194 34796
rect 39194 34756 39234 34796
rect 39234 34756 39255 34796
rect 39337 34756 39358 34796
rect 39358 34756 39398 34796
rect 39398 34756 39423 34796
rect 39169 34733 39255 34756
rect 39337 34733 39423 34756
rect 43169 34796 43255 34819
rect 43337 34796 43423 34819
rect 43169 34756 43194 34796
rect 43194 34756 43234 34796
rect 43234 34756 43255 34796
rect 43337 34756 43358 34796
rect 43358 34756 43398 34796
rect 43398 34756 43423 34796
rect 43169 34733 43255 34756
rect 43337 34733 43423 34756
rect 47169 34796 47255 34819
rect 47337 34796 47423 34819
rect 47169 34756 47194 34796
rect 47194 34756 47234 34796
rect 47234 34756 47255 34796
rect 47337 34756 47358 34796
rect 47358 34756 47398 34796
rect 47398 34756 47423 34796
rect 47169 34733 47255 34756
rect 47337 34733 47423 34756
rect 51169 34796 51255 34819
rect 51337 34796 51423 34819
rect 51169 34756 51194 34796
rect 51194 34756 51234 34796
rect 51234 34756 51255 34796
rect 51337 34756 51358 34796
rect 51358 34756 51398 34796
rect 51398 34756 51423 34796
rect 51169 34733 51255 34756
rect 51337 34733 51423 34756
rect 55169 34796 55255 34819
rect 55337 34796 55423 34819
rect 55169 34756 55194 34796
rect 55194 34756 55234 34796
rect 55234 34756 55255 34796
rect 55337 34756 55358 34796
rect 55358 34756 55398 34796
rect 55398 34756 55423 34796
rect 55169 34733 55255 34756
rect 55337 34733 55423 34756
rect 59169 34796 59255 34819
rect 59337 34796 59423 34819
rect 59169 34756 59194 34796
rect 59194 34756 59234 34796
rect 59234 34756 59255 34796
rect 59337 34756 59358 34796
rect 59358 34756 59398 34796
rect 59398 34756 59423 34796
rect 59169 34733 59255 34756
rect 59337 34733 59423 34756
rect 63169 34796 63255 34819
rect 63337 34796 63423 34819
rect 63169 34756 63194 34796
rect 63194 34756 63234 34796
rect 63234 34756 63255 34796
rect 63337 34756 63358 34796
rect 63358 34756 63398 34796
rect 63398 34756 63423 34796
rect 63169 34733 63255 34756
rect 63337 34733 63423 34756
rect 67169 34796 67255 34819
rect 67337 34796 67423 34819
rect 67169 34756 67194 34796
rect 67194 34756 67234 34796
rect 67234 34756 67255 34796
rect 67337 34756 67358 34796
rect 67358 34756 67398 34796
rect 67398 34756 67423 34796
rect 67169 34733 67255 34756
rect 67337 34733 67423 34756
rect 71169 34796 71255 34819
rect 71337 34796 71423 34819
rect 71169 34756 71194 34796
rect 71194 34756 71234 34796
rect 71234 34756 71255 34796
rect 71337 34756 71358 34796
rect 71358 34756 71398 34796
rect 71398 34756 71423 34796
rect 71169 34733 71255 34756
rect 71337 34733 71423 34756
rect 75169 34796 75255 34819
rect 75337 34796 75423 34819
rect 75169 34756 75194 34796
rect 75194 34756 75234 34796
rect 75234 34756 75255 34796
rect 75337 34756 75358 34796
rect 75358 34756 75398 34796
rect 75398 34756 75423 34796
rect 75169 34733 75255 34756
rect 75337 34733 75423 34756
rect 79169 34796 79255 34819
rect 79337 34796 79423 34819
rect 79169 34756 79194 34796
rect 79194 34756 79234 34796
rect 79234 34756 79255 34796
rect 79337 34756 79358 34796
rect 79358 34756 79398 34796
rect 79398 34756 79423 34796
rect 79169 34733 79255 34756
rect 79337 34733 79423 34756
rect 83169 34796 83255 34819
rect 83337 34796 83423 34819
rect 83169 34756 83194 34796
rect 83194 34756 83234 34796
rect 83234 34756 83255 34796
rect 83337 34756 83358 34796
rect 83358 34756 83398 34796
rect 83398 34756 83423 34796
rect 83169 34733 83255 34756
rect 83337 34733 83423 34756
rect 87169 34796 87255 34819
rect 87337 34796 87423 34819
rect 87169 34756 87194 34796
rect 87194 34756 87234 34796
rect 87234 34756 87255 34796
rect 87337 34756 87358 34796
rect 87358 34756 87398 34796
rect 87398 34756 87423 34796
rect 87169 34733 87255 34756
rect 87337 34733 87423 34756
rect 91169 34796 91255 34819
rect 91337 34796 91423 34819
rect 91169 34756 91194 34796
rect 91194 34756 91234 34796
rect 91234 34756 91255 34796
rect 91337 34756 91358 34796
rect 91358 34756 91398 34796
rect 91398 34756 91423 34796
rect 91169 34733 91255 34756
rect 91337 34733 91423 34756
rect 95169 34796 95255 34819
rect 95337 34796 95423 34819
rect 95169 34756 95194 34796
rect 95194 34756 95234 34796
rect 95234 34756 95255 34796
rect 95337 34756 95358 34796
rect 95358 34756 95398 34796
rect 95398 34756 95423 34796
rect 95169 34733 95255 34756
rect 95337 34733 95423 34756
rect 99169 34796 99255 34819
rect 99337 34796 99423 34819
rect 99169 34756 99194 34796
rect 99194 34756 99234 34796
rect 99234 34756 99255 34796
rect 99337 34756 99358 34796
rect 99358 34756 99398 34796
rect 99398 34756 99423 34796
rect 99169 34733 99255 34756
rect 99337 34733 99423 34756
rect 4409 34040 4495 34063
rect 4577 34040 4663 34063
rect 4409 34000 4434 34040
rect 4434 34000 4474 34040
rect 4474 34000 4495 34040
rect 4577 34000 4598 34040
rect 4598 34000 4638 34040
rect 4638 34000 4663 34040
rect 4409 33977 4495 34000
rect 4577 33977 4663 34000
rect 8409 34040 8495 34063
rect 8577 34040 8663 34063
rect 8409 34000 8434 34040
rect 8434 34000 8474 34040
rect 8474 34000 8495 34040
rect 8577 34000 8598 34040
rect 8598 34000 8638 34040
rect 8638 34000 8663 34040
rect 8409 33977 8495 34000
rect 8577 33977 8663 34000
rect 12409 34040 12495 34063
rect 12577 34040 12663 34063
rect 12409 34000 12434 34040
rect 12434 34000 12474 34040
rect 12474 34000 12495 34040
rect 12577 34000 12598 34040
rect 12598 34000 12638 34040
rect 12638 34000 12663 34040
rect 12409 33977 12495 34000
rect 12577 33977 12663 34000
rect 16409 34040 16495 34063
rect 16577 34040 16663 34063
rect 16409 34000 16434 34040
rect 16434 34000 16474 34040
rect 16474 34000 16495 34040
rect 16577 34000 16598 34040
rect 16598 34000 16638 34040
rect 16638 34000 16663 34040
rect 16409 33977 16495 34000
rect 16577 33977 16663 34000
rect 20409 34040 20495 34063
rect 20577 34040 20663 34063
rect 20409 34000 20434 34040
rect 20434 34000 20474 34040
rect 20474 34000 20495 34040
rect 20577 34000 20598 34040
rect 20598 34000 20638 34040
rect 20638 34000 20663 34040
rect 20409 33977 20495 34000
rect 20577 33977 20663 34000
rect 24409 34040 24495 34063
rect 24577 34040 24663 34063
rect 24409 34000 24434 34040
rect 24434 34000 24474 34040
rect 24474 34000 24495 34040
rect 24577 34000 24598 34040
rect 24598 34000 24638 34040
rect 24638 34000 24663 34040
rect 24409 33977 24495 34000
rect 24577 33977 24663 34000
rect 28409 34040 28495 34063
rect 28577 34040 28663 34063
rect 28409 34000 28434 34040
rect 28434 34000 28474 34040
rect 28474 34000 28495 34040
rect 28577 34000 28598 34040
rect 28598 34000 28638 34040
rect 28638 34000 28663 34040
rect 28409 33977 28495 34000
rect 28577 33977 28663 34000
rect 32409 34040 32495 34063
rect 32577 34040 32663 34063
rect 32409 34000 32434 34040
rect 32434 34000 32474 34040
rect 32474 34000 32495 34040
rect 32577 34000 32598 34040
rect 32598 34000 32638 34040
rect 32638 34000 32663 34040
rect 32409 33977 32495 34000
rect 32577 33977 32663 34000
rect 36409 34040 36495 34063
rect 36577 34040 36663 34063
rect 36409 34000 36434 34040
rect 36434 34000 36474 34040
rect 36474 34000 36495 34040
rect 36577 34000 36598 34040
rect 36598 34000 36638 34040
rect 36638 34000 36663 34040
rect 36409 33977 36495 34000
rect 36577 33977 36663 34000
rect 40409 34040 40495 34063
rect 40577 34040 40663 34063
rect 40409 34000 40434 34040
rect 40434 34000 40474 34040
rect 40474 34000 40495 34040
rect 40577 34000 40598 34040
rect 40598 34000 40638 34040
rect 40638 34000 40663 34040
rect 40409 33977 40495 34000
rect 40577 33977 40663 34000
rect 44409 34040 44495 34063
rect 44577 34040 44663 34063
rect 44409 34000 44434 34040
rect 44434 34000 44474 34040
rect 44474 34000 44495 34040
rect 44577 34000 44598 34040
rect 44598 34000 44638 34040
rect 44638 34000 44663 34040
rect 44409 33977 44495 34000
rect 44577 33977 44663 34000
rect 48409 34040 48495 34063
rect 48577 34040 48663 34063
rect 48409 34000 48434 34040
rect 48434 34000 48474 34040
rect 48474 34000 48495 34040
rect 48577 34000 48598 34040
rect 48598 34000 48638 34040
rect 48638 34000 48663 34040
rect 48409 33977 48495 34000
rect 48577 33977 48663 34000
rect 52409 34040 52495 34063
rect 52577 34040 52663 34063
rect 52409 34000 52434 34040
rect 52434 34000 52474 34040
rect 52474 34000 52495 34040
rect 52577 34000 52598 34040
rect 52598 34000 52638 34040
rect 52638 34000 52663 34040
rect 52409 33977 52495 34000
rect 52577 33977 52663 34000
rect 56409 34040 56495 34063
rect 56577 34040 56663 34063
rect 56409 34000 56434 34040
rect 56434 34000 56474 34040
rect 56474 34000 56495 34040
rect 56577 34000 56598 34040
rect 56598 34000 56638 34040
rect 56638 34000 56663 34040
rect 56409 33977 56495 34000
rect 56577 33977 56663 34000
rect 60409 34040 60495 34063
rect 60577 34040 60663 34063
rect 60409 34000 60434 34040
rect 60434 34000 60474 34040
rect 60474 34000 60495 34040
rect 60577 34000 60598 34040
rect 60598 34000 60638 34040
rect 60638 34000 60663 34040
rect 60409 33977 60495 34000
rect 60577 33977 60663 34000
rect 64409 34040 64495 34063
rect 64577 34040 64663 34063
rect 64409 34000 64434 34040
rect 64434 34000 64474 34040
rect 64474 34000 64495 34040
rect 64577 34000 64598 34040
rect 64598 34000 64638 34040
rect 64638 34000 64663 34040
rect 64409 33977 64495 34000
rect 64577 33977 64663 34000
rect 68409 34040 68495 34063
rect 68577 34040 68663 34063
rect 68409 34000 68434 34040
rect 68434 34000 68474 34040
rect 68474 34000 68495 34040
rect 68577 34000 68598 34040
rect 68598 34000 68638 34040
rect 68638 34000 68663 34040
rect 68409 33977 68495 34000
rect 68577 33977 68663 34000
rect 86469 33389 86555 33475
rect 3169 33284 3255 33307
rect 3337 33284 3423 33307
rect 3169 33244 3194 33284
rect 3194 33244 3234 33284
rect 3234 33244 3255 33284
rect 3337 33244 3358 33284
rect 3358 33244 3398 33284
rect 3398 33244 3423 33284
rect 3169 33221 3255 33244
rect 3337 33221 3423 33244
rect 7169 33284 7255 33307
rect 7337 33284 7423 33307
rect 7169 33244 7194 33284
rect 7194 33244 7234 33284
rect 7234 33244 7255 33284
rect 7337 33244 7358 33284
rect 7358 33244 7398 33284
rect 7398 33244 7423 33284
rect 7169 33221 7255 33244
rect 7337 33221 7423 33244
rect 11169 33284 11255 33307
rect 11337 33284 11423 33307
rect 11169 33244 11194 33284
rect 11194 33244 11234 33284
rect 11234 33244 11255 33284
rect 11337 33244 11358 33284
rect 11358 33244 11398 33284
rect 11398 33244 11423 33284
rect 11169 33221 11255 33244
rect 11337 33221 11423 33244
rect 15169 33284 15255 33307
rect 15337 33284 15423 33307
rect 15169 33244 15194 33284
rect 15194 33244 15234 33284
rect 15234 33244 15255 33284
rect 15337 33244 15358 33284
rect 15358 33244 15398 33284
rect 15398 33244 15423 33284
rect 15169 33221 15255 33244
rect 15337 33221 15423 33244
rect 19169 33284 19255 33307
rect 19337 33284 19423 33307
rect 19169 33244 19194 33284
rect 19194 33244 19234 33284
rect 19234 33244 19255 33284
rect 19337 33244 19358 33284
rect 19358 33244 19398 33284
rect 19398 33244 19423 33284
rect 19169 33221 19255 33244
rect 19337 33221 19423 33244
rect 23169 33284 23255 33307
rect 23337 33284 23423 33307
rect 23169 33244 23194 33284
rect 23194 33244 23234 33284
rect 23234 33244 23255 33284
rect 23337 33244 23358 33284
rect 23358 33244 23398 33284
rect 23398 33244 23423 33284
rect 23169 33221 23255 33244
rect 23337 33221 23423 33244
rect 27169 33284 27255 33307
rect 27337 33284 27423 33307
rect 27169 33244 27194 33284
rect 27194 33244 27234 33284
rect 27234 33244 27255 33284
rect 27337 33244 27358 33284
rect 27358 33244 27398 33284
rect 27398 33244 27423 33284
rect 27169 33221 27255 33244
rect 27337 33221 27423 33244
rect 31169 33284 31255 33307
rect 31337 33284 31423 33307
rect 31169 33244 31194 33284
rect 31194 33244 31234 33284
rect 31234 33244 31255 33284
rect 31337 33244 31358 33284
rect 31358 33244 31398 33284
rect 31398 33244 31423 33284
rect 31169 33221 31255 33244
rect 31337 33221 31423 33244
rect 35169 33284 35255 33307
rect 35337 33284 35423 33307
rect 35169 33244 35194 33284
rect 35194 33244 35234 33284
rect 35234 33244 35255 33284
rect 35337 33244 35358 33284
rect 35358 33244 35398 33284
rect 35398 33244 35423 33284
rect 35169 33221 35255 33244
rect 35337 33221 35423 33244
rect 39169 33284 39255 33307
rect 39337 33284 39423 33307
rect 39169 33244 39194 33284
rect 39194 33244 39234 33284
rect 39234 33244 39255 33284
rect 39337 33244 39358 33284
rect 39358 33244 39398 33284
rect 39398 33244 39423 33284
rect 39169 33221 39255 33244
rect 39337 33221 39423 33244
rect 43169 33284 43255 33307
rect 43337 33284 43423 33307
rect 43169 33244 43194 33284
rect 43194 33244 43234 33284
rect 43234 33244 43255 33284
rect 43337 33244 43358 33284
rect 43358 33244 43398 33284
rect 43398 33244 43423 33284
rect 43169 33221 43255 33244
rect 43337 33221 43423 33244
rect 47169 33284 47255 33307
rect 47337 33284 47423 33307
rect 47169 33244 47194 33284
rect 47194 33244 47234 33284
rect 47234 33244 47255 33284
rect 47337 33244 47358 33284
rect 47358 33244 47398 33284
rect 47398 33244 47423 33284
rect 47169 33221 47255 33244
rect 47337 33221 47423 33244
rect 51169 33284 51255 33307
rect 51337 33284 51423 33307
rect 51169 33244 51194 33284
rect 51194 33244 51234 33284
rect 51234 33244 51255 33284
rect 51337 33244 51358 33284
rect 51358 33244 51398 33284
rect 51398 33244 51423 33284
rect 51169 33221 51255 33244
rect 51337 33221 51423 33244
rect 55169 33284 55255 33307
rect 55337 33284 55423 33307
rect 55169 33244 55194 33284
rect 55194 33244 55234 33284
rect 55234 33244 55255 33284
rect 55337 33244 55358 33284
rect 55358 33244 55398 33284
rect 55398 33244 55423 33284
rect 55169 33221 55255 33244
rect 55337 33221 55423 33244
rect 59169 33284 59255 33307
rect 59337 33284 59423 33307
rect 59169 33244 59194 33284
rect 59194 33244 59234 33284
rect 59234 33244 59255 33284
rect 59337 33244 59358 33284
rect 59358 33244 59398 33284
rect 59398 33244 59423 33284
rect 59169 33221 59255 33244
rect 59337 33221 59423 33244
rect 63169 33284 63255 33307
rect 63337 33284 63423 33307
rect 63169 33244 63194 33284
rect 63194 33244 63234 33284
rect 63234 33244 63255 33284
rect 63337 33244 63358 33284
rect 63358 33244 63398 33284
rect 63398 33244 63423 33284
rect 63169 33221 63255 33244
rect 63337 33221 63423 33244
rect 67169 33284 67255 33307
rect 67337 33284 67423 33307
rect 67169 33244 67194 33284
rect 67194 33244 67234 33284
rect 67234 33244 67255 33284
rect 67337 33244 67358 33284
rect 67358 33244 67398 33284
rect 67398 33244 67423 33284
rect 67169 33221 67255 33244
rect 67337 33221 67423 33244
rect 73245 32801 73331 32887
rect 4409 32528 4495 32551
rect 4577 32528 4663 32551
rect 4409 32488 4434 32528
rect 4434 32488 4474 32528
rect 4474 32488 4495 32528
rect 4577 32488 4598 32528
rect 4598 32488 4638 32528
rect 4638 32488 4663 32528
rect 4409 32465 4495 32488
rect 4577 32465 4663 32488
rect 8409 32528 8495 32551
rect 8577 32528 8663 32551
rect 8409 32488 8434 32528
rect 8434 32488 8474 32528
rect 8474 32488 8495 32528
rect 8577 32488 8598 32528
rect 8598 32488 8638 32528
rect 8638 32488 8663 32528
rect 8409 32465 8495 32488
rect 8577 32465 8663 32488
rect 12409 32528 12495 32551
rect 12577 32528 12663 32551
rect 12409 32488 12434 32528
rect 12434 32488 12474 32528
rect 12474 32488 12495 32528
rect 12577 32488 12598 32528
rect 12598 32488 12638 32528
rect 12638 32488 12663 32528
rect 12409 32465 12495 32488
rect 12577 32465 12663 32488
rect 16409 32528 16495 32551
rect 16577 32528 16663 32551
rect 16409 32488 16434 32528
rect 16434 32488 16474 32528
rect 16474 32488 16495 32528
rect 16577 32488 16598 32528
rect 16598 32488 16638 32528
rect 16638 32488 16663 32528
rect 16409 32465 16495 32488
rect 16577 32465 16663 32488
rect 20409 32528 20495 32551
rect 20577 32528 20663 32551
rect 20409 32488 20434 32528
rect 20434 32488 20474 32528
rect 20474 32488 20495 32528
rect 20577 32488 20598 32528
rect 20598 32488 20638 32528
rect 20638 32488 20663 32528
rect 20409 32465 20495 32488
rect 20577 32465 20663 32488
rect 24409 32528 24495 32551
rect 24577 32528 24663 32551
rect 24409 32488 24434 32528
rect 24434 32488 24474 32528
rect 24474 32488 24495 32528
rect 24577 32488 24598 32528
rect 24598 32488 24638 32528
rect 24638 32488 24663 32528
rect 24409 32465 24495 32488
rect 24577 32465 24663 32488
rect 28409 32528 28495 32551
rect 28577 32528 28663 32551
rect 28409 32488 28434 32528
rect 28434 32488 28474 32528
rect 28474 32488 28495 32528
rect 28577 32488 28598 32528
rect 28598 32488 28638 32528
rect 28638 32488 28663 32528
rect 28409 32465 28495 32488
rect 28577 32465 28663 32488
rect 32409 32528 32495 32551
rect 32577 32528 32663 32551
rect 32409 32488 32434 32528
rect 32434 32488 32474 32528
rect 32474 32488 32495 32528
rect 32577 32488 32598 32528
rect 32598 32488 32638 32528
rect 32638 32488 32663 32528
rect 32409 32465 32495 32488
rect 32577 32465 32663 32488
rect 36409 32528 36495 32551
rect 36577 32528 36663 32551
rect 36409 32488 36434 32528
rect 36434 32488 36474 32528
rect 36474 32488 36495 32528
rect 36577 32488 36598 32528
rect 36598 32488 36638 32528
rect 36638 32488 36663 32528
rect 36409 32465 36495 32488
rect 36577 32465 36663 32488
rect 40409 32528 40495 32551
rect 40577 32528 40663 32551
rect 40409 32488 40434 32528
rect 40434 32488 40474 32528
rect 40474 32488 40495 32528
rect 40577 32488 40598 32528
rect 40598 32488 40638 32528
rect 40638 32488 40663 32528
rect 40409 32465 40495 32488
rect 40577 32465 40663 32488
rect 44409 32528 44495 32551
rect 44577 32528 44663 32551
rect 44409 32488 44434 32528
rect 44434 32488 44474 32528
rect 44474 32488 44495 32528
rect 44577 32488 44598 32528
rect 44598 32488 44638 32528
rect 44638 32488 44663 32528
rect 44409 32465 44495 32488
rect 44577 32465 44663 32488
rect 48409 32528 48495 32551
rect 48577 32528 48663 32551
rect 48409 32488 48434 32528
rect 48434 32488 48474 32528
rect 48474 32488 48495 32528
rect 48577 32488 48598 32528
rect 48598 32488 48638 32528
rect 48638 32488 48663 32528
rect 48409 32465 48495 32488
rect 48577 32465 48663 32488
rect 52409 32528 52495 32551
rect 52577 32528 52663 32551
rect 52409 32488 52434 32528
rect 52434 32488 52474 32528
rect 52474 32488 52495 32528
rect 52577 32488 52598 32528
rect 52598 32488 52638 32528
rect 52638 32488 52663 32528
rect 52409 32465 52495 32488
rect 52577 32465 52663 32488
rect 56409 32528 56495 32551
rect 56577 32528 56663 32551
rect 56409 32488 56434 32528
rect 56434 32488 56474 32528
rect 56474 32488 56495 32528
rect 56577 32488 56598 32528
rect 56598 32488 56638 32528
rect 56638 32488 56663 32528
rect 56409 32465 56495 32488
rect 56577 32465 56663 32488
rect 60409 32528 60495 32551
rect 60577 32528 60663 32551
rect 60409 32488 60434 32528
rect 60434 32488 60474 32528
rect 60474 32488 60495 32528
rect 60577 32488 60598 32528
rect 60598 32488 60638 32528
rect 60638 32488 60663 32528
rect 60409 32465 60495 32488
rect 60577 32465 60663 32488
rect 64409 32528 64495 32551
rect 64577 32528 64663 32551
rect 64409 32488 64434 32528
rect 64434 32488 64474 32528
rect 64474 32488 64495 32528
rect 64577 32488 64598 32528
rect 64598 32488 64638 32528
rect 64638 32488 64663 32528
rect 64409 32465 64495 32488
rect 64577 32465 64663 32488
rect 68409 32528 68495 32551
rect 68577 32528 68663 32551
rect 68409 32488 68434 32528
rect 68434 32488 68474 32528
rect 68474 32488 68495 32528
rect 68577 32488 68598 32528
rect 68598 32488 68638 32528
rect 68638 32488 68663 32528
rect 68409 32465 68495 32488
rect 68577 32465 68663 32488
rect 3169 31772 3255 31795
rect 3337 31772 3423 31795
rect 3169 31732 3194 31772
rect 3194 31732 3234 31772
rect 3234 31732 3255 31772
rect 3337 31732 3358 31772
rect 3358 31732 3398 31772
rect 3398 31732 3423 31772
rect 3169 31709 3255 31732
rect 3337 31709 3423 31732
rect 7169 31772 7255 31795
rect 7337 31772 7423 31795
rect 7169 31732 7194 31772
rect 7194 31732 7234 31772
rect 7234 31732 7255 31772
rect 7337 31732 7358 31772
rect 7358 31732 7398 31772
rect 7398 31732 7423 31772
rect 7169 31709 7255 31732
rect 7337 31709 7423 31732
rect 11169 31772 11255 31795
rect 11337 31772 11423 31795
rect 11169 31732 11194 31772
rect 11194 31732 11234 31772
rect 11234 31732 11255 31772
rect 11337 31732 11358 31772
rect 11358 31732 11398 31772
rect 11398 31732 11423 31772
rect 11169 31709 11255 31732
rect 11337 31709 11423 31732
rect 15169 31772 15255 31795
rect 15337 31772 15423 31795
rect 15169 31732 15194 31772
rect 15194 31732 15234 31772
rect 15234 31732 15255 31772
rect 15337 31732 15358 31772
rect 15358 31732 15398 31772
rect 15398 31732 15423 31772
rect 15169 31709 15255 31732
rect 15337 31709 15423 31732
rect 19169 31772 19255 31795
rect 19337 31772 19423 31795
rect 19169 31732 19194 31772
rect 19194 31732 19234 31772
rect 19234 31732 19255 31772
rect 19337 31732 19358 31772
rect 19358 31732 19398 31772
rect 19398 31732 19423 31772
rect 19169 31709 19255 31732
rect 19337 31709 19423 31732
rect 23169 31772 23255 31795
rect 23337 31772 23423 31795
rect 23169 31732 23194 31772
rect 23194 31732 23234 31772
rect 23234 31732 23255 31772
rect 23337 31732 23358 31772
rect 23358 31732 23398 31772
rect 23398 31732 23423 31772
rect 23169 31709 23255 31732
rect 23337 31709 23423 31732
rect 27169 31772 27255 31795
rect 27337 31772 27423 31795
rect 27169 31732 27194 31772
rect 27194 31732 27234 31772
rect 27234 31732 27255 31772
rect 27337 31732 27358 31772
rect 27358 31732 27398 31772
rect 27398 31732 27423 31772
rect 27169 31709 27255 31732
rect 27337 31709 27423 31732
rect 31169 31772 31255 31795
rect 31337 31772 31423 31795
rect 31169 31732 31194 31772
rect 31194 31732 31234 31772
rect 31234 31732 31255 31772
rect 31337 31732 31358 31772
rect 31358 31732 31398 31772
rect 31398 31732 31423 31772
rect 31169 31709 31255 31732
rect 31337 31709 31423 31732
rect 35169 31772 35255 31795
rect 35337 31772 35423 31795
rect 35169 31732 35194 31772
rect 35194 31732 35234 31772
rect 35234 31732 35255 31772
rect 35337 31732 35358 31772
rect 35358 31732 35398 31772
rect 35398 31732 35423 31772
rect 35169 31709 35255 31732
rect 35337 31709 35423 31732
rect 39169 31772 39255 31795
rect 39337 31772 39423 31795
rect 39169 31732 39194 31772
rect 39194 31732 39234 31772
rect 39234 31732 39255 31772
rect 39337 31732 39358 31772
rect 39358 31732 39398 31772
rect 39398 31732 39423 31772
rect 39169 31709 39255 31732
rect 39337 31709 39423 31732
rect 43169 31772 43255 31795
rect 43337 31772 43423 31795
rect 43169 31732 43194 31772
rect 43194 31732 43234 31772
rect 43234 31732 43255 31772
rect 43337 31732 43358 31772
rect 43358 31732 43398 31772
rect 43398 31732 43423 31772
rect 43169 31709 43255 31732
rect 43337 31709 43423 31732
rect 47169 31772 47255 31795
rect 47337 31772 47423 31795
rect 47169 31732 47194 31772
rect 47194 31732 47234 31772
rect 47234 31732 47255 31772
rect 47337 31732 47358 31772
rect 47358 31732 47398 31772
rect 47398 31732 47423 31772
rect 47169 31709 47255 31732
rect 47337 31709 47423 31732
rect 51169 31772 51255 31795
rect 51337 31772 51423 31795
rect 51169 31732 51194 31772
rect 51194 31732 51234 31772
rect 51234 31732 51255 31772
rect 51337 31732 51358 31772
rect 51358 31732 51398 31772
rect 51398 31732 51423 31772
rect 51169 31709 51255 31732
rect 51337 31709 51423 31732
rect 55169 31772 55255 31795
rect 55337 31772 55423 31795
rect 55169 31732 55194 31772
rect 55194 31732 55234 31772
rect 55234 31732 55255 31772
rect 55337 31732 55358 31772
rect 55358 31732 55398 31772
rect 55398 31732 55423 31772
rect 55169 31709 55255 31732
rect 55337 31709 55423 31732
rect 59169 31772 59255 31795
rect 59337 31772 59423 31795
rect 59169 31732 59194 31772
rect 59194 31732 59234 31772
rect 59234 31732 59255 31772
rect 59337 31732 59358 31772
rect 59358 31732 59398 31772
rect 59398 31732 59423 31772
rect 59169 31709 59255 31732
rect 59337 31709 59423 31732
rect 63169 31772 63255 31795
rect 63337 31772 63423 31795
rect 63169 31732 63194 31772
rect 63194 31732 63234 31772
rect 63234 31732 63255 31772
rect 63337 31732 63358 31772
rect 63358 31732 63398 31772
rect 63398 31732 63423 31772
rect 63169 31709 63255 31732
rect 63337 31709 63423 31732
rect 67169 31772 67255 31795
rect 67337 31772 67423 31795
rect 67169 31732 67194 31772
rect 67194 31732 67234 31772
rect 67234 31732 67255 31772
rect 67337 31732 67358 31772
rect 67358 31732 67398 31772
rect 67398 31732 67423 31772
rect 67169 31709 67255 31732
rect 67337 31709 67423 31732
rect 72409 31770 72495 31856
rect 72577 31770 72663 31856
rect 72409 31602 72495 31688
rect 72577 31602 72663 31688
rect 72409 31434 72495 31520
rect 72577 31434 72663 31520
rect 72409 31266 72495 31352
rect 72577 31266 72663 31352
rect 72409 31098 72495 31184
rect 72577 31098 72663 31184
rect 4409 31016 4495 31039
rect 4577 31016 4663 31039
rect 4409 30976 4434 31016
rect 4434 30976 4474 31016
rect 4474 30976 4495 31016
rect 4577 30976 4598 31016
rect 4598 30976 4638 31016
rect 4638 30976 4663 31016
rect 4409 30953 4495 30976
rect 4577 30953 4663 30976
rect 8409 31016 8495 31039
rect 8577 31016 8663 31039
rect 8409 30976 8434 31016
rect 8434 30976 8474 31016
rect 8474 30976 8495 31016
rect 8577 30976 8598 31016
rect 8598 30976 8638 31016
rect 8638 30976 8663 31016
rect 8409 30953 8495 30976
rect 8577 30953 8663 30976
rect 12409 31016 12495 31039
rect 12577 31016 12663 31039
rect 12409 30976 12434 31016
rect 12434 30976 12474 31016
rect 12474 30976 12495 31016
rect 12577 30976 12598 31016
rect 12598 30976 12638 31016
rect 12638 30976 12663 31016
rect 12409 30953 12495 30976
rect 12577 30953 12663 30976
rect 16409 31016 16495 31039
rect 16577 31016 16663 31039
rect 16409 30976 16434 31016
rect 16434 30976 16474 31016
rect 16474 30976 16495 31016
rect 16577 30976 16598 31016
rect 16598 30976 16638 31016
rect 16638 30976 16663 31016
rect 16409 30953 16495 30976
rect 16577 30953 16663 30976
rect 20409 31016 20495 31039
rect 20577 31016 20663 31039
rect 20409 30976 20434 31016
rect 20434 30976 20474 31016
rect 20474 30976 20495 31016
rect 20577 30976 20598 31016
rect 20598 30976 20638 31016
rect 20638 30976 20663 31016
rect 20409 30953 20495 30976
rect 20577 30953 20663 30976
rect 24409 31016 24495 31039
rect 24577 31016 24663 31039
rect 24409 30976 24434 31016
rect 24434 30976 24474 31016
rect 24474 30976 24495 31016
rect 24577 30976 24598 31016
rect 24598 30976 24638 31016
rect 24638 30976 24663 31016
rect 24409 30953 24495 30976
rect 24577 30953 24663 30976
rect 28409 31016 28495 31039
rect 28577 31016 28663 31039
rect 28409 30976 28434 31016
rect 28434 30976 28474 31016
rect 28474 30976 28495 31016
rect 28577 30976 28598 31016
rect 28598 30976 28638 31016
rect 28638 30976 28663 31016
rect 28409 30953 28495 30976
rect 28577 30953 28663 30976
rect 32409 31016 32495 31039
rect 32577 31016 32663 31039
rect 32409 30976 32434 31016
rect 32434 30976 32474 31016
rect 32474 30976 32495 31016
rect 32577 30976 32598 31016
rect 32598 30976 32638 31016
rect 32638 30976 32663 31016
rect 32409 30953 32495 30976
rect 32577 30953 32663 30976
rect 36409 31016 36495 31039
rect 36577 31016 36663 31039
rect 36409 30976 36434 31016
rect 36434 30976 36474 31016
rect 36474 30976 36495 31016
rect 36577 30976 36598 31016
rect 36598 30976 36638 31016
rect 36638 30976 36663 31016
rect 36409 30953 36495 30976
rect 36577 30953 36663 30976
rect 40409 31016 40495 31039
rect 40577 31016 40663 31039
rect 40409 30976 40434 31016
rect 40434 30976 40474 31016
rect 40474 30976 40495 31016
rect 40577 30976 40598 31016
rect 40598 30976 40638 31016
rect 40638 30976 40663 31016
rect 40409 30953 40495 30976
rect 40577 30953 40663 30976
rect 44409 31016 44495 31039
rect 44577 31016 44663 31039
rect 44409 30976 44434 31016
rect 44434 30976 44474 31016
rect 44474 30976 44495 31016
rect 44577 30976 44598 31016
rect 44598 30976 44638 31016
rect 44638 30976 44663 31016
rect 44409 30953 44495 30976
rect 44577 30953 44663 30976
rect 48409 31016 48495 31039
rect 48577 31016 48663 31039
rect 48409 30976 48434 31016
rect 48434 30976 48474 31016
rect 48474 30976 48495 31016
rect 48577 30976 48598 31016
rect 48598 30976 48638 31016
rect 48638 30976 48663 31016
rect 48409 30953 48495 30976
rect 48577 30953 48663 30976
rect 52409 31016 52495 31039
rect 52577 31016 52663 31039
rect 52409 30976 52434 31016
rect 52434 30976 52474 31016
rect 52474 30976 52495 31016
rect 52577 30976 52598 31016
rect 52598 30976 52638 31016
rect 52638 30976 52663 31016
rect 52409 30953 52495 30976
rect 52577 30953 52663 30976
rect 56409 31016 56495 31039
rect 56577 31016 56663 31039
rect 56409 30976 56434 31016
rect 56434 30976 56474 31016
rect 56474 30976 56495 31016
rect 56577 30976 56598 31016
rect 56598 30976 56638 31016
rect 56638 30976 56663 31016
rect 56409 30953 56495 30976
rect 56577 30953 56663 30976
rect 60409 31016 60495 31039
rect 60577 31016 60663 31039
rect 60409 30976 60434 31016
rect 60434 30976 60474 31016
rect 60474 30976 60495 31016
rect 60577 30976 60598 31016
rect 60598 30976 60638 31016
rect 60638 30976 60663 31016
rect 60409 30953 60495 30976
rect 60577 30953 60663 30976
rect 64409 31016 64495 31039
rect 64577 31016 64663 31039
rect 64409 30976 64434 31016
rect 64434 30976 64474 31016
rect 64474 30976 64495 31016
rect 64577 30976 64598 31016
rect 64598 30976 64638 31016
rect 64638 30976 64663 31016
rect 64409 30953 64495 30976
rect 64577 30953 64663 30976
rect 68409 31016 68495 31039
rect 68577 31016 68663 31039
rect 68409 30976 68434 31016
rect 68434 30976 68474 31016
rect 68474 30976 68495 31016
rect 68577 30976 68598 31016
rect 68598 30976 68638 31016
rect 68638 30976 68663 31016
rect 68409 30953 68495 30976
rect 68577 30953 68663 30976
rect 72409 30930 72495 31016
rect 72577 30930 72663 31016
rect 72409 30762 72495 30848
rect 72577 30762 72663 30848
rect 72409 30594 72495 30680
rect 72577 30594 72663 30680
rect 72409 30426 72495 30512
rect 72577 30426 72663 30512
rect 3169 30260 3255 30283
rect 3337 30260 3423 30283
rect 3169 30220 3194 30260
rect 3194 30220 3234 30260
rect 3234 30220 3255 30260
rect 3337 30220 3358 30260
rect 3358 30220 3398 30260
rect 3398 30220 3423 30260
rect 3169 30197 3255 30220
rect 3337 30197 3423 30220
rect 7169 30260 7255 30283
rect 7337 30260 7423 30283
rect 7169 30220 7194 30260
rect 7194 30220 7234 30260
rect 7234 30220 7255 30260
rect 7337 30220 7358 30260
rect 7358 30220 7398 30260
rect 7398 30220 7423 30260
rect 7169 30197 7255 30220
rect 7337 30197 7423 30220
rect 11169 30260 11255 30283
rect 11337 30260 11423 30283
rect 11169 30220 11194 30260
rect 11194 30220 11234 30260
rect 11234 30220 11255 30260
rect 11337 30220 11358 30260
rect 11358 30220 11398 30260
rect 11398 30220 11423 30260
rect 11169 30197 11255 30220
rect 11337 30197 11423 30220
rect 15169 30260 15255 30283
rect 15337 30260 15423 30283
rect 15169 30220 15194 30260
rect 15194 30220 15234 30260
rect 15234 30220 15255 30260
rect 15337 30220 15358 30260
rect 15358 30220 15398 30260
rect 15398 30220 15423 30260
rect 15169 30197 15255 30220
rect 15337 30197 15423 30220
rect 19169 30260 19255 30283
rect 19337 30260 19423 30283
rect 19169 30220 19194 30260
rect 19194 30220 19234 30260
rect 19234 30220 19255 30260
rect 19337 30220 19358 30260
rect 19358 30220 19398 30260
rect 19398 30220 19423 30260
rect 19169 30197 19255 30220
rect 19337 30197 19423 30220
rect 23169 30260 23255 30283
rect 23337 30260 23423 30283
rect 23169 30220 23194 30260
rect 23194 30220 23234 30260
rect 23234 30220 23255 30260
rect 23337 30220 23358 30260
rect 23358 30220 23398 30260
rect 23398 30220 23423 30260
rect 23169 30197 23255 30220
rect 23337 30197 23423 30220
rect 27169 30260 27255 30283
rect 27337 30260 27423 30283
rect 27169 30220 27194 30260
rect 27194 30220 27234 30260
rect 27234 30220 27255 30260
rect 27337 30220 27358 30260
rect 27358 30220 27398 30260
rect 27398 30220 27423 30260
rect 27169 30197 27255 30220
rect 27337 30197 27423 30220
rect 31169 30260 31255 30283
rect 31337 30260 31423 30283
rect 31169 30220 31194 30260
rect 31194 30220 31234 30260
rect 31234 30220 31255 30260
rect 31337 30220 31358 30260
rect 31358 30220 31398 30260
rect 31398 30220 31423 30260
rect 31169 30197 31255 30220
rect 31337 30197 31423 30220
rect 35169 30260 35255 30283
rect 35337 30260 35423 30283
rect 35169 30220 35194 30260
rect 35194 30220 35234 30260
rect 35234 30220 35255 30260
rect 35337 30220 35358 30260
rect 35358 30220 35398 30260
rect 35398 30220 35423 30260
rect 35169 30197 35255 30220
rect 35337 30197 35423 30220
rect 39169 30260 39255 30283
rect 39337 30260 39423 30283
rect 39169 30220 39194 30260
rect 39194 30220 39234 30260
rect 39234 30220 39255 30260
rect 39337 30220 39358 30260
rect 39358 30220 39398 30260
rect 39398 30220 39423 30260
rect 39169 30197 39255 30220
rect 39337 30197 39423 30220
rect 43169 30260 43255 30283
rect 43337 30260 43423 30283
rect 43169 30220 43194 30260
rect 43194 30220 43234 30260
rect 43234 30220 43255 30260
rect 43337 30220 43358 30260
rect 43358 30220 43398 30260
rect 43398 30220 43423 30260
rect 43169 30197 43255 30220
rect 43337 30197 43423 30220
rect 47169 30260 47255 30283
rect 47337 30260 47423 30283
rect 47169 30220 47194 30260
rect 47194 30220 47234 30260
rect 47234 30220 47255 30260
rect 47337 30220 47358 30260
rect 47358 30220 47398 30260
rect 47398 30220 47423 30260
rect 47169 30197 47255 30220
rect 47337 30197 47423 30220
rect 51169 30260 51255 30283
rect 51337 30260 51423 30283
rect 51169 30220 51194 30260
rect 51194 30220 51234 30260
rect 51234 30220 51255 30260
rect 51337 30220 51358 30260
rect 51358 30220 51398 30260
rect 51398 30220 51423 30260
rect 51169 30197 51255 30220
rect 51337 30197 51423 30220
rect 55169 30260 55255 30283
rect 55337 30260 55423 30283
rect 55169 30220 55194 30260
rect 55194 30220 55234 30260
rect 55234 30220 55255 30260
rect 55337 30220 55358 30260
rect 55358 30220 55398 30260
rect 55398 30220 55423 30260
rect 55169 30197 55255 30220
rect 55337 30197 55423 30220
rect 59169 30260 59255 30283
rect 59337 30260 59423 30283
rect 59169 30220 59194 30260
rect 59194 30220 59234 30260
rect 59234 30220 59255 30260
rect 59337 30220 59358 30260
rect 59358 30220 59398 30260
rect 59398 30220 59423 30260
rect 59169 30197 59255 30220
rect 59337 30197 59423 30220
rect 63169 30260 63255 30283
rect 63337 30260 63423 30283
rect 63169 30220 63194 30260
rect 63194 30220 63234 30260
rect 63234 30220 63255 30260
rect 63337 30220 63358 30260
rect 63358 30220 63398 30260
rect 63398 30220 63423 30260
rect 63169 30197 63255 30220
rect 63337 30197 63423 30220
rect 67169 30260 67255 30283
rect 67337 30260 67423 30283
rect 67169 30220 67194 30260
rect 67194 30220 67234 30260
rect 67234 30220 67255 30260
rect 67337 30220 67358 30260
rect 67358 30220 67398 30260
rect 67398 30220 67423 30260
rect 67169 30197 67255 30220
rect 67337 30197 67423 30220
rect 72409 30258 72495 30344
rect 72577 30258 72663 30344
rect 72409 30090 72495 30176
rect 72577 30090 72663 30176
rect 72409 29922 72495 30008
rect 72577 29922 72663 30008
rect 72409 29754 72495 29840
rect 72577 29754 72663 29840
rect 76409 31770 76495 31856
rect 76577 31770 76663 31856
rect 76409 31602 76495 31688
rect 76577 31602 76663 31688
rect 76409 31434 76495 31520
rect 76577 31434 76663 31520
rect 76409 31266 76495 31352
rect 76577 31266 76663 31352
rect 76409 31098 76495 31184
rect 76577 31098 76663 31184
rect 76409 30930 76495 31016
rect 76577 30930 76663 31016
rect 76409 30762 76495 30848
rect 76577 30762 76663 30848
rect 76409 30594 76495 30680
rect 76577 30594 76663 30680
rect 76409 30426 76495 30512
rect 76577 30426 76663 30512
rect 76409 30258 76495 30344
rect 76577 30258 76663 30344
rect 76409 30090 76495 30176
rect 76577 30090 76663 30176
rect 76409 29922 76495 30008
rect 76577 29922 76663 30008
rect 76409 29754 76495 29840
rect 76577 29754 76663 29840
rect 80409 31770 80495 31856
rect 80577 31770 80663 31856
rect 80409 31602 80495 31688
rect 80577 31602 80663 31688
rect 80409 31434 80495 31520
rect 80577 31434 80663 31520
rect 80409 31266 80495 31352
rect 80577 31266 80663 31352
rect 80409 31098 80495 31184
rect 80577 31098 80663 31184
rect 80409 30930 80495 31016
rect 80577 30930 80663 31016
rect 80409 30762 80495 30848
rect 80577 30762 80663 30848
rect 80409 30594 80495 30680
rect 80577 30594 80663 30680
rect 80409 30426 80495 30512
rect 80577 30426 80663 30512
rect 80409 30258 80495 30344
rect 80577 30258 80663 30344
rect 80409 30090 80495 30176
rect 80577 30090 80663 30176
rect 80409 29922 80495 30008
rect 80577 29922 80663 30008
rect 80409 29754 80495 29840
rect 80577 29754 80663 29840
rect 84409 31770 84495 31856
rect 84577 31770 84663 31856
rect 84409 31602 84495 31688
rect 84577 31602 84663 31688
rect 84409 31434 84495 31520
rect 84577 31434 84663 31520
rect 84409 31266 84495 31352
rect 84577 31266 84663 31352
rect 84409 31098 84495 31184
rect 84577 31098 84663 31184
rect 84409 30930 84495 31016
rect 84577 30930 84663 31016
rect 84409 30762 84495 30848
rect 84577 30762 84663 30848
rect 84409 30594 84495 30680
rect 84577 30594 84663 30680
rect 84409 30426 84495 30512
rect 84577 30426 84663 30512
rect 84409 30258 84495 30344
rect 84577 30258 84663 30344
rect 84409 30090 84495 30176
rect 84577 30090 84663 30176
rect 84409 29922 84495 30008
rect 84577 29922 84663 30008
rect 84409 29754 84495 29840
rect 84577 29754 84663 29840
rect 88409 31770 88495 31856
rect 88577 31770 88663 31856
rect 88409 31602 88495 31688
rect 88577 31602 88663 31688
rect 88409 31434 88495 31520
rect 88577 31434 88663 31520
rect 88409 31266 88495 31352
rect 88577 31266 88663 31352
rect 88409 31098 88495 31184
rect 88577 31098 88663 31184
rect 88409 30930 88495 31016
rect 88577 30930 88663 31016
rect 88409 30762 88495 30848
rect 88577 30762 88663 30848
rect 88409 30594 88495 30680
rect 88577 30594 88663 30680
rect 88409 30426 88495 30512
rect 88577 30426 88663 30512
rect 88409 30258 88495 30344
rect 88577 30258 88663 30344
rect 88409 30090 88495 30176
rect 88577 30090 88663 30176
rect 88409 29922 88495 30008
rect 88577 29922 88663 30008
rect 88409 29754 88495 29840
rect 88577 29754 88663 29840
rect 92409 31770 92495 31856
rect 92577 31770 92663 31856
rect 92409 31602 92495 31688
rect 92577 31602 92663 31688
rect 92409 31434 92495 31520
rect 92577 31434 92663 31520
rect 92409 31266 92495 31352
rect 92577 31266 92663 31352
rect 92409 31098 92495 31184
rect 92577 31098 92663 31184
rect 92409 30930 92495 31016
rect 92577 30930 92663 31016
rect 92409 30762 92495 30848
rect 92577 30762 92663 30848
rect 92409 30594 92495 30680
rect 92577 30594 92663 30680
rect 92409 30426 92495 30512
rect 92577 30426 92663 30512
rect 92409 30258 92495 30344
rect 92577 30258 92663 30344
rect 92409 30090 92495 30176
rect 92577 30090 92663 30176
rect 92409 29922 92495 30008
rect 92577 29922 92663 30008
rect 92409 29754 92495 29840
rect 92577 29754 92663 29840
rect 96409 31770 96495 31856
rect 96577 31770 96663 31856
rect 96409 31602 96495 31688
rect 96577 31602 96663 31688
rect 96409 31434 96495 31520
rect 96577 31434 96663 31520
rect 96409 31266 96495 31352
rect 96577 31266 96663 31352
rect 96409 31098 96495 31184
rect 96577 31098 96663 31184
rect 96409 30930 96495 31016
rect 96577 30930 96663 31016
rect 96409 30762 96495 30848
rect 96577 30762 96663 30848
rect 96409 30594 96495 30680
rect 96577 30594 96663 30680
rect 96409 30426 96495 30512
rect 96577 30426 96663 30512
rect 96409 30258 96495 30344
rect 96577 30258 96663 30344
rect 96409 30090 96495 30176
rect 96577 30090 96663 30176
rect 96409 29922 96495 30008
rect 96577 29922 96663 30008
rect 96409 29754 96495 29840
rect 96577 29754 96663 29840
rect 4409 29504 4495 29527
rect 4577 29504 4663 29527
rect 4409 29464 4434 29504
rect 4434 29464 4474 29504
rect 4474 29464 4495 29504
rect 4577 29464 4598 29504
rect 4598 29464 4638 29504
rect 4638 29464 4663 29504
rect 4409 29441 4495 29464
rect 4577 29441 4663 29464
rect 8409 29504 8495 29527
rect 8577 29504 8663 29527
rect 8409 29464 8434 29504
rect 8434 29464 8474 29504
rect 8474 29464 8495 29504
rect 8577 29464 8598 29504
rect 8598 29464 8638 29504
rect 8638 29464 8663 29504
rect 8409 29441 8495 29464
rect 8577 29441 8663 29464
rect 12409 29504 12495 29527
rect 12577 29504 12663 29527
rect 12409 29464 12434 29504
rect 12434 29464 12474 29504
rect 12474 29464 12495 29504
rect 12577 29464 12598 29504
rect 12598 29464 12638 29504
rect 12638 29464 12663 29504
rect 12409 29441 12495 29464
rect 12577 29441 12663 29464
rect 16409 29504 16495 29527
rect 16577 29504 16663 29527
rect 16409 29464 16434 29504
rect 16434 29464 16474 29504
rect 16474 29464 16495 29504
rect 16577 29464 16598 29504
rect 16598 29464 16638 29504
rect 16638 29464 16663 29504
rect 16409 29441 16495 29464
rect 16577 29441 16663 29464
rect 20409 29504 20495 29527
rect 20577 29504 20663 29527
rect 20409 29464 20434 29504
rect 20434 29464 20474 29504
rect 20474 29464 20495 29504
rect 20577 29464 20598 29504
rect 20598 29464 20638 29504
rect 20638 29464 20663 29504
rect 20409 29441 20495 29464
rect 20577 29441 20663 29464
rect 24409 29504 24495 29527
rect 24577 29504 24663 29527
rect 24409 29464 24434 29504
rect 24434 29464 24474 29504
rect 24474 29464 24495 29504
rect 24577 29464 24598 29504
rect 24598 29464 24638 29504
rect 24638 29464 24663 29504
rect 24409 29441 24495 29464
rect 24577 29441 24663 29464
rect 28409 29504 28495 29527
rect 28577 29504 28663 29527
rect 28409 29464 28434 29504
rect 28434 29464 28474 29504
rect 28474 29464 28495 29504
rect 28577 29464 28598 29504
rect 28598 29464 28638 29504
rect 28638 29464 28663 29504
rect 28409 29441 28495 29464
rect 28577 29441 28663 29464
rect 32409 29504 32495 29527
rect 32577 29504 32663 29527
rect 32409 29464 32434 29504
rect 32434 29464 32474 29504
rect 32474 29464 32495 29504
rect 32577 29464 32598 29504
rect 32598 29464 32638 29504
rect 32638 29464 32663 29504
rect 32409 29441 32495 29464
rect 32577 29441 32663 29464
rect 36409 29504 36495 29527
rect 36577 29504 36663 29527
rect 36409 29464 36434 29504
rect 36434 29464 36474 29504
rect 36474 29464 36495 29504
rect 36577 29464 36598 29504
rect 36598 29464 36638 29504
rect 36638 29464 36663 29504
rect 36409 29441 36495 29464
rect 36577 29441 36663 29464
rect 40409 29504 40495 29527
rect 40577 29504 40663 29527
rect 40409 29464 40434 29504
rect 40434 29464 40474 29504
rect 40474 29464 40495 29504
rect 40577 29464 40598 29504
rect 40598 29464 40638 29504
rect 40638 29464 40663 29504
rect 40409 29441 40495 29464
rect 40577 29441 40663 29464
rect 44409 29504 44495 29527
rect 44577 29504 44663 29527
rect 44409 29464 44434 29504
rect 44434 29464 44474 29504
rect 44474 29464 44495 29504
rect 44577 29464 44598 29504
rect 44598 29464 44638 29504
rect 44638 29464 44663 29504
rect 44409 29441 44495 29464
rect 44577 29441 44663 29464
rect 48409 29504 48495 29527
rect 48577 29504 48663 29527
rect 48409 29464 48434 29504
rect 48434 29464 48474 29504
rect 48474 29464 48495 29504
rect 48577 29464 48598 29504
rect 48598 29464 48638 29504
rect 48638 29464 48663 29504
rect 48409 29441 48495 29464
rect 48577 29441 48663 29464
rect 52409 29504 52495 29527
rect 52577 29504 52663 29527
rect 52409 29464 52434 29504
rect 52434 29464 52474 29504
rect 52474 29464 52495 29504
rect 52577 29464 52598 29504
rect 52598 29464 52638 29504
rect 52638 29464 52663 29504
rect 52409 29441 52495 29464
rect 52577 29441 52663 29464
rect 56409 29504 56495 29527
rect 56577 29504 56663 29527
rect 56409 29464 56434 29504
rect 56434 29464 56474 29504
rect 56474 29464 56495 29504
rect 56577 29464 56598 29504
rect 56598 29464 56638 29504
rect 56638 29464 56663 29504
rect 56409 29441 56495 29464
rect 56577 29441 56663 29464
rect 60409 29504 60495 29527
rect 60577 29504 60663 29527
rect 60409 29464 60434 29504
rect 60434 29464 60474 29504
rect 60474 29464 60495 29504
rect 60577 29464 60598 29504
rect 60598 29464 60638 29504
rect 60638 29464 60663 29504
rect 60409 29441 60495 29464
rect 60577 29441 60663 29464
rect 64409 29504 64495 29527
rect 64577 29504 64663 29527
rect 64409 29464 64434 29504
rect 64434 29464 64474 29504
rect 64474 29464 64495 29504
rect 64577 29464 64598 29504
rect 64598 29464 64638 29504
rect 64638 29464 64663 29504
rect 64409 29441 64495 29464
rect 64577 29441 64663 29464
rect 68409 29504 68495 29527
rect 68577 29504 68663 29527
rect 68409 29464 68434 29504
rect 68434 29464 68474 29504
rect 68474 29464 68495 29504
rect 68577 29464 68598 29504
rect 68598 29464 68638 29504
rect 68638 29464 68663 29504
rect 68409 29441 68495 29464
rect 68577 29441 68663 29464
rect 75169 28894 75255 28980
rect 75337 28894 75423 28980
rect 3169 28748 3255 28771
rect 3337 28748 3423 28771
rect 3169 28708 3194 28748
rect 3194 28708 3234 28748
rect 3234 28708 3255 28748
rect 3337 28708 3358 28748
rect 3358 28708 3398 28748
rect 3398 28708 3423 28748
rect 3169 28685 3255 28708
rect 3337 28685 3423 28708
rect 7169 28748 7255 28771
rect 7337 28748 7423 28771
rect 7169 28708 7194 28748
rect 7194 28708 7234 28748
rect 7234 28708 7255 28748
rect 7337 28708 7358 28748
rect 7358 28708 7398 28748
rect 7398 28708 7423 28748
rect 7169 28685 7255 28708
rect 7337 28685 7423 28708
rect 11169 28748 11255 28771
rect 11337 28748 11423 28771
rect 11169 28708 11194 28748
rect 11194 28708 11234 28748
rect 11234 28708 11255 28748
rect 11337 28708 11358 28748
rect 11358 28708 11398 28748
rect 11398 28708 11423 28748
rect 11169 28685 11255 28708
rect 11337 28685 11423 28708
rect 15169 28748 15255 28771
rect 15337 28748 15423 28771
rect 15169 28708 15194 28748
rect 15194 28708 15234 28748
rect 15234 28708 15255 28748
rect 15337 28708 15358 28748
rect 15358 28708 15398 28748
rect 15398 28708 15423 28748
rect 15169 28685 15255 28708
rect 15337 28685 15423 28708
rect 19169 28748 19255 28771
rect 19337 28748 19423 28771
rect 19169 28708 19194 28748
rect 19194 28708 19234 28748
rect 19234 28708 19255 28748
rect 19337 28708 19358 28748
rect 19358 28708 19398 28748
rect 19398 28708 19423 28748
rect 19169 28685 19255 28708
rect 19337 28685 19423 28708
rect 23169 28748 23255 28771
rect 23337 28748 23423 28771
rect 23169 28708 23194 28748
rect 23194 28708 23234 28748
rect 23234 28708 23255 28748
rect 23337 28708 23358 28748
rect 23358 28708 23398 28748
rect 23398 28708 23423 28748
rect 23169 28685 23255 28708
rect 23337 28685 23423 28708
rect 27169 28748 27255 28771
rect 27337 28748 27423 28771
rect 27169 28708 27194 28748
rect 27194 28708 27234 28748
rect 27234 28708 27255 28748
rect 27337 28708 27358 28748
rect 27358 28708 27398 28748
rect 27398 28708 27423 28748
rect 27169 28685 27255 28708
rect 27337 28685 27423 28708
rect 31169 28748 31255 28771
rect 31337 28748 31423 28771
rect 31169 28708 31194 28748
rect 31194 28708 31234 28748
rect 31234 28708 31255 28748
rect 31337 28708 31358 28748
rect 31358 28708 31398 28748
rect 31398 28708 31423 28748
rect 31169 28685 31255 28708
rect 31337 28685 31423 28708
rect 35169 28748 35255 28771
rect 35337 28748 35423 28771
rect 35169 28708 35194 28748
rect 35194 28708 35234 28748
rect 35234 28708 35255 28748
rect 35337 28708 35358 28748
rect 35358 28708 35398 28748
rect 35398 28708 35423 28748
rect 35169 28685 35255 28708
rect 35337 28685 35423 28708
rect 39169 28748 39255 28771
rect 39337 28748 39423 28771
rect 39169 28708 39194 28748
rect 39194 28708 39234 28748
rect 39234 28708 39255 28748
rect 39337 28708 39358 28748
rect 39358 28708 39398 28748
rect 39398 28708 39423 28748
rect 39169 28685 39255 28708
rect 39337 28685 39423 28708
rect 43169 28748 43255 28771
rect 43337 28748 43423 28771
rect 43169 28708 43194 28748
rect 43194 28708 43234 28748
rect 43234 28708 43255 28748
rect 43337 28708 43358 28748
rect 43358 28708 43398 28748
rect 43398 28708 43423 28748
rect 43169 28685 43255 28708
rect 43337 28685 43423 28708
rect 47169 28748 47255 28771
rect 47337 28748 47423 28771
rect 47169 28708 47194 28748
rect 47194 28708 47234 28748
rect 47234 28708 47255 28748
rect 47337 28708 47358 28748
rect 47358 28708 47398 28748
rect 47398 28708 47423 28748
rect 47169 28685 47255 28708
rect 47337 28685 47423 28708
rect 51169 28748 51255 28771
rect 51337 28748 51423 28771
rect 51169 28708 51194 28748
rect 51194 28708 51234 28748
rect 51234 28708 51255 28748
rect 51337 28708 51358 28748
rect 51358 28708 51398 28748
rect 51398 28708 51423 28748
rect 51169 28685 51255 28708
rect 51337 28685 51423 28708
rect 55169 28748 55255 28771
rect 55337 28748 55423 28771
rect 55169 28708 55194 28748
rect 55194 28708 55234 28748
rect 55234 28708 55255 28748
rect 55337 28708 55358 28748
rect 55358 28708 55398 28748
rect 55398 28708 55423 28748
rect 55169 28685 55255 28708
rect 55337 28685 55423 28708
rect 59169 28748 59255 28771
rect 59337 28748 59423 28771
rect 59169 28708 59194 28748
rect 59194 28708 59234 28748
rect 59234 28708 59255 28748
rect 59337 28708 59358 28748
rect 59358 28708 59398 28748
rect 59398 28708 59423 28748
rect 59169 28685 59255 28708
rect 59337 28685 59423 28708
rect 63169 28748 63255 28771
rect 63337 28748 63423 28771
rect 63169 28708 63194 28748
rect 63194 28708 63234 28748
rect 63234 28708 63255 28748
rect 63337 28708 63358 28748
rect 63358 28708 63398 28748
rect 63398 28708 63423 28748
rect 63169 28685 63255 28708
rect 63337 28685 63423 28708
rect 67169 28748 67255 28771
rect 67337 28748 67423 28771
rect 67169 28708 67194 28748
rect 67194 28708 67234 28748
rect 67234 28708 67255 28748
rect 67337 28708 67358 28748
rect 67358 28708 67398 28748
rect 67398 28708 67423 28748
rect 67169 28685 67255 28708
rect 67337 28685 67423 28708
rect 75169 28726 75255 28812
rect 75337 28726 75423 28812
rect 75169 28558 75255 28644
rect 75337 28558 75423 28644
rect 75169 28390 75255 28476
rect 75337 28390 75423 28476
rect 75169 28222 75255 28308
rect 75337 28222 75423 28308
rect 75169 28054 75255 28140
rect 75337 28054 75423 28140
rect 4409 27992 4495 28015
rect 4577 27992 4663 28015
rect 4409 27952 4434 27992
rect 4434 27952 4474 27992
rect 4474 27952 4495 27992
rect 4577 27952 4598 27992
rect 4598 27952 4638 27992
rect 4638 27952 4663 27992
rect 4409 27929 4495 27952
rect 4577 27929 4663 27952
rect 8409 27992 8495 28015
rect 8577 27992 8663 28015
rect 8409 27952 8434 27992
rect 8434 27952 8474 27992
rect 8474 27952 8495 27992
rect 8577 27952 8598 27992
rect 8598 27952 8638 27992
rect 8638 27952 8663 27992
rect 8409 27929 8495 27952
rect 8577 27929 8663 27952
rect 12409 27992 12495 28015
rect 12577 27992 12663 28015
rect 12409 27952 12434 27992
rect 12434 27952 12474 27992
rect 12474 27952 12495 27992
rect 12577 27952 12598 27992
rect 12598 27952 12638 27992
rect 12638 27952 12663 27992
rect 12409 27929 12495 27952
rect 12577 27929 12663 27952
rect 16409 27992 16495 28015
rect 16577 27992 16663 28015
rect 16409 27952 16434 27992
rect 16434 27952 16474 27992
rect 16474 27952 16495 27992
rect 16577 27952 16598 27992
rect 16598 27952 16638 27992
rect 16638 27952 16663 27992
rect 16409 27929 16495 27952
rect 16577 27929 16663 27952
rect 20409 27992 20495 28015
rect 20577 27992 20663 28015
rect 20409 27952 20434 27992
rect 20434 27952 20474 27992
rect 20474 27952 20495 27992
rect 20577 27952 20598 27992
rect 20598 27952 20638 27992
rect 20638 27952 20663 27992
rect 20409 27929 20495 27952
rect 20577 27929 20663 27952
rect 24409 27992 24495 28015
rect 24577 27992 24663 28015
rect 24409 27952 24434 27992
rect 24434 27952 24474 27992
rect 24474 27952 24495 27992
rect 24577 27952 24598 27992
rect 24598 27952 24638 27992
rect 24638 27952 24663 27992
rect 24409 27929 24495 27952
rect 24577 27929 24663 27952
rect 28409 27992 28495 28015
rect 28577 27992 28663 28015
rect 28409 27952 28434 27992
rect 28434 27952 28474 27992
rect 28474 27952 28495 27992
rect 28577 27952 28598 27992
rect 28598 27952 28638 27992
rect 28638 27952 28663 27992
rect 28409 27929 28495 27952
rect 28577 27929 28663 27952
rect 32409 27992 32495 28015
rect 32577 27992 32663 28015
rect 32409 27952 32434 27992
rect 32434 27952 32474 27992
rect 32474 27952 32495 27992
rect 32577 27952 32598 27992
rect 32598 27952 32638 27992
rect 32638 27952 32663 27992
rect 32409 27929 32495 27952
rect 32577 27929 32663 27952
rect 36409 27992 36495 28015
rect 36577 27992 36663 28015
rect 36409 27952 36434 27992
rect 36434 27952 36474 27992
rect 36474 27952 36495 27992
rect 36577 27952 36598 27992
rect 36598 27952 36638 27992
rect 36638 27952 36663 27992
rect 36409 27929 36495 27952
rect 36577 27929 36663 27952
rect 40409 27992 40495 28015
rect 40577 27992 40663 28015
rect 40409 27952 40434 27992
rect 40434 27952 40474 27992
rect 40474 27952 40495 27992
rect 40577 27952 40598 27992
rect 40598 27952 40638 27992
rect 40638 27952 40663 27992
rect 40409 27929 40495 27952
rect 40577 27929 40663 27952
rect 44409 27992 44495 28015
rect 44577 27992 44663 28015
rect 44409 27952 44434 27992
rect 44434 27952 44474 27992
rect 44474 27952 44495 27992
rect 44577 27952 44598 27992
rect 44598 27952 44638 27992
rect 44638 27952 44663 27992
rect 44409 27929 44495 27952
rect 44577 27929 44663 27952
rect 48409 27992 48495 28015
rect 48577 27992 48663 28015
rect 48409 27952 48434 27992
rect 48434 27952 48474 27992
rect 48474 27952 48495 27992
rect 48577 27952 48598 27992
rect 48598 27952 48638 27992
rect 48638 27952 48663 27992
rect 48409 27929 48495 27952
rect 48577 27929 48663 27952
rect 52409 27992 52495 28015
rect 52577 27992 52663 28015
rect 52409 27952 52434 27992
rect 52434 27952 52474 27992
rect 52474 27952 52495 27992
rect 52577 27952 52598 27992
rect 52598 27952 52638 27992
rect 52638 27952 52663 27992
rect 52409 27929 52495 27952
rect 52577 27929 52663 27952
rect 56409 27992 56495 28015
rect 56577 27992 56663 28015
rect 56409 27952 56434 27992
rect 56434 27952 56474 27992
rect 56474 27952 56495 27992
rect 56577 27952 56598 27992
rect 56598 27952 56638 27992
rect 56638 27952 56663 27992
rect 56409 27929 56495 27952
rect 56577 27929 56663 27952
rect 60409 27992 60495 28015
rect 60577 27992 60663 28015
rect 60409 27952 60434 27992
rect 60434 27952 60474 27992
rect 60474 27952 60495 27992
rect 60577 27952 60598 27992
rect 60598 27952 60638 27992
rect 60638 27952 60663 27992
rect 60409 27929 60495 27952
rect 60577 27929 60663 27952
rect 64409 27992 64495 28015
rect 64577 27992 64663 28015
rect 64409 27952 64434 27992
rect 64434 27952 64474 27992
rect 64474 27952 64495 27992
rect 64577 27952 64598 27992
rect 64598 27952 64638 27992
rect 64638 27952 64663 27992
rect 64409 27929 64495 27952
rect 64577 27929 64663 27952
rect 68409 27992 68495 28015
rect 68577 27992 68663 28015
rect 68409 27952 68434 27992
rect 68434 27952 68474 27992
rect 68474 27952 68495 27992
rect 68577 27952 68598 27992
rect 68598 27952 68638 27992
rect 68638 27952 68663 27992
rect 68409 27929 68495 27952
rect 68577 27929 68663 27952
rect 75169 27886 75255 27972
rect 75337 27886 75423 27972
rect 75169 27718 75255 27804
rect 75337 27718 75423 27804
rect 75169 27550 75255 27636
rect 75337 27550 75423 27636
rect 75169 27382 75255 27468
rect 75337 27382 75423 27468
rect 3169 27236 3255 27259
rect 3337 27236 3423 27259
rect 3169 27196 3194 27236
rect 3194 27196 3234 27236
rect 3234 27196 3255 27236
rect 3337 27196 3358 27236
rect 3358 27196 3398 27236
rect 3398 27196 3423 27236
rect 3169 27173 3255 27196
rect 3337 27173 3423 27196
rect 7169 27236 7255 27259
rect 7337 27236 7423 27259
rect 7169 27196 7194 27236
rect 7194 27196 7234 27236
rect 7234 27196 7255 27236
rect 7337 27196 7358 27236
rect 7358 27196 7398 27236
rect 7398 27196 7423 27236
rect 7169 27173 7255 27196
rect 7337 27173 7423 27196
rect 11169 27236 11255 27259
rect 11337 27236 11423 27259
rect 11169 27196 11194 27236
rect 11194 27196 11234 27236
rect 11234 27196 11255 27236
rect 11337 27196 11358 27236
rect 11358 27196 11398 27236
rect 11398 27196 11423 27236
rect 11169 27173 11255 27196
rect 11337 27173 11423 27196
rect 15169 27236 15255 27259
rect 15337 27236 15423 27259
rect 15169 27196 15194 27236
rect 15194 27196 15234 27236
rect 15234 27196 15255 27236
rect 15337 27196 15358 27236
rect 15358 27196 15398 27236
rect 15398 27196 15423 27236
rect 15169 27173 15255 27196
rect 15337 27173 15423 27196
rect 19169 27236 19255 27259
rect 19337 27236 19423 27259
rect 19169 27196 19194 27236
rect 19194 27196 19234 27236
rect 19234 27196 19255 27236
rect 19337 27196 19358 27236
rect 19358 27196 19398 27236
rect 19398 27196 19423 27236
rect 19169 27173 19255 27196
rect 19337 27173 19423 27196
rect 23169 27236 23255 27259
rect 23337 27236 23423 27259
rect 23169 27196 23194 27236
rect 23194 27196 23234 27236
rect 23234 27196 23255 27236
rect 23337 27196 23358 27236
rect 23358 27196 23398 27236
rect 23398 27196 23423 27236
rect 23169 27173 23255 27196
rect 23337 27173 23423 27196
rect 27169 27236 27255 27259
rect 27337 27236 27423 27259
rect 27169 27196 27194 27236
rect 27194 27196 27234 27236
rect 27234 27196 27255 27236
rect 27337 27196 27358 27236
rect 27358 27196 27398 27236
rect 27398 27196 27423 27236
rect 27169 27173 27255 27196
rect 27337 27173 27423 27196
rect 31169 27236 31255 27259
rect 31337 27236 31423 27259
rect 31169 27196 31194 27236
rect 31194 27196 31234 27236
rect 31234 27196 31255 27236
rect 31337 27196 31358 27236
rect 31358 27196 31398 27236
rect 31398 27196 31423 27236
rect 31169 27173 31255 27196
rect 31337 27173 31423 27196
rect 35169 27236 35255 27259
rect 35337 27236 35423 27259
rect 35169 27196 35194 27236
rect 35194 27196 35234 27236
rect 35234 27196 35255 27236
rect 35337 27196 35358 27236
rect 35358 27196 35398 27236
rect 35398 27196 35423 27236
rect 35169 27173 35255 27196
rect 35337 27173 35423 27196
rect 39169 27236 39255 27259
rect 39337 27236 39423 27259
rect 39169 27196 39194 27236
rect 39194 27196 39234 27236
rect 39234 27196 39255 27236
rect 39337 27196 39358 27236
rect 39358 27196 39398 27236
rect 39398 27196 39423 27236
rect 39169 27173 39255 27196
rect 39337 27173 39423 27196
rect 43169 27236 43255 27259
rect 43337 27236 43423 27259
rect 43169 27196 43194 27236
rect 43194 27196 43234 27236
rect 43234 27196 43255 27236
rect 43337 27196 43358 27236
rect 43358 27196 43398 27236
rect 43398 27196 43423 27236
rect 43169 27173 43255 27196
rect 43337 27173 43423 27196
rect 47169 27236 47255 27259
rect 47337 27236 47423 27259
rect 47169 27196 47194 27236
rect 47194 27196 47234 27236
rect 47234 27196 47255 27236
rect 47337 27196 47358 27236
rect 47358 27196 47398 27236
rect 47398 27196 47423 27236
rect 47169 27173 47255 27196
rect 47337 27173 47423 27196
rect 51169 27236 51255 27259
rect 51337 27236 51423 27259
rect 51169 27196 51194 27236
rect 51194 27196 51234 27236
rect 51234 27196 51255 27236
rect 51337 27196 51358 27236
rect 51358 27196 51398 27236
rect 51398 27196 51423 27236
rect 51169 27173 51255 27196
rect 51337 27173 51423 27196
rect 55169 27236 55255 27259
rect 55337 27236 55423 27259
rect 55169 27196 55194 27236
rect 55194 27196 55234 27236
rect 55234 27196 55255 27236
rect 55337 27196 55358 27236
rect 55358 27196 55398 27236
rect 55398 27196 55423 27236
rect 55169 27173 55255 27196
rect 55337 27173 55423 27196
rect 59169 27236 59255 27259
rect 59337 27236 59423 27259
rect 59169 27196 59194 27236
rect 59194 27196 59234 27236
rect 59234 27196 59255 27236
rect 59337 27196 59358 27236
rect 59358 27196 59398 27236
rect 59398 27196 59423 27236
rect 59169 27173 59255 27196
rect 59337 27173 59423 27196
rect 63169 27236 63255 27259
rect 63337 27236 63423 27259
rect 63169 27196 63194 27236
rect 63194 27196 63234 27236
rect 63234 27196 63255 27236
rect 63337 27196 63358 27236
rect 63358 27196 63398 27236
rect 63398 27196 63423 27236
rect 63169 27173 63255 27196
rect 63337 27173 63423 27196
rect 67169 27236 67255 27259
rect 67337 27236 67423 27259
rect 67169 27196 67194 27236
rect 67194 27196 67234 27236
rect 67234 27196 67255 27236
rect 67337 27196 67358 27236
rect 67358 27196 67398 27236
rect 67398 27196 67423 27236
rect 67169 27173 67255 27196
rect 67337 27173 67423 27196
rect 75169 27214 75255 27300
rect 75337 27214 75423 27300
rect 75169 27046 75255 27132
rect 75337 27046 75423 27132
rect 75169 26878 75255 26964
rect 75337 26878 75423 26964
rect 79169 28894 79255 28980
rect 79337 28894 79423 28980
rect 79169 28726 79255 28812
rect 79337 28726 79423 28812
rect 79169 28558 79255 28644
rect 79337 28558 79423 28644
rect 79169 28390 79255 28476
rect 79337 28390 79423 28476
rect 79169 28222 79255 28308
rect 79337 28222 79423 28308
rect 79169 28054 79255 28140
rect 79337 28054 79423 28140
rect 79169 27886 79255 27972
rect 79337 27886 79423 27972
rect 79169 27718 79255 27804
rect 79337 27718 79423 27804
rect 79169 27550 79255 27636
rect 79337 27550 79423 27636
rect 79169 27382 79255 27468
rect 79337 27382 79423 27468
rect 79169 27214 79255 27300
rect 79337 27214 79423 27300
rect 79169 27046 79255 27132
rect 79337 27046 79423 27132
rect 79169 26878 79255 26964
rect 79337 26878 79423 26964
rect 83169 28894 83255 28980
rect 83337 28894 83423 28980
rect 83169 28726 83255 28812
rect 83337 28726 83423 28812
rect 83169 28558 83255 28644
rect 83337 28558 83423 28644
rect 83169 28390 83255 28476
rect 83337 28390 83423 28476
rect 83169 28222 83255 28308
rect 83337 28222 83423 28308
rect 83169 28054 83255 28140
rect 83337 28054 83423 28140
rect 83169 27886 83255 27972
rect 83337 27886 83423 27972
rect 83169 27718 83255 27804
rect 83337 27718 83423 27804
rect 83169 27550 83255 27636
rect 83337 27550 83423 27636
rect 83169 27382 83255 27468
rect 83337 27382 83423 27468
rect 83169 27214 83255 27300
rect 83337 27214 83423 27300
rect 83169 27046 83255 27132
rect 83337 27046 83423 27132
rect 83169 26878 83255 26964
rect 83337 26878 83423 26964
rect 87169 28894 87255 28980
rect 87337 28894 87423 28980
rect 87169 28726 87255 28812
rect 87337 28726 87423 28812
rect 87169 28558 87255 28644
rect 87337 28558 87423 28644
rect 87169 28390 87255 28476
rect 87337 28390 87423 28476
rect 87169 28222 87255 28308
rect 87337 28222 87423 28308
rect 87169 28054 87255 28140
rect 87337 28054 87423 28140
rect 87169 27886 87255 27972
rect 87337 27886 87423 27972
rect 87169 27718 87255 27804
rect 87337 27718 87423 27804
rect 87169 27550 87255 27636
rect 87337 27550 87423 27636
rect 87169 27382 87255 27468
rect 87337 27382 87423 27468
rect 87169 27214 87255 27300
rect 87337 27214 87423 27300
rect 87169 27046 87255 27132
rect 87337 27046 87423 27132
rect 87169 26878 87255 26964
rect 87337 26878 87423 26964
rect 91169 28894 91255 28980
rect 91337 28894 91423 28980
rect 91169 28726 91255 28812
rect 91337 28726 91423 28812
rect 91169 28558 91255 28644
rect 91337 28558 91423 28644
rect 91169 28390 91255 28476
rect 91337 28390 91423 28476
rect 91169 28222 91255 28308
rect 91337 28222 91423 28308
rect 91169 28054 91255 28140
rect 91337 28054 91423 28140
rect 91169 27886 91255 27972
rect 91337 27886 91423 27972
rect 91169 27718 91255 27804
rect 91337 27718 91423 27804
rect 91169 27550 91255 27636
rect 91337 27550 91423 27636
rect 91169 27382 91255 27468
rect 91337 27382 91423 27468
rect 91169 27214 91255 27300
rect 91337 27214 91423 27300
rect 91169 27046 91255 27132
rect 91337 27046 91423 27132
rect 91169 26878 91255 26964
rect 91337 26878 91423 26964
rect 95169 28894 95255 28980
rect 95337 28894 95423 28980
rect 95169 28726 95255 28812
rect 95337 28726 95423 28812
rect 95169 28558 95255 28644
rect 95337 28558 95423 28644
rect 95169 28390 95255 28476
rect 95337 28390 95423 28476
rect 95169 28222 95255 28308
rect 95337 28222 95423 28308
rect 95169 28054 95255 28140
rect 95337 28054 95423 28140
rect 95169 27886 95255 27972
rect 95337 27886 95423 27972
rect 95169 27718 95255 27804
rect 95337 27718 95423 27804
rect 95169 27550 95255 27636
rect 95337 27550 95423 27636
rect 95169 27382 95255 27468
rect 95337 27382 95423 27468
rect 95169 27214 95255 27300
rect 95337 27214 95423 27300
rect 95169 27046 95255 27132
rect 95337 27046 95423 27132
rect 95169 26878 95255 26964
rect 95337 26878 95423 26964
rect 73245 26564 73331 26587
rect 73245 26524 73268 26564
rect 73268 26524 73331 26564
rect 4409 26480 4495 26503
rect 4577 26480 4663 26503
rect 4409 26440 4434 26480
rect 4434 26440 4474 26480
rect 4474 26440 4495 26480
rect 4577 26440 4598 26480
rect 4598 26440 4638 26480
rect 4638 26440 4663 26480
rect 4409 26417 4495 26440
rect 4577 26417 4663 26440
rect 8409 26480 8495 26503
rect 8577 26480 8663 26503
rect 8409 26440 8434 26480
rect 8434 26440 8474 26480
rect 8474 26440 8495 26480
rect 8577 26440 8598 26480
rect 8598 26440 8638 26480
rect 8638 26440 8663 26480
rect 8409 26417 8495 26440
rect 8577 26417 8663 26440
rect 12409 26480 12495 26503
rect 12577 26480 12663 26503
rect 12409 26440 12434 26480
rect 12434 26440 12474 26480
rect 12474 26440 12495 26480
rect 12577 26440 12598 26480
rect 12598 26440 12638 26480
rect 12638 26440 12663 26480
rect 12409 26417 12495 26440
rect 12577 26417 12663 26440
rect 16409 26480 16495 26503
rect 16577 26480 16663 26503
rect 16409 26440 16434 26480
rect 16434 26440 16474 26480
rect 16474 26440 16495 26480
rect 16577 26440 16598 26480
rect 16598 26440 16638 26480
rect 16638 26440 16663 26480
rect 16409 26417 16495 26440
rect 16577 26417 16663 26440
rect 20409 26480 20495 26503
rect 20577 26480 20663 26503
rect 20409 26440 20434 26480
rect 20434 26440 20474 26480
rect 20474 26440 20495 26480
rect 20577 26440 20598 26480
rect 20598 26440 20638 26480
rect 20638 26440 20663 26480
rect 20409 26417 20495 26440
rect 20577 26417 20663 26440
rect 24409 26480 24495 26503
rect 24577 26480 24663 26503
rect 24409 26440 24434 26480
rect 24434 26440 24474 26480
rect 24474 26440 24495 26480
rect 24577 26440 24598 26480
rect 24598 26440 24638 26480
rect 24638 26440 24663 26480
rect 24409 26417 24495 26440
rect 24577 26417 24663 26440
rect 28409 26480 28495 26503
rect 28577 26480 28663 26503
rect 28409 26440 28434 26480
rect 28434 26440 28474 26480
rect 28474 26440 28495 26480
rect 28577 26440 28598 26480
rect 28598 26440 28638 26480
rect 28638 26440 28663 26480
rect 28409 26417 28495 26440
rect 28577 26417 28663 26440
rect 32409 26480 32495 26503
rect 32577 26480 32663 26503
rect 32409 26440 32434 26480
rect 32434 26440 32474 26480
rect 32474 26440 32495 26480
rect 32577 26440 32598 26480
rect 32598 26440 32638 26480
rect 32638 26440 32663 26480
rect 32409 26417 32495 26440
rect 32577 26417 32663 26440
rect 36409 26480 36495 26503
rect 36577 26480 36663 26503
rect 36409 26440 36434 26480
rect 36434 26440 36474 26480
rect 36474 26440 36495 26480
rect 36577 26440 36598 26480
rect 36598 26440 36638 26480
rect 36638 26440 36663 26480
rect 36409 26417 36495 26440
rect 36577 26417 36663 26440
rect 40409 26480 40495 26503
rect 40577 26480 40663 26503
rect 40409 26440 40434 26480
rect 40434 26440 40474 26480
rect 40474 26440 40495 26480
rect 40577 26440 40598 26480
rect 40598 26440 40638 26480
rect 40638 26440 40663 26480
rect 40409 26417 40495 26440
rect 40577 26417 40663 26440
rect 44409 26480 44495 26503
rect 44577 26480 44663 26503
rect 44409 26440 44434 26480
rect 44434 26440 44474 26480
rect 44474 26440 44495 26480
rect 44577 26440 44598 26480
rect 44598 26440 44638 26480
rect 44638 26440 44663 26480
rect 44409 26417 44495 26440
rect 44577 26417 44663 26440
rect 48409 26480 48495 26503
rect 48577 26480 48663 26503
rect 48409 26440 48434 26480
rect 48434 26440 48474 26480
rect 48474 26440 48495 26480
rect 48577 26440 48598 26480
rect 48598 26440 48638 26480
rect 48638 26440 48663 26480
rect 48409 26417 48495 26440
rect 48577 26417 48663 26440
rect 52409 26480 52495 26503
rect 52577 26480 52663 26503
rect 52409 26440 52434 26480
rect 52434 26440 52474 26480
rect 52474 26440 52495 26480
rect 52577 26440 52598 26480
rect 52598 26440 52638 26480
rect 52638 26440 52663 26480
rect 52409 26417 52495 26440
rect 52577 26417 52663 26440
rect 56409 26480 56495 26503
rect 56577 26480 56663 26503
rect 56409 26440 56434 26480
rect 56434 26440 56474 26480
rect 56474 26440 56495 26480
rect 56577 26440 56598 26480
rect 56598 26440 56638 26480
rect 56638 26440 56663 26480
rect 56409 26417 56495 26440
rect 56577 26417 56663 26440
rect 60409 26480 60495 26503
rect 60577 26480 60663 26503
rect 60409 26440 60434 26480
rect 60434 26440 60474 26480
rect 60474 26440 60495 26480
rect 60577 26440 60598 26480
rect 60598 26440 60638 26480
rect 60638 26440 60663 26480
rect 60409 26417 60495 26440
rect 60577 26417 60663 26440
rect 64409 26480 64495 26503
rect 64577 26480 64663 26503
rect 64409 26440 64434 26480
rect 64434 26440 64474 26480
rect 64474 26440 64495 26480
rect 64577 26440 64598 26480
rect 64598 26440 64638 26480
rect 64638 26440 64663 26480
rect 64409 26417 64495 26440
rect 64577 26417 64663 26440
rect 68409 26480 68495 26503
rect 68577 26480 68663 26503
rect 73245 26501 73331 26524
rect 68409 26440 68434 26480
rect 68434 26440 68474 26480
rect 68474 26440 68495 26480
rect 68577 26440 68598 26480
rect 68598 26440 68638 26480
rect 68638 26440 68663 26480
rect 68409 26417 68495 26440
rect 68577 26417 68663 26440
rect 3169 25724 3255 25747
rect 3337 25724 3423 25747
rect 3169 25684 3194 25724
rect 3194 25684 3234 25724
rect 3234 25684 3255 25724
rect 3337 25684 3358 25724
rect 3358 25684 3398 25724
rect 3398 25684 3423 25724
rect 3169 25661 3255 25684
rect 3337 25661 3423 25684
rect 7169 25724 7255 25747
rect 7337 25724 7423 25747
rect 7169 25684 7194 25724
rect 7194 25684 7234 25724
rect 7234 25684 7255 25724
rect 7337 25684 7358 25724
rect 7358 25684 7398 25724
rect 7398 25684 7423 25724
rect 7169 25661 7255 25684
rect 7337 25661 7423 25684
rect 11169 25724 11255 25747
rect 11337 25724 11423 25747
rect 11169 25684 11194 25724
rect 11194 25684 11234 25724
rect 11234 25684 11255 25724
rect 11337 25684 11358 25724
rect 11358 25684 11398 25724
rect 11398 25684 11423 25724
rect 11169 25661 11255 25684
rect 11337 25661 11423 25684
rect 15169 25724 15255 25747
rect 15337 25724 15423 25747
rect 15169 25684 15194 25724
rect 15194 25684 15234 25724
rect 15234 25684 15255 25724
rect 15337 25684 15358 25724
rect 15358 25684 15398 25724
rect 15398 25684 15423 25724
rect 15169 25661 15255 25684
rect 15337 25661 15423 25684
rect 19169 25724 19255 25747
rect 19337 25724 19423 25747
rect 19169 25684 19194 25724
rect 19194 25684 19234 25724
rect 19234 25684 19255 25724
rect 19337 25684 19358 25724
rect 19358 25684 19398 25724
rect 19398 25684 19423 25724
rect 19169 25661 19255 25684
rect 19337 25661 19423 25684
rect 23169 25724 23255 25747
rect 23337 25724 23423 25747
rect 23169 25684 23194 25724
rect 23194 25684 23234 25724
rect 23234 25684 23255 25724
rect 23337 25684 23358 25724
rect 23358 25684 23398 25724
rect 23398 25684 23423 25724
rect 23169 25661 23255 25684
rect 23337 25661 23423 25684
rect 27169 25724 27255 25747
rect 27337 25724 27423 25747
rect 27169 25684 27194 25724
rect 27194 25684 27234 25724
rect 27234 25684 27255 25724
rect 27337 25684 27358 25724
rect 27358 25684 27398 25724
rect 27398 25684 27423 25724
rect 27169 25661 27255 25684
rect 27337 25661 27423 25684
rect 31169 25724 31255 25747
rect 31337 25724 31423 25747
rect 31169 25684 31194 25724
rect 31194 25684 31234 25724
rect 31234 25684 31255 25724
rect 31337 25684 31358 25724
rect 31358 25684 31398 25724
rect 31398 25684 31423 25724
rect 31169 25661 31255 25684
rect 31337 25661 31423 25684
rect 35169 25724 35255 25747
rect 35337 25724 35423 25747
rect 35169 25684 35194 25724
rect 35194 25684 35234 25724
rect 35234 25684 35255 25724
rect 35337 25684 35358 25724
rect 35358 25684 35398 25724
rect 35398 25684 35423 25724
rect 35169 25661 35255 25684
rect 35337 25661 35423 25684
rect 39169 25724 39255 25747
rect 39337 25724 39423 25747
rect 39169 25684 39194 25724
rect 39194 25684 39234 25724
rect 39234 25684 39255 25724
rect 39337 25684 39358 25724
rect 39358 25684 39398 25724
rect 39398 25684 39423 25724
rect 39169 25661 39255 25684
rect 39337 25661 39423 25684
rect 43169 25724 43255 25747
rect 43337 25724 43423 25747
rect 43169 25684 43194 25724
rect 43194 25684 43234 25724
rect 43234 25684 43255 25724
rect 43337 25684 43358 25724
rect 43358 25684 43398 25724
rect 43398 25684 43423 25724
rect 43169 25661 43255 25684
rect 43337 25661 43423 25684
rect 47169 25724 47255 25747
rect 47337 25724 47423 25747
rect 47169 25684 47194 25724
rect 47194 25684 47234 25724
rect 47234 25684 47255 25724
rect 47337 25684 47358 25724
rect 47358 25684 47398 25724
rect 47398 25684 47423 25724
rect 47169 25661 47255 25684
rect 47337 25661 47423 25684
rect 51169 25724 51255 25747
rect 51337 25724 51423 25747
rect 51169 25684 51194 25724
rect 51194 25684 51234 25724
rect 51234 25684 51255 25724
rect 51337 25684 51358 25724
rect 51358 25684 51398 25724
rect 51398 25684 51423 25724
rect 51169 25661 51255 25684
rect 51337 25661 51423 25684
rect 55169 25724 55255 25747
rect 55337 25724 55423 25747
rect 55169 25684 55194 25724
rect 55194 25684 55234 25724
rect 55234 25684 55255 25724
rect 55337 25684 55358 25724
rect 55358 25684 55398 25724
rect 55398 25684 55423 25724
rect 55169 25661 55255 25684
rect 55337 25661 55423 25684
rect 59169 25724 59255 25747
rect 59337 25724 59423 25747
rect 59169 25684 59194 25724
rect 59194 25684 59234 25724
rect 59234 25684 59255 25724
rect 59337 25684 59358 25724
rect 59358 25684 59398 25724
rect 59398 25684 59423 25724
rect 59169 25661 59255 25684
rect 59337 25661 59423 25684
rect 63169 25724 63255 25747
rect 63337 25724 63423 25747
rect 63169 25684 63194 25724
rect 63194 25684 63234 25724
rect 63234 25684 63255 25724
rect 63337 25684 63358 25724
rect 63358 25684 63398 25724
rect 63398 25684 63423 25724
rect 63169 25661 63255 25684
rect 63337 25661 63423 25684
rect 67169 25724 67255 25747
rect 67337 25724 67423 25747
rect 67169 25684 67194 25724
rect 67194 25684 67234 25724
rect 67234 25684 67255 25724
rect 67337 25684 67358 25724
rect 67358 25684 67398 25724
rect 67398 25684 67423 25724
rect 67169 25661 67255 25684
rect 67337 25661 67423 25684
rect 86469 25325 86555 25411
rect 4409 24968 4495 24991
rect 4577 24968 4663 24991
rect 4409 24928 4434 24968
rect 4434 24928 4474 24968
rect 4474 24928 4495 24968
rect 4577 24928 4598 24968
rect 4598 24928 4638 24968
rect 4638 24928 4663 24968
rect 4409 24905 4495 24928
rect 4577 24905 4663 24928
rect 8409 24968 8495 24991
rect 8577 24968 8663 24991
rect 8409 24928 8434 24968
rect 8434 24928 8474 24968
rect 8474 24928 8495 24968
rect 8577 24928 8598 24968
rect 8598 24928 8638 24968
rect 8638 24928 8663 24968
rect 8409 24905 8495 24928
rect 8577 24905 8663 24928
rect 12409 24968 12495 24991
rect 12577 24968 12663 24991
rect 12409 24928 12434 24968
rect 12434 24928 12474 24968
rect 12474 24928 12495 24968
rect 12577 24928 12598 24968
rect 12598 24928 12638 24968
rect 12638 24928 12663 24968
rect 12409 24905 12495 24928
rect 12577 24905 12663 24928
rect 16409 24968 16495 24991
rect 16577 24968 16663 24991
rect 16409 24928 16434 24968
rect 16434 24928 16474 24968
rect 16474 24928 16495 24968
rect 16577 24928 16598 24968
rect 16598 24928 16638 24968
rect 16638 24928 16663 24968
rect 16409 24905 16495 24928
rect 16577 24905 16663 24928
rect 20409 24968 20495 24991
rect 20577 24968 20663 24991
rect 20409 24928 20434 24968
rect 20434 24928 20474 24968
rect 20474 24928 20495 24968
rect 20577 24928 20598 24968
rect 20598 24928 20638 24968
rect 20638 24928 20663 24968
rect 20409 24905 20495 24928
rect 20577 24905 20663 24928
rect 24409 24968 24495 24991
rect 24577 24968 24663 24991
rect 24409 24928 24434 24968
rect 24434 24928 24474 24968
rect 24474 24928 24495 24968
rect 24577 24928 24598 24968
rect 24598 24928 24638 24968
rect 24638 24928 24663 24968
rect 24409 24905 24495 24928
rect 24577 24905 24663 24928
rect 28409 24968 28495 24991
rect 28577 24968 28663 24991
rect 28409 24928 28434 24968
rect 28434 24928 28474 24968
rect 28474 24928 28495 24968
rect 28577 24928 28598 24968
rect 28598 24928 28638 24968
rect 28638 24928 28663 24968
rect 28409 24905 28495 24928
rect 28577 24905 28663 24928
rect 32409 24968 32495 24991
rect 32577 24968 32663 24991
rect 32409 24928 32434 24968
rect 32434 24928 32474 24968
rect 32474 24928 32495 24968
rect 32577 24928 32598 24968
rect 32598 24928 32638 24968
rect 32638 24928 32663 24968
rect 32409 24905 32495 24928
rect 32577 24905 32663 24928
rect 36409 24968 36495 24991
rect 36577 24968 36663 24991
rect 36409 24928 36434 24968
rect 36434 24928 36474 24968
rect 36474 24928 36495 24968
rect 36577 24928 36598 24968
rect 36598 24928 36638 24968
rect 36638 24928 36663 24968
rect 36409 24905 36495 24928
rect 36577 24905 36663 24928
rect 40409 24968 40495 24991
rect 40577 24968 40663 24991
rect 40409 24928 40434 24968
rect 40434 24928 40474 24968
rect 40474 24928 40495 24968
rect 40577 24928 40598 24968
rect 40598 24928 40638 24968
rect 40638 24928 40663 24968
rect 40409 24905 40495 24928
rect 40577 24905 40663 24928
rect 44409 24968 44495 24991
rect 44577 24968 44663 24991
rect 44409 24928 44434 24968
rect 44434 24928 44474 24968
rect 44474 24928 44495 24968
rect 44577 24928 44598 24968
rect 44598 24928 44638 24968
rect 44638 24928 44663 24968
rect 44409 24905 44495 24928
rect 44577 24905 44663 24928
rect 48409 24968 48495 24991
rect 48577 24968 48663 24991
rect 48409 24928 48434 24968
rect 48434 24928 48474 24968
rect 48474 24928 48495 24968
rect 48577 24928 48598 24968
rect 48598 24928 48638 24968
rect 48638 24928 48663 24968
rect 48409 24905 48495 24928
rect 48577 24905 48663 24928
rect 52409 24968 52495 24991
rect 52577 24968 52663 24991
rect 52409 24928 52434 24968
rect 52434 24928 52474 24968
rect 52474 24928 52495 24968
rect 52577 24928 52598 24968
rect 52598 24928 52638 24968
rect 52638 24928 52663 24968
rect 52409 24905 52495 24928
rect 52577 24905 52663 24928
rect 56409 24968 56495 24991
rect 56577 24968 56663 24991
rect 56409 24928 56434 24968
rect 56434 24928 56474 24968
rect 56474 24928 56495 24968
rect 56577 24928 56598 24968
rect 56598 24928 56638 24968
rect 56638 24928 56663 24968
rect 56409 24905 56495 24928
rect 56577 24905 56663 24928
rect 60409 24968 60495 24991
rect 60577 24968 60663 24991
rect 60409 24928 60434 24968
rect 60434 24928 60474 24968
rect 60474 24928 60495 24968
rect 60577 24928 60598 24968
rect 60598 24928 60638 24968
rect 60638 24928 60663 24968
rect 60409 24905 60495 24928
rect 60577 24905 60663 24928
rect 64409 24968 64495 24991
rect 64577 24968 64663 24991
rect 64409 24928 64434 24968
rect 64434 24928 64474 24968
rect 64474 24928 64495 24968
rect 64577 24928 64598 24968
rect 64598 24928 64638 24968
rect 64638 24928 64663 24968
rect 64409 24905 64495 24928
rect 64577 24905 64663 24928
rect 68409 24968 68495 24991
rect 68577 24968 68663 24991
rect 68409 24928 68434 24968
rect 68434 24928 68474 24968
rect 68474 24928 68495 24968
rect 68577 24928 68598 24968
rect 68598 24928 68638 24968
rect 68638 24928 68663 24968
rect 68409 24905 68495 24928
rect 68577 24905 68663 24928
rect 3169 24212 3255 24235
rect 3337 24212 3423 24235
rect 3169 24172 3194 24212
rect 3194 24172 3234 24212
rect 3234 24172 3255 24212
rect 3337 24172 3358 24212
rect 3358 24172 3398 24212
rect 3398 24172 3423 24212
rect 3169 24149 3255 24172
rect 3337 24149 3423 24172
rect 7169 24212 7255 24235
rect 7337 24212 7423 24235
rect 7169 24172 7194 24212
rect 7194 24172 7234 24212
rect 7234 24172 7255 24212
rect 7337 24172 7358 24212
rect 7358 24172 7398 24212
rect 7398 24172 7423 24212
rect 7169 24149 7255 24172
rect 7337 24149 7423 24172
rect 11169 24212 11255 24235
rect 11337 24212 11423 24235
rect 11169 24172 11194 24212
rect 11194 24172 11234 24212
rect 11234 24172 11255 24212
rect 11337 24172 11358 24212
rect 11358 24172 11398 24212
rect 11398 24172 11423 24212
rect 11169 24149 11255 24172
rect 11337 24149 11423 24172
rect 15169 24212 15255 24235
rect 15337 24212 15423 24235
rect 15169 24172 15194 24212
rect 15194 24172 15234 24212
rect 15234 24172 15255 24212
rect 15337 24172 15358 24212
rect 15358 24172 15398 24212
rect 15398 24172 15423 24212
rect 15169 24149 15255 24172
rect 15337 24149 15423 24172
rect 19169 24212 19255 24235
rect 19337 24212 19423 24235
rect 19169 24172 19194 24212
rect 19194 24172 19234 24212
rect 19234 24172 19255 24212
rect 19337 24172 19358 24212
rect 19358 24172 19398 24212
rect 19398 24172 19423 24212
rect 19169 24149 19255 24172
rect 19337 24149 19423 24172
rect 23169 24212 23255 24235
rect 23337 24212 23423 24235
rect 23169 24172 23194 24212
rect 23194 24172 23234 24212
rect 23234 24172 23255 24212
rect 23337 24172 23358 24212
rect 23358 24172 23398 24212
rect 23398 24172 23423 24212
rect 23169 24149 23255 24172
rect 23337 24149 23423 24172
rect 27169 24212 27255 24235
rect 27337 24212 27423 24235
rect 27169 24172 27194 24212
rect 27194 24172 27234 24212
rect 27234 24172 27255 24212
rect 27337 24172 27358 24212
rect 27358 24172 27398 24212
rect 27398 24172 27423 24212
rect 27169 24149 27255 24172
rect 27337 24149 27423 24172
rect 31169 24212 31255 24235
rect 31337 24212 31423 24235
rect 31169 24172 31194 24212
rect 31194 24172 31234 24212
rect 31234 24172 31255 24212
rect 31337 24172 31358 24212
rect 31358 24172 31398 24212
rect 31398 24172 31423 24212
rect 31169 24149 31255 24172
rect 31337 24149 31423 24172
rect 35169 24212 35255 24235
rect 35337 24212 35423 24235
rect 35169 24172 35194 24212
rect 35194 24172 35234 24212
rect 35234 24172 35255 24212
rect 35337 24172 35358 24212
rect 35358 24172 35398 24212
rect 35398 24172 35423 24212
rect 35169 24149 35255 24172
rect 35337 24149 35423 24172
rect 39169 24212 39255 24235
rect 39337 24212 39423 24235
rect 39169 24172 39194 24212
rect 39194 24172 39234 24212
rect 39234 24172 39255 24212
rect 39337 24172 39358 24212
rect 39358 24172 39398 24212
rect 39398 24172 39423 24212
rect 39169 24149 39255 24172
rect 39337 24149 39423 24172
rect 43169 24212 43255 24235
rect 43337 24212 43423 24235
rect 43169 24172 43194 24212
rect 43194 24172 43234 24212
rect 43234 24172 43255 24212
rect 43337 24172 43358 24212
rect 43358 24172 43398 24212
rect 43398 24172 43423 24212
rect 43169 24149 43255 24172
rect 43337 24149 43423 24172
rect 47169 24212 47255 24235
rect 47337 24212 47423 24235
rect 47169 24172 47194 24212
rect 47194 24172 47234 24212
rect 47234 24172 47255 24212
rect 47337 24172 47358 24212
rect 47358 24172 47398 24212
rect 47398 24172 47423 24212
rect 47169 24149 47255 24172
rect 47337 24149 47423 24172
rect 51169 24212 51255 24235
rect 51337 24212 51423 24235
rect 51169 24172 51194 24212
rect 51194 24172 51234 24212
rect 51234 24172 51255 24212
rect 51337 24172 51358 24212
rect 51358 24172 51398 24212
rect 51398 24172 51423 24212
rect 51169 24149 51255 24172
rect 51337 24149 51423 24172
rect 55169 24212 55255 24235
rect 55337 24212 55423 24235
rect 55169 24172 55194 24212
rect 55194 24172 55234 24212
rect 55234 24172 55255 24212
rect 55337 24172 55358 24212
rect 55358 24172 55398 24212
rect 55398 24172 55423 24212
rect 55169 24149 55255 24172
rect 55337 24149 55423 24172
rect 59169 24212 59255 24235
rect 59337 24212 59423 24235
rect 59169 24172 59194 24212
rect 59194 24172 59234 24212
rect 59234 24172 59255 24212
rect 59337 24172 59358 24212
rect 59358 24172 59398 24212
rect 59398 24172 59423 24212
rect 59169 24149 59255 24172
rect 59337 24149 59423 24172
rect 63169 24212 63255 24235
rect 63337 24212 63423 24235
rect 63169 24172 63194 24212
rect 63194 24172 63234 24212
rect 63234 24172 63255 24212
rect 63337 24172 63358 24212
rect 63358 24172 63398 24212
rect 63398 24172 63423 24212
rect 63169 24149 63255 24172
rect 63337 24149 63423 24172
rect 67169 24212 67255 24235
rect 67337 24212 67423 24235
rect 67169 24172 67194 24212
rect 67194 24172 67234 24212
rect 67234 24172 67255 24212
rect 67337 24172 67358 24212
rect 67358 24172 67398 24212
rect 67398 24172 67423 24212
rect 67169 24149 67255 24172
rect 67337 24149 67423 24172
rect 71169 24212 71255 24235
rect 71337 24212 71423 24235
rect 71169 24172 71194 24212
rect 71194 24172 71234 24212
rect 71234 24172 71255 24212
rect 71337 24172 71358 24212
rect 71358 24172 71398 24212
rect 71398 24172 71423 24212
rect 71169 24149 71255 24172
rect 71337 24149 71423 24172
rect 75169 24212 75255 24235
rect 75337 24212 75423 24235
rect 75169 24172 75194 24212
rect 75194 24172 75234 24212
rect 75234 24172 75255 24212
rect 75337 24172 75358 24212
rect 75358 24172 75398 24212
rect 75398 24172 75423 24212
rect 75169 24149 75255 24172
rect 75337 24149 75423 24172
rect 79169 24212 79255 24235
rect 79337 24212 79423 24235
rect 79169 24172 79194 24212
rect 79194 24172 79234 24212
rect 79234 24172 79255 24212
rect 79337 24172 79358 24212
rect 79358 24172 79398 24212
rect 79398 24172 79423 24212
rect 79169 24149 79255 24172
rect 79337 24149 79423 24172
rect 83169 24212 83255 24235
rect 83337 24212 83423 24235
rect 83169 24172 83194 24212
rect 83194 24172 83234 24212
rect 83234 24172 83255 24212
rect 83337 24172 83358 24212
rect 83358 24172 83398 24212
rect 83398 24172 83423 24212
rect 83169 24149 83255 24172
rect 83337 24149 83423 24172
rect 87169 24212 87255 24235
rect 87337 24212 87423 24235
rect 87169 24172 87194 24212
rect 87194 24172 87234 24212
rect 87234 24172 87255 24212
rect 87337 24172 87358 24212
rect 87358 24172 87398 24212
rect 87398 24172 87423 24212
rect 87169 24149 87255 24172
rect 87337 24149 87423 24172
rect 91169 24212 91255 24235
rect 91337 24212 91423 24235
rect 91169 24172 91194 24212
rect 91194 24172 91234 24212
rect 91234 24172 91255 24212
rect 91337 24172 91358 24212
rect 91358 24172 91398 24212
rect 91398 24172 91423 24212
rect 91169 24149 91255 24172
rect 91337 24149 91423 24172
rect 95169 24212 95255 24235
rect 95337 24212 95423 24235
rect 95169 24172 95194 24212
rect 95194 24172 95234 24212
rect 95234 24172 95255 24212
rect 95337 24172 95358 24212
rect 95358 24172 95398 24212
rect 95398 24172 95423 24212
rect 95169 24149 95255 24172
rect 95337 24149 95423 24172
rect 99169 24212 99255 24235
rect 99337 24212 99423 24235
rect 99169 24172 99194 24212
rect 99194 24172 99234 24212
rect 99234 24172 99255 24212
rect 99337 24172 99358 24212
rect 99358 24172 99398 24212
rect 99398 24172 99423 24212
rect 99169 24149 99255 24172
rect 99337 24149 99423 24172
rect 4409 23456 4495 23479
rect 4577 23456 4663 23479
rect 4409 23416 4434 23456
rect 4434 23416 4474 23456
rect 4474 23416 4495 23456
rect 4577 23416 4598 23456
rect 4598 23416 4638 23456
rect 4638 23416 4663 23456
rect 4409 23393 4495 23416
rect 4577 23393 4663 23416
rect 8409 23456 8495 23479
rect 8577 23456 8663 23479
rect 8409 23416 8434 23456
rect 8434 23416 8474 23456
rect 8474 23416 8495 23456
rect 8577 23416 8598 23456
rect 8598 23416 8638 23456
rect 8638 23416 8663 23456
rect 8409 23393 8495 23416
rect 8577 23393 8663 23416
rect 12409 23456 12495 23479
rect 12577 23456 12663 23479
rect 12409 23416 12434 23456
rect 12434 23416 12474 23456
rect 12474 23416 12495 23456
rect 12577 23416 12598 23456
rect 12598 23416 12638 23456
rect 12638 23416 12663 23456
rect 12409 23393 12495 23416
rect 12577 23393 12663 23416
rect 16409 23456 16495 23479
rect 16577 23456 16663 23479
rect 16409 23416 16434 23456
rect 16434 23416 16474 23456
rect 16474 23416 16495 23456
rect 16577 23416 16598 23456
rect 16598 23416 16638 23456
rect 16638 23416 16663 23456
rect 16409 23393 16495 23416
rect 16577 23393 16663 23416
rect 20409 23456 20495 23479
rect 20577 23456 20663 23479
rect 20409 23416 20434 23456
rect 20434 23416 20474 23456
rect 20474 23416 20495 23456
rect 20577 23416 20598 23456
rect 20598 23416 20638 23456
rect 20638 23416 20663 23456
rect 20409 23393 20495 23416
rect 20577 23393 20663 23416
rect 24409 23456 24495 23479
rect 24577 23456 24663 23479
rect 24409 23416 24434 23456
rect 24434 23416 24474 23456
rect 24474 23416 24495 23456
rect 24577 23416 24598 23456
rect 24598 23416 24638 23456
rect 24638 23416 24663 23456
rect 24409 23393 24495 23416
rect 24577 23393 24663 23416
rect 28409 23456 28495 23479
rect 28577 23456 28663 23479
rect 28409 23416 28434 23456
rect 28434 23416 28474 23456
rect 28474 23416 28495 23456
rect 28577 23416 28598 23456
rect 28598 23416 28638 23456
rect 28638 23416 28663 23456
rect 28409 23393 28495 23416
rect 28577 23393 28663 23416
rect 32409 23456 32495 23479
rect 32577 23456 32663 23479
rect 32409 23416 32434 23456
rect 32434 23416 32474 23456
rect 32474 23416 32495 23456
rect 32577 23416 32598 23456
rect 32598 23416 32638 23456
rect 32638 23416 32663 23456
rect 32409 23393 32495 23416
rect 32577 23393 32663 23416
rect 36409 23456 36495 23479
rect 36577 23456 36663 23479
rect 36409 23416 36434 23456
rect 36434 23416 36474 23456
rect 36474 23416 36495 23456
rect 36577 23416 36598 23456
rect 36598 23416 36638 23456
rect 36638 23416 36663 23456
rect 36409 23393 36495 23416
rect 36577 23393 36663 23416
rect 40409 23456 40495 23479
rect 40577 23456 40663 23479
rect 40409 23416 40434 23456
rect 40434 23416 40474 23456
rect 40474 23416 40495 23456
rect 40577 23416 40598 23456
rect 40598 23416 40638 23456
rect 40638 23416 40663 23456
rect 40409 23393 40495 23416
rect 40577 23393 40663 23416
rect 44409 23456 44495 23479
rect 44577 23456 44663 23479
rect 44409 23416 44434 23456
rect 44434 23416 44474 23456
rect 44474 23416 44495 23456
rect 44577 23416 44598 23456
rect 44598 23416 44638 23456
rect 44638 23416 44663 23456
rect 44409 23393 44495 23416
rect 44577 23393 44663 23416
rect 48409 23456 48495 23479
rect 48577 23456 48663 23479
rect 48409 23416 48434 23456
rect 48434 23416 48474 23456
rect 48474 23416 48495 23456
rect 48577 23416 48598 23456
rect 48598 23416 48638 23456
rect 48638 23416 48663 23456
rect 48409 23393 48495 23416
rect 48577 23393 48663 23416
rect 52409 23456 52495 23479
rect 52577 23456 52663 23479
rect 52409 23416 52434 23456
rect 52434 23416 52474 23456
rect 52474 23416 52495 23456
rect 52577 23416 52598 23456
rect 52598 23416 52638 23456
rect 52638 23416 52663 23456
rect 52409 23393 52495 23416
rect 52577 23393 52663 23416
rect 56409 23456 56495 23479
rect 56577 23456 56663 23479
rect 56409 23416 56434 23456
rect 56434 23416 56474 23456
rect 56474 23416 56495 23456
rect 56577 23416 56598 23456
rect 56598 23416 56638 23456
rect 56638 23416 56663 23456
rect 56409 23393 56495 23416
rect 56577 23393 56663 23416
rect 60409 23456 60495 23479
rect 60577 23456 60663 23479
rect 60409 23416 60434 23456
rect 60434 23416 60474 23456
rect 60474 23416 60495 23456
rect 60577 23416 60598 23456
rect 60598 23416 60638 23456
rect 60638 23416 60663 23456
rect 60409 23393 60495 23416
rect 60577 23393 60663 23416
rect 64409 23456 64495 23479
rect 64577 23456 64663 23479
rect 64409 23416 64434 23456
rect 64434 23416 64474 23456
rect 64474 23416 64495 23456
rect 64577 23416 64598 23456
rect 64598 23416 64638 23456
rect 64638 23416 64663 23456
rect 64409 23393 64495 23416
rect 64577 23393 64663 23416
rect 68409 23456 68495 23479
rect 68577 23456 68663 23479
rect 68409 23416 68434 23456
rect 68434 23416 68474 23456
rect 68474 23416 68495 23456
rect 68577 23416 68598 23456
rect 68598 23416 68638 23456
rect 68638 23416 68663 23456
rect 68409 23393 68495 23416
rect 68577 23393 68663 23416
rect 72409 23456 72495 23479
rect 72577 23456 72663 23479
rect 72409 23416 72434 23456
rect 72434 23416 72474 23456
rect 72474 23416 72495 23456
rect 72577 23416 72598 23456
rect 72598 23416 72638 23456
rect 72638 23416 72663 23456
rect 72409 23393 72495 23416
rect 72577 23393 72663 23416
rect 76409 23456 76495 23479
rect 76577 23456 76663 23479
rect 76409 23416 76434 23456
rect 76434 23416 76474 23456
rect 76474 23416 76495 23456
rect 76577 23416 76598 23456
rect 76598 23416 76638 23456
rect 76638 23416 76663 23456
rect 76409 23393 76495 23416
rect 76577 23393 76663 23416
rect 80409 23456 80495 23479
rect 80577 23456 80663 23479
rect 80409 23416 80434 23456
rect 80434 23416 80474 23456
rect 80474 23416 80495 23456
rect 80577 23416 80598 23456
rect 80598 23416 80638 23456
rect 80638 23416 80663 23456
rect 80409 23393 80495 23416
rect 80577 23393 80663 23416
rect 84409 23456 84495 23479
rect 84577 23456 84663 23479
rect 84409 23416 84434 23456
rect 84434 23416 84474 23456
rect 84474 23416 84495 23456
rect 84577 23416 84598 23456
rect 84598 23416 84638 23456
rect 84638 23416 84663 23456
rect 84409 23393 84495 23416
rect 84577 23393 84663 23416
rect 88409 23456 88495 23479
rect 88577 23456 88663 23479
rect 88409 23416 88434 23456
rect 88434 23416 88474 23456
rect 88474 23416 88495 23456
rect 88577 23416 88598 23456
rect 88598 23416 88638 23456
rect 88638 23416 88663 23456
rect 88409 23393 88495 23416
rect 88577 23393 88663 23416
rect 92409 23456 92495 23479
rect 92577 23456 92663 23479
rect 92409 23416 92434 23456
rect 92434 23416 92474 23456
rect 92474 23416 92495 23456
rect 92577 23416 92598 23456
rect 92598 23416 92638 23456
rect 92638 23416 92663 23456
rect 92409 23393 92495 23416
rect 92577 23393 92663 23416
rect 96409 23456 96495 23479
rect 96577 23456 96663 23479
rect 96409 23416 96434 23456
rect 96434 23416 96474 23456
rect 96474 23416 96495 23456
rect 96577 23416 96598 23456
rect 96598 23416 96638 23456
rect 96638 23416 96663 23456
rect 96409 23393 96495 23416
rect 96577 23393 96663 23416
rect 3169 22700 3255 22723
rect 3337 22700 3423 22723
rect 3169 22660 3194 22700
rect 3194 22660 3234 22700
rect 3234 22660 3255 22700
rect 3337 22660 3358 22700
rect 3358 22660 3398 22700
rect 3398 22660 3423 22700
rect 3169 22637 3255 22660
rect 3337 22637 3423 22660
rect 7169 22700 7255 22723
rect 7337 22700 7423 22723
rect 7169 22660 7194 22700
rect 7194 22660 7234 22700
rect 7234 22660 7255 22700
rect 7337 22660 7358 22700
rect 7358 22660 7398 22700
rect 7398 22660 7423 22700
rect 7169 22637 7255 22660
rect 7337 22637 7423 22660
rect 11169 22700 11255 22723
rect 11337 22700 11423 22723
rect 11169 22660 11194 22700
rect 11194 22660 11234 22700
rect 11234 22660 11255 22700
rect 11337 22660 11358 22700
rect 11358 22660 11398 22700
rect 11398 22660 11423 22700
rect 11169 22637 11255 22660
rect 11337 22637 11423 22660
rect 15169 22700 15255 22723
rect 15337 22700 15423 22723
rect 15169 22660 15194 22700
rect 15194 22660 15234 22700
rect 15234 22660 15255 22700
rect 15337 22660 15358 22700
rect 15358 22660 15398 22700
rect 15398 22660 15423 22700
rect 15169 22637 15255 22660
rect 15337 22637 15423 22660
rect 19169 22700 19255 22723
rect 19337 22700 19423 22723
rect 19169 22660 19194 22700
rect 19194 22660 19234 22700
rect 19234 22660 19255 22700
rect 19337 22660 19358 22700
rect 19358 22660 19398 22700
rect 19398 22660 19423 22700
rect 19169 22637 19255 22660
rect 19337 22637 19423 22660
rect 23169 22700 23255 22723
rect 23337 22700 23423 22723
rect 23169 22660 23194 22700
rect 23194 22660 23234 22700
rect 23234 22660 23255 22700
rect 23337 22660 23358 22700
rect 23358 22660 23398 22700
rect 23398 22660 23423 22700
rect 23169 22637 23255 22660
rect 23337 22637 23423 22660
rect 27169 22700 27255 22723
rect 27337 22700 27423 22723
rect 27169 22660 27194 22700
rect 27194 22660 27234 22700
rect 27234 22660 27255 22700
rect 27337 22660 27358 22700
rect 27358 22660 27398 22700
rect 27398 22660 27423 22700
rect 27169 22637 27255 22660
rect 27337 22637 27423 22660
rect 31169 22700 31255 22723
rect 31337 22700 31423 22723
rect 31169 22660 31194 22700
rect 31194 22660 31234 22700
rect 31234 22660 31255 22700
rect 31337 22660 31358 22700
rect 31358 22660 31398 22700
rect 31398 22660 31423 22700
rect 31169 22637 31255 22660
rect 31337 22637 31423 22660
rect 35169 22700 35255 22723
rect 35337 22700 35423 22723
rect 35169 22660 35194 22700
rect 35194 22660 35234 22700
rect 35234 22660 35255 22700
rect 35337 22660 35358 22700
rect 35358 22660 35398 22700
rect 35398 22660 35423 22700
rect 35169 22637 35255 22660
rect 35337 22637 35423 22660
rect 39169 22700 39255 22723
rect 39337 22700 39423 22723
rect 39169 22660 39194 22700
rect 39194 22660 39234 22700
rect 39234 22660 39255 22700
rect 39337 22660 39358 22700
rect 39358 22660 39398 22700
rect 39398 22660 39423 22700
rect 39169 22637 39255 22660
rect 39337 22637 39423 22660
rect 43169 22700 43255 22723
rect 43337 22700 43423 22723
rect 43169 22660 43194 22700
rect 43194 22660 43234 22700
rect 43234 22660 43255 22700
rect 43337 22660 43358 22700
rect 43358 22660 43398 22700
rect 43398 22660 43423 22700
rect 43169 22637 43255 22660
rect 43337 22637 43423 22660
rect 47169 22700 47255 22723
rect 47337 22700 47423 22723
rect 47169 22660 47194 22700
rect 47194 22660 47234 22700
rect 47234 22660 47255 22700
rect 47337 22660 47358 22700
rect 47358 22660 47398 22700
rect 47398 22660 47423 22700
rect 47169 22637 47255 22660
rect 47337 22637 47423 22660
rect 51169 22700 51255 22723
rect 51337 22700 51423 22723
rect 51169 22660 51194 22700
rect 51194 22660 51234 22700
rect 51234 22660 51255 22700
rect 51337 22660 51358 22700
rect 51358 22660 51398 22700
rect 51398 22660 51423 22700
rect 51169 22637 51255 22660
rect 51337 22637 51423 22660
rect 55169 22700 55255 22723
rect 55337 22700 55423 22723
rect 55169 22660 55194 22700
rect 55194 22660 55234 22700
rect 55234 22660 55255 22700
rect 55337 22660 55358 22700
rect 55358 22660 55398 22700
rect 55398 22660 55423 22700
rect 55169 22637 55255 22660
rect 55337 22637 55423 22660
rect 59169 22700 59255 22723
rect 59337 22700 59423 22723
rect 59169 22660 59194 22700
rect 59194 22660 59234 22700
rect 59234 22660 59255 22700
rect 59337 22660 59358 22700
rect 59358 22660 59398 22700
rect 59398 22660 59423 22700
rect 59169 22637 59255 22660
rect 59337 22637 59423 22660
rect 63169 22700 63255 22723
rect 63337 22700 63423 22723
rect 63169 22660 63194 22700
rect 63194 22660 63234 22700
rect 63234 22660 63255 22700
rect 63337 22660 63358 22700
rect 63358 22660 63398 22700
rect 63398 22660 63423 22700
rect 63169 22637 63255 22660
rect 63337 22637 63423 22660
rect 67169 22700 67255 22723
rect 67337 22700 67423 22723
rect 67169 22660 67194 22700
rect 67194 22660 67234 22700
rect 67234 22660 67255 22700
rect 67337 22660 67358 22700
rect 67358 22660 67398 22700
rect 67398 22660 67423 22700
rect 67169 22637 67255 22660
rect 67337 22637 67423 22660
rect 71169 22700 71255 22723
rect 71337 22700 71423 22723
rect 71169 22660 71194 22700
rect 71194 22660 71234 22700
rect 71234 22660 71255 22700
rect 71337 22660 71358 22700
rect 71358 22660 71398 22700
rect 71398 22660 71423 22700
rect 71169 22637 71255 22660
rect 71337 22637 71423 22660
rect 75169 22700 75255 22723
rect 75337 22700 75423 22723
rect 75169 22660 75194 22700
rect 75194 22660 75234 22700
rect 75234 22660 75255 22700
rect 75337 22660 75358 22700
rect 75358 22660 75398 22700
rect 75398 22660 75423 22700
rect 75169 22637 75255 22660
rect 75337 22637 75423 22660
rect 79169 22700 79255 22723
rect 79337 22700 79423 22723
rect 79169 22660 79194 22700
rect 79194 22660 79234 22700
rect 79234 22660 79255 22700
rect 79337 22660 79358 22700
rect 79358 22660 79398 22700
rect 79398 22660 79423 22700
rect 79169 22637 79255 22660
rect 79337 22637 79423 22660
rect 83169 22700 83255 22723
rect 83337 22700 83423 22723
rect 83169 22660 83194 22700
rect 83194 22660 83234 22700
rect 83234 22660 83255 22700
rect 83337 22660 83358 22700
rect 83358 22660 83398 22700
rect 83398 22660 83423 22700
rect 83169 22637 83255 22660
rect 83337 22637 83423 22660
rect 87169 22700 87255 22723
rect 87337 22700 87423 22723
rect 87169 22660 87194 22700
rect 87194 22660 87234 22700
rect 87234 22660 87255 22700
rect 87337 22660 87358 22700
rect 87358 22660 87398 22700
rect 87398 22660 87423 22700
rect 87169 22637 87255 22660
rect 87337 22637 87423 22660
rect 91169 22700 91255 22723
rect 91337 22700 91423 22723
rect 91169 22660 91194 22700
rect 91194 22660 91234 22700
rect 91234 22660 91255 22700
rect 91337 22660 91358 22700
rect 91358 22660 91398 22700
rect 91398 22660 91423 22700
rect 91169 22637 91255 22660
rect 91337 22637 91423 22660
rect 95169 22700 95255 22723
rect 95337 22700 95423 22723
rect 95169 22660 95194 22700
rect 95194 22660 95234 22700
rect 95234 22660 95255 22700
rect 95337 22660 95358 22700
rect 95358 22660 95398 22700
rect 95398 22660 95423 22700
rect 95169 22637 95255 22660
rect 95337 22637 95423 22660
rect 99169 22700 99255 22723
rect 99337 22700 99423 22723
rect 99169 22660 99194 22700
rect 99194 22660 99234 22700
rect 99234 22660 99255 22700
rect 99337 22660 99358 22700
rect 99358 22660 99398 22700
rect 99398 22660 99423 22700
rect 99169 22637 99255 22660
rect 99337 22637 99423 22660
rect 4409 21944 4495 21967
rect 4577 21944 4663 21967
rect 4409 21904 4434 21944
rect 4434 21904 4474 21944
rect 4474 21904 4495 21944
rect 4577 21904 4598 21944
rect 4598 21904 4638 21944
rect 4638 21904 4663 21944
rect 4409 21881 4495 21904
rect 4577 21881 4663 21904
rect 8409 21944 8495 21967
rect 8577 21944 8663 21967
rect 8409 21904 8434 21944
rect 8434 21904 8474 21944
rect 8474 21904 8495 21944
rect 8577 21904 8598 21944
rect 8598 21904 8638 21944
rect 8638 21904 8663 21944
rect 8409 21881 8495 21904
rect 8577 21881 8663 21904
rect 12409 21944 12495 21967
rect 12577 21944 12663 21967
rect 12409 21904 12434 21944
rect 12434 21904 12474 21944
rect 12474 21904 12495 21944
rect 12577 21904 12598 21944
rect 12598 21904 12638 21944
rect 12638 21904 12663 21944
rect 12409 21881 12495 21904
rect 12577 21881 12663 21904
rect 16409 21944 16495 21967
rect 16577 21944 16663 21967
rect 16409 21904 16434 21944
rect 16434 21904 16474 21944
rect 16474 21904 16495 21944
rect 16577 21904 16598 21944
rect 16598 21904 16638 21944
rect 16638 21904 16663 21944
rect 16409 21881 16495 21904
rect 16577 21881 16663 21904
rect 20409 21944 20495 21967
rect 20577 21944 20663 21967
rect 20409 21904 20434 21944
rect 20434 21904 20474 21944
rect 20474 21904 20495 21944
rect 20577 21904 20598 21944
rect 20598 21904 20638 21944
rect 20638 21904 20663 21944
rect 20409 21881 20495 21904
rect 20577 21881 20663 21904
rect 24409 21944 24495 21967
rect 24577 21944 24663 21967
rect 24409 21904 24434 21944
rect 24434 21904 24474 21944
rect 24474 21904 24495 21944
rect 24577 21904 24598 21944
rect 24598 21904 24638 21944
rect 24638 21904 24663 21944
rect 24409 21881 24495 21904
rect 24577 21881 24663 21904
rect 28409 21944 28495 21967
rect 28577 21944 28663 21967
rect 28409 21904 28434 21944
rect 28434 21904 28474 21944
rect 28474 21904 28495 21944
rect 28577 21904 28598 21944
rect 28598 21904 28638 21944
rect 28638 21904 28663 21944
rect 28409 21881 28495 21904
rect 28577 21881 28663 21904
rect 32409 21944 32495 21967
rect 32577 21944 32663 21967
rect 32409 21904 32434 21944
rect 32434 21904 32474 21944
rect 32474 21904 32495 21944
rect 32577 21904 32598 21944
rect 32598 21904 32638 21944
rect 32638 21904 32663 21944
rect 32409 21881 32495 21904
rect 32577 21881 32663 21904
rect 36409 21944 36495 21967
rect 36577 21944 36663 21967
rect 36409 21904 36434 21944
rect 36434 21904 36474 21944
rect 36474 21904 36495 21944
rect 36577 21904 36598 21944
rect 36598 21904 36638 21944
rect 36638 21904 36663 21944
rect 36409 21881 36495 21904
rect 36577 21881 36663 21904
rect 40409 21944 40495 21967
rect 40577 21944 40663 21967
rect 40409 21904 40434 21944
rect 40434 21904 40474 21944
rect 40474 21904 40495 21944
rect 40577 21904 40598 21944
rect 40598 21904 40638 21944
rect 40638 21904 40663 21944
rect 40409 21881 40495 21904
rect 40577 21881 40663 21904
rect 44409 21944 44495 21967
rect 44577 21944 44663 21967
rect 44409 21904 44434 21944
rect 44434 21904 44474 21944
rect 44474 21904 44495 21944
rect 44577 21904 44598 21944
rect 44598 21904 44638 21944
rect 44638 21904 44663 21944
rect 44409 21881 44495 21904
rect 44577 21881 44663 21904
rect 48409 21944 48495 21967
rect 48577 21944 48663 21967
rect 48409 21904 48434 21944
rect 48434 21904 48474 21944
rect 48474 21904 48495 21944
rect 48577 21904 48598 21944
rect 48598 21904 48638 21944
rect 48638 21904 48663 21944
rect 48409 21881 48495 21904
rect 48577 21881 48663 21904
rect 52409 21944 52495 21967
rect 52577 21944 52663 21967
rect 52409 21904 52434 21944
rect 52434 21904 52474 21944
rect 52474 21904 52495 21944
rect 52577 21904 52598 21944
rect 52598 21904 52638 21944
rect 52638 21904 52663 21944
rect 52409 21881 52495 21904
rect 52577 21881 52663 21904
rect 56409 21944 56495 21967
rect 56577 21944 56663 21967
rect 56409 21904 56434 21944
rect 56434 21904 56474 21944
rect 56474 21904 56495 21944
rect 56577 21904 56598 21944
rect 56598 21904 56638 21944
rect 56638 21904 56663 21944
rect 56409 21881 56495 21904
rect 56577 21881 56663 21904
rect 60409 21944 60495 21967
rect 60577 21944 60663 21967
rect 60409 21904 60434 21944
rect 60434 21904 60474 21944
rect 60474 21904 60495 21944
rect 60577 21904 60598 21944
rect 60598 21904 60638 21944
rect 60638 21904 60663 21944
rect 60409 21881 60495 21904
rect 60577 21881 60663 21904
rect 64409 21944 64495 21967
rect 64577 21944 64663 21967
rect 64409 21904 64434 21944
rect 64434 21904 64474 21944
rect 64474 21904 64495 21944
rect 64577 21904 64598 21944
rect 64598 21904 64638 21944
rect 64638 21904 64663 21944
rect 64409 21881 64495 21904
rect 64577 21881 64663 21904
rect 68409 21944 68495 21967
rect 68577 21944 68663 21967
rect 68409 21904 68434 21944
rect 68434 21904 68474 21944
rect 68474 21904 68495 21944
rect 68577 21904 68598 21944
rect 68598 21904 68638 21944
rect 68638 21904 68663 21944
rect 68409 21881 68495 21904
rect 68577 21881 68663 21904
rect 72409 21944 72495 21967
rect 72577 21944 72663 21967
rect 72409 21904 72434 21944
rect 72434 21904 72474 21944
rect 72474 21904 72495 21944
rect 72577 21904 72598 21944
rect 72598 21904 72638 21944
rect 72638 21904 72663 21944
rect 72409 21881 72495 21904
rect 72577 21881 72663 21904
rect 76409 21944 76495 21967
rect 76577 21944 76663 21967
rect 76409 21904 76434 21944
rect 76434 21904 76474 21944
rect 76474 21904 76495 21944
rect 76577 21904 76598 21944
rect 76598 21904 76638 21944
rect 76638 21904 76663 21944
rect 76409 21881 76495 21904
rect 76577 21881 76663 21904
rect 80409 21944 80495 21967
rect 80577 21944 80663 21967
rect 80409 21904 80434 21944
rect 80434 21904 80474 21944
rect 80474 21904 80495 21944
rect 80577 21904 80598 21944
rect 80598 21904 80638 21944
rect 80638 21904 80663 21944
rect 80409 21881 80495 21904
rect 80577 21881 80663 21904
rect 84409 21944 84495 21967
rect 84577 21944 84663 21967
rect 84409 21904 84434 21944
rect 84434 21904 84474 21944
rect 84474 21904 84495 21944
rect 84577 21904 84598 21944
rect 84598 21904 84638 21944
rect 84638 21904 84663 21944
rect 84409 21881 84495 21904
rect 84577 21881 84663 21904
rect 88409 21944 88495 21967
rect 88577 21944 88663 21967
rect 88409 21904 88434 21944
rect 88434 21904 88474 21944
rect 88474 21904 88495 21944
rect 88577 21904 88598 21944
rect 88598 21904 88638 21944
rect 88638 21904 88663 21944
rect 88409 21881 88495 21904
rect 88577 21881 88663 21904
rect 92409 21944 92495 21967
rect 92577 21944 92663 21967
rect 92409 21904 92434 21944
rect 92434 21904 92474 21944
rect 92474 21904 92495 21944
rect 92577 21904 92598 21944
rect 92598 21904 92638 21944
rect 92638 21904 92663 21944
rect 92409 21881 92495 21904
rect 92577 21881 92663 21904
rect 96409 21944 96495 21967
rect 96577 21944 96663 21967
rect 96409 21904 96434 21944
rect 96434 21904 96474 21944
rect 96474 21904 96495 21944
rect 96577 21904 96598 21944
rect 96598 21904 96638 21944
rect 96638 21904 96663 21944
rect 96409 21881 96495 21904
rect 96577 21881 96663 21904
rect 3169 21188 3255 21211
rect 3337 21188 3423 21211
rect 3169 21148 3194 21188
rect 3194 21148 3234 21188
rect 3234 21148 3255 21188
rect 3337 21148 3358 21188
rect 3358 21148 3398 21188
rect 3398 21148 3423 21188
rect 3169 21125 3255 21148
rect 3337 21125 3423 21148
rect 7169 21188 7255 21211
rect 7337 21188 7423 21211
rect 7169 21148 7194 21188
rect 7194 21148 7234 21188
rect 7234 21148 7255 21188
rect 7337 21148 7358 21188
rect 7358 21148 7398 21188
rect 7398 21148 7423 21188
rect 7169 21125 7255 21148
rect 7337 21125 7423 21148
rect 11169 21188 11255 21211
rect 11337 21188 11423 21211
rect 11169 21148 11194 21188
rect 11194 21148 11234 21188
rect 11234 21148 11255 21188
rect 11337 21148 11358 21188
rect 11358 21148 11398 21188
rect 11398 21148 11423 21188
rect 11169 21125 11255 21148
rect 11337 21125 11423 21148
rect 15169 21188 15255 21211
rect 15337 21188 15423 21211
rect 15169 21148 15194 21188
rect 15194 21148 15234 21188
rect 15234 21148 15255 21188
rect 15337 21148 15358 21188
rect 15358 21148 15398 21188
rect 15398 21148 15423 21188
rect 15169 21125 15255 21148
rect 15337 21125 15423 21148
rect 19169 21188 19255 21211
rect 19337 21188 19423 21211
rect 19169 21148 19194 21188
rect 19194 21148 19234 21188
rect 19234 21148 19255 21188
rect 19337 21148 19358 21188
rect 19358 21148 19398 21188
rect 19398 21148 19423 21188
rect 19169 21125 19255 21148
rect 19337 21125 19423 21148
rect 23169 21188 23255 21211
rect 23337 21188 23423 21211
rect 23169 21148 23194 21188
rect 23194 21148 23234 21188
rect 23234 21148 23255 21188
rect 23337 21148 23358 21188
rect 23358 21148 23398 21188
rect 23398 21148 23423 21188
rect 23169 21125 23255 21148
rect 23337 21125 23423 21148
rect 27169 21188 27255 21211
rect 27337 21188 27423 21211
rect 27169 21148 27194 21188
rect 27194 21148 27234 21188
rect 27234 21148 27255 21188
rect 27337 21148 27358 21188
rect 27358 21148 27398 21188
rect 27398 21148 27423 21188
rect 27169 21125 27255 21148
rect 27337 21125 27423 21148
rect 31169 21188 31255 21211
rect 31337 21188 31423 21211
rect 31169 21148 31194 21188
rect 31194 21148 31234 21188
rect 31234 21148 31255 21188
rect 31337 21148 31358 21188
rect 31358 21148 31398 21188
rect 31398 21148 31423 21188
rect 31169 21125 31255 21148
rect 31337 21125 31423 21148
rect 35169 21188 35255 21211
rect 35337 21188 35423 21211
rect 35169 21148 35194 21188
rect 35194 21148 35234 21188
rect 35234 21148 35255 21188
rect 35337 21148 35358 21188
rect 35358 21148 35398 21188
rect 35398 21148 35423 21188
rect 35169 21125 35255 21148
rect 35337 21125 35423 21148
rect 39169 21188 39255 21211
rect 39337 21188 39423 21211
rect 39169 21148 39194 21188
rect 39194 21148 39234 21188
rect 39234 21148 39255 21188
rect 39337 21148 39358 21188
rect 39358 21148 39398 21188
rect 39398 21148 39423 21188
rect 39169 21125 39255 21148
rect 39337 21125 39423 21148
rect 43169 21188 43255 21211
rect 43337 21188 43423 21211
rect 43169 21148 43194 21188
rect 43194 21148 43234 21188
rect 43234 21148 43255 21188
rect 43337 21148 43358 21188
rect 43358 21148 43398 21188
rect 43398 21148 43423 21188
rect 43169 21125 43255 21148
rect 43337 21125 43423 21148
rect 47169 21188 47255 21211
rect 47337 21188 47423 21211
rect 47169 21148 47194 21188
rect 47194 21148 47234 21188
rect 47234 21148 47255 21188
rect 47337 21148 47358 21188
rect 47358 21148 47398 21188
rect 47398 21148 47423 21188
rect 47169 21125 47255 21148
rect 47337 21125 47423 21148
rect 51169 21188 51255 21211
rect 51337 21188 51423 21211
rect 51169 21148 51194 21188
rect 51194 21148 51234 21188
rect 51234 21148 51255 21188
rect 51337 21148 51358 21188
rect 51358 21148 51398 21188
rect 51398 21148 51423 21188
rect 51169 21125 51255 21148
rect 51337 21125 51423 21148
rect 55169 21188 55255 21211
rect 55337 21188 55423 21211
rect 55169 21148 55194 21188
rect 55194 21148 55234 21188
rect 55234 21148 55255 21188
rect 55337 21148 55358 21188
rect 55358 21148 55398 21188
rect 55398 21148 55423 21188
rect 55169 21125 55255 21148
rect 55337 21125 55423 21148
rect 59169 21188 59255 21211
rect 59337 21188 59423 21211
rect 59169 21148 59194 21188
rect 59194 21148 59234 21188
rect 59234 21148 59255 21188
rect 59337 21148 59358 21188
rect 59358 21148 59398 21188
rect 59398 21148 59423 21188
rect 59169 21125 59255 21148
rect 59337 21125 59423 21148
rect 63169 21188 63255 21211
rect 63337 21188 63423 21211
rect 63169 21148 63194 21188
rect 63194 21148 63234 21188
rect 63234 21148 63255 21188
rect 63337 21148 63358 21188
rect 63358 21148 63398 21188
rect 63398 21148 63423 21188
rect 63169 21125 63255 21148
rect 63337 21125 63423 21148
rect 67169 21188 67255 21211
rect 67337 21188 67423 21211
rect 67169 21148 67194 21188
rect 67194 21148 67234 21188
rect 67234 21148 67255 21188
rect 67337 21148 67358 21188
rect 67358 21148 67398 21188
rect 67398 21148 67423 21188
rect 67169 21125 67255 21148
rect 67337 21125 67423 21148
rect 71169 21188 71255 21211
rect 71337 21188 71423 21211
rect 71169 21148 71194 21188
rect 71194 21148 71234 21188
rect 71234 21148 71255 21188
rect 71337 21148 71358 21188
rect 71358 21148 71398 21188
rect 71398 21148 71423 21188
rect 71169 21125 71255 21148
rect 71337 21125 71423 21148
rect 75169 21188 75255 21211
rect 75337 21188 75423 21211
rect 75169 21148 75194 21188
rect 75194 21148 75234 21188
rect 75234 21148 75255 21188
rect 75337 21148 75358 21188
rect 75358 21148 75398 21188
rect 75398 21148 75423 21188
rect 75169 21125 75255 21148
rect 75337 21125 75423 21148
rect 79169 21188 79255 21211
rect 79337 21188 79423 21211
rect 79169 21148 79194 21188
rect 79194 21148 79234 21188
rect 79234 21148 79255 21188
rect 79337 21148 79358 21188
rect 79358 21148 79398 21188
rect 79398 21148 79423 21188
rect 79169 21125 79255 21148
rect 79337 21125 79423 21148
rect 83169 21188 83255 21211
rect 83337 21188 83423 21211
rect 83169 21148 83194 21188
rect 83194 21148 83234 21188
rect 83234 21148 83255 21188
rect 83337 21148 83358 21188
rect 83358 21148 83398 21188
rect 83398 21148 83423 21188
rect 83169 21125 83255 21148
rect 83337 21125 83423 21148
rect 87169 21188 87255 21211
rect 87337 21188 87423 21211
rect 87169 21148 87194 21188
rect 87194 21148 87234 21188
rect 87234 21148 87255 21188
rect 87337 21148 87358 21188
rect 87358 21148 87398 21188
rect 87398 21148 87423 21188
rect 87169 21125 87255 21148
rect 87337 21125 87423 21148
rect 91169 21188 91255 21211
rect 91337 21188 91423 21211
rect 91169 21148 91194 21188
rect 91194 21148 91234 21188
rect 91234 21148 91255 21188
rect 91337 21148 91358 21188
rect 91358 21148 91398 21188
rect 91398 21148 91423 21188
rect 91169 21125 91255 21148
rect 91337 21125 91423 21148
rect 95169 21188 95255 21211
rect 95337 21188 95423 21211
rect 95169 21148 95194 21188
rect 95194 21148 95234 21188
rect 95234 21148 95255 21188
rect 95337 21148 95358 21188
rect 95358 21148 95398 21188
rect 95398 21148 95423 21188
rect 95169 21125 95255 21148
rect 95337 21125 95423 21148
rect 99169 21188 99255 21211
rect 99337 21188 99423 21211
rect 99169 21148 99194 21188
rect 99194 21148 99234 21188
rect 99234 21148 99255 21188
rect 99337 21148 99358 21188
rect 99358 21148 99398 21188
rect 99398 21148 99423 21188
rect 99169 21125 99255 21148
rect 99337 21125 99423 21148
rect 4409 20432 4495 20455
rect 4577 20432 4663 20455
rect 4409 20392 4434 20432
rect 4434 20392 4474 20432
rect 4474 20392 4495 20432
rect 4577 20392 4598 20432
rect 4598 20392 4638 20432
rect 4638 20392 4663 20432
rect 4409 20369 4495 20392
rect 4577 20369 4663 20392
rect 8409 20432 8495 20455
rect 8577 20432 8663 20455
rect 8409 20392 8434 20432
rect 8434 20392 8474 20432
rect 8474 20392 8495 20432
rect 8577 20392 8598 20432
rect 8598 20392 8638 20432
rect 8638 20392 8663 20432
rect 8409 20369 8495 20392
rect 8577 20369 8663 20392
rect 12409 20432 12495 20455
rect 12577 20432 12663 20455
rect 12409 20392 12434 20432
rect 12434 20392 12474 20432
rect 12474 20392 12495 20432
rect 12577 20392 12598 20432
rect 12598 20392 12638 20432
rect 12638 20392 12663 20432
rect 12409 20369 12495 20392
rect 12577 20369 12663 20392
rect 16409 20432 16495 20455
rect 16577 20432 16663 20455
rect 16409 20392 16434 20432
rect 16434 20392 16474 20432
rect 16474 20392 16495 20432
rect 16577 20392 16598 20432
rect 16598 20392 16638 20432
rect 16638 20392 16663 20432
rect 16409 20369 16495 20392
rect 16577 20369 16663 20392
rect 20409 20432 20495 20455
rect 20577 20432 20663 20455
rect 20409 20392 20434 20432
rect 20434 20392 20474 20432
rect 20474 20392 20495 20432
rect 20577 20392 20598 20432
rect 20598 20392 20638 20432
rect 20638 20392 20663 20432
rect 20409 20369 20495 20392
rect 20577 20369 20663 20392
rect 24409 20432 24495 20455
rect 24577 20432 24663 20455
rect 24409 20392 24434 20432
rect 24434 20392 24474 20432
rect 24474 20392 24495 20432
rect 24577 20392 24598 20432
rect 24598 20392 24638 20432
rect 24638 20392 24663 20432
rect 24409 20369 24495 20392
rect 24577 20369 24663 20392
rect 28409 20432 28495 20455
rect 28577 20432 28663 20455
rect 28409 20392 28434 20432
rect 28434 20392 28474 20432
rect 28474 20392 28495 20432
rect 28577 20392 28598 20432
rect 28598 20392 28638 20432
rect 28638 20392 28663 20432
rect 28409 20369 28495 20392
rect 28577 20369 28663 20392
rect 32409 20432 32495 20455
rect 32577 20432 32663 20455
rect 32409 20392 32434 20432
rect 32434 20392 32474 20432
rect 32474 20392 32495 20432
rect 32577 20392 32598 20432
rect 32598 20392 32638 20432
rect 32638 20392 32663 20432
rect 32409 20369 32495 20392
rect 32577 20369 32663 20392
rect 36409 20432 36495 20455
rect 36577 20432 36663 20455
rect 36409 20392 36434 20432
rect 36434 20392 36474 20432
rect 36474 20392 36495 20432
rect 36577 20392 36598 20432
rect 36598 20392 36638 20432
rect 36638 20392 36663 20432
rect 36409 20369 36495 20392
rect 36577 20369 36663 20392
rect 40409 20432 40495 20455
rect 40577 20432 40663 20455
rect 40409 20392 40434 20432
rect 40434 20392 40474 20432
rect 40474 20392 40495 20432
rect 40577 20392 40598 20432
rect 40598 20392 40638 20432
rect 40638 20392 40663 20432
rect 40409 20369 40495 20392
rect 40577 20369 40663 20392
rect 44409 20432 44495 20455
rect 44577 20432 44663 20455
rect 44409 20392 44434 20432
rect 44434 20392 44474 20432
rect 44474 20392 44495 20432
rect 44577 20392 44598 20432
rect 44598 20392 44638 20432
rect 44638 20392 44663 20432
rect 44409 20369 44495 20392
rect 44577 20369 44663 20392
rect 48409 20432 48495 20455
rect 48577 20432 48663 20455
rect 48409 20392 48434 20432
rect 48434 20392 48474 20432
rect 48474 20392 48495 20432
rect 48577 20392 48598 20432
rect 48598 20392 48638 20432
rect 48638 20392 48663 20432
rect 48409 20369 48495 20392
rect 48577 20369 48663 20392
rect 52409 20432 52495 20455
rect 52577 20432 52663 20455
rect 52409 20392 52434 20432
rect 52434 20392 52474 20432
rect 52474 20392 52495 20432
rect 52577 20392 52598 20432
rect 52598 20392 52638 20432
rect 52638 20392 52663 20432
rect 52409 20369 52495 20392
rect 52577 20369 52663 20392
rect 56409 20432 56495 20455
rect 56577 20432 56663 20455
rect 56409 20392 56434 20432
rect 56434 20392 56474 20432
rect 56474 20392 56495 20432
rect 56577 20392 56598 20432
rect 56598 20392 56638 20432
rect 56638 20392 56663 20432
rect 56409 20369 56495 20392
rect 56577 20369 56663 20392
rect 60409 20432 60495 20455
rect 60577 20432 60663 20455
rect 60409 20392 60434 20432
rect 60434 20392 60474 20432
rect 60474 20392 60495 20432
rect 60577 20392 60598 20432
rect 60598 20392 60638 20432
rect 60638 20392 60663 20432
rect 60409 20369 60495 20392
rect 60577 20369 60663 20392
rect 64409 20432 64495 20455
rect 64577 20432 64663 20455
rect 64409 20392 64434 20432
rect 64434 20392 64474 20432
rect 64474 20392 64495 20432
rect 64577 20392 64598 20432
rect 64598 20392 64638 20432
rect 64638 20392 64663 20432
rect 64409 20369 64495 20392
rect 64577 20369 64663 20392
rect 68409 20432 68495 20455
rect 68577 20432 68663 20455
rect 68409 20392 68434 20432
rect 68434 20392 68474 20432
rect 68474 20392 68495 20432
rect 68577 20392 68598 20432
rect 68598 20392 68638 20432
rect 68638 20392 68663 20432
rect 68409 20369 68495 20392
rect 68577 20369 68663 20392
rect 72409 20432 72495 20455
rect 72577 20432 72663 20455
rect 72409 20392 72434 20432
rect 72434 20392 72474 20432
rect 72474 20392 72495 20432
rect 72577 20392 72598 20432
rect 72598 20392 72638 20432
rect 72638 20392 72663 20432
rect 72409 20369 72495 20392
rect 72577 20369 72663 20392
rect 76409 20432 76495 20455
rect 76577 20432 76663 20455
rect 76409 20392 76434 20432
rect 76434 20392 76474 20432
rect 76474 20392 76495 20432
rect 76577 20392 76598 20432
rect 76598 20392 76638 20432
rect 76638 20392 76663 20432
rect 76409 20369 76495 20392
rect 76577 20369 76663 20392
rect 80409 20432 80495 20455
rect 80577 20432 80663 20455
rect 80409 20392 80434 20432
rect 80434 20392 80474 20432
rect 80474 20392 80495 20432
rect 80577 20392 80598 20432
rect 80598 20392 80638 20432
rect 80638 20392 80663 20432
rect 80409 20369 80495 20392
rect 80577 20369 80663 20392
rect 84409 20432 84495 20455
rect 84577 20432 84663 20455
rect 84409 20392 84434 20432
rect 84434 20392 84474 20432
rect 84474 20392 84495 20432
rect 84577 20392 84598 20432
rect 84598 20392 84638 20432
rect 84638 20392 84663 20432
rect 84409 20369 84495 20392
rect 84577 20369 84663 20392
rect 88409 20432 88495 20455
rect 88577 20432 88663 20455
rect 88409 20392 88434 20432
rect 88434 20392 88474 20432
rect 88474 20392 88495 20432
rect 88577 20392 88598 20432
rect 88598 20392 88638 20432
rect 88638 20392 88663 20432
rect 88409 20369 88495 20392
rect 88577 20369 88663 20392
rect 92409 20432 92495 20455
rect 92577 20432 92663 20455
rect 92409 20392 92434 20432
rect 92434 20392 92474 20432
rect 92474 20392 92495 20432
rect 92577 20392 92598 20432
rect 92598 20392 92638 20432
rect 92638 20392 92663 20432
rect 92409 20369 92495 20392
rect 92577 20369 92663 20392
rect 96409 20432 96495 20455
rect 96577 20432 96663 20455
rect 96409 20392 96434 20432
rect 96434 20392 96474 20432
rect 96474 20392 96495 20432
rect 96577 20392 96598 20432
rect 96598 20392 96638 20432
rect 96638 20392 96663 20432
rect 96409 20369 96495 20392
rect 96577 20369 96663 20392
rect 3169 19676 3255 19699
rect 3337 19676 3423 19699
rect 3169 19636 3194 19676
rect 3194 19636 3234 19676
rect 3234 19636 3255 19676
rect 3337 19636 3358 19676
rect 3358 19636 3398 19676
rect 3398 19636 3423 19676
rect 3169 19613 3255 19636
rect 3337 19613 3423 19636
rect 7169 19676 7255 19699
rect 7337 19676 7423 19699
rect 7169 19636 7194 19676
rect 7194 19636 7234 19676
rect 7234 19636 7255 19676
rect 7337 19636 7358 19676
rect 7358 19636 7398 19676
rect 7398 19636 7423 19676
rect 7169 19613 7255 19636
rect 7337 19613 7423 19636
rect 11169 19676 11255 19699
rect 11337 19676 11423 19699
rect 11169 19636 11194 19676
rect 11194 19636 11234 19676
rect 11234 19636 11255 19676
rect 11337 19636 11358 19676
rect 11358 19636 11398 19676
rect 11398 19636 11423 19676
rect 11169 19613 11255 19636
rect 11337 19613 11423 19636
rect 15169 19676 15255 19699
rect 15337 19676 15423 19699
rect 15169 19636 15194 19676
rect 15194 19636 15234 19676
rect 15234 19636 15255 19676
rect 15337 19636 15358 19676
rect 15358 19636 15398 19676
rect 15398 19636 15423 19676
rect 15169 19613 15255 19636
rect 15337 19613 15423 19636
rect 19169 19676 19255 19699
rect 19337 19676 19423 19699
rect 19169 19636 19194 19676
rect 19194 19636 19234 19676
rect 19234 19636 19255 19676
rect 19337 19636 19358 19676
rect 19358 19636 19398 19676
rect 19398 19636 19423 19676
rect 19169 19613 19255 19636
rect 19337 19613 19423 19636
rect 23169 19676 23255 19699
rect 23337 19676 23423 19699
rect 23169 19636 23194 19676
rect 23194 19636 23234 19676
rect 23234 19636 23255 19676
rect 23337 19636 23358 19676
rect 23358 19636 23398 19676
rect 23398 19636 23423 19676
rect 23169 19613 23255 19636
rect 23337 19613 23423 19636
rect 27169 19676 27255 19699
rect 27337 19676 27423 19699
rect 27169 19636 27194 19676
rect 27194 19636 27234 19676
rect 27234 19636 27255 19676
rect 27337 19636 27358 19676
rect 27358 19636 27398 19676
rect 27398 19636 27423 19676
rect 27169 19613 27255 19636
rect 27337 19613 27423 19636
rect 31169 19676 31255 19699
rect 31337 19676 31423 19699
rect 31169 19636 31194 19676
rect 31194 19636 31234 19676
rect 31234 19636 31255 19676
rect 31337 19636 31358 19676
rect 31358 19636 31398 19676
rect 31398 19636 31423 19676
rect 31169 19613 31255 19636
rect 31337 19613 31423 19636
rect 35169 19676 35255 19699
rect 35337 19676 35423 19699
rect 35169 19636 35194 19676
rect 35194 19636 35234 19676
rect 35234 19636 35255 19676
rect 35337 19636 35358 19676
rect 35358 19636 35398 19676
rect 35398 19636 35423 19676
rect 35169 19613 35255 19636
rect 35337 19613 35423 19636
rect 39169 19676 39255 19699
rect 39337 19676 39423 19699
rect 39169 19636 39194 19676
rect 39194 19636 39234 19676
rect 39234 19636 39255 19676
rect 39337 19636 39358 19676
rect 39358 19636 39398 19676
rect 39398 19636 39423 19676
rect 39169 19613 39255 19636
rect 39337 19613 39423 19636
rect 43169 19676 43255 19699
rect 43337 19676 43423 19699
rect 43169 19636 43194 19676
rect 43194 19636 43234 19676
rect 43234 19636 43255 19676
rect 43337 19636 43358 19676
rect 43358 19636 43398 19676
rect 43398 19636 43423 19676
rect 43169 19613 43255 19636
rect 43337 19613 43423 19636
rect 47169 19676 47255 19699
rect 47337 19676 47423 19699
rect 47169 19636 47194 19676
rect 47194 19636 47234 19676
rect 47234 19636 47255 19676
rect 47337 19636 47358 19676
rect 47358 19636 47398 19676
rect 47398 19636 47423 19676
rect 47169 19613 47255 19636
rect 47337 19613 47423 19636
rect 51169 19676 51255 19699
rect 51337 19676 51423 19699
rect 51169 19636 51194 19676
rect 51194 19636 51234 19676
rect 51234 19636 51255 19676
rect 51337 19636 51358 19676
rect 51358 19636 51398 19676
rect 51398 19636 51423 19676
rect 51169 19613 51255 19636
rect 51337 19613 51423 19636
rect 55169 19676 55255 19699
rect 55337 19676 55423 19699
rect 55169 19636 55194 19676
rect 55194 19636 55234 19676
rect 55234 19636 55255 19676
rect 55337 19636 55358 19676
rect 55358 19636 55398 19676
rect 55398 19636 55423 19676
rect 55169 19613 55255 19636
rect 55337 19613 55423 19636
rect 59169 19676 59255 19699
rect 59337 19676 59423 19699
rect 59169 19636 59194 19676
rect 59194 19636 59234 19676
rect 59234 19636 59255 19676
rect 59337 19636 59358 19676
rect 59358 19636 59398 19676
rect 59398 19636 59423 19676
rect 59169 19613 59255 19636
rect 59337 19613 59423 19636
rect 63169 19676 63255 19699
rect 63337 19676 63423 19699
rect 63169 19636 63194 19676
rect 63194 19636 63234 19676
rect 63234 19636 63255 19676
rect 63337 19636 63358 19676
rect 63358 19636 63398 19676
rect 63398 19636 63423 19676
rect 63169 19613 63255 19636
rect 63337 19613 63423 19636
rect 67169 19676 67255 19699
rect 67337 19676 67423 19699
rect 67169 19636 67194 19676
rect 67194 19636 67234 19676
rect 67234 19636 67255 19676
rect 67337 19636 67358 19676
rect 67358 19636 67398 19676
rect 67398 19636 67423 19676
rect 67169 19613 67255 19636
rect 67337 19613 67423 19636
rect 71169 19676 71255 19699
rect 71337 19676 71423 19699
rect 71169 19636 71194 19676
rect 71194 19636 71234 19676
rect 71234 19636 71255 19676
rect 71337 19636 71358 19676
rect 71358 19636 71398 19676
rect 71398 19636 71423 19676
rect 71169 19613 71255 19636
rect 71337 19613 71423 19636
rect 75169 19676 75255 19699
rect 75337 19676 75423 19699
rect 75169 19636 75194 19676
rect 75194 19636 75234 19676
rect 75234 19636 75255 19676
rect 75337 19636 75358 19676
rect 75358 19636 75398 19676
rect 75398 19636 75423 19676
rect 75169 19613 75255 19636
rect 75337 19613 75423 19636
rect 79169 19676 79255 19699
rect 79337 19676 79423 19699
rect 79169 19636 79194 19676
rect 79194 19636 79234 19676
rect 79234 19636 79255 19676
rect 79337 19636 79358 19676
rect 79358 19636 79398 19676
rect 79398 19636 79423 19676
rect 79169 19613 79255 19636
rect 79337 19613 79423 19636
rect 83169 19676 83255 19699
rect 83337 19676 83423 19699
rect 83169 19636 83194 19676
rect 83194 19636 83234 19676
rect 83234 19636 83255 19676
rect 83337 19636 83358 19676
rect 83358 19636 83398 19676
rect 83398 19636 83423 19676
rect 83169 19613 83255 19636
rect 83337 19613 83423 19636
rect 87169 19676 87255 19699
rect 87337 19676 87423 19699
rect 87169 19636 87194 19676
rect 87194 19636 87234 19676
rect 87234 19636 87255 19676
rect 87337 19636 87358 19676
rect 87358 19636 87398 19676
rect 87398 19636 87423 19676
rect 87169 19613 87255 19636
rect 87337 19613 87423 19636
rect 91169 19676 91255 19699
rect 91337 19676 91423 19699
rect 91169 19636 91194 19676
rect 91194 19636 91234 19676
rect 91234 19636 91255 19676
rect 91337 19636 91358 19676
rect 91358 19636 91398 19676
rect 91398 19636 91423 19676
rect 91169 19613 91255 19636
rect 91337 19613 91423 19636
rect 95169 19676 95255 19699
rect 95337 19676 95423 19699
rect 95169 19636 95194 19676
rect 95194 19636 95234 19676
rect 95234 19636 95255 19676
rect 95337 19636 95358 19676
rect 95358 19636 95398 19676
rect 95398 19636 95423 19676
rect 95169 19613 95255 19636
rect 95337 19613 95423 19636
rect 99169 19676 99255 19699
rect 99337 19676 99423 19699
rect 99169 19636 99194 19676
rect 99194 19636 99234 19676
rect 99234 19636 99255 19676
rect 99337 19636 99358 19676
rect 99358 19636 99398 19676
rect 99398 19636 99423 19676
rect 99169 19613 99255 19636
rect 99337 19613 99423 19636
rect 4409 18920 4495 18943
rect 4577 18920 4663 18943
rect 4409 18880 4434 18920
rect 4434 18880 4474 18920
rect 4474 18880 4495 18920
rect 4577 18880 4598 18920
rect 4598 18880 4638 18920
rect 4638 18880 4663 18920
rect 4409 18857 4495 18880
rect 4577 18857 4663 18880
rect 8409 18920 8495 18943
rect 8577 18920 8663 18943
rect 8409 18880 8434 18920
rect 8434 18880 8474 18920
rect 8474 18880 8495 18920
rect 8577 18880 8598 18920
rect 8598 18880 8638 18920
rect 8638 18880 8663 18920
rect 8409 18857 8495 18880
rect 8577 18857 8663 18880
rect 12409 18920 12495 18943
rect 12577 18920 12663 18943
rect 12409 18880 12434 18920
rect 12434 18880 12474 18920
rect 12474 18880 12495 18920
rect 12577 18880 12598 18920
rect 12598 18880 12638 18920
rect 12638 18880 12663 18920
rect 12409 18857 12495 18880
rect 12577 18857 12663 18880
rect 16409 18920 16495 18943
rect 16577 18920 16663 18943
rect 16409 18880 16434 18920
rect 16434 18880 16474 18920
rect 16474 18880 16495 18920
rect 16577 18880 16598 18920
rect 16598 18880 16638 18920
rect 16638 18880 16663 18920
rect 16409 18857 16495 18880
rect 16577 18857 16663 18880
rect 20409 18920 20495 18943
rect 20577 18920 20663 18943
rect 20409 18880 20434 18920
rect 20434 18880 20474 18920
rect 20474 18880 20495 18920
rect 20577 18880 20598 18920
rect 20598 18880 20638 18920
rect 20638 18880 20663 18920
rect 20409 18857 20495 18880
rect 20577 18857 20663 18880
rect 24409 18920 24495 18943
rect 24577 18920 24663 18943
rect 24409 18880 24434 18920
rect 24434 18880 24474 18920
rect 24474 18880 24495 18920
rect 24577 18880 24598 18920
rect 24598 18880 24638 18920
rect 24638 18880 24663 18920
rect 24409 18857 24495 18880
rect 24577 18857 24663 18880
rect 28409 18920 28495 18943
rect 28577 18920 28663 18943
rect 28409 18880 28434 18920
rect 28434 18880 28474 18920
rect 28474 18880 28495 18920
rect 28577 18880 28598 18920
rect 28598 18880 28638 18920
rect 28638 18880 28663 18920
rect 28409 18857 28495 18880
rect 28577 18857 28663 18880
rect 32409 18920 32495 18943
rect 32577 18920 32663 18943
rect 32409 18880 32434 18920
rect 32434 18880 32474 18920
rect 32474 18880 32495 18920
rect 32577 18880 32598 18920
rect 32598 18880 32638 18920
rect 32638 18880 32663 18920
rect 32409 18857 32495 18880
rect 32577 18857 32663 18880
rect 36409 18920 36495 18943
rect 36577 18920 36663 18943
rect 36409 18880 36434 18920
rect 36434 18880 36474 18920
rect 36474 18880 36495 18920
rect 36577 18880 36598 18920
rect 36598 18880 36638 18920
rect 36638 18880 36663 18920
rect 36409 18857 36495 18880
rect 36577 18857 36663 18880
rect 40409 18920 40495 18943
rect 40577 18920 40663 18943
rect 40409 18880 40434 18920
rect 40434 18880 40474 18920
rect 40474 18880 40495 18920
rect 40577 18880 40598 18920
rect 40598 18880 40638 18920
rect 40638 18880 40663 18920
rect 40409 18857 40495 18880
rect 40577 18857 40663 18880
rect 44409 18920 44495 18943
rect 44577 18920 44663 18943
rect 44409 18880 44434 18920
rect 44434 18880 44474 18920
rect 44474 18880 44495 18920
rect 44577 18880 44598 18920
rect 44598 18880 44638 18920
rect 44638 18880 44663 18920
rect 44409 18857 44495 18880
rect 44577 18857 44663 18880
rect 48409 18920 48495 18943
rect 48577 18920 48663 18943
rect 48409 18880 48434 18920
rect 48434 18880 48474 18920
rect 48474 18880 48495 18920
rect 48577 18880 48598 18920
rect 48598 18880 48638 18920
rect 48638 18880 48663 18920
rect 48409 18857 48495 18880
rect 48577 18857 48663 18880
rect 52409 18920 52495 18943
rect 52577 18920 52663 18943
rect 52409 18880 52434 18920
rect 52434 18880 52474 18920
rect 52474 18880 52495 18920
rect 52577 18880 52598 18920
rect 52598 18880 52638 18920
rect 52638 18880 52663 18920
rect 52409 18857 52495 18880
rect 52577 18857 52663 18880
rect 56409 18920 56495 18943
rect 56577 18920 56663 18943
rect 56409 18880 56434 18920
rect 56434 18880 56474 18920
rect 56474 18880 56495 18920
rect 56577 18880 56598 18920
rect 56598 18880 56638 18920
rect 56638 18880 56663 18920
rect 56409 18857 56495 18880
rect 56577 18857 56663 18880
rect 60409 18920 60495 18943
rect 60577 18920 60663 18943
rect 60409 18880 60434 18920
rect 60434 18880 60474 18920
rect 60474 18880 60495 18920
rect 60577 18880 60598 18920
rect 60598 18880 60638 18920
rect 60638 18880 60663 18920
rect 60409 18857 60495 18880
rect 60577 18857 60663 18880
rect 64409 18920 64495 18943
rect 64577 18920 64663 18943
rect 64409 18880 64434 18920
rect 64434 18880 64474 18920
rect 64474 18880 64495 18920
rect 64577 18880 64598 18920
rect 64598 18880 64638 18920
rect 64638 18880 64663 18920
rect 64409 18857 64495 18880
rect 64577 18857 64663 18880
rect 68409 18920 68495 18943
rect 68577 18920 68663 18943
rect 68409 18880 68434 18920
rect 68434 18880 68474 18920
rect 68474 18880 68495 18920
rect 68577 18880 68598 18920
rect 68598 18880 68638 18920
rect 68638 18880 68663 18920
rect 68409 18857 68495 18880
rect 68577 18857 68663 18880
rect 72409 18920 72495 18943
rect 72577 18920 72663 18943
rect 72409 18880 72434 18920
rect 72434 18880 72474 18920
rect 72474 18880 72495 18920
rect 72577 18880 72598 18920
rect 72598 18880 72638 18920
rect 72638 18880 72663 18920
rect 72409 18857 72495 18880
rect 72577 18857 72663 18880
rect 76409 18920 76495 18943
rect 76577 18920 76663 18943
rect 76409 18880 76434 18920
rect 76434 18880 76474 18920
rect 76474 18880 76495 18920
rect 76577 18880 76598 18920
rect 76598 18880 76638 18920
rect 76638 18880 76663 18920
rect 76409 18857 76495 18880
rect 76577 18857 76663 18880
rect 80409 18920 80495 18943
rect 80577 18920 80663 18943
rect 80409 18880 80434 18920
rect 80434 18880 80474 18920
rect 80474 18880 80495 18920
rect 80577 18880 80598 18920
rect 80598 18880 80638 18920
rect 80638 18880 80663 18920
rect 80409 18857 80495 18880
rect 80577 18857 80663 18880
rect 84409 18920 84495 18943
rect 84577 18920 84663 18943
rect 84409 18880 84434 18920
rect 84434 18880 84474 18920
rect 84474 18880 84495 18920
rect 84577 18880 84598 18920
rect 84598 18880 84638 18920
rect 84638 18880 84663 18920
rect 84409 18857 84495 18880
rect 84577 18857 84663 18880
rect 88409 18920 88495 18943
rect 88577 18920 88663 18943
rect 88409 18880 88434 18920
rect 88434 18880 88474 18920
rect 88474 18880 88495 18920
rect 88577 18880 88598 18920
rect 88598 18880 88638 18920
rect 88638 18880 88663 18920
rect 88409 18857 88495 18880
rect 88577 18857 88663 18880
rect 92409 18920 92495 18943
rect 92577 18920 92663 18943
rect 92409 18880 92434 18920
rect 92434 18880 92474 18920
rect 92474 18880 92495 18920
rect 92577 18880 92598 18920
rect 92598 18880 92638 18920
rect 92638 18880 92663 18920
rect 92409 18857 92495 18880
rect 92577 18857 92663 18880
rect 96409 18920 96495 18943
rect 96577 18920 96663 18943
rect 96409 18880 96434 18920
rect 96434 18880 96474 18920
rect 96474 18880 96495 18920
rect 96577 18880 96598 18920
rect 96598 18880 96638 18920
rect 96638 18880 96663 18920
rect 96409 18857 96495 18880
rect 96577 18857 96663 18880
rect 3169 18164 3255 18187
rect 3337 18164 3423 18187
rect 3169 18124 3194 18164
rect 3194 18124 3234 18164
rect 3234 18124 3255 18164
rect 3337 18124 3358 18164
rect 3358 18124 3398 18164
rect 3398 18124 3423 18164
rect 3169 18101 3255 18124
rect 3337 18101 3423 18124
rect 7169 18164 7255 18187
rect 7337 18164 7423 18187
rect 7169 18124 7194 18164
rect 7194 18124 7234 18164
rect 7234 18124 7255 18164
rect 7337 18124 7358 18164
rect 7358 18124 7398 18164
rect 7398 18124 7423 18164
rect 7169 18101 7255 18124
rect 7337 18101 7423 18124
rect 11169 18164 11255 18187
rect 11337 18164 11423 18187
rect 11169 18124 11194 18164
rect 11194 18124 11234 18164
rect 11234 18124 11255 18164
rect 11337 18124 11358 18164
rect 11358 18124 11398 18164
rect 11398 18124 11423 18164
rect 11169 18101 11255 18124
rect 11337 18101 11423 18124
rect 15169 18164 15255 18187
rect 15337 18164 15423 18187
rect 15169 18124 15194 18164
rect 15194 18124 15234 18164
rect 15234 18124 15255 18164
rect 15337 18124 15358 18164
rect 15358 18124 15398 18164
rect 15398 18124 15423 18164
rect 15169 18101 15255 18124
rect 15337 18101 15423 18124
rect 19169 18164 19255 18187
rect 19337 18164 19423 18187
rect 19169 18124 19194 18164
rect 19194 18124 19234 18164
rect 19234 18124 19255 18164
rect 19337 18124 19358 18164
rect 19358 18124 19398 18164
rect 19398 18124 19423 18164
rect 19169 18101 19255 18124
rect 19337 18101 19423 18124
rect 23169 18164 23255 18187
rect 23337 18164 23423 18187
rect 23169 18124 23194 18164
rect 23194 18124 23234 18164
rect 23234 18124 23255 18164
rect 23337 18124 23358 18164
rect 23358 18124 23398 18164
rect 23398 18124 23423 18164
rect 23169 18101 23255 18124
rect 23337 18101 23423 18124
rect 27169 18164 27255 18187
rect 27337 18164 27423 18187
rect 27169 18124 27194 18164
rect 27194 18124 27234 18164
rect 27234 18124 27255 18164
rect 27337 18124 27358 18164
rect 27358 18124 27398 18164
rect 27398 18124 27423 18164
rect 27169 18101 27255 18124
rect 27337 18101 27423 18124
rect 31169 18164 31255 18187
rect 31337 18164 31423 18187
rect 31169 18124 31194 18164
rect 31194 18124 31234 18164
rect 31234 18124 31255 18164
rect 31337 18124 31358 18164
rect 31358 18124 31398 18164
rect 31398 18124 31423 18164
rect 31169 18101 31255 18124
rect 31337 18101 31423 18124
rect 35169 18164 35255 18187
rect 35337 18164 35423 18187
rect 35169 18124 35194 18164
rect 35194 18124 35234 18164
rect 35234 18124 35255 18164
rect 35337 18124 35358 18164
rect 35358 18124 35398 18164
rect 35398 18124 35423 18164
rect 35169 18101 35255 18124
rect 35337 18101 35423 18124
rect 39169 18164 39255 18187
rect 39337 18164 39423 18187
rect 39169 18124 39194 18164
rect 39194 18124 39234 18164
rect 39234 18124 39255 18164
rect 39337 18124 39358 18164
rect 39358 18124 39398 18164
rect 39398 18124 39423 18164
rect 39169 18101 39255 18124
rect 39337 18101 39423 18124
rect 43169 18164 43255 18187
rect 43337 18164 43423 18187
rect 43169 18124 43194 18164
rect 43194 18124 43234 18164
rect 43234 18124 43255 18164
rect 43337 18124 43358 18164
rect 43358 18124 43398 18164
rect 43398 18124 43423 18164
rect 43169 18101 43255 18124
rect 43337 18101 43423 18124
rect 47169 18164 47255 18187
rect 47337 18164 47423 18187
rect 47169 18124 47194 18164
rect 47194 18124 47234 18164
rect 47234 18124 47255 18164
rect 47337 18124 47358 18164
rect 47358 18124 47398 18164
rect 47398 18124 47423 18164
rect 47169 18101 47255 18124
rect 47337 18101 47423 18124
rect 51169 18164 51255 18187
rect 51337 18164 51423 18187
rect 51169 18124 51194 18164
rect 51194 18124 51234 18164
rect 51234 18124 51255 18164
rect 51337 18124 51358 18164
rect 51358 18124 51398 18164
rect 51398 18124 51423 18164
rect 51169 18101 51255 18124
rect 51337 18101 51423 18124
rect 55169 18164 55255 18187
rect 55337 18164 55423 18187
rect 55169 18124 55194 18164
rect 55194 18124 55234 18164
rect 55234 18124 55255 18164
rect 55337 18124 55358 18164
rect 55358 18124 55398 18164
rect 55398 18124 55423 18164
rect 55169 18101 55255 18124
rect 55337 18101 55423 18124
rect 59169 18164 59255 18187
rect 59337 18164 59423 18187
rect 59169 18124 59194 18164
rect 59194 18124 59234 18164
rect 59234 18124 59255 18164
rect 59337 18124 59358 18164
rect 59358 18124 59398 18164
rect 59398 18124 59423 18164
rect 59169 18101 59255 18124
rect 59337 18101 59423 18124
rect 63169 18164 63255 18187
rect 63337 18164 63423 18187
rect 63169 18124 63194 18164
rect 63194 18124 63234 18164
rect 63234 18124 63255 18164
rect 63337 18124 63358 18164
rect 63358 18124 63398 18164
rect 63398 18124 63423 18164
rect 63169 18101 63255 18124
rect 63337 18101 63423 18124
rect 67169 18164 67255 18187
rect 67337 18164 67423 18187
rect 67169 18124 67194 18164
rect 67194 18124 67234 18164
rect 67234 18124 67255 18164
rect 67337 18124 67358 18164
rect 67358 18124 67398 18164
rect 67398 18124 67423 18164
rect 67169 18101 67255 18124
rect 67337 18101 67423 18124
rect 71169 18164 71255 18187
rect 71337 18164 71423 18187
rect 71169 18124 71194 18164
rect 71194 18124 71234 18164
rect 71234 18124 71255 18164
rect 71337 18124 71358 18164
rect 71358 18124 71398 18164
rect 71398 18124 71423 18164
rect 71169 18101 71255 18124
rect 71337 18101 71423 18124
rect 75169 18164 75255 18187
rect 75337 18164 75423 18187
rect 75169 18124 75194 18164
rect 75194 18124 75234 18164
rect 75234 18124 75255 18164
rect 75337 18124 75358 18164
rect 75358 18124 75398 18164
rect 75398 18124 75423 18164
rect 75169 18101 75255 18124
rect 75337 18101 75423 18124
rect 79169 18164 79255 18187
rect 79337 18164 79423 18187
rect 79169 18124 79194 18164
rect 79194 18124 79234 18164
rect 79234 18124 79255 18164
rect 79337 18124 79358 18164
rect 79358 18124 79398 18164
rect 79398 18124 79423 18164
rect 79169 18101 79255 18124
rect 79337 18101 79423 18124
rect 83169 18164 83255 18187
rect 83337 18164 83423 18187
rect 83169 18124 83194 18164
rect 83194 18124 83234 18164
rect 83234 18124 83255 18164
rect 83337 18124 83358 18164
rect 83358 18124 83398 18164
rect 83398 18124 83423 18164
rect 83169 18101 83255 18124
rect 83337 18101 83423 18124
rect 87169 18164 87255 18187
rect 87337 18164 87423 18187
rect 87169 18124 87194 18164
rect 87194 18124 87234 18164
rect 87234 18124 87255 18164
rect 87337 18124 87358 18164
rect 87358 18124 87398 18164
rect 87398 18124 87423 18164
rect 87169 18101 87255 18124
rect 87337 18101 87423 18124
rect 91169 18164 91255 18187
rect 91337 18164 91423 18187
rect 91169 18124 91194 18164
rect 91194 18124 91234 18164
rect 91234 18124 91255 18164
rect 91337 18124 91358 18164
rect 91358 18124 91398 18164
rect 91398 18124 91423 18164
rect 91169 18101 91255 18124
rect 91337 18101 91423 18124
rect 95169 18164 95255 18187
rect 95337 18164 95423 18187
rect 95169 18124 95194 18164
rect 95194 18124 95234 18164
rect 95234 18124 95255 18164
rect 95337 18124 95358 18164
rect 95358 18124 95398 18164
rect 95398 18124 95423 18164
rect 95169 18101 95255 18124
rect 95337 18101 95423 18124
rect 99169 18164 99255 18187
rect 99337 18164 99423 18187
rect 99169 18124 99194 18164
rect 99194 18124 99234 18164
rect 99234 18124 99255 18164
rect 99337 18124 99358 18164
rect 99358 18124 99398 18164
rect 99398 18124 99423 18164
rect 99169 18101 99255 18124
rect 99337 18101 99423 18124
rect 4409 17408 4495 17431
rect 4577 17408 4663 17431
rect 4409 17368 4434 17408
rect 4434 17368 4474 17408
rect 4474 17368 4495 17408
rect 4577 17368 4598 17408
rect 4598 17368 4638 17408
rect 4638 17368 4663 17408
rect 4409 17345 4495 17368
rect 4577 17345 4663 17368
rect 8409 17408 8495 17431
rect 8577 17408 8663 17431
rect 8409 17368 8434 17408
rect 8434 17368 8474 17408
rect 8474 17368 8495 17408
rect 8577 17368 8598 17408
rect 8598 17368 8638 17408
rect 8638 17368 8663 17408
rect 8409 17345 8495 17368
rect 8577 17345 8663 17368
rect 12409 17408 12495 17431
rect 12577 17408 12663 17431
rect 12409 17368 12434 17408
rect 12434 17368 12474 17408
rect 12474 17368 12495 17408
rect 12577 17368 12598 17408
rect 12598 17368 12638 17408
rect 12638 17368 12663 17408
rect 12409 17345 12495 17368
rect 12577 17345 12663 17368
rect 16409 17408 16495 17431
rect 16577 17408 16663 17431
rect 16409 17368 16434 17408
rect 16434 17368 16474 17408
rect 16474 17368 16495 17408
rect 16577 17368 16598 17408
rect 16598 17368 16638 17408
rect 16638 17368 16663 17408
rect 16409 17345 16495 17368
rect 16577 17345 16663 17368
rect 20409 17408 20495 17431
rect 20577 17408 20663 17431
rect 20409 17368 20434 17408
rect 20434 17368 20474 17408
rect 20474 17368 20495 17408
rect 20577 17368 20598 17408
rect 20598 17368 20638 17408
rect 20638 17368 20663 17408
rect 20409 17345 20495 17368
rect 20577 17345 20663 17368
rect 24409 17408 24495 17431
rect 24577 17408 24663 17431
rect 24409 17368 24434 17408
rect 24434 17368 24474 17408
rect 24474 17368 24495 17408
rect 24577 17368 24598 17408
rect 24598 17368 24638 17408
rect 24638 17368 24663 17408
rect 24409 17345 24495 17368
rect 24577 17345 24663 17368
rect 28409 17408 28495 17431
rect 28577 17408 28663 17431
rect 28409 17368 28434 17408
rect 28434 17368 28474 17408
rect 28474 17368 28495 17408
rect 28577 17368 28598 17408
rect 28598 17368 28638 17408
rect 28638 17368 28663 17408
rect 28409 17345 28495 17368
rect 28577 17345 28663 17368
rect 32409 17408 32495 17431
rect 32577 17408 32663 17431
rect 32409 17368 32434 17408
rect 32434 17368 32474 17408
rect 32474 17368 32495 17408
rect 32577 17368 32598 17408
rect 32598 17368 32638 17408
rect 32638 17368 32663 17408
rect 32409 17345 32495 17368
rect 32577 17345 32663 17368
rect 36409 17408 36495 17431
rect 36577 17408 36663 17431
rect 36409 17368 36434 17408
rect 36434 17368 36474 17408
rect 36474 17368 36495 17408
rect 36577 17368 36598 17408
rect 36598 17368 36638 17408
rect 36638 17368 36663 17408
rect 36409 17345 36495 17368
rect 36577 17345 36663 17368
rect 40409 17408 40495 17431
rect 40577 17408 40663 17431
rect 40409 17368 40434 17408
rect 40434 17368 40474 17408
rect 40474 17368 40495 17408
rect 40577 17368 40598 17408
rect 40598 17368 40638 17408
rect 40638 17368 40663 17408
rect 40409 17345 40495 17368
rect 40577 17345 40663 17368
rect 44409 17408 44495 17431
rect 44577 17408 44663 17431
rect 44409 17368 44434 17408
rect 44434 17368 44474 17408
rect 44474 17368 44495 17408
rect 44577 17368 44598 17408
rect 44598 17368 44638 17408
rect 44638 17368 44663 17408
rect 44409 17345 44495 17368
rect 44577 17345 44663 17368
rect 48409 17408 48495 17431
rect 48577 17408 48663 17431
rect 48409 17368 48434 17408
rect 48434 17368 48474 17408
rect 48474 17368 48495 17408
rect 48577 17368 48598 17408
rect 48598 17368 48638 17408
rect 48638 17368 48663 17408
rect 48409 17345 48495 17368
rect 48577 17345 48663 17368
rect 52409 17408 52495 17431
rect 52577 17408 52663 17431
rect 52409 17368 52434 17408
rect 52434 17368 52474 17408
rect 52474 17368 52495 17408
rect 52577 17368 52598 17408
rect 52598 17368 52638 17408
rect 52638 17368 52663 17408
rect 52409 17345 52495 17368
rect 52577 17345 52663 17368
rect 56409 17408 56495 17431
rect 56577 17408 56663 17431
rect 56409 17368 56434 17408
rect 56434 17368 56474 17408
rect 56474 17368 56495 17408
rect 56577 17368 56598 17408
rect 56598 17368 56638 17408
rect 56638 17368 56663 17408
rect 56409 17345 56495 17368
rect 56577 17345 56663 17368
rect 60409 17408 60495 17431
rect 60577 17408 60663 17431
rect 60409 17368 60434 17408
rect 60434 17368 60474 17408
rect 60474 17368 60495 17408
rect 60577 17368 60598 17408
rect 60598 17368 60638 17408
rect 60638 17368 60663 17408
rect 60409 17345 60495 17368
rect 60577 17345 60663 17368
rect 64409 17408 64495 17431
rect 64577 17408 64663 17431
rect 64409 17368 64434 17408
rect 64434 17368 64474 17408
rect 64474 17368 64495 17408
rect 64577 17368 64598 17408
rect 64598 17368 64638 17408
rect 64638 17368 64663 17408
rect 64409 17345 64495 17368
rect 64577 17345 64663 17368
rect 68409 17408 68495 17431
rect 68577 17408 68663 17431
rect 68409 17368 68434 17408
rect 68434 17368 68474 17408
rect 68474 17368 68495 17408
rect 68577 17368 68598 17408
rect 68598 17368 68638 17408
rect 68638 17368 68663 17408
rect 68409 17345 68495 17368
rect 68577 17345 68663 17368
rect 72409 17408 72495 17431
rect 72577 17408 72663 17431
rect 72409 17368 72434 17408
rect 72434 17368 72474 17408
rect 72474 17368 72495 17408
rect 72577 17368 72598 17408
rect 72598 17368 72638 17408
rect 72638 17368 72663 17408
rect 72409 17345 72495 17368
rect 72577 17345 72663 17368
rect 76409 17408 76495 17431
rect 76577 17408 76663 17431
rect 76409 17368 76434 17408
rect 76434 17368 76474 17408
rect 76474 17368 76495 17408
rect 76577 17368 76598 17408
rect 76598 17368 76638 17408
rect 76638 17368 76663 17408
rect 76409 17345 76495 17368
rect 76577 17345 76663 17368
rect 80409 17408 80495 17431
rect 80577 17408 80663 17431
rect 80409 17368 80434 17408
rect 80434 17368 80474 17408
rect 80474 17368 80495 17408
rect 80577 17368 80598 17408
rect 80598 17368 80638 17408
rect 80638 17368 80663 17408
rect 80409 17345 80495 17368
rect 80577 17345 80663 17368
rect 84409 17408 84495 17431
rect 84577 17408 84663 17431
rect 84409 17368 84434 17408
rect 84434 17368 84474 17408
rect 84474 17368 84495 17408
rect 84577 17368 84598 17408
rect 84598 17368 84638 17408
rect 84638 17368 84663 17408
rect 84409 17345 84495 17368
rect 84577 17345 84663 17368
rect 88409 17408 88495 17431
rect 88577 17408 88663 17431
rect 88409 17368 88434 17408
rect 88434 17368 88474 17408
rect 88474 17368 88495 17408
rect 88577 17368 88598 17408
rect 88598 17368 88638 17408
rect 88638 17368 88663 17408
rect 88409 17345 88495 17368
rect 88577 17345 88663 17368
rect 92409 17408 92495 17431
rect 92577 17408 92663 17431
rect 92409 17368 92434 17408
rect 92434 17368 92474 17408
rect 92474 17368 92495 17408
rect 92577 17368 92598 17408
rect 92598 17368 92638 17408
rect 92638 17368 92663 17408
rect 92409 17345 92495 17368
rect 92577 17345 92663 17368
rect 96409 17408 96495 17431
rect 96577 17408 96663 17431
rect 96409 17368 96434 17408
rect 96434 17368 96474 17408
rect 96474 17368 96495 17408
rect 96577 17368 96598 17408
rect 96598 17368 96638 17408
rect 96638 17368 96663 17408
rect 96409 17345 96495 17368
rect 96577 17345 96663 17368
rect 3169 16652 3255 16675
rect 3337 16652 3423 16675
rect 3169 16612 3194 16652
rect 3194 16612 3234 16652
rect 3234 16612 3255 16652
rect 3337 16612 3358 16652
rect 3358 16612 3398 16652
rect 3398 16612 3423 16652
rect 3169 16589 3255 16612
rect 3337 16589 3423 16612
rect 7169 16652 7255 16675
rect 7337 16652 7423 16675
rect 7169 16612 7194 16652
rect 7194 16612 7234 16652
rect 7234 16612 7255 16652
rect 7337 16612 7358 16652
rect 7358 16612 7398 16652
rect 7398 16612 7423 16652
rect 7169 16589 7255 16612
rect 7337 16589 7423 16612
rect 11169 16652 11255 16675
rect 11337 16652 11423 16675
rect 11169 16612 11194 16652
rect 11194 16612 11234 16652
rect 11234 16612 11255 16652
rect 11337 16612 11358 16652
rect 11358 16612 11398 16652
rect 11398 16612 11423 16652
rect 11169 16589 11255 16612
rect 11337 16589 11423 16612
rect 15169 16652 15255 16675
rect 15337 16652 15423 16675
rect 15169 16612 15194 16652
rect 15194 16612 15234 16652
rect 15234 16612 15255 16652
rect 15337 16612 15358 16652
rect 15358 16612 15398 16652
rect 15398 16612 15423 16652
rect 15169 16589 15255 16612
rect 15337 16589 15423 16612
rect 19169 16652 19255 16675
rect 19337 16652 19423 16675
rect 19169 16612 19194 16652
rect 19194 16612 19234 16652
rect 19234 16612 19255 16652
rect 19337 16612 19358 16652
rect 19358 16612 19398 16652
rect 19398 16612 19423 16652
rect 19169 16589 19255 16612
rect 19337 16589 19423 16612
rect 23169 16652 23255 16675
rect 23337 16652 23423 16675
rect 23169 16612 23194 16652
rect 23194 16612 23234 16652
rect 23234 16612 23255 16652
rect 23337 16612 23358 16652
rect 23358 16612 23398 16652
rect 23398 16612 23423 16652
rect 23169 16589 23255 16612
rect 23337 16589 23423 16612
rect 27169 16652 27255 16675
rect 27337 16652 27423 16675
rect 27169 16612 27194 16652
rect 27194 16612 27234 16652
rect 27234 16612 27255 16652
rect 27337 16612 27358 16652
rect 27358 16612 27398 16652
rect 27398 16612 27423 16652
rect 27169 16589 27255 16612
rect 27337 16589 27423 16612
rect 31169 16652 31255 16675
rect 31337 16652 31423 16675
rect 31169 16612 31194 16652
rect 31194 16612 31234 16652
rect 31234 16612 31255 16652
rect 31337 16612 31358 16652
rect 31358 16612 31398 16652
rect 31398 16612 31423 16652
rect 31169 16589 31255 16612
rect 31337 16589 31423 16612
rect 35169 16652 35255 16675
rect 35337 16652 35423 16675
rect 35169 16612 35194 16652
rect 35194 16612 35234 16652
rect 35234 16612 35255 16652
rect 35337 16612 35358 16652
rect 35358 16612 35398 16652
rect 35398 16612 35423 16652
rect 35169 16589 35255 16612
rect 35337 16589 35423 16612
rect 39169 16652 39255 16675
rect 39337 16652 39423 16675
rect 39169 16612 39194 16652
rect 39194 16612 39234 16652
rect 39234 16612 39255 16652
rect 39337 16612 39358 16652
rect 39358 16612 39398 16652
rect 39398 16612 39423 16652
rect 39169 16589 39255 16612
rect 39337 16589 39423 16612
rect 43169 16652 43255 16675
rect 43337 16652 43423 16675
rect 43169 16612 43194 16652
rect 43194 16612 43234 16652
rect 43234 16612 43255 16652
rect 43337 16612 43358 16652
rect 43358 16612 43398 16652
rect 43398 16612 43423 16652
rect 43169 16589 43255 16612
rect 43337 16589 43423 16612
rect 47169 16652 47255 16675
rect 47337 16652 47423 16675
rect 47169 16612 47194 16652
rect 47194 16612 47234 16652
rect 47234 16612 47255 16652
rect 47337 16612 47358 16652
rect 47358 16612 47398 16652
rect 47398 16612 47423 16652
rect 47169 16589 47255 16612
rect 47337 16589 47423 16612
rect 51169 16652 51255 16675
rect 51337 16652 51423 16675
rect 51169 16612 51194 16652
rect 51194 16612 51234 16652
rect 51234 16612 51255 16652
rect 51337 16612 51358 16652
rect 51358 16612 51398 16652
rect 51398 16612 51423 16652
rect 51169 16589 51255 16612
rect 51337 16589 51423 16612
rect 55169 16652 55255 16675
rect 55337 16652 55423 16675
rect 55169 16612 55194 16652
rect 55194 16612 55234 16652
rect 55234 16612 55255 16652
rect 55337 16612 55358 16652
rect 55358 16612 55398 16652
rect 55398 16612 55423 16652
rect 55169 16589 55255 16612
rect 55337 16589 55423 16612
rect 59169 16652 59255 16675
rect 59337 16652 59423 16675
rect 59169 16612 59194 16652
rect 59194 16612 59234 16652
rect 59234 16612 59255 16652
rect 59337 16612 59358 16652
rect 59358 16612 59398 16652
rect 59398 16612 59423 16652
rect 59169 16589 59255 16612
rect 59337 16589 59423 16612
rect 63169 16652 63255 16675
rect 63337 16652 63423 16675
rect 63169 16612 63194 16652
rect 63194 16612 63234 16652
rect 63234 16612 63255 16652
rect 63337 16612 63358 16652
rect 63358 16612 63398 16652
rect 63398 16612 63423 16652
rect 63169 16589 63255 16612
rect 63337 16589 63423 16612
rect 67169 16652 67255 16675
rect 67337 16652 67423 16675
rect 67169 16612 67194 16652
rect 67194 16612 67234 16652
rect 67234 16612 67255 16652
rect 67337 16612 67358 16652
rect 67358 16612 67398 16652
rect 67398 16612 67423 16652
rect 67169 16589 67255 16612
rect 67337 16589 67423 16612
rect 71169 16652 71255 16675
rect 71337 16652 71423 16675
rect 71169 16612 71194 16652
rect 71194 16612 71234 16652
rect 71234 16612 71255 16652
rect 71337 16612 71358 16652
rect 71358 16612 71398 16652
rect 71398 16612 71423 16652
rect 71169 16589 71255 16612
rect 71337 16589 71423 16612
rect 75169 16652 75255 16675
rect 75337 16652 75423 16675
rect 75169 16612 75194 16652
rect 75194 16612 75234 16652
rect 75234 16612 75255 16652
rect 75337 16612 75358 16652
rect 75358 16612 75398 16652
rect 75398 16612 75423 16652
rect 75169 16589 75255 16612
rect 75337 16589 75423 16612
rect 79169 16652 79255 16675
rect 79337 16652 79423 16675
rect 79169 16612 79194 16652
rect 79194 16612 79234 16652
rect 79234 16612 79255 16652
rect 79337 16612 79358 16652
rect 79358 16612 79398 16652
rect 79398 16612 79423 16652
rect 79169 16589 79255 16612
rect 79337 16589 79423 16612
rect 83169 16652 83255 16675
rect 83337 16652 83423 16675
rect 83169 16612 83194 16652
rect 83194 16612 83234 16652
rect 83234 16612 83255 16652
rect 83337 16612 83358 16652
rect 83358 16612 83398 16652
rect 83398 16612 83423 16652
rect 83169 16589 83255 16612
rect 83337 16589 83423 16612
rect 87169 16652 87255 16675
rect 87337 16652 87423 16675
rect 87169 16612 87194 16652
rect 87194 16612 87234 16652
rect 87234 16612 87255 16652
rect 87337 16612 87358 16652
rect 87358 16612 87398 16652
rect 87398 16612 87423 16652
rect 87169 16589 87255 16612
rect 87337 16589 87423 16612
rect 91169 16652 91255 16675
rect 91337 16652 91423 16675
rect 91169 16612 91194 16652
rect 91194 16612 91234 16652
rect 91234 16612 91255 16652
rect 91337 16612 91358 16652
rect 91358 16612 91398 16652
rect 91398 16612 91423 16652
rect 91169 16589 91255 16612
rect 91337 16589 91423 16612
rect 95169 16652 95255 16675
rect 95337 16652 95423 16675
rect 95169 16612 95194 16652
rect 95194 16612 95234 16652
rect 95234 16612 95255 16652
rect 95337 16612 95358 16652
rect 95358 16612 95398 16652
rect 95398 16612 95423 16652
rect 95169 16589 95255 16612
rect 95337 16589 95423 16612
rect 99169 16652 99255 16675
rect 99337 16652 99423 16675
rect 99169 16612 99194 16652
rect 99194 16612 99234 16652
rect 99234 16612 99255 16652
rect 99337 16612 99358 16652
rect 99358 16612 99398 16652
rect 99398 16612 99423 16652
rect 99169 16589 99255 16612
rect 99337 16589 99423 16612
rect 86469 16337 86555 16423
rect 4409 15896 4495 15919
rect 4577 15896 4663 15919
rect 4409 15856 4434 15896
rect 4434 15856 4474 15896
rect 4474 15856 4495 15896
rect 4577 15856 4598 15896
rect 4598 15856 4638 15896
rect 4638 15856 4663 15896
rect 4409 15833 4495 15856
rect 4577 15833 4663 15856
rect 8409 15896 8495 15919
rect 8577 15896 8663 15919
rect 8409 15856 8434 15896
rect 8434 15856 8474 15896
rect 8474 15856 8495 15896
rect 8577 15856 8598 15896
rect 8598 15856 8638 15896
rect 8638 15856 8663 15896
rect 8409 15833 8495 15856
rect 8577 15833 8663 15856
rect 12409 15896 12495 15919
rect 12577 15896 12663 15919
rect 12409 15856 12434 15896
rect 12434 15856 12474 15896
rect 12474 15856 12495 15896
rect 12577 15856 12598 15896
rect 12598 15856 12638 15896
rect 12638 15856 12663 15896
rect 12409 15833 12495 15856
rect 12577 15833 12663 15856
rect 16409 15896 16495 15919
rect 16577 15896 16663 15919
rect 16409 15856 16434 15896
rect 16434 15856 16474 15896
rect 16474 15856 16495 15896
rect 16577 15856 16598 15896
rect 16598 15856 16638 15896
rect 16638 15856 16663 15896
rect 16409 15833 16495 15856
rect 16577 15833 16663 15856
rect 20409 15896 20495 15919
rect 20577 15896 20663 15919
rect 20409 15856 20434 15896
rect 20434 15856 20474 15896
rect 20474 15856 20495 15896
rect 20577 15856 20598 15896
rect 20598 15856 20638 15896
rect 20638 15856 20663 15896
rect 20409 15833 20495 15856
rect 20577 15833 20663 15856
rect 24409 15896 24495 15919
rect 24577 15896 24663 15919
rect 24409 15856 24434 15896
rect 24434 15856 24474 15896
rect 24474 15856 24495 15896
rect 24577 15856 24598 15896
rect 24598 15856 24638 15896
rect 24638 15856 24663 15896
rect 24409 15833 24495 15856
rect 24577 15833 24663 15856
rect 28409 15896 28495 15919
rect 28577 15896 28663 15919
rect 28409 15856 28434 15896
rect 28434 15856 28474 15896
rect 28474 15856 28495 15896
rect 28577 15856 28598 15896
rect 28598 15856 28638 15896
rect 28638 15856 28663 15896
rect 28409 15833 28495 15856
rect 28577 15833 28663 15856
rect 32409 15896 32495 15919
rect 32577 15896 32663 15919
rect 32409 15856 32434 15896
rect 32434 15856 32474 15896
rect 32474 15856 32495 15896
rect 32577 15856 32598 15896
rect 32598 15856 32638 15896
rect 32638 15856 32663 15896
rect 32409 15833 32495 15856
rect 32577 15833 32663 15856
rect 36409 15896 36495 15919
rect 36577 15896 36663 15919
rect 36409 15856 36434 15896
rect 36434 15856 36474 15896
rect 36474 15856 36495 15896
rect 36577 15856 36598 15896
rect 36598 15856 36638 15896
rect 36638 15856 36663 15896
rect 36409 15833 36495 15856
rect 36577 15833 36663 15856
rect 40409 15896 40495 15919
rect 40577 15896 40663 15919
rect 40409 15856 40434 15896
rect 40434 15856 40474 15896
rect 40474 15856 40495 15896
rect 40577 15856 40598 15896
rect 40598 15856 40638 15896
rect 40638 15856 40663 15896
rect 40409 15833 40495 15856
rect 40577 15833 40663 15856
rect 44409 15896 44495 15919
rect 44577 15896 44663 15919
rect 44409 15856 44434 15896
rect 44434 15856 44474 15896
rect 44474 15856 44495 15896
rect 44577 15856 44598 15896
rect 44598 15856 44638 15896
rect 44638 15856 44663 15896
rect 44409 15833 44495 15856
rect 44577 15833 44663 15856
rect 48409 15896 48495 15919
rect 48577 15896 48663 15919
rect 48409 15856 48434 15896
rect 48434 15856 48474 15896
rect 48474 15856 48495 15896
rect 48577 15856 48598 15896
rect 48598 15856 48638 15896
rect 48638 15856 48663 15896
rect 48409 15833 48495 15856
rect 48577 15833 48663 15856
rect 52409 15896 52495 15919
rect 52577 15896 52663 15919
rect 52409 15856 52434 15896
rect 52434 15856 52474 15896
rect 52474 15856 52495 15896
rect 52577 15856 52598 15896
rect 52598 15856 52638 15896
rect 52638 15856 52663 15896
rect 52409 15833 52495 15856
rect 52577 15833 52663 15856
rect 56409 15896 56495 15919
rect 56577 15896 56663 15919
rect 56409 15856 56434 15896
rect 56434 15856 56474 15896
rect 56474 15856 56495 15896
rect 56577 15856 56598 15896
rect 56598 15856 56638 15896
rect 56638 15856 56663 15896
rect 56409 15833 56495 15856
rect 56577 15833 56663 15856
rect 60409 15896 60495 15919
rect 60577 15896 60663 15919
rect 60409 15856 60434 15896
rect 60434 15856 60474 15896
rect 60474 15856 60495 15896
rect 60577 15856 60598 15896
rect 60598 15856 60638 15896
rect 60638 15856 60663 15896
rect 60409 15833 60495 15856
rect 60577 15833 60663 15856
rect 64409 15896 64495 15919
rect 64577 15896 64663 15919
rect 64409 15856 64434 15896
rect 64434 15856 64474 15896
rect 64474 15856 64495 15896
rect 64577 15856 64598 15896
rect 64598 15856 64638 15896
rect 64638 15856 64663 15896
rect 64409 15833 64495 15856
rect 64577 15833 64663 15856
rect 68409 15896 68495 15919
rect 68577 15896 68663 15919
rect 68409 15856 68434 15896
rect 68434 15856 68474 15896
rect 68474 15856 68495 15896
rect 68577 15856 68598 15896
rect 68598 15856 68638 15896
rect 68638 15856 68663 15896
rect 68409 15833 68495 15856
rect 68577 15833 68663 15856
rect 72409 15896 72495 15919
rect 72577 15896 72663 15919
rect 72409 15856 72434 15896
rect 72434 15856 72474 15896
rect 72474 15856 72495 15896
rect 72577 15856 72598 15896
rect 72598 15856 72638 15896
rect 72638 15856 72663 15896
rect 72409 15833 72495 15856
rect 72577 15833 72663 15856
rect 76409 15896 76495 15919
rect 76577 15896 76663 15919
rect 76409 15856 76434 15896
rect 76434 15856 76474 15896
rect 76474 15856 76495 15896
rect 76577 15856 76598 15896
rect 76598 15856 76638 15896
rect 76638 15856 76663 15896
rect 76409 15833 76495 15856
rect 76577 15833 76663 15856
rect 80409 15896 80495 15919
rect 80577 15896 80663 15919
rect 80409 15856 80434 15896
rect 80434 15856 80474 15896
rect 80474 15856 80495 15896
rect 80577 15856 80598 15896
rect 80598 15856 80638 15896
rect 80638 15856 80663 15896
rect 80409 15833 80495 15856
rect 80577 15833 80663 15856
rect 84409 15896 84495 15919
rect 84577 15896 84663 15919
rect 84409 15856 84434 15896
rect 84434 15856 84474 15896
rect 84474 15856 84495 15896
rect 84577 15856 84598 15896
rect 84598 15856 84638 15896
rect 84638 15856 84663 15896
rect 84409 15833 84495 15856
rect 84577 15833 84663 15856
rect 88409 15896 88495 15919
rect 88577 15896 88663 15919
rect 88409 15856 88434 15896
rect 88434 15856 88474 15896
rect 88474 15856 88495 15896
rect 88577 15856 88598 15896
rect 88598 15856 88638 15896
rect 88638 15856 88663 15896
rect 88409 15833 88495 15856
rect 88577 15833 88663 15856
rect 92409 15896 92495 15919
rect 92577 15896 92663 15919
rect 92409 15856 92434 15896
rect 92434 15856 92474 15896
rect 92474 15856 92495 15896
rect 92577 15856 92598 15896
rect 92598 15856 92638 15896
rect 92638 15856 92663 15896
rect 92409 15833 92495 15856
rect 92577 15833 92663 15856
rect 96409 15896 96495 15919
rect 96577 15896 96663 15919
rect 96409 15856 96434 15896
rect 96434 15856 96474 15896
rect 96474 15856 96495 15896
rect 96577 15856 96598 15896
rect 96598 15856 96638 15896
rect 96638 15856 96663 15896
rect 96409 15833 96495 15856
rect 96577 15833 96663 15856
rect 3169 15140 3255 15163
rect 3337 15140 3423 15163
rect 3169 15100 3194 15140
rect 3194 15100 3234 15140
rect 3234 15100 3255 15140
rect 3337 15100 3358 15140
rect 3358 15100 3398 15140
rect 3398 15100 3423 15140
rect 3169 15077 3255 15100
rect 3337 15077 3423 15100
rect 7169 15140 7255 15163
rect 7337 15140 7423 15163
rect 7169 15100 7194 15140
rect 7194 15100 7234 15140
rect 7234 15100 7255 15140
rect 7337 15100 7358 15140
rect 7358 15100 7398 15140
rect 7398 15100 7423 15140
rect 7169 15077 7255 15100
rect 7337 15077 7423 15100
rect 11169 15140 11255 15163
rect 11337 15140 11423 15163
rect 11169 15100 11194 15140
rect 11194 15100 11234 15140
rect 11234 15100 11255 15140
rect 11337 15100 11358 15140
rect 11358 15100 11398 15140
rect 11398 15100 11423 15140
rect 11169 15077 11255 15100
rect 11337 15077 11423 15100
rect 15169 15140 15255 15163
rect 15337 15140 15423 15163
rect 15169 15100 15194 15140
rect 15194 15100 15234 15140
rect 15234 15100 15255 15140
rect 15337 15100 15358 15140
rect 15358 15100 15398 15140
rect 15398 15100 15423 15140
rect 15169 15077 15255 15100
rect 15337 15077 15423 15100
rect 19169 15140 19255 15163
rect 19337 15140 19423 15163
rect 19169 15100 19194 15140
rect 19194 15100 19234 15140
rect 19234 15100 19255 15140
rect 19337 15100 19358 15140
rect 19358 15100 19398 15140
rect 19398 15100 19423 15140
rect 19169 15077 19255 15100
rect 19337 15077 19423 15100
rect 23169 15140 23255 15163
rect 23337 15140 23423 15163
rect 23169 15100 23194 15140
rect 23194 15100 23234 15140
rect 23234 15100 23255 15140
rect 23337 15100 23358 15140
rect 23358 15100 23398 15140
rect 23398 15100 23423 15140
rect 23169 15077 23255 15100
rect 23337 15077 23423 15100
rect 27169 15140 27255 15163
rect 27337 15140 27423 15163
rect 27169 15100 27194 15140
rect 27194 15100 27234 15140
rect 27234 15100 27255 15140
rect 27337 15100 27358 15140
rect 27358 15100 27398 15140
rect 27398 15100 27423 15140
rect 27169 15077 27255 15100
rect 27337 15077 27423 15100
rect 31169 15140 31255 15163
rect 31337 15140 31423 15163
rect 31169 15100 31194 15140
rect 31194 15100 31234 15140
rect 31234 15100 31255 15140
rect 31337 15100 31358 15140
rect 31358 15100 31398 15140
rect 31398 15100 31423 15140
rect 31169 15077 31255 15100
rect 31337 15077 31423 15100
rect 35169 15140 35255 15163
rect 35337 15140 35423 15163
rect 35169 15100 35194 15140
rect 35194 15100 35234 15140
rect 35234 15100 35255 15140
rect 35337 15100 35358 15140
rect 35358 15100 35398 15140
rect 35398 15100 35423 15140
rect 35169 15077 35255 15100
rect 35337 15077 35423 15100
rect 39169 15140 39255 15163
rect 39337 15140 39423 15163
rect 39169 15100 39194 15140
rect 39194 15100 39234 15140
rect 39234 15100 39255 15140
rect 39337 15100 39358 15140
rect 39358 15100 39398 15140
rect 39398 15100 39423 15140
rect 39169 15077 39255 15100
rect 39337 15077 39423 15100
rect 43169 15140 43255 15163
rect 43337 15140 43423 15163
rect 43169 15100 43194 15140
rect 43194 15100 43234 15140
rect 43234 15100 43255 15140
rect 43337 15100 43358 15140
rect 43358 15100 43398 15140
rect 43398 15100 43423 15140
rect 43169 15077 43255 15100
rect 43337 15077 43423 15100
rect 47169 15140 47255 15163
rect 47337 15140 47423 15163
rect 47169 15100 47194 15140
rect 47194 15100 47234 15140
rect 47234 15100 47255 15140
rect 47337 15100 47358 15140
rect 47358 15100 47398 15140
rect 47398 15100 47423 15140
rect 47169 15077 47255 15100
rect 47337 15077 47423 15100
rect 51169 15140 51255 15163
rect 51337 15140 51423 15163
rect 51169 15100 51194 15140
rect 51194 15100 51234 15140
rect 51234 15100 51255 15140
rect 51337 15100 51358 15140
rect 51358 15100 51398 15140
rect 51398 15100 51423 15140
rect 51169 15077 51255 15100
rect 51337 15077 51423 15100
rect 55169 15140 55255 15163
rect 55337 15140 55423 15163
rect 55169 15100 55194 15140
rect 55194 15100 55234 15140
rect 55234 15100 55255 15140
rect 55337 15100 55358 15140
rect 55358 15100 55398 15140
rect 55398 15100 55423 15140
rect 55169 15077 55255 15100
rect 55337 15077 55423 15100
rect 59169 15140 59255 15163
rect 59337 15140 59423 15163
rect 59169 15100 59194 15140
rect 59194 15100 59234 15140
rect 59234 15100 59255 15140
rect 59337 15100 59358 15140
rect 59358 15100 59398 15140
rect 59398 15100 59423 15140
rect 59169 15077 59255 15100
rect 59337 15077 59423 15100
rect 63169 15140 63255 15163
rect 63337 15140 63423 15163
rect 63169 15100 63194 15140
rect 63194 15100 63234 15140
rect 63234 15100 63255 15140
rect 63337 15100 63358 15140
rect 63358 15100 63398 15140
rect 63398 15100 63423 15140
rect 63169 15077 63255 15100
rect 63337 15077 63423 15100
rect 67169 15140 67255 15163
rect 67337 15140 67423 15163
rect 67169 15100 67194 15140
rect 67194 15100 67234 15140
rect 67234 15100 67255 15140
rect 67337 15100 67358 15140
rect 67358 15100 67398 15140
rect 67398 15100 67423 15140
rect 67169 15077 67255 15100
rect 67337 15077 67423 15100
rect 4409 14384 4495 14407
rect 4577 14384 4663 14407
rect 4409 14344 4434 14384
rect 4434 14344 4474 14384
rect 4474 14344 4495 14384
rect 4577 14344 4598 14384
rect 4598 14344 4638 14384
rect 4638 14344 4663 14384
rect 4409 14321 4495 14344
rect 4577 14321 4663 14344
rect 8409 14384 8495 14407
rect 8577 14384 8663 14407
rect 8409 14344 8434 14384
rect 8434 14344 8474 14384
rect 8474 14344 8495 14384
rect 8577 14344 8598 14384
rect 8598 14344 8638 14384
rect 8638 14344 8663 14384
rect 8409 14321 8495 14344
rect 8577 14321 8663 14344
rect 12409 14384 12495 14407
rect 12577 14384 12663 14407
rect 12409 14344 12434 14384
rect 12434 14344 12474 14384
rect 12474 14344 12495 14384
rect 12577 14344 12598 14384
rect 12598 14344 12638 14384
rect 12638 14344 12663 14384
rect 12409 14321 12495 14344
rect 12577 14321 12663 14344
rect 16409 14384 16495 14407
rect 16577 14384 16663 14407
rect 16409 14344 16434 14384
rect 16434 14344 16474 14384
rect 16474 14344 16495 14384
rect 16577 14344 16598 14384
rect 16598 14344 16638 14384
rect 16638 14344 16663 14384
rect 16409 14321 16495 14344
rect 16577 14321 16663 14344
rect 20409 14384 20495 14407
rect 20577 14384 20663 14407
rect 20409 14344 20434 14384
rect 20434 14344 20474 14384
rect 20474 14344 20495 14384
rect 20577 14344 20598 14384
rect 20598 14344 20638 14384
rect 20638 14344 20663 14384
rect 20409 14321 20495 14344
rect 20577 14321 20663 14344
rect 24409 14384 24495 14407
rect 24577 14384 24663 14407
rect 24409 14344 24434 14384
rect 24434 14344 24474 14384
rect 24474 14344 24495 14384
rect 24577 14344 24598 14384
rect 24598 14344 24638 14384
rect 24638 14344 24663 14384
rect 24409 14321 24495 14344
rect 24577 14321 24663 14344
rect 28409 14384 28495 14407
rect 28577 14384 28663 14407
rect 28409 14344 28434 14384
rect 28434 14344 28474 14384
rect 28474 14344 28495 14384
rect 28577 14344 28598 14384
rect 28598 14344 28638 14384
rect 28638 14344 28663 14384
rect 28409 14321 28495 14344
rect 28577 14321 28663 14344
rect 32409 14384 32495 14407
rect 32577 14384 32663 14407
rect 32409 14344 32434 14384
rect 32434 14344 32474 14384
rect 32474 14344 32495 14384
rect 32577 14344 32598 14384
rect 32598 14344 32638 14384
rect 32638 14344 32663 14384
rect 32409 14321 32495 14344
rect 32577 14321 32663 14344
rect 36409 14384 36495 14407
rect 36577 14384 36663 14407
rect 36409 14344 36434 14384
rect 36434 14344 36474 14384
rect 36474 14344 36495 14384
rect 36577 14344 36598 14384
rect 36598 14344 36638 14384
rect 36638 14344 36663 14384
rect 36409 14321 36495 14344
rect 36577 14321 36663 14344
rect 40409 14384 40495 14407
rect 40577 14384 40663 14407
rect 40409 14344 40434 14384
rect 40434 14344 40474 14384
rect 40474 14344 40495 14384
rect 40577 14344 40598 14384
rect 40598 14344 40638 14384
rect 40638 14344 40663 14384
rect 40409 14321 40495 14344
rect 40577 14321 40663 14344
rect 44409 14384 44495 14407
rect 44577 14384 44663 14407
rect 44409 14344 44434 14384
rect 44434 14344 44474 14384
rect 44474 14344 44495 14384
rect 44577 14344 44598 14384
rect 44598 14344 44638 14384
rect 44638 14344 44663 14384
rect 44409 14321 44495 14344
rect 44577 14321 44663 14344
rect 48409 14384 48495 14407
rect 48577 14384 48663 14407
rect 48409 14344 48434 14384
rect 48434 14344 48474 14384
rect 48474 14344 48495 14384
rect 48577 14344 48598 14384
rect 48598 14344 48638 14384
rect 48638 14344 48663 14384
rect 48409 14321 48495 14344
rect 48577 14321 48663 14344
rect 52409 14384 52495 14407
rect 52577 14384 52663 14407
rect 52409 14344 52434 14384
rect 52434 14344 52474 14384
rect 52474 14344 52495 14384
rect 52577 14344 52598 14384
rect 52598 14344 52638 14384
rect 52638 14344 52663 14384
rect 52409 14321 52495 14344
rect 52577 14321 52663 14344
rect 56409 14384 56495 14407
rect 56577 14384 56663 14407
rect 56409 14344 56434 14384
rect 56434 14344 56474 14384
rect 56474 14344 56495 14384
rect 56577 14344 56598 14384
rect 56598 14344 56638 14384
rect 56638 14344 56663 14384
rect 56409 14321 56495 14344
rect 56577 14321 56663 14344
rect 60409 14384 60495 14407
rect 60577 14384 60663 14407
rect 60409 14344 60434 14384
rect 60434 14344 60474 14384
rect 60474 14344 60495 14384
rect 60577 14344 60598 14384
rect 60598 14344 60638 14384
rect 60638 14344 60663 14384
rect 60409 14321 60495 14344
rect 60577 14321 60663 14344
rect 64409 14384 64495 14407
rect 64577 14384 64663 14407
rect 64409 14344 64434 14384
rect 64434 14344 64474 14384
rect 64474 14344 64495 14384
rect 64577 14344 64598 14384
rect 64598 14344 64638 14384
rect 64638 14344 64663 14384
rect 64409 14321 64495 14344
rect 64577 14321 64663 14344
rect 68409 14384 68495 14407
rect 68577 14384 68663 14407
rect 68409 14344 68434 14384
rect 68434 14344 68474 14384
rect 68474 14344 68495 14384
rect 68577 14344 68598 14384
rect 68598 14344 68638 14384
rect 68638 14344 68663 14384
rect 68409 14321 68495 14344
rect 68577 14321 68663 14344
rect 3169 13628 3255 13651
rect 3337 13628 3423 13651
rect 3169 13588 3194 13628
rect 3194 13588 3234 13628
rect 3234 13588 3255 13628
rect 3337 13588 3358 13628
rect 3358 13588 3398 13628
rect 3398 13588 3423 13628
rect 3169 13565 3255 13588
rect 3337 13565 3423 13588
rect 7169 13628 7255 13651
rect 7337 13628 7423 13651
rect 7169 13588 7194 13628
rect 7194 13588 7234 13628
rect 7234 13588 7255 13628
rect 7337 13588 7358 13628
rect 7358 13588 7398 13628
rect 7398 13588 7423 13628
rect 7169 13565 7255 13588
rect 7337 13565 7423 13588
rect 11169 13628 11255 13651
rect 11337 13628 11423 13651
rect 11169 13588 11194 13628
rect 11194 13588 11234 13628
rect 11234 13588 11255 13628
rect 11337 13588 11358 13628
rect 11358 13588 11398 13628
rect 11398 13588 11423 13628
rect 11169 13565 11255 13588
rect 11337 13565 11423 13588
rect 15169 13628 15255 13651
rect 15337 13628 15423 13651
rect 15169 13588 15194 13628
rect 15194 13588 15234 13628
rect 15234 13588 15255 13628
rect 15337 13588 15358 13628
rect 15358 13588 15398 13628
rect 15398 13588 15423 13628
rect 15169 13565 15255 13588
rect 15337 13565 15423 13588
rect 19169 13628 19255 13651
rect 19337 13628 19423 13651
rect 19169 13588 19194 13628
rect 19194 13588 19234 13628
rect 19234 13588 19255 13628
rect 19337 13588 19358 13628
rect 19358 13588 19398 13628
rect 19398 13588 19423 13628
rect 19169 13565 19255 13588
rect 19337 13565 19423 13588
rect 23169 13628 23255 13651
rect 23337 13628 23423 13651
rect 23169 13588 23194 13628
rect 23194 13588 23234 13628
rect 23234 13588 23255 13628
rect 23337 13588 23358 13628
rect 23358 13588 23398 13628
rect 23398 13588 23423 13628
rect 23169 13565 23255 13588
rect 23337 13565 23423 13588
rect 27169 13628 27255 13651
rect 27337 13628 27423 13651
rect 27169 13588 27194 13628
rect 27194 13588 27234 13628
rect 27234 13588 27255 13628
rect 27337 13588 27358 13628
rect 27358 13588 27398 13628
rect 27398 13588 27423 13628
rect 27169 13565 27255 13588
rect 27337 13565 27423 13588
rect 31169 13628 31255 13651
rect 31337 13628 31423 13651
rect 31169 13588 31194 13628
rect 31194 13588 31234 13628
rect 31234 13588 31255 13628
rect 31337 13588 31358 13628
rect 31358 13588 31398 13628
rect 31398 13588 31423 13628
rect 31169 13565 31255 13588
rect 31337 13565 31423 13588
rect 35169 13628 35255 13651
rect 35337 13628 35423 13651
rect 35169 13588 35194 13628
rect 35194 13588 35234 13628
rect 35234 13588 35255 13628
rect 35337 13588 35358 13628
rect 35358 13588 35398 13628
rect 35398 13588 35423 13628
rect 35169 13565 35255 13588
rect 35337 13565 35423 13588
rect 39169 13628 39255 13651
rect 39337 13628 39423 13651
rect 39169 13588 39194 13628
rect 39194 13588 39234 13628
rect 39234 13588 39255 13628
rect 39337 13588 39358 13628
rect 39358 13588 39398 13628
rect 39398 13588 39423 13628
rect 39169 13565 39255 13588
rect 39337 13565 39423 13588
rect 43169 13628 43255 13651
rect 43337 13628 43423 13651
rect 43169 13588 43194 13628
rect 43194 13588 43234 13628
rect 43234 13588 43255 13628
rect 43337 13588 43358 13628
rect 43358 13588 43398 13628
rect 43398 13588 43423 13628
rect 43169 13565 43255 13588
rect 43337 13565 43423 13588
rect 47169 13628 47255 13651
rect 47337 13628 47423 13651
rect 47169 13588 47194 13628
rect 47194 13588 47234 13628
rect 47234 13588 47255 13628
rect 47337 13588 47358 13628
rect 47358 13588 47398 13628
rect 47398 13588 47423 13628
rect 47169 13565 47255 13588
rect 47337 13565 47423 13588
rect 51169 13628 51255 13651
rect 51337 13628 51423 13651
rect 51169 13588 51194 13628
rect 51194 13588 51234 13628
rect 51234 13588 51255 13628
rect 51337 13588 51358 13628
rect 51358 13588 51398 13628
rect 51398 13588 51423 13628
rect 51169 13565 51255 13588
rect 51337 13565 51423 13588
rect 55169 13628 55255 13651
rect 55337 13628 55423 13651
rect 55169 13588 55194 13628
rect 55194 13588 55234 13628
rect 55234 13588 55255 13628
rect 55337 13588 55358 13628
rect 55358 13588 55398 13628
rect 55398 13588 55423 13628
rect 55169 13565 55255 13588
rect 55337 13565 55423 13588
rect 59169 13628 59255 13651
rect 59337 13628 59423 13651
rect 59169 13588 59194 13628
rect 59194 13588 59234 13628
rect 59234 13588 59255 13628
rect 59337 13588 59358 13628
rect 59358 13588 59398 13628
rect 59398 13588 59423 13628
rect 59169 13565 59255 13588
rect 59337 13565 59423 13588
rect 63169 13628 63255 13651
rect 63337 13628 63423 13651
rect 63169 13588 63194 13628
rect 63194 13588 63234 13628
rect 63234 13588 63255 13628
rect 63337 13588 63358 13628
rect 63358 13588 63398 13628
rect 63398 13588 63423 13628
rect 63169 13565 63255 13588
rect 63337 13565 63423 13588
rect 67169 13628 67255 13651
rect 67337 13628 67423 13651
rect 67169 13588 67194 13628
rect 67194 13588 67234 13628
rect 67234 13588 67255 13628
rect 67337 13588 67358 13628
rect 67358 13588 67398 13628
rect 67398 13588 67423 13628
rect 67169 13565 67255 13588
rect 67337 13565 67423 13588
rect 72409 13036 72495 13122
rect 72577 13036 72663 13122
rect 4409 12872 4495 12895
rect 4577 12872 4663 12895
rect 4409 12832 4434 12872
rect 4434 12832 4474 12872
rect 4474 12832 4495 12872
rect 4577 12832 4598 12872
rect 4598 12832 4638 12872
rect 4638 12832 4663 12872
rect 4409 12809 4495 12832
rect 4577 12809 4663 12832
rect 8409 12872 8495 12895
rect 8577 12872 8663 12895
rect 8409 12832 8434 12872
rect 8434 12832 8474 12872
rect 8474 12832 8495 12872
rect 8577 12832 8598 12872
rect 8598 12832 8638 12872
rect 8638 12832 8663 12872
rect 8409 12809 8495 12832
rect 8577 12809 8663 12832
rect 12409 12872 12495 12895
rect 12577 12872 12663 12895
rect 12409 12832 12434 12872
rect 12434 12832 12474 12872
rect 12474 12832 12495 12872
rect 12577 12832 12598 12872
rect 12598 12832 12638 12872
rect 12638 12832 12663 12872
rect 12409 12809 12495 12832
rect 12577 12809 12663 12832
rect 16409 12872 16495 12895
rect 16577 12872 16663 12895
rect 16409 12832 16434 12872
rect 16434 12832 16474 12872
rect 16474 12832 16495 12872
rect 16577 12832 16598 12872
rect 16598 12832 16638 12872
rect 16638 12832 16663 12872
rect 16409 12809 16495 12832
rect 16577 12809 16663 12832
rect 20409 12872 20495 12895
rect 20577 12872 20663 12895
rect 20409 12832 20434 12872
rect 20434 12832 20474 12872
rect 20474 12832 20495 12872
rect 20577 12832 20598 12872
rect 20598 12832 20638 12872
rect 20638 12832 20663 12872
rect 20409 12809 20495 12832
rect 20577 12809 20663 12832
rect 24409 12872 24495 12895
rect 24577 12872 24663 12895
rect 24409 12832 24434 12872
rect 24434 12832 24474 12872
rect 24474 12832 24495 12872
rect 24577 12832 24598 12872
rect 24598 12832 24638 12872
rect 24638 12832 24663 12872
rect 24409 12809 24495 12832
rect 24577 12809 24663 12832
rect 28409 12872 28495 12895
rect 28577 12872 28663 12895
rect 28409 12832 28434 12872
rect 28434 12832 28474 12872
rect 28474 12832 28495 12872
rect 28577 12832 28598 12872
rect 28598 12832 28638 12872
rect 28638 12832 28663 12872
rect 28409 12809 28495 12832
rect 28577 12809 28663 12832
rect 32409 12872 32495 12895
rect 32577 12872 32663 12895
rect 32409 12832 32434 12872
rect 32434 12832 32474 12872
rect 32474 12832 32495 12872
rect 32577 12832 32598 12872
rect 32598 12832 32638 12872
rect 32638 12832 32663 12872
rect 32409 12809 32495 12832
rect 32577 12809 32663 12832
rect 36409 12872 36495 12895
rect 36577 12872 36663 12895
rect 36409 12832 36434 12872
rect 36434 12832 36474 12872
rect 36474 12832 36495 12872
rect 36577 12832 36598 12872
rect 36598 12832 36638 12872
rect 36638 12832 36663 12872
rect 36409 12809 36495 12832
rect 36577 12809 36663 12832
rect 40409 12872 40495 12895
rect 40577 12872 40663 12895
rect 40409 12832 40434 12872
rect 40434 12832 40474 12872
rect 40474 12832 40495 12872
rect 40577 12832 40598 12872
rect 40598 12832 40638 12872
rect 40638 12832 40663 12872
rect 40409 12809 40495 12832
rect 40577 12809 40663 12832
rect 44409 12872 44495 12895
rect 44577 12872 44663 12895
rect 44409 12832 44434 12872
rect 44434 12832 44474 12872
rect 44474 12832 44495 12872
rect 44577 12832 44598 12872
rect 44598 12832 44638 12872
rect 44638 12832 44663 12872
rect 44409 12809 44495 12832
rect 44577 12809 44663 12832
rect 48409 12872 48495 12895
rect 48577 12872 48663 12895
rect 48409 12832 48434 12872
rect 48434 12832 48474 12872
rect 48474 12832 48495 12872
rect 48577 12832 48598 12872
rect 48598 12832 48638 12872
rect 48638 12832 48663 12872
rect 48409 12809 48495 12832
rect 48577 12809 48663 12832
rect 52409 12872 52495 12895
rect 52577 12872 52663 12895
rect 52409 12832 52434 12872
rect 52434 12832 52474 12872
rect 52474 12832 52495 12872
rect 52577 12832 52598 12872
rect 52598 12832 52638 12872
rect 52638 12832 52663 12872
rect 52409 12809 52495 12832
rect 52577 12809 52663 12832
rect 56409 12872 56495 12895
rect 56577 12872 56663 12895
rect 56409 12832 56434 12872
rect 56434 12832 56474 12872
rect 56474 12832 56495 12872
rect 56577 12832 56598 12872
rect 56598 12832 56638 12872
rect 56638 12832 56663 12872
rect 56409 12809 56495 12832
rect 56577 12809 56663 12832
rect 60409 12872 60495 12895
rect 60577 12872 60663 12895
rect 60409 12832 60434 12872
rect 60434 12832 60474 12872
rect 60474 12832 60495 12872
rect 60577 12832 60598 12872
rect 60598 12832 60638 12872
rect 60638 12832 60663 12872
rect 60409 12809 60495 12832
rect 60577 12809 60663 12832
rect 64409 12872 64495 12895
rect 64577 12872 64663 12895
rect 64409 12832 64434 12872
rect 64434 12832 64474 12872
rect 64474 12832 64495 12872
rect 64577 12832 64598 12872
rect 64598 12832 64638 12872
rect 64638 12832 64663 12872
rect 64409 12809 64495 12832
rect 64577 12809 64663 12832
rect 68409 12872 68495 12895
rect 68577 12872 68663 12895
rect 68409 12832 68434 12872
rect 68434 12832 68474 12872
rect 68474 12832 68495 12872
rect 68577 12832 68598 12872
rect 68598 12832 68638 12872
rect 68638 12832 68663 12872
rect 68409 12809 68495 12832
rect 68577 12809 68663 12832
rect 72409 12868 72495 12954
rect 72577 12868 72663 12954
rect 72409 12700 72495 12786
rect 72577 12700 72663 12786
rect 72409 12532 72495 12618
rect 72577 12532 72663 12618
rect 72409 12364 72495 12450
rect 72577 12364 72663 12450
rect 72409 12196 72495 12282
rect 72577 12196 72663 12282
rect 3169 12116 3255 12139
rect 3337 12116 3423 12139
rect 3169 12076 3194 12116
rect 3194 12076 3234 12116
rect 3234 12076 3255 12116
rect 3337 12076 3358 12116
rect 3358 12076 3398 12116
rect 3398 12076 3423 12116
rect 3169 12053 3255 12076
rect 3337 12053 3423 12076
rect 7169 12116 7255 12139
rect 7337 12116 7423 12139
rect 7169 12076 7194 12116
rect 7194 12076 7234 12116
rect 7234 12076 7255 12116
rect 7337 12076 7358 12116
rect 7358 12076 7398 12116
rect 7398 12076 7423 12116
rect 7169 12053 7255 12076
rect 7337 12053 7423 12076
rect 11169 12116 11255 12139
rect 11337 12116 11423 12139
rect 11169 12076 11194 12116
rect 11194 12076 11234 12116
rect 11234 12076 11255 12116
rect 11337 12076 11358 12116
rect 11358 12076 11398 12116
rect 11398 12076 11423 12116
rect 11169 12053 11255 12076
rect 11337 12053 11423 12076
rect 15169 12116 15255 12139
rect 15337 12116 15423 12139
rect 15169 12076 15194 12116
rect 15194 12076 15234 12116
rect 15234 12076 15255 12116
rect 15337 12076 15358 12116
rect 15358 12076 15398 12116
rect 15398 12076 15423 12116
rect 15169 12053 15255 12076
rect 15337 12053 15423 12076
rect 19169 12116 19255 12139
rect 19337 12116 19423 12139
rect 19169 12076 19194 12116
rect 19194 12076 19234 12116
rect 19234 12076 19255 12116
rect 19337 12076 19358 12116
rect 19358 12076 19398 12116
rect 19398 12076 19423 12116
rect 19169 12053 19255 12076
rect 19337 12053 19423 12076
rect 23169 12116 23255 12139
rect 23337 12116 23423 12139
rect 23169 12076 23194 12116
rect 23194 12076 23234 12116
rect 23234 12076 23255 12116
rect 23337 12076 23358 12116
rect 23358 12076 23398 12116
rect 23398 12076 23423 12116
rect 23169 12053 23255 12076
rect 23337 12053 23423 12076
rect 27169 12116 27255 12139
rect 27337 12116 27423 12139
rect 27169 12076 27194 12116
rect 27194 12076 27234 12116
rect 27234 12076 27255 12116
rect 27337 12076 27358 12116
rect 27358 12076 27398 12116
rect 27398 12076 27423 12116
rect 27169 12053 27255 12076
rect 27337 12053 27423 12076
rect 31169 12116 31255 12139
rect 31337 12116 31423 12139
rect 31169 12076 31194 12116
rect 31194 12076 31234 12116
rect 31234 12076 31255 12116
rect 31337 12076 31358 12116
rect 31358 12076 31398 12116
rect 31398 12076 31423 12116
rect 31169 12053 31255 12076
rect 31337 12053 31423 12076
rect 35169 12116 35255 12139
rect 35337 12116 35423 12139
rect 35169 12076 35194 12116
rect 35194 12076 35234 12116
rect 35234 12076 35255 12116
rect 35337 12076 35358 12116
rect 35358 12076 35398 12116
rect 35398 12076 35423 12116
rect 35169 12053 35255 12076
rect 35337 12053 35423 12076
rect 39169 12116 39255 12139
rect 39337 12116 39423 12139
rect 39169 12076 39194 12116
rect 39194 12076 39234 12116
rect 39234 12076 39255 12116
rect 39337 12076 39358 12116
rect 39358 12076 39398 12116
rect 39398 12076 39423 12116
rect 39169 12053 39255 12076
rect 39337 12053 39423 12076
rect 43169 12116 43255 12139
rect 43337 12116 43423 12139
rect 43169 12076 43194 12116
rect 43194 12076 43234 12116
rect 43234 12076 43255 12116
rect 43337 12076 43358 12116
rect 43358 12076 43398 12116
rect 43398 12076 43423 12116
rect 43169 12053 43255 12076
rect 43337 12053 43423 12076
rect 47169 12116 47255 12139
rect 47337 12116 47423 12139
rect 47169 12076 47194 12116
rect 47194 12076 47234 12116
rect 47234 12076 47255 12116
rect 47337 12076 47358 12116
rect 47358 12076 47398 12116
rect 47398 12076 47423 12116
rect 47169 12053 47255 12076
rect 47337 12053 47423 12076
rect 51169 12116 51255 12139
rect 51337 12116 51423 12139
rect 51169 12076 51194 12116
rect 51194 12076 51234 12116
rect 51234 12076 51255 12116
rect 51337 12076 51358 12116
rect 51358 12076 51398 12116
rect 51398 12076 51423 12116
rect 51169 12053 51255 12076
rect 51337 12053 51423 12076
rect 55169 12116 55255 12139
rect 55337 12116 55423 12139
rect 55169 12076 55194 12116
rect 55194 12076 55234 12116
rect 55234 12076 55255 12116
rect 55337 12076 55358 12116
rect 55358 12076 55398 12116
rect 55398 12076 55423 12116
rect 55169 12053 55255 12076
rect 55337 12053 55423 12076
rect 59169 12116 59255 12139
rect 59337 12116 59423 12139
rect 59169 12076 59194 12116
rect 59194 12076 59234 12116
rect 59234 12076 59255 12116
rect 59337 12076 59358 12116
rect 59358 12076 59398 12116
rect 59398 12076 59423 12116
rect 59169 12053 59255 12076
rect 59337 12053 59423 12076
rect 63169 12116 63255 12139
rect 63337 12116 63423 12139
rect 63169 12076 63194 12116
rect 63194 12076 63234 12116
rect 63234 12076 63255 12116
rect 63337 12076 63358 12116
rect 63358 12076 63398 12116
rect 63398 12076 63423 12116
rect 63169 12053 63255 12076
rect 63337 12053 63423 12076
rect 67169 12116 67255 12139
rect 67337 12116 67423 12139
rect 67169 12076 67194 12116
rect 67194 12076 67234 12116
rect 67234 12076 67255 12116
rect 67337 12076 67358 12116
rect 67358 12076 67398 12116
rect 67398 12076 67423 12116
rect 67169 12053 67255 12076
rect 67337 12053 67423 12076
rect 72409 12028 72495 12114
rect 72577 12028 72663 12114
rect 72409 11860 72495 11946
rect 72577 11860 72663 11946
rect 72409 11692 72495 11778
rect 72577 11692 72663 11778
rect 72409 11524 72495 11610
rect 72577 11524 72663 11610
rect 4409 11360 4495 11383
rect 4577 11360 4663 11383
rect 4409 11320 4434 11360
rect 4434 11320 4474 11360
rect 4474 11320 4495 11360
rect 4577 11320 4598 11360
rect 4598 11320 4638 11360
rect 4638 11320 4663 11360
rect 4409 11297 4495 11320
rect 4577 11297 4663 11320
rect 8409 11360 8495 11383
rect 8577 11360 8663 11383
rect 8409 11320 8434 11360
rect 8434 11320 8474 11360
rect 8474 11320 8495 11360
rect 8577 11320 8598 11360
rect 8598 11320 8638 11360
rect 8638 11320 8663 11360
rect 8409 11297 8495 11320
rect 8577 11297 8663 11320
rect 12409 11360 12495 11383
rect 12577 11360 12663 11383
rect 12409 11320 12434 11360
rect 12434 11320 12474 11360
rect 12474 11320 12495 11360
rect 12577 11320 12598 11360
rect 12598 11320 12638 11360
rect 12638 11320 12663 11360
rect 12409 11297 12495 11320
rect 12577 11297 12663 11320
rect 16409 11360 16495 11383
rect 16577 11360 16663 11383
rect 16409 11320 16434 11360
rect 16434 11320 16474 11360
rect 16474 11320 16495 11360
rect 16577 11320 16598 11360
rect 16598 11320 16638 11360
rect 16638 11320 16663 11360
rect 16409 11297 16495 11320
rect 16577 11297 16663 11320
rect 20409 11360 20495 11383
rect 20577 11360 20663 11383
rect 20409 11320 20434 11360
rect 20434 11320 20474 11360
rect 20474 11320 20495 11360
rect 20577 11320 20598 11360
rect 20598 11320 20638 11360
rect 20638 11320 20663 11360
rect 20409 11297 20495 11320
rect 20577 11297 20663 11320
rect 24409 11360 24495 11383
rect 24577 11360 24663 11383
rect 24409 11320 24434 11360
rect 24434 11320 24474 11360
rect 24474 11320 24495 11360
rect 24577 11320 24598 11360
rect 24598 11320 24638 11360
rect 24638 11320 24663 11360
rect 24409 11297 24495 11320
rect 24577 11297 24663 11320
rect 28409 11360 28495 11383
rect 28577 11360 28663 11383
rect 28409 11320 28434 11360
rect 28434 11320 28474 11360
rect 28474 11320 28495 11360
rect 28577 11320 28598 11360
rect 28598 11320 28638 11360
rect 28638 11320 28663 11360
rect 28409 11297 28495 11320
rect 28577 11297 28663 11320
rect 32409 11360 32495 11383
rect 32577 11360 32663 11383
rect 32409 11320 32434 11360
rect 32434 11320 32474 11360
rect 32474 11320 32495 11360
rect 32577 11320 32598 11360
rect 32598 11320 32638 11360
rect 32638 11320 32663 11360
rect 32409 11297 32495 11320
rect 32577 11297 32663 11320
rect 36409 11360 36495 11383
rect 36577 11360 36663 11383
rect 36409 11320 36434 11360
rect 36434 11320 36474 11360
rect 36474 11320 36495 11360
rect 36577 11320 36598 11360
rect 36598 11320 36638 11360
rect 36638 11320 36663 11360
rect 36409 11297 36495 11320
rect 36577 11297 36663 11320
rect 40409 11360 40495 11383
rect 40577 11360 40663 11383
rect 40409 11320 40434 11360
rect 40434 11320 40474 11360
rect 40474 11320 40495 11360
rect 40577 11320 40598 11360
rect 40598 11320 40638 11360
rect 40638 11320 40663 11360
rect 40409 11297 40495 11320
rect 40577 11297 40663 11320
rect 44409 11360 44495 11383
rect 44577 11360 44663 11383
rect 44409 11320 44434 11360
rect 44434 11320 44474 11360
rect 44474 11320 44495 11360
rect 44577 11320 44598 11360
rect 44598 11320 44638 11360
rect 44638 11320 44663 11360
rect 44409 11297 44495 11320
rect 44577 11297 44663 11320
rect 48409 11360 48495 11383
rect 48577 11360 48663 11383
rect 48409 11320 48434 11360
rect 48434 11320 48474 11360
rect 48474 11320 48495 11360
rect 48577 11320 48598 11360
rect 48598 11320 48638 11360
rect 48638 11320 48663 11360
rect 48409 11297 48495 11320
rect 48577 11297 48663 11320
rect 52409 11360 52495 11383
rect 52577 11360 52663 11383
rect 52409 11320 52434 11360
rect 52434 11320 52474 11360
rect 52474 11320 52495 11360
rect 52577 11320 52598 11360
rect 52598 11320 52638 11360
rect 52638 11320 52663 11360
rect 52409 11297 52495 11320
rect 52577 11297 52663 11320
rect 56409 11360 56495 11383
rect 56577 11360 56663 11383
rect 56409 11320 56434 11360
rect 56434 11320 56474 11360
rect 56474 11320 56495 11360
rect 56577 11320 56598 11360
rect 56598 11320 56638 11360
rect 56638 11320 56663 11360
rect 56409 11297 56495 11320
rect 56577 11297 56663 11320
rect 60409 11360 60495 11383
rect 60577 11360 60663 11383
rect 60409 11320 60434 11360
rect 60434 11320 60474 11360
rect 60474 11320 60495 11360
rect 60577 11320 60598 11360
rect 60598 11320 60638 11360
rect 60638 11320 60663 11360
rect 60409 11297 60495 11320
rect 60577 11297 60663 11320
rect 64409 11360 64495 11383
rect 64577 11360 64663 11383
rect 64409 11320 64434 11360
rect 64434 11320 64474 11360
rect 64474 11320 64495 11360
rect 64577 11320 64598 11360
rect 64598 11320 64638 11360
rect 64638 11320 64663 11360
rect 64409 11297 64495 11320
rect 64577 11297 64663 11320
rect 68409 11360 68495 11383
rect 68577 11360 68663 11383
rect 68409 11320 68434 11360
rect 68434 11320 68474 11360
rect 68474 11320 68495 11360
rect 68577 11320 68598 11360
rect 68598 11320 68638 11360
rect 68638 11320 68663 11360
rect 68409 11297 68495 11320
rect 68577 11297 68663 11320
rect 72409 11356 72495 11442
rect 72577 11356 72663 11442
rect 72409 11188 72495 11274
rect 72577 11188 72663 11274
rect 72409 11020 72495 11106
rect 72577 11020 72663 11106
rect 76409 13036 76495 13122
rect 76577 13036 76663 13122
rect 76409 12868 76495 12954
rect 76577 12868 76663 12954
rect 76409 12700 76495 12786
rect 76577 12700 76663 12786
rect 76409 12532 76495 12618
rect 76577 12532 76663 12618
rect 76409 12364 76495 12450
rect 76577 12364 76663 12450
rect 76409 12196 76495 12282
rect 76577 12196 76663 12282
rect 76409 12028 76495 12114
rect 76577 12028 76663 12114
rect 76409 11860 76495 11946
rect 76577 11860 76663 11946
rect 76409 11692 76495 11778
rect 76577 11692 76663 11778
rect 76409 11524 76495 11610
rect 76577 11524 76663 11610
rect 76409 11356 76495 11442
rect 76577 11356 76663 11442
rect 76409 11188 76495 11274
rect 76577 11188 76663 11274
rect 76409 11020 76495 11106
rect 76577 11020 76663 11106
rect 80409 13036 80495 13122
rect 80577 13036 80663 13122
rect 80409 12868 80495 12954
rect 80577 12868 80663 12954
rect 80409 12700 80495 12786
rect 80577 12700 80663 12786
rect 80409 12532 80495 12618
rect 80577 12532 80663 12618
rect 80409 12364 80495 12450
rect 80577 12364 80663 12450
rect 80409 12196 80495 12282
rect 80577 12196 80663 12282
rect 80409 12028 80495 12114
rect 80577 12028 80663 12114
rect 80409 11860 80495 11946
rect 80577 11860 80663 11946
rect 80409 11692 80495 11778
rect 80577 11692 80663 11778
rect 80409 11524 80495 11610
rect 80577 11524 80663 11610
rect 80409 11356 80495 11442
rect 80577 11356 80663 11442
rect 80409 11188 80495 11274
rect 80577 11188 80663 11274
rect 80409 11020 80495 11106
rect 80577 11020 80663 11106
rect 84409 13036 84495 13122
rect 84577 13036 84663 13122
rect 84409 12868 84495 12954
rect 84577 12868 84663 12954
rect 84409 12700 84495 12786
rect 84577 12700 84663 12786
rect 84409 12532 84495 12618
rect 84577 12532 84663 12618
rect 84409 12364 84495 12450
rect 84577 12364 84663 12450
rect 84409 12196 84495 12282
rect 84577 12196 84663 12282
rect 84409 12028 84495 12114
rect 84577 12028 84663 12114
rect 84409 11860 84495 11946
rect 84577 11860 84663 11946
rect 84409 11692 84495 11778
rect 84577 11692 84663 11778
rect 84409 11524 84495 11610
rect 84577 11524 84663 11610
rect 84409 11356 84495 11442
rect 84577 11356 84663 11442
rect 84409 11188 84495 11274
rect 84577 11188 84663 11274
rect 84409 11020 84495 11106
rect 84577 11020 84663 11106
rect 88409 13036 88495 13122
rect 88577 13036 88663 13122
rect 88409 12868 88495 12954
rect 88577 12868 88663 12954
rect 88409 12700 88495 12786
rect 88577 12700 88663 12786
rect 88409 12532 88495 12618
rect 88577 12532 88663 12618
rect 88409 12364 88495 12450
rect 88577 12364 88663 12450
rect 88409 12196 88495 12282
rect 88577 12196 88663 12282
rect 88409 12028 88495 12114
rect 88577 12028 88663 12114
rect 88409 11860 88495 11946
rect 88577 11860 88663 11946
rect 88409 11692 88495 11778
rect 88577 11692 88663 11778
rect 88409 11524 88495 11610
rect 88577 11524 88663 11610
rect 88409 11356 88495 11442
rect 88577 11356 88663 11442
rect 88409 11188 88495 11274
rect 88577 11188 88663 11274
rect 88409 11020 88495 11106
rect 88577 11020 88663 11106
rect 92409 13036 92495 13122
rect 92577 13036 92663 13122
rect 92409 12868 92495 12954
rect 92577 12868 92663 12954
rect 92409 12700 92495 12786
rect 92577 12700 92663 12786
rect 92409 12532 92495 12618
rect 92577 12532 92663 12618
rect 92409 12364 92495 12450
rect 92577 12364 92663 12450
rect 92409 12196 92495 12282
rect 92577 12196 92663 12282
rect 92409 12028 92495 12114
rect 92577 12028 92663 12114
rect 92409 11860 92495 11946
rect 92577 11860 92663 11946
rect 92409 11692 92495 11778
rect 92577 11692 92663 11778
rect 92409 11524 92495 11610
rect 92577 11524 92663 11610
rect 92409 11356 92495 11442
rect 92577 11356 92663 11442
rect 92409 11188 92495 11274
rect 92577 11188 92663 11274
rect 92409 11020 92495 11106
rect 92577 11020 92663 11106
rect 96409 13036 96495 13122
rect 96577 13036 96663 13122
rect 96409 12868 96495 12954
rect 96577 12868 96663 12954
rect 96409 12700 96495 12786
rect 96577 12700 96663 12786
rect 96409 12532 96495 12618
rect 96577 12532 96663 12618
rect 96409 12364 96495 12450
rect 96577 12364 96663 12450
rect 96409 12196 96495 12282
rect 96577 12196 96663 12282
rect 96409 12028 96495 12114
rect 96577 12028 96663 12114
rect 96409 11860 96495 11946
rect 96577 11860 96663 11946
rect 96409 11692 96495 11778
rect 96577 11692 96663 11778
rect 96409 11524 96495 11610
rect 96577 11524 96663 11610
rect 96409 11356 96495 11442
rect 96577 11356 96663 11442
rect 96409 11188 96495 11274
rect 96577 11188 96663 11274
rect 96409 11020 96495 11106
rect 96577 11020 96663 11106
rect 3169 10604 3255 10627
rect 3337 10604 3423 10627
rect 3169 10564 3194 10604
rect 3194 10564 3234 10604
rect 3234 10564 3255 10604
rect 3337 10564 3358 10604
rect 3358 10564 3398 10604
rect 3398 10564 3423 10604
rect 3169 10541 3255 10564
rect 3337 10541 3423 10564
rect 7169 10604 7255 10627
rect 7337 10604 7423 10627
rect 7169 10564 7194 10604
rect 7194 10564 7234 10604
rect 7234 10564 7255 10604
rect 7337 10564 7358 10604
rect 7358 10564 7398 10604
rect 7398 10564 7423 10604
rect 7169 10541 7255 10564
rect 7337 10541 7423 10564
rect 11169 10604 11255 10627
rect 11337 10604 11423 10627
rect 11169 10564 11194 10604
rect 11194 10564 11234 10604
rect 11234 10564 11255 10604
rect 11337 10564 11358 10604
rect 11358 10564 11398 10604
rect 11398 10564 11423 10604
rect 11169 10541 11255 10564
rect 11337 10541 11423 10564
rect 15169 10604 15255 10627
rect 15337 10604 15423 10627
rect 15169 10564 15194 10604
rect 15194 10564 15234 10604
rect 15234 10564 15255 10604
rect 15337 10564 15358 10604
rect 15358 10564 15398 10604
rect 15398 10564 15423 10604
rect 15169 10541 15255 10564
rect 15337 10541 15423 10564
rect 19169 10604 19255 10627
rect 19337 10604 19423 10627
rect 19169 10564 19194 10604
rect 19194 10564 19234 10604
rect 19234 10564 19255 10604
rect 19337 10564 19358 10604
rect 19358 10564 19398 10604
rect 19398 10564 19423 10604
rect 19169 10541 19255 10564
rect 19337 10541 19423 10564
rect 23169 10604 23255 10627
rect 23337 10604 23423 10627
rect 23169 10564 23194 10604
rect 23194 10564 23234 10604
rect 23234 10564 23255 10604
rect 23337 10564 23358 10604
rect 23358 10564 23398 10604
rect 23398 10564 23423 10604
rect 23169 10541 23255 10564
rect 23337 10541 23423 10564
rect 27169 10604 27255 10627
rect 27337 10604 27423 10627
rect 27169 10564 27194 10604
rect 27194 10564 27234 10604
rect 27234 10564 27255 10604
rect 27337 10564 27358 10604
rect 27358 10564 27398 10604
rect 27398 10564 27423 10604
rect 27169 10541 27255 10564
rect 27337 10541 27423 10564
rect 31169 10604 31255 10627
rect 31337 10604 31423 10627
rect 31169 10564 31194 10604
rect 31194 10564 31234 10604
rect 31234 10564 31255 10604
rect 31337 10564 31358 10604
rect 31358 10564 31398 10604
rect 31398 10564 31423 10604
rect 31169 10541 31255 10564
rect 31337 10541 31423 10564
rect 35169 10604 35255 10627
rect 35337 10604 35423 10627
rect 35169 10564 35194 10604
rect 35194 10564 35234 10604
rect 35234 10564 35255 10604
rect 35337 10564 35358 10604
rect 35358 10564 35398 10604
rect 35398 10564 35423 10604
rect 35169 10541 35255 10564
rect 35337 10541 35423 10564
rect 39169 10604 39255 10627
rect 39337 10604 39423 10627
rect 39169 10564 39194 10604
rect 39194 10564 39234 10604
rect 39234 10564 39255 10604
rect 39337 10564 39358 10604
rect 39358 10564 39398 10604
rect 39398 10564 39423 10604
rect 39169 10541 39255 10564
rect 39337 10541 39423 10564
rect 43169 10604 43255 10627
rect 43337 10604 43423 10627
rect 43169 10564 43194 10604
rect 43194 10564 43234 10604
rect 43234 10564 43255 10604
rect 43337 10564 43358 10604
rect 43358 10564 43398 10604
rect 43398 10564 43423 10604
rect 43169 10541 43255 10564
rect 43337 10541 43423 10564
rect 47169 10604 47255 10627
rect 47337 10604 47423 10627
rect 47169 10564 47194 10604
rect 47194 10564 47234 10604
rect 47234 10564 47255 10604
rect 47337 10564 47358 10604
rect 47358 10564 47398 10604
rect 47398 10564 47423 10604
rect 47169 10541 47255 10564
rect 47337 10541 47423 10564
rect 51169 10604 51255 10627
rect 51337 10604 51423 10627
rect 51169 10564 51194 10604
rect 51194 10564 51234 10604
rect 51234 10564 51255 10604
rect 51337 10564 51358 10604
rect 51358 10564 51398 10604
rect 51398 10564 51423 10604
rect 51169 10541 51255 10564
rect 51337 10541 51423 10564
rect 55169 10604 55255 10627
rect 55337 10604 55423 10627
rect 55169 10564 55194 10604
rect 55194 10564 55234 10604
rect 55234 10564 55255 10604
rect 55337 10564 55358 10604
rect 55358 10564 55398 10604
rect 55398 10564 55423 10604
rect 55169 10541 55255 10564
rect 55337 10541 55423 10564
rect 59169 10604 59255 10627
rect 59337 10604 59423 10627
rect 59169 10564 59194 10604
rect 59194 10564 59234 10604
rect 59234 10564 59255 10604
rect 59337 10564 59358 10604
rect 59358 10564 59398 10604
rect 59398 10564 59423 10604
rect 59169 10541 59255 10564
rect 59337 10541 59423 10564
rect 63169 10604 63255 10627
rect 63337 10604 63423 10627
rect 63169 10564 63194 10604
rect 63194 10564 63234 10604
rect 63234 10564 63255 10604
rect 63337 10564 63358 10604
rect 63358 10564 63398 10604
rect 63398 10564 63423 10604
rect 63169 10541 63255 10564
rect 63337 10541 63423 10564
rect 67169 10604 67255 10627
rect 67337 10604 67423 10627
rect 67169 10564 67194 10604
rect 67194 10564 67234 10604
rect 67234 10564 67255 10604
rect 67337 10564 67358 10604
rect 67358 10564 67398 10604
rect 67398 10564 67423 10604
rect 67169 10541 67255 10564
rect 67337 10541 67423 10564
rect 75169 10160 75255 10246
rect 75337 10160 75423 10246
rect 75169 9992 75255 10078
rect 75337 9992 75423 10078
rect 4409 9848 4495 9871
rect 4577 9848 4663 9871
rect 4409 9808 4434 9848
rect 4434 9808 4474 9848
rect 4474 9808 4495 9848
rect 4577 9808 4598 9848
rect 4598 9808 4638 9848
rect 4638 9808 4663 9848
rect 4409 9785 4495 9808
rect 4577 9785 4663 9808
rect 8409 9848 8495 9871
rect 8577 9848 8663 9871
rect 8409 9808 8434 9848
rect 8434 9808 8474 9848
rect 8474 9808 8495 9848
rect 8577 9808 8598 9848
rect 8598 9808 8638 9848
rect 8638 9808 8663 9848
rect 8409 9785 8495 9808
rect 8577 9785 8663 9808
rect 12409 9848 12495 9871
rect 12577 9848 12663 9871
rect 12409 9808 12434 9848
rect 12434 9808 12474 9848
rect 12474 9808 12495 9848
rect 12577 9808 12598 9848
rect 12598 9808 12638 9848
rect 12638 9808 12663 9848
rect 12409 9785 12495 9808
rect 12577 9785 12663 9808
rect 16409 9848 16495 9871
rect 16577 9848 16663 9871
rect 16409 9808 16434 9848
rect 16434 9808 16474 9848
rect 16474 9808 16495 9848
rect 16577 9808 16598 9848
rect 16598 9808 16638 9848
rect 16638 9808 16663 9848
rect 16409 9785 16495 9808
rect 16577 9785 16663 9808
rect 20409 9848 20495 9871
rect 20577 9848 20663 9871
rect 20409 9808 20434 9848
rect 20434 9808 20474 9848
rect 20474 9808 20495 9848
rect 20577 9808 20598 9848
rect 20598 9808 20638 9848
rect 20638 9808 20663 9848
rect 20409 9785 20495 9808
rect 20577 9785 20663 9808
rect 24409 9848 24495 9871
rect 24577 9848 24663 9871
rect 24409 9808 24434 9848
rect 24434 9808 24474 9848
rect 24474 9808 24495 9848
rect 24577 9808 24598 9848
rect 24598 9808 24638 9848
rect 24638 9808 24663 9848
rect 24409 9785 24495 9808
rect 24577 9785 24663 9808
rect 28409 9848 28495 9871
rect 28577 9848 28663 9871
rect 28409 9808 28434 9848
rect 28434 9808 28474 9848
rect 28474 9808 28495 9848
rect 28577 9808 28598 9848
rect 28598 9808 28638 9848
rect 28638 9808 28663 9848
rect 28409 9785 28495 9808
rect 28577 9785 28663 9808
rect 32409 9848 32495 9871
rect 32577 9848 32663 9871
rect 32409 9808 32434 9848
rect 32434 9808 32474 9848
rect 32474 9808 32495 9848
rect 32577 9808 32598 9848
rect 32598 9808 32638 9848
rect 32638 9808 32663 9848
rect 32409 9785 32495 9808
rect 32577 9785 32663 9808
rect 36409 9848 36495 9871
rect 36577 9848 36663 9871
rect 36409 9808 36434 9848
rect 36434 9808 36474 9848
rect 36474 9808 36495 9848
rect 36577 9808 36598 9848
rect 36598 9808 36638 9848
rect 36638 9808 36663 9848
rect 36409 9785 36495 9808
rect 36577 9785 36663 9808
rect 40409 9848 40495 9871
rect 40577 9848 40663 9871
rect 40409 9808 40434 9848
rect 40434 9808 40474 9848
rect 40474 9808 40495 9848
rect 40577 9808 40598 9848
rect 40598 9808 40638 9848
rect 40638 9808 40663 9848
rect 40409 9785 40495 9808
rect 40577 9785 40663 9808
rect 44409 9848 44495 9871
rect 44577 9848 44663 9871
rect 44409 9808 44434 9848
rect 44434 9808 44474 9848
rect 44474 9808 44495 9848
rect 44577 9808 44598 9848
rect 44598 9808 44638 9848
rect 44638 9808 44663 9848
rect 44409 9785 44495 9808
rect 44577 9785 44663 9808
rect 48409 9848 48495 9871
rect 48577 9848 48663 9871
rect 48409 9808 48434 9848
rect 48434 9808 48474 9848
rect 48474 9808 48495 9848
rect 48577 9808 48598 9848
rect 48598 9808 48638 9848
rect 48638 9808 48663 9848
rect 48409 9785 48495 9808
rect 48577 9785 48663 9808
rect 52409 9848 52495 9871
rect 52577 9848 52663 9871
rect 52409 9808 52434 9848
rect 52434 9808 52474 9848
rect 52474 9808 52495 9848
rect 52577 9808 52598 9848
rect 52598 9808 52638 9848
rect 52638 9808 52663 9848
rect 52409 9785 52495 9808
rect 52577 9785 52663 9808
rect 56409 9848 56495 9871
rect 56577 9848 56663 9871
rect 56409 9808 56434 9848
rect 56434 9808 56474 9848
rect 56474 9808 56495 9848
rect 56577 9808 56598 9848
rect 56598 9808 56638 9848
rect 56638 9808 56663 9848
rect 56409 9785 56495 9808
rect 56577 9785 56663 9808
rect 60409 9848 60495 9871
rect 60577 9848 60663 9871
rect 60409 9808 60434 9848
rect 60434 9808 60474 9848
rect 60474 9808 60495 9848
rect 60577 9808 60598 9848
rect 60598 9808 60638 9848
rect 60638 9808 60663 9848
rect 60409 9785 60495 9808
rect 60577 9785 60663 9808
rect 64409 9848 64495 9871
rect 64577 9848 64663 9871
rect 64409 9808 64434 9848
rect 64434 9808 64474 9848
rect 64474 9808 64495 9848
rect 64577 9808 64598 9848
rect 64598 9808 64638 9848
rect 64638 9808 64663 9848
rect 64409 9785 64495 9808
rect 64577 9785 64663 9808
rect 68409 9848 68495 9871
rect 68577 9848 68663 9871
rect 68409 9808 68434 9848
rect 68434 9808 68474 9848
rect 68474 9808 68495 9848
rect 68577 9808 68598 9848
rect 68598 9808 68638 9848
rect 68638 9808 68663 9848
rect 68409 9785 68495 9808
rect 68577 9785 68663 9808
rect 75169 9824 75255 9910
rect 75337 9824 75423 9910
rect 75169 9656 75255 9742
rect 75337 9656 75423 9742
rect 75169 9488 75255 9574
rect 75337 9488 75423 9574
rect 75169 9320 75255 9406
rect 75337 9320 75423 9406
rect 75169 9152 75255 9238
rect 75337 9152 75423 9238
rect 3169 9092 3255 9115
rect 3337 9092 3423 9115
rect 3169 9052 3194 9092
rect 3194 9052 3234 9092
rect 3234 9052 3255 9092
rect 3337 9052 3358 9092
rect 3358 9052 3398 9092
rect 3398 9052 3423 9092
rect 3169 9029 3255 9052
rect 3337 9029 3423 9052
rect 7169 9092 7255 9115
rect 7337 9092 7423 9115
rect 7169 9052 7194 9092
rect 7194 9052 7234 9092
rect 7234 9052 7255 9092
rect 7337 9052 7358 9092
rect 7358 9052 7398 9092
rect 7398 9052 7423 9092
rect 7169 9029 7255 9052
rect 7337 9029 7423 9052
rect 11169 9092 11255 9115
rect 11337 9092 11423 9115
rect 11169 9052 11194 9092
rect 11194 9052 11234 9092
rect 11234 9052 11255 9092
rect 11337 9052 11358 9092
rect 11358 9052 11398 9092
rect 11398 9052 11423 9092
rect 11169 9029 11255 9052
rect 11337 9029 11423 9052
rect 15169 9092 15255 9115
rect 15337 9092 15423 9115
rect 15169 9052 15194 9092
rect 15194 9052 15234 9092
rect 15234 9052 15255 9092
rect 15337 9052 15358 9092
rect 15358 9052 15398 9092
rect 15398 9052 15423 9092
rect 15169 9029 15255 9052
rect 15337 9029 15423 9052
rect 19169 9092 19255 9115
rect 19337 9092 19423 9115
rect 19169 9052 19194 9092
rect 19194 9052 19234 9092
rect 19234 9052 19255 9092
rect 19337 9052 19358 9092
rect 19358 9052 19398 9092
rect 19398 9052 19423 9092
rect 19169 9029 19255 9052
rect 19337 9029 19423 9052
rect 23169 9092 23255 9115
rect 23337 9092 23423 9115
rect 23169 9052 23194 9092
rect 23194 9052 23234 9092
rect 23234 9052 23255 9092
rect 23337 9052 23358 9092
rect 23358 9052 23398 9092
rect 23398 9052 23423 9092
rect 23169 9029 23255 9052
rect 23337 9029 23423 9052
rect 27169 9092 27255 9115
rect 27337 9092 27423 9115
rect 27169 9052 27194 9092
rect 27194 9052 27234 9092
rect 27234 9052 27255 9092
rect 27337 9052 27358 9092
rect 27358 9052 27398 9092
rect 27398 9052 27423 9092
rect 27169 9029 27255 9052
rect 27337 9029 27423 9052
rect 31169 9092 31255 9115
rect 31337 9092 31423 9115
rect 31169 9052 31194 9092
rect 31194 9052 31234 9092
rect 31234 9052 31255 9092
rect 31337 9052 31358 9092
rect 31358 9052 31398 9092
rect 31398 9052 31423 9092
rect 31169 9029 31255 9052
rect 31337 9029 31423 9052
rect 35169 9092 35255 9115
rect 35337 9092 35423 9115
rect 35169 9052 35194 9092
rect 35194 9052 35234 9092
rect 35234 9052 35255 9092
rect 35337 9052 35358 9092
rect 35358 9052 35398 9092
rect 35398 9052 35423 9092
rect 35169 9029 35255 9052
rect 35337 9029 35423 9052
rect 39169 9092 39255 9115
rect 39337 9092 39423 9115
rect 39169 9052 39194 9092
rect 39194 9052 39234 9092
rect 39234 9052 39255 9092
rect 39337 9052 39358 9092
rect 39358 9052 39398 9092
rect 39398 9052 39423 9092
rect 39169 9029 39255 9052
rect 39337 9029 39423 9052
rect 43169 9092 43255 9115
rect 43337 9092 43423 9115
rect 43169 9052 43194 9092
rect 43194 9052 43234 9092
rect 43234 9052 43255 9092
rect 43337 9052 43358 9092
rect 43358 9052 43398 9092
rect 43398 9052 43423 9092
rect 43169 9029 43255 9052
rect 43337 9029 43423 9052
rect 47169 9092 47255 9115
rect 47337 9092 47423 9115
rect 47169 9052 47194 9092
rect 47194 9052 47234 9092
rect 47234 9052 47255 9092
rect 47337 9052 47358 9092
rect 47358 9052 47398 9092
rect 47398 9052 47423 9092
rect 47169 9029 47255 9052
rect 47337 9029 47423 9052
rect 51169 9092 51255 9115
rect 51337 9092 51423 9115
rect 51169 9052 51194 9092
rect 51194 9052 51234 9092
rect 51234 9052 51255 9092
rect 51337 9052 51358 9092
rect 51358 9052 51398 9092
rect 51398 9052 51423 9092
rect 51169 9029 51255 9052
rect 51337 9029 51423 9052
rect 55169 9092 55255 9115
rect 55337 9092 55423 9115
rect 55169 9052 55194 9092
rect 55194 9052 55234 9092
rect 55234 9052 55255 9092
rect 55337 9052 55358 9092
rect 55358 9052 55398 9092
rect 55398 9052 55423 9092
rect 55169 9029 55255 9052
rect 55337 9029 55423 9052
rect 59169 9092 59255 9115
rect 59337 9092 59423 9115
rect 59169 9052 59194 9092
rect 59194 9052 59234 9092
rect 59234 9052 59255 9092
rect 59337 9052 59358 9092
rect 59358 9052 59398 9092
rect 59398 9052 59423 9092
rect 59169 9029 59255 9052
rect 59337 9029 59423 9052
rect 63169 9092 63255 9115
rect 63337 9092 63423 9115
rect 63169 9052 63194 9092
rect 63194 9052 63234 9092
rect 63234 9052 63255 9092
rect 63337 9052 63358 9092
rect 63358 9052 63398 9092
rect 63398 9052 63423 9092
rect 63169 9029 63255 9052
rect 63337 9029 63423 9052
rect 67169 9092 67255 9115
rect 67337 9092 67423 9115
rect 67169 9052 67194 9092
rect 67194 9052 67234 9092
rect 67234 9052 67255 9092
rect 67337 9052 67358 9092
rect 67358 9052 67398 9092
rect 67398 9052 67423 9092
rect 67169 9029 67255 9052
rect 67337 9029 67423 9052
rect 75169 8984 75255 9070
rect 75337 8984 75423 9070
rect 75169 8816 75255 8902
rect 75337 8816 75423 8902
rect 75169 8648 75255 8734
rect 75337 8648 75423 8734
rect 75169 8480 75255 8566
rect 75337 8480 75423 8566
rect 4409 8336 4495 8359
rect 4577 8336 4663 8359
rect 4409 8296 4434 8336
rect 4434 8296 4474 8336
rect 4474 8296 4495 8336
rect 4577 8296 4598 8336
rect 4598 8296 4638 8336
rect 4638 8296 4663 8336
rect 4409 8273 4495 8296
rect 4577 8273 4663 8296
rect 8409 8336 8495 8359
rect 8577 8336 8663 8359
rect 8409 8296 8434 8336
rect 8434 8296 8474 8336
rect 8474 8296 8495 8336
rect 8577 8296 8598 8336
rect 8598 8296 8638 8336
rect 8638 8296 8663 8336
rect 8409 8273 8495 8296
rect 8577 8273 8663 8296
rect 12409 8336 12495 8359
rect 12577 8336 12663 8359
rect 12409 8296 12434 8336
rect 12434 8296 12474 8336
rect 12474 8296 12495 8336
rect 12577 8296 12598 8336
rect 12598 8296 12638 8336
rect 12638 8296 12663 8336
rect 12409 8273 12495 8296
rect 12577 8273 12663 8296
rect 16409 8336 16495 8359
rect 16577 8336 16663 8359
rect 16409 8296 16434 8336
rect 16434 8296 16474 8336
rect 16474 8296 16495 8336
rect 16577 8296 16598 8336
rect 16598 8296 16638 8336
rect 16638 8296 16663 8336
rect 16409 8273 16495 8296
rect 16577 8273 16663 8296
rect 20409 8336 20495 8359
rect 20577 8336 20663 8359
rect 20409 8296 20434 8336
rect 20434 8296 20474 8336
rect 20474 8296 20495 8336
rect 20577 8296 20598 8336
rect 20598 8296 20638 8336
rect 20638 8296 20663 8336
rect 20409 8273 20495 8296
rect 20577 8273 20663 8296
rect 24409 8336 24495 8359
rect 24577 8336 24663 8359
rect 24409 8296 24434 8336
rect 24434 8296 24474 8336
rect 24474 8296 24495 8336
rect 24577 8296 24598 8336
rect 24598 8296 24638 8336
rect 24638 8296 24663 8336
rect 24409 8273 24495 8296
rect 24577 8273 24663 8296
rect 28409 8336 28495 8359
rect 28577 8336 28663 8359
rect 28409 8296 28434 8336
rect 28434 8296 28474 8336
rect 28474 8296 28495 8336
rect 28577 8296 28598 8336
rect 28598 8296 28638 8336
rect 28638 8296 28663 8336
rect 28409 8273 28495 8296
rect 28577 8273 28663 8296
rect 32409 8336 32495 8359
rect 32577 8336 32663 8359
rect 32409 8296 32434 8336
rect 32434 8296 32474 8336
rect 32474 8296 32495 8336
rect 32577 8296 32598 8336
rect 32598 8296 32638 8336
rect 32638 8296 32663 8336
rect 32409 8273 32495 8296
rect 32577 8273 32663 8296
rect 36409 8336 36495 8359
rect 36577 8336 36663 8359
rect 36409 8296 36434 8336
rect 36434 8296 36474 8336
rect 36474 8296 36495 8336
rect 36577 8296 36598 8336
rect 36598 8296 36638 8336
rect 36638 8296 36663 8336
rect 36409 8273 36495 8296
rect 36577 8273 36663 8296
rect 40409 8336 40495 8359
rect 40577 8336 40663 8359
rect 40409 8296 40434 8336
rect 40434 8296 40474 8336
rect 40474 8296 40495 8336
rect 40577 8296 40598 8336
rect 40598 8296 40638 8336
rect 40638 8296 40663 8336
rect 40409 8273 40495 8296
rect 40577 8273 40663 8296
rect 44409 8336 44495 8359
rect 44577 8336 44663 8359
rect 44409 8296 44434 8336
rect 44434 8296 44474 8336
rect 44474 8296 44495 8336
rect 44577 8296 44598 8336
rect 44598 8296 44638 8336
rect 44638 8296 44663 8336
rect 44409 8273 44495 8296
rect 44577 8273 44663 8296
rect 48409 8336 48495 8359
rect 48577 8336 48663 8359
rect 48409 8296 48434 8336
rect 48434 8296 48474 8336
rect 48474 8296 48495 8336
rect 48577 8296 48598 8336
rect 48598 8296 48638 8336
rect 48638 8296 48663 8336
rect 48409 8273 48495 8296
rect 48577 8273 48663 8296
rect 52409 8336 52495 8359
rect 52577 8336 52663 8359
rect 52409 8296 52434 8336
rect 52434 8296 52474 8336
rect 52474 8296 52495 8336
rect 52577 8296 52598 8336
rect 52598 8296 52638 8336
rect 52638 8296 52663 8336
rect 52409 8273 52495 8296
rect 52577 8273 52663 8296
rect 56409 8336 56495 8359
rect 56577 8336 56663 8359
rect 56409 8296 56434 8336
rect 56434 8296 56474 8336
rect 56474 8296 56495 8336
rect 56577 8296 56598 8336
rect 56598 8296 56638 8336
rect 56638 8296 56663 8336
rect 56409 8273 56495 8296
rect 56577 8273 56663 8296
rect 60409 8336 60495 8359
rect 60577 8336 60663 8359
rect 60409 8296 60434 8336
rect 60434 8296 60474 8336
rect 60474 8296 60495 8336
rect 60577 8296 60598 8336
rect 60598 8296 60638 8336
rect 60638 8296 60663 8336
rect 60409 8273 60495 8296
rect 60577 8273 60663 8296
rect 64409 8336 64495 8359
rect 64577 8336 64663 8359
rect 64409 8296 64434 8336
rect 64434 8296 64474 8336
rect 64474 8296 64495 8336
rect 64577 8296 64598 8336
rect 64598 8296 64638 8336
rect 64638 8296 64663 8336
rect 64409 8273 64495 8296
rect 64577 8273 64663 8296
rect 68409 8336 68495 8359
rect 68577 8336 68663 8359
rect 68409 8296 68434 8336
rect 68434 8296 68474 8336
rect 68474 8296 68495 8336
rect 68577 8296 68598 8336
rect 68598 8296 68638 8336
rect 68638 8296 68663 8336
rect 68409 8273 68495 8296
rect 68577 8273 68663 8296
rect 75169 8312 75255 8398
rect 75337 8312 75423 8398
rect 75169 8144 75255 8230
rect 75337 8144 75423 8230
rect 79169 10160 79255 10246
rect 79337 10160 79423 10246
rect 79169 9992 79255 10078
rect 79337 9992 79423 10078
rect 79169 9824 79255 9910
rect 79337 9824 79423 9910
rect 79169 9656 79255 9742
rect 79337 9656 79423 9742
rect 79169 9488 79255 9574
rect 79337 9488 79423 9574
rect 79169 9320 79255 9406
rect 79337 9320 79423 9406
rect 79169 9152 79255 9238
rect 79337 9152 79423 9238
rect 79169 8984 79255 9070
rect 79337 8984 79423 9070
rect 79169 8816 79255 8902
rect 79337 8816 79423 8902
rect 79169 8648 79255 8734
rect 79337 8648 79423 8734
rect 79169 8480 79255 8566
rect 79337 8480 79423 8566
rect 79169 8312 79255 8398
rect 79337 8312 79423 8398
rect 79169 8144 79255 8230
rect 79337 8144 79423 8230
rect 83169 10160 83255 10246
rect 83337 10160 83423 10246
rect 83169 9992 83255 10078
rect 83337 9992 83423 10078
rect 83169 9824 83255 9910
rect 83337 9824 83423 9910
rect 83169 9656 83255 9742
rect 83337 9656 83423 9742
rect 83169 9488 83255 9574
rect 83337 9488 83423 9574
rect 83169 9320 83255 9406
rect 83337 9320 83423 9406
rect 83169 9152 83255 9238
rect 83337 9152 83423 9238
rect 83169 8984 83255 9070
rect 83337 8984 83423 9070
rect 83169 8816 83255 8902
rect 83337 8816 83423 8902
rect 83169 8648 83255 8734
rect 83337 8648 83423 8734
rect 83169 8480 83255 8566
rect 83337 8480 83423 8566
rect 83169 8312 83255 8398
rect 83337 8312 83423 8398
rect 83169 8144 83255 8230
rect 83337 8144 83423 8230
rect 87169 10160 87255 10246
rect 87337 10160 87423 10246
rect 87169 9992 87255 10078
rect 87337 9992 87423 10078
rect 87169 9824 87255 9910
rect 87337 9824 87423 9910
rect 87169 9656 87255 9742
rect 87337 9656 87423 9742
rect 87169 9488 87255 9574
rect 87337 9488 87423 9574
rect 87169 9320 87255 9406
rect 87337 9320 87423 9406
rect 87169 9152 87255 9238
rect 87337 9152 87423 9238
rect 87169 8984 87255 9070
rect 87337 8984 87423 9070
rect 87169 8816 87255 8902
rect 87337 8816 87423 8902
rect 87169 8648 87255 8734
rect 87337 8648 87423 8734
rect 87169 8480 87255 8566
rect 87337 8480 87423 8566
rect 87169 8312 87255 8398
rect 87337 8312 87423 8398
rect 87169 8144 87255 8230
rect 87337 8144 87423 8230
rect 91169 10160 91255 10246
rect 91337 10160 91423 10246
rect 91169 9992 91255 10078
rect 91337 9992 91423 10078
rect 91169 9824 91255 9910
rect 91337 9824 91423 9910
rect 91169 9656 91255 9742
rect 91337 9656 91423 9742
rect 91169 9488 91255 9574
rect 91337 9488 91423 9574
rect 91169 9320 91255 9406
rect 91337 9320 91423 9406
rect 91169 9152 91255 9238
rect 91337 9152 91423 9238
rect 91169 8984 91255 9070
rect 91337 8984 91423 9070
rect 91169 8816 91255 8902
rect 91337 8816 91423 8902
rect 91169 8648 91255 8734
rect 91337 8648 91423 8734
rect 91169 8480 91255 8566
rect 91337 8480 91423 8566
rect 91169 8312 91255 8398
rect 91337 8312 91423 8398
rect 91169 8144 91255 8230
rect 91337 8144 91423 8230
rect 95169 10160 95255 10246
rect 95337 10160 95423 10246
rect 95169 9992 95255 10078
rect 95337 9992 95423 10078
rect 95169 9824 95255 9910
rect 95337 9824 95423 9910
rect 95169 9656 95255 9742
rect 95337 9656 95423 9742
rect 95169 9488 95255 9574
rect 95337 9488 95423 9574
rect 95169 9320 95255 9406
rect 95337 9320 95423 9406
rect 95169 9152 95255 9238
rect 95337 9152 95423 9238
rect 95169 8984 95255 9070
rect 95337 8984 95423 9070
rect 95169 8816 95255 8902
rect 95337 8816 95423 8902
rect 95169 8648 95255 8734
rect 95337 8648 95423 8734
rect 95169 8480 95255 8566
rect 95337 8480 95423 8566
rect 95169 8312 95255 8398
rect 95337 8312 95423 8398
rect 95169 8144 95255 8230
rect 95337 8144 95423 8230
rect 3169 7580 3255 7603
rect 3337 7580 3423 7603
rect 3169 7540 3194 7580
rect 3194 7540 3234 7580
rect 3234 7540 3255 7580
rect 3337 7540 3358 7580
rect 3358 7540 3398 7580
rect 3398 7540 3423 7580
rect 3169 7517 3255 7540
rect 3337 7517 3423 7540
rect 7169 7580 7255 7603
rect 7337 7580 7423 7603
rect 7169 7540 7194 7580
rect 7194 7540 7234 7580
rect 7234 7540 7255 7580
rect 7337 7540 7358 7580
rect 7358 7540 7398 7580
rect 7398 7540 7423 7580
rect 7169 7517 7255 7540
rect 7337 7517 7423 7540
rect 11169 7580 11255 7603
rect 11337 7580 11423 7603
rect 11169 7540 11194 7580
rect 11194 7540 11234 7580
rect 11234 7540 11255 7580
rect 11337 7540 11358 7580
rect 11358 7540 11398 7580
rect 11398 7540 11423 7580
rect 11169 7517 11255 7540
rect 11337 7517 11423 7540
rect 15169 7580 15255 7603
rect 15337 7580 15423 7603
rect 15169 7540 15194 7580
rect 15194 7540 15234 7580
rect 15234 7540 15255 7580
rect 15337 7540 15358 7580
rect 15358 7540 15398 7580
rect 15398 7540 15423 7580
rect 15169 7517 15255 7540
rect 15337 7517 15423 7540
rect 19169 7580 19255 7603
rect 19337 7580 19423 7603
rect 19169 7540 19194 7580
rect 19194 7540 19234 7580
rect 19234 7540 19255 7580
rect 19337 7540 19358 7580
rect 19358 7540 19398 7580
rect 19398 7540 19423 7580
rect 19169 7517 19255 7540
rect 19337 7517 19423 7540
rect 23169 7580 23255 7603
rect 23337 7580 23423 7603
rect 23169 7540 23194 7580
rect 23194 7540 23234 7580
rect 23234 7540 23255 7580
rect 23337 7540 23358 7580
rect 23358 7540 23398 7580
rect 23398 7540 23423 7580
rect 23169 7517 23255 7540
rect 23337 7517 23423 7540
rect 27169 7580 27255 7603
rect 27337 7580 27423 7603
rect 27169 7540 27194 7580
rect 27194 7540 27234 7580
rect 27234 7540 27255 7580
rect 27337 7540 27358 7580
rect 27358 7540 27398 7580
rect 27398 7540 27423 7580
rect 27169 7517 27255 7540
rect 27337 7517 27423 7540
rect 31169 7580 31255 7603
rect 31337 7580 31423 7603
rect 31169 7540 31194 7580
rect 31194 7540 31234 7580
rect 31234 7540 31255 7580
rect 31337 7540 31358 7580
rect 31358 7540 31398 7580
rect 31398 7540 31423 7580
rect 31169 7517 31255 7540
rect 31337 7517 31423 7540
rect 35169 7580 35255 7603
rect 35337 7580 35423 7603
rect 35169 7540 35194 7580
rect 35194 7540 35234 7580
rect 35234 7540 35255 7580
rect 35337 7540 35358 7580
rect 35358 7540 35398 7580
rect 35398 7540 35423 7580
rect 35169 7517 35255 7540
rect 35337 7517 35423 7540
rect 39169 7580 39255 7603
rect 39337 7580 39423 7603
rect 39169 7540 39194 7580
rect 39194 7540 39234 7580
rect 39234 7540 39255 7580
rect 39337 7540 39358 7580
rect 39358 7540 39398 7580
rect 39398 7540 39423 7580
rect 39169 7517 39255 7540
rect 39337 7517 39423 7540
rect 43169 7580 43255 7603
rect 43337 7580 43423 7603
rect 43169 7540 43194 7580
rect 43194 7540 43234 7580
rect 43234 7540 43255 7580
rect 43337 7540 43358 7580
rect 43358 7540 43398 7580
rect 43398 7540 43423 7580
rect 43169 7517 43255 7540
rect 43337 7517 43423 7540
rect 47169 7580 47255 7603
rect 47337 7580 47423 7603
rect 47169 7540 47194 7580
rect 47194 7540 47234 7580
rect 47234 7540 47255 7580
rect 47337 7540 47358 7580
rect 47358 7540 47398 7580
rect 47398 7540 47423 7580
rect 47169 7517 47255 7540
rect 47337 7517 47423 7540
rect 51169 7580 51255 7603
rect 51337 7580 51423 7603
rect 51169 7540 51194 7580
rect 51194 7540 51234 7580
rect 51234 7540 51255 7580
rect 51337 7540 51358 7580
rect 51358 7540 51398 7580
rect 51398 7540 51423 7580
rect 51169 7517 51255 7540
rect 51337 7517 51423 7540
rect 55169 7580 55255 7603
rect 55337 7580 55423 7603
rect 55169 7540 55194 7580
rect 55194 7540 55234 7580
rect 55234 7540 55255 7580
rect 55337 7540 55358 7580
rect 55358 7540 55398 7580
rect 55398 7540 55423 7580
rect 55169 7517 55255 7540
rect 55337 7517 55423 7540
rect 59169 7580 59255 7603
rect 59337 7580 59423 7603
rect 59169 7540 59194 7580
rect 59194 7540 59234 7580
rect 59234 7540 59255 7580
rect 59337 7540 59358 7580
rect 59358 7540 59398 7580
rect 59398 7540 59423 7580
rect 59169 7517 59255 7540
rect 59337 7517 59423 7540
rect 63169 7580 63255 7603
rect 63337 7580 63423 7603
rect 63169 7540 63194 7580
rect 63194 7540 63234 7580
rect 63234 7540 63255 7580
rect 63337 7540 63358 7580
rect 63358 7540 63398 7580
rect 63398 7540 63423 7580
rect 63169 7517 63255 7540
rect 63337 7517 63423 7540
rect 67169 7580 67255 7603
rect 67337 7580 67423 7603
rect 67169 7540 67194 7580
rect 67194 7540 67234 7580
rect 67234 7540 67255 7580
rect 67337 7540 67358 7580
rect 67358 7540 67398 7580
rect 67398 7540 67423 7580
rect 67169 7517 67255 7540
rect 67337 7517 67423 7540
rect 86469 7433 86555 7519
rect 4409 6824 4495 6847
rect 4577 6824 4663 6847
rect 4409 6784 4434 6824
rect 4434 6784 4474 6824
rect 4474 6784 4495 6824
rect 4577 6784 4598 6824
rect 4598 6784 4638 6824
rect 4638 6784 4663 6824
rect 4409 6761 4495 6784
rect 4577 6761 4663 6784
rect 8409 6824 8495 6847
rect 8577 6824 8663 6847
rect 8409 6784 8434 6824
rect 8434 6784 8474 6824
rect 8474 6784 8495 6824
rect 8577 6784 8598 6824
rect 8598 6784 8638 6824
rect 8638 6784 8663 6824
rect 8409 6761 8495 6784
rect 8577 6761 8663 6784
rect 12409 6824 12495 6847
rect 12577 6824 12663 6847
rect 12409 6784 12434 6824
rect 12434 6784 12474 6824
rect 12474 6784 12495 6824
rect 12577 6784 12598 6824
rect 12598 6784 12638 6824
rect 12638 6784 12663 6824
rect 12409 6761 12495 6784
rect 12577 6761 12663 6784
rect 16409 6824 16495 6847
rect 16577 6824 16663 6847
rect 16409 6784 16434 6824
rect 16434 6784 16474 6824
rect 16474 6784 16495 6824
rect 16577 6784 16598 6824
rect 16598 6784 16638 6824
rect 16638 6784 16663 6824
rect 16409 6761 16495 6784
rect 16577 6761 16663 6784
rect 20409 6824 20495 6847
rect 20577 6824 20663 6847
rect 20409 6784 20434 6824
rect 20434 6784 20474 6824
rect 20474 6784 20495 6824
rect 20577 6784 20598 6824
rect 20598 6784 20638 6824
rect 20638 6784 20663 6824
rect 20409 6761 20495 6784
rect 20577 6761 20663 6784
rect 24409 6824 24495 6847
rect 24577 6824 24663 6847
rect 24409 6784 24434 6824
rect 24434 6784 24474 6824
rect 24474 6784 24495 6824
rect 24577 6784 24598 6824
rect 24598 6784 24638 6824
rect 24638 6784 24663 6824
rect 24409 6761 24495 6784
rect 24577 6761 24663 6784
rect 28409 6824 28495 6847
rect 28577 6824 28663 6847
rect 28409 6784 28434 6824
rect 28434 6784 28474 6824
rect 28474 6784 28495 6824
rect 28577 6784 28598 6824
rect 28598 6784 28638 6824
rect 28638 6784 28663 6824
rect 28409 6761 28495 6784
rect 28577 6761 28663 6784
rect 32409 6824 32495 6847
rect 32577 6824 32663 6847
rect 32409 6784 32434 6824
rect 32434 6784 32474 6824
rect 32474 6784 32495 6824
rect 32577 6784 32598 6824
rect 32598 6784 32638 6824
rect 32638 6784 32663 6824
rect 32409 6761 32495 6784
rect 32577 6761 32663 6784
rect 36409 6824 36495 6847
rect 36577 6824 36663 6847
rect 36409 6784 36434 6824
rect 36434 6784 36474 6824
rect 36474 6784 36495 6824
rect 36577 6784 36598 6824
rect 36598 6784 36638 6824
rect 36638 6784 36663 6824
rect 36409 6761 36495 6784
rect 36577 6761 36663 6784
rect 40409 6824 40495 6847
rect 40577 6824 40663 6847
rect 40409 6784 40434 6824
rect 40434 6784 40474 6824
rect 40474 6784 40495 6824
rect 40577 6784 40598 6824
rect 40598 6784 40638 6824
rect 40638 6784 40663 6824
rect 40409 6761 40495 6784
rect 40577 6761 40663 6784
rect 44409 6824 44495 6847
rect 44577 6824 44663 6847
rect 44409 6784 44434 6824
rect 44434 6784 44474 6824
rect 44474 6784 44495 6824
rect 44577 6784 44598 6824
rect 44598 6784 44638 6824
rect 44638 6784 44663 6824
rect 44409 6761 44495 6784
rect 44577 6761 44663 6784
rect 48409 6824 48495 6847
rect 48577 6824 48663 6847
rect 48409 6784 48434 6824
rect 48434 6784 48474 6824
rect 48474 6784 48495 6824
rect 48577 6784 48598 6824
rect 48598 6784 48638 6824
rect 48638 6784 48663 6824
rect 48409 6761 48495 6784
rect 48577 6761 48663 6784
rect 52409 6824 52495 6847
rect 52577 6824 52663 6847
rect 52409 6784 52434 6824
rect 52434 6784 52474 6824
rect 52474 6784 52495 6824
rect 52577 6784 52598 6824
rect 52598 6784 52638 6824
rect 52638 6784 52663 6824
rect 52409 6761 52495 6784
rect 52577 6761 52663 6784
rect 56409 6824 56495 6847
rect 56577 6824 56663 6847
rect 56409 6784 56434 6824
rect 56434 6784 56474 6824
rect 56474 6784 56495 6824
rect 56577 6784 56598 6824
rect 56598 6784 56638 6824
rect 56638 6784 56663 6824
rect 56409 6761 56495 6784
rect 56577 6761 56663 6784
rect 60409 6824 60495 6847
rect 60577 6824 60663 6847
rect 60409 6784 60434 6824
rect 60434 6784 60474 6824
rect 60474 6784 60495 6824
rect 60577 6784 60598 6824
rect 60598 6784 60638 6824
rect 60638 6784 60663 6824
rect 60409 6761 60495 6784
rect 60577 6761 60663 6784
rect 64409 6824 64495 6847
rect 64577 6824 64663 6847
rect 64409 6784 64434 6824
rect 64434 6784 64474 6824
rect 64474 6784 64495 6824
rect 64577 6784 64598 6824
rect 64598 6784 64638 6824
rect 64638 6784 64663 6824
rect 64409 6761 64495 6784
rect 64577 6761 64663 6784
rect 68409 6824 68495 6847
rect 68577 6824 68663 6847
rect 68409 6784 68434 6824
rect 68434 6784 68474 6824
rect 68474 6784 68495 6824
rect 68577 6784 68598 6824
rect 68598 6784 68638 6824
rect 68638 6784 68663 6824
rect 68409 6761 68495 6784
rect 68577 6761 68663 6784
rect 3169 6068 3255 6091
rect 3337 6068 3423 6091
rect 3169 6028 3194 6068
rect 3194 6028 3234 6068
rect 3234 6028 3255 6068
rect 3337 6028 3358 6068
rect 3358 6028 3398 6068
rect 3398 6028 3423 6068
rect 3169 6005 3255 6028
rect 3337 6005 3423 6028
rect 7169 6068 7255 6091
rect 7337 6068 7423 6091
rect 7169 6028 7194 6068
rect 7194 6028 7234 6068
rect 7234 6028 7255 6068
rect 7337 6028 7358 6068
rect 7358 6028 7398 6068
rect 7398 6028 7423 6068
rect 7169 6005 7255 6028
rect 7337 6005 7423 6028
rect 11169 6068 11255 6091
rect 11337 6068 11423 6091
rect 11169 6028 11194 6068
rect 11194 6028 11234 6068
rect 11234 6028 11255 6068
rect 11337 6028 11358 6068
rect 11358 6028 11398 6068
rect 11398 6028 11423 6068
rect 11169 6005 11255 6028
rect 11337 6005 11423 6028
rect 15169 6068 15255 6091
rect 15337 6068 15423 6091
rect 15169 6028 15194 6068
rect 15194 6028 15234 6068
rect 15234 6028 15255 6068
rect 15337 6028 15358 6068
rect 15358 6028 15398 6068
rect 15398 6028 15423 6068
rect 15169 6005 15255 6028
rect 15337 6005 15423 6028
rect 19169 6068 19255 6091
rect 19337 6068 19423 6091
rect 19169 6028 19194 6068
rect 19194 6028 19234 6068
rect 19234 6028 19255 6068
rect 19337 6028 19358 6068
rect 19358 6028 19398 6068
rect 19398 6028 19423 6068
rect 19169 6005 19255 6028
rect 19337 6005 19423 6028
rect 23169 6068 23255 6091
rect 23337 6068 23423 6091
rect 23169 6028 23194 6068
rect 23194 6028 23234 6068
rect 23234 6028 23255 6068
rect 23337 6028 23358 6068
rect 23358 6028 23398 6068
rect 23398 6028 23423 6068
rect 23169 6005 23255 6028
rect 23337 6005 23423 6028
rect 27169 6068 27255 6091
rect 27337 6068 27423 6091
rect 27169 6028 27194 6068
rect 27194 6028 27234 6068
rect 27234 6028 27255 6068
rect 27337 6028 27358 6068
rect 27358 6028 27398 6068
rect 27398 6028 27423 6068
rect 27169 6005 27255 6028
rect 27337 6005 27423 6028
rect 31169 6068 31255 6091
rect 31337 6068 31423 6091
rect 31169 6028 31194 6068
rect 31194 6028 31234 6068
rect 31234 6028 31255 6068
rect 31337 6028 31358 6068
rect 31358 6028 31398 6068
rect 31398 6028 31423 6068
rect 31169 6005 31255 6028
rect 31337 6005 31423 6028
rect 35169 6068 35255 6091
rect 35337 6068 35423 6091
rect 35169 6028 35194 6068
rect 35194 6028 35234 6068
rect 35234 6028 35255 6068
rect 35337 6028 35358 6068
rect 35358 6028 35398 6068
rect 35398 6028 35423 6068
rect 35169 6005 35255 6028
rect 35337 6005 35423 6028
rect 39169 6068 39255 6091
rect 39337 6068 39423 6091
rect 39169 6028 39194 6068
rect 39194 6028 39234 6068
rect 39234 6028 39255 6068
rect 39337 6028 39358 6068
rect 39358 6028 39398 6068
rect 39398 6028 39423 6068
rect 39169 6005 39255 6028
rect 39337 6005 39423 6028
rect 43169 6068 43255 6091
rect 43337 6068 43423 6091
rect 43169 6028 43194 6068
rect 43194 6028 43234 6068
rect 43234 6028 43255 6068
rect 43337 6028 43358 6068
rect 43358 6028 43398 6068
rect 43398 6028 43423 6068
rect 43169 6005 43255 6028
rect 43337 6005 43423 6028
rect 47169 6068 47255 6091
rect 47337 6068 47423 6091
rect 47169 6028 47194 6068
rect 47194 6028 47234 6068
rect 47234 6028 47255 6068
rect 47337 6028 47358 6068
rect 47358 6028 47398 6068
rect 47398 6028 47423 6068
rect 47169 6005 47255 6028
rect 47337 6005 47423 6028
rect 51169 6068 51255 6091
rect 51337 6068 51423 6091
rect 51169 6028 51194 6068
rect 51194 6028 51234 6068
rect 51234 6028 51255 6068
rect 51337 6028 51358 6068
rect 51358 6028 51398 6068
rect 51398 6028 51423 6068
rect 51169 6005 51255 6028
rect 51337 6005 51423 6028
rect 55169 6068 55255 6091
rect 55337 6068 55423 6091
rect 55169 6028 55194 6068
rect 55194 6028 55234 6068
rect 55234 6028 55255 6068
rect 55337 6028 55358 6068
rect 55358 6028 55398 6068
rect 55398 6028 55423 6068
rect 55169 6005 55255 6028
rect 55337 6005 55423 6028
rect 59169 6068 59255 6091
rect 59337 6068 59423 6091
rect 59169 6028 59194 6068
rect 59194 6028 59234 6068
rect 59234 6028 59255 6068
rect 59337 6028 59358 6068
rect 59358 6028 59398 6068
rect 59398 6028 59423 6068
rect 59169 6005 59255 6028
rect 59337 6005 59423 6028
rect 63169 6068 63255 6091
rect 63337 6068 63423 6091
rect 63169 6028 63194 6068
rect 63194 6028 63234 6068
rect 63234 6028 63255 6068
rect 63337 6028 63358 6068
rect 63358 6028 63398 6068
rect 63398 6028 63423 6068
rect 63169 6005 63255 6028
rect 63337 6005 63423 6028
rect 67169 6068 67255 6091
rect 67337 6068 67423 6091
rect 67169 6028 67194 6068
rect 67194 6028 67234 6068
rect 67234 6028 67255 6068
rect 67337 6028 67358 6068
rect 67358 6028 67398 6068
rect 67398 6028 67423 6068
rect 67169 6005 67255 6028
rect 67337 6005 67423 6028
rect 4409 5312 4495 5335
rect 4577 5312 4663 5335
rect 4409 5272 4434 5312
rect 4434 5272 4474 5312
rect 4474 5272 4495 5312
rect 4577 5272 4598 5312
rect 4598 5272 4638 5312
rect 4638 5272 4663 5312
rect 4409 5249 4495 5272
rect 4577 5249 4663 5272
rect 8409 5312 8495 5335
rect 8577 5312 8663 5335
rect 8409 5272 8434 5312
rect 8434 5272 8474 5312
rect 8474 5272 8495 5312
rect 8577 5272 8598 5312
rect 8598 5272 8638 5312
rect 8638 5272 8663 5312
rect 8409 5249 8495 5272
rect 8577 5249 8663 5272
rect 12409 5312 12495 5335
rect 12577 5312 12663 5335
rect 12409 5272 12434 5312
rect 12434 5272 12474 5312
rect 12474 5272 12495 5312
rect 12577 5272 12598 5312
rect 12598 5272 12638 5312
rect 12638 5272 12663 5312
rect 12409 5249 12495 5272
rect 12577 5249 12663 5272
rect 16409 5312 16495 5335
rect 16577 5312 16663 5335
rect 16409 5272 16434 5312
rect 16434 5272 16474 5312
rect 16474 5272 16495 5312
rect 16577 5272 16598 5312
rect 16598 5272 16638 5312
rect 16638 5272 16663 5312
rect 16409 5249 16495 5272
rect 16577 5249 16663 5272
rect 20409 5312 20495 5335
rect 20577 5312 20663 5335
rect 20409 5272 20434 5312
rect 20434 5272 20474 5312
rect 20474 5272 20495 5312
rect 20577 5272 20598 5312
rect 20598 5272 20638 5312
rect 20638 5272 20663 5312
rect 20409 5249 20495 5272
rect 20577 5249 20663 5272
rect 24409 5312 24495 5335
rect 24577 5312 24663 5335
rect 24409 5272 24434 5312
rect 24434 5272 24474 5312
rect 24474 5272 24495 5312
rect 24577 5272 24598 5312
rect 24598 5272 24638 5312
rect 24638 5272 24663 5312
rect 24409 5249 24495 5272
rect 24577 5249 24663 5272
rect 28409 5312 28495 5335
rect 28577 5312 28663 5335
rect 28409 5272 28434 5312
rect 28434 5272 28474 5312
rect 28474 5272 28495 5312
rect 28577 5272 28598 5312
rect 28598 5272 28638 5312
rect 28638 5272 28663 5312
rect 28409 5249 28495 5272
rect 28577 5249 28663 5272
rect 32409 5312 32495 5335
rect 32577 5312 32663 5335
rect 32409 5272 32434 5312
rect 32434 5272 32474 5312
rect 32474 5272 32495 5312
rect 32577 5272 32598 5312
rect 32598 5272 32638 5312
rect 32638 5272 32663 5312
rect 32409 5249 32495 5272
rect 32577 5249 32663 5272
rect 36409 5312 36495 5335
rect 36577 5312 36663 5335
rect 36409 5272 36434 5312
rect 36434 5272 36474 5312
rect 36474 5272 36495 5312
rect 36577 5272 36598 5312
rect 36598 5272 36638 5312
rect 36638 5272 36663 5312
rect 36409 5249 36495 5272
rect 36577 5249 36663 5272
rect 40409 5312 40495 5335
rect 40577 5312 40663 5335
rect 40409 5272 40434 5312
rect 40434 5272 40474 5312
rect 40474 5272 40495 5312
rect 40577 5272 40598 5312
rect 40598 5272 40638 5312
rect 40638 5272 40663 5312
rect 40409 5249 40495 5272
rect 40577 5249 40663 5272
rect 44409 5312 44495 5335
rect 44577 5312 44663 5335
rect 44409 5272 44434 5312
rect 44434 5272 44474 5312
rect 44474 5272 44495 5312
rect 44577 5272 44598 5312
rect 44598 5272 44638 5312
rect 44638 5272 44663 5312
rect 44409 5249 44495 5272
rect 44577 5249 44663 5272
rect 48409 5312 48495 5335
rect 48577 5312 48663 5335
rect 48409 5272 48434 5312
rect 48434 5272 48474 5312
rect 48474 5272 48495 5312
rect 48577 5272 48598 5312
rect 48598 5272 48638 5312
rect 48638 5272 48663 5312
rect 48409 5249 48495 5272
rect 48577 5249 48663 5272
rect 52409 5312 52495 5335
rect 52577 5312 52663 5335
rect 52409 5272 52434 5312
rect 52434 5272 52474 5312
rect 52474 5272 52495 5312
rect 52577 5272 52598 5312
rect 52598 5272 52638 5312
rect 52638 5272 52663 5312
rect 52409 5249 52495 5272
rect 52577 5249 52663 5272
rect 56409 5312 56495 5335
rect 56577 5312 56663 5335
rect 56409 5272 56434 5312
rect 56434 5272 56474 5312
rect 56474 5272 56495 5312
rect 56577 5272 56598 5312
rect 56598 5272 56638 5312
rect 56638 5272 56663 5312
rect 56409 5249 56495 5272
rect 56577 5249 56663 5272
rect 60409 5312 60495 5335
rect 60577 5312 60663 5335
rect 60409 5272 60434 5312
rect 60434 5272 60474 5312
rect 60474 5272 60495 5312
rect 60577 5272 60598 5312
rect 60598 5272 60638 5312
rect 60638 5272 60663 5312
rect 60409 5249 60495 5272
rect 60577 5249 60663 5272
rect 64409 5312 64495 5335
rect 64577 5312 64663 5335
rect 64409 5272 64434 5312
rect 64434 5272 64474 5312
rect 64474 5272 64495 5312
rect 64577 5272 64598 5312
rect 64598 5272 64638 5312
rect 64638 5272 64663 5312
rect 64409 5249 64495 5272
rect 64577 5249 64663 5272
rect 68409 5312 68495 5335
rect 68577 5312 68663 5335
rect 68409 5272 68434 5312
rect 68434 5272 68474 5312
rect 68474 5272 68495 5312
rect 68577 5272 68598 5312
rect 68598 5272 68638 5312
rect 68638 5272 68663 5312
rect 68409 5249 68495 5272
rect 68577 5249 68663 5272
rect 72409 5312 72495 5335
rect 72577 5312 72663 5335
rect 72409 5272 72434 5312
rect 72434 5272 72474 5312
rect 72474 5272 72495 5312
rect 72577 5272 72598 5312
rect 72598 5272 72638 5312
rect 72638 5272 72663 5312
rect 72409 5249 72495 5272
rect 72577 5249 72663 5272
rect 76409 5312 76495 5335
rect 76577 5312 76663 5335
rect 76409 5272 76434 5312
rect 76434 5272 76474 5312
rect 76474 5272 76495 5312
rect 76577 5272 76598 5312
rect 76598 5272 76638 5312
rect 76638 5272 76663 5312
rect 76409 5249 76495 5272
rect 76577 5249 76663 5272
rect 80409 5312 80495 5335
rect 80577 5312 80663 5335
rect 80409 5272 80434 5312
rect 80434 5272 80474 5312
rect 80474 5272 80495 5312
rect 80577 5272 80598 5312
rect 80598 5272 80638 5312
rect 80638 5272 80663 5312
rect 80409 5249 80495 5272
rect 80577 5249 80663 5272
rect 84409 5312 84495 5335
rect 84577 5312 84663 5335
rect 84409 5272 84434 5312
rect 84434 5272 84474 5312
rect 84474 5272 84495 5312
rect 84577 5272 84598 5312
rect 84598 5272 84638 5312
rect 84638 5272 84663 5312
rect 84409 5249 84495 5272
rect 84577 5249 84663 5272
rect 88409 5312 88495 5335
rect 88577 5312 88663 5335
rect 88409 5272 88434 5312
rect 88434 5272 88474 5312
rect 88474 5272 88495 5312
rect 88577 5272 88598 5312
rect 88598 5272 88638 5312
rect 88638 5272 88663 5312
rect 88409 5249 88495 5272
rect 88577 5249 88663 5272
rect 92409 5312 92495 5335
rect 92577 5312 92663 5335
rect 92409 5272 92434 5312
rect 92434 5272 92474 5312
rect 92474 5272 92495 5312
rect 92577 5272 92598 5312
rect 92598 5272 92638 5312
rect 92638 5272 92663 5312
rect 92409 5249 92495 5272
rect 92577 5249 92663 5272
rect 96409 5312 96495 5335
rect 96577 5312 96663 5335
rect 96409 5272 96434 5312
rect 96434 5272 96474 5312
rect 96474 5272 96495 5312
rect 96577 5272 96598 5312
rect 96598 5272 96638 5312
rect 96638 5272 96663 5312
rect 96409 5249 96495 5272
rect 96577 5249 96663 5272
rect 3169 4556 3255 4579
rect 3337 4556 3423 4579
rect 3169 4516 3194 4556
rect 3194 4516 3234 4556
rect 3234 4516 3255 4556
rect 3337 4516 3358 4556
rect 3358 4516 3398 4556
rect 3398 4516 3423 4556
rect 3169 4493 3255 4516
rect 3337 4493 3423 4516
rect 7169 4556 7255 4579
rect 7337 4556 7423 4579
rect 7169 4516 7194 4556
rect 7194 4516 7234 4556
rect 7234 4516 7255 4556
rect 7337 4516 7358 4556
rect 7358 4516 7398 4556
rect 7398 4516 7423 4556
rect 7169 4493 7255 4516
rect 7337 4493 7423 4516
rect 11169 4556 11255 4579
rect 11337 4556 11423 4579
rect 11169 4516 11194 4556
rect 11194 4516 11234 4556
rect 11234 4516 11255 4556
rect 11337 4516 11358 4556
rect 11358 4516 11398 4556
rect 11398 4516 11423 4556
rect 11169 4493 11255 4516
rect 11337 4493 11423 4516
rect 15169 4556 15255 4579
rect 15337 4556 15423 4579
rect 15169 4516 15194 4556
rect 15194 4516 15234 4556
rect 15234 4516 15255 4556
rect 15337 4516 15358 4556
rect 15358 4516 15398 4556
rect 15398 4516 15423 4556
rect 15169 4493 15255 4516
rect 15337 4493 15423 4516
rect 19169 4556 19255 4579
rect 19337 4556 19423 4579
rect 19169 4516 19194 4556
rect 19194 4516 19234 4556
rect 19234 4516 19255 4556
rect 19337 4516 19358 4556
rect 19358 4516 19398 4556
rect 19398 4516 19423 4556
rect 19169 4493 19255 4516
rect 19337 4493 19423 4516
rect 23169 4556 23255 4579
rect 23337 4556 23423 4579
rect 23169 4516 23194 4556
rect 23194 4516 23234 4556
rect 23234 4516 23255 4556
rect 23337 4516 23358 4556
rect 23358 4516 23398 4556
rect 23398 4516 23423 4556
rect 23169 4493 23255 4516
rect 23337 4493 23423 4516
rect 27169 4556 27255 4579
rect 27337 4556 27423 4579
rect 27169 4516 27194 4556
rect 27194 4516 27234 4556
rect 27234 4516 27255 4556
rect 27337 4516 27358 4556
rect 27358 4516 27398 4556
rect 27398 4516 27423 4556
rect 27169 4493 27255 4516
rect 27337 4493 27423 4516
rect 31169 4556 31255 4579
rect 31337 4556 31423 4579
rect 31169 4516 31194 4556
rect 31194 4516 31234 4556
rect 31234 4516 31255 4556
rect 31337 4516 31358 4556
rect 31358 4516 31398 4556
rect 31398 4516 31423 4556
rect 31169 4493 31255 4516
rect 31337 4493 31423 4516
rect 35169 4556 35255 4579
rect 35337 4556 35423 4579
rect 35169 4516 35194 4556
rect 35194 4516 35234 4556
rect 35234 4516 35255 4556
rect 35337 4516 35358 4556
rect 35358 4516 35398 4556
rect 35398 4516 35423 4556
rect 35169 4493 35255 4516
rect 35337 4493 35423 4516
rect 39169 4556 39255 4579
rect 39337 4556 39423 4579
rect 39169 4516 39194 4556
rect 39194 4516 39234 4556
rect 39234 4516 39255 4556
rect 39337 4516 39358 4556
rect 39358 4516 39398 4556
rect 39398 4516 39423 4556
rect 39169 4493 39255 4516
rect 39337 4493 39423 4516
rect 43169 4556 43255 4579
rect 43337 4556 43423 4579
rect 43169 4516 43194 4556
rect 43194 4516 43234 4556
rect 43234 4516 43255 4556
rect 43337 4516 43358 4556
rect 43358 4516 43398 4556
rect 43398 4516 43423 4556
rect 43169 4493 43255 4516
rect 43337 4493 43423 4516
rect 47169 4556 47255 4579
rect 47337 4556 47423 4579
rect 47169 4516 47194 4556
rect 47194 4516 47234 4556
rect 47234 4516 47255 4556
rect 47337 4516 47358 4556
rect 47358 4516 47398 4556
rect 47398 4516 47423 4556
rect 47169 4493 47255 4516
rect 47337 4493 47423 4516
rect 51169 4556 51255 4579
rect 51337 4556 51423 4579
rect 51169 4516 51194 4556
rect 51194 4516 51234 4556
rect 51234 4516 51255 4556
rect 51337 4516 51358 4556
rect 51358 4516 51398 4556
rect 51398 4516 51423 4556
rect 51169 4493 51255 4516
rect 51337 4493 51423 4516
rect 55169 4556 55255 4579
rect 55337 4556 55423 4579
rect 55169 4516 55194 4556
rect 55194 4516 55234 4556
rect 55234 4516 55255 4556
rect 55337 4516 55358 4556
rect 55358 4516 55398 4556
rect 55398 4516 55423 4556
rect 55169 4493 55255 4516
rect 55337 4493 55423 4516
rect 59169 4556 59255 4579
rect 59337 4556 59423 4579
rect 59169 4516 59194 4556
rect 59194 4516 59234 4556
rect 59234 4516 59255 4556
rect 59337 4516 59358 4556
rect 59358 4516 59398 4556
rect 59398 4516 59423 4556
rect 59169 4493 59255 4516
rect 59337 4493 59423 4516
rect 63169 4556 63255 4579
rect 63337 4556 63423 4579
rect 63169 4516 63194 4556
rect 63194 4516 63234 4556
rect 63234 4516 63255 4556
rect 63337 4516 63358 4556
rect 63358 4516 63398 4556
rect 63398 4516 63423 4556
rect 63169 4493 63255 4516
rect 63337 4493 63423 4516
rect 67169 4556 67255 4579
rect 67337 4556 67423 4579
rect 67169 4516 67194 4556
rect 67194 4516 67234 4556
rect 67234 4516 67255 4556
rect 67337 4516 67358 4556
rect 67358 4516 67398 4556
rect 67398 4516 67423 4556
rect 67169 4493 67255 4516
rect 67337 4493 67423 4516
rect 71169 4556 71255 4579
rect 71337 4556 71423 4579
rect 71169 4516 71194 4556
rect 71194 4516 71234 4556
rect 71234 4516 71255 4556
rect 71337 4516 71358 4556
rect 71358 4516 71398 4556
rect 71398 4516 71423 4556
rect 71169 4493 71255 4516
rect 71337 4493 71423 4516
rect 75169 4556 75255 4579
rect 75337 4556 75423 4579
rect 75169 4516 75194 4556
rect 75194 4516 75234 4556
rect 75234 4516 75255 4556
rect 75337 4516 75358 4556
rect 75358 4516 75398 4556
rect 75398 4516 75423 4556
rect 75169 4493 75255 4516
rect 75337 4493 75423 4516
rect 79169 4556 79255 4579
rect 79337 4556 79423 4579
rect 79169 4516 79194 4556
rect 79194 4516 79234 4556
rect 79234 4516 79255 4556
rect 79337 4516 79358 4556
rect 79358 4516 79398 4556
rect 79398 4516 79423 4556
rect 79169 4493 79255 4516
rect 79337 4493 79423 4516
rect 83169 4556 83255 4579
rect 83337 4556 83423 4579
rect 83169 4516 83194 4556
rect 83194 4516 83234 4556
rect 83234 4516 83255 4556
rect 83337 4516 83358 4556
rect 83358 4516 83398 4556
rect 83398 4516 83423 4556
rect 83169 4493 83255 4516
rect 83337 4493 83423 4516
rect 87169 4556 87255 4579
rect 87337 4556 87423 4579
rect 87169 4516 87194 4556
rect 87194 4516 87234 4556
rect 87234 4516 87255 4556
rect 87337 4516 87358 4556
rect 87358 4516 87398 4556
rect 87398 4516 87423 4556
rect 87169 4493 87255 4516
rect 87337 4493 87423 4516
rect 91169 4556 91255 4579
rect 91337 4556 91423 4579
rect 91169 4516 91194 4556
rect 91194 4516 91234 4556
rect 91234 4516 91255 4556
rect 91337 4516 91358 4556
rect 91358 4516 91398 4556
rect 91398 4516 91423 4556
rect 91169 4493 91255 4516
rect 91337 4493 91423 4516
rect 95169 4556 95255 4579
rect 95337 4556 95423 4579
rect 95169 4516 95194 4556
rect 95194 4516 95234 4556
rect 95234 4516 95255 4556
rect 95337 4516 95358 4556
rect 95358 4516 95398 4556
rect 95398 4516 95423 4556
rect 95169 4493 95255 4516
rect 95337 4493 95423 4516
rect 99169 4556 99255 4579
rect 99337 4556 99423 4579
rect 99169 4516 99194 4556
rect 99194 4516 99234 4556
rect 99234 4516 99255 4556
rect 99337 4516 99358 4556
rect 99358 4516 99398 4556
rect 99398 4516 99423 4556
rect 99169 4493 99255 4516
rect 99337 4493 99423 4516
rect 4409 3800 4495 3823
rect 4577 3800 4663 3823
rect 4409 3760 4434 3800
rect 4434 3760 4474 3800
rect 4474 3760 4495 3800
rect 4577 3760 4598 3800
rect 4598 3760 4638 3800
rect 4638 3760 4663 3800
rect 4409 3737 4495 3760
rect 4577 3737 4663 3760
rect 8409 3800 8495 3823
rect 8577 3800 8663 3823
rect 8409 3760 8434 3800
rect 8434 3760 8474 3800
rect 8474 3760 8495 3800
rect 8577 3760 8598 3800
rect 8598 3760 8638 3800
rect 8638 3760 8663 3800
rect 8409 3737 8495 3760
rect 8577 3737 8663 3760
rect 12409 3800 12495 3823
rect 12577 3800 12663 3823
rect 12409 3760 12434 3800
rect 12434 3760 12474 3800
rect 12474 3760 12495 3800
rect 12577 3760 12598 3800
rect 12598 3760 12638 3800
rect 12638 3760 12663 3800
rect 12409 3737 12495 3760
rect 12577 3737 12663 3760
rect 16409 3800 16495 3823
rect 16577 3800 16663 3823
rect 16409 3760 16434 3800
rect 16434 3760 16474 3800
rect 16474 3760 16495 3800
rect 16577 3760 16598 3800
rect 16598 3760 16638 3800
rect 16638 3760 16663 3800
rect 16409 3737 16495 3760
rect 16577 3737 16663 3760
rect 20409 3800 20495 3823
rect 20577 3800 20663 3823
rect 20409 3760 20434 3800
rect 20434 3760 20474 3800
rect 20474 3760 20495 3800
rect 20577 3760 20598 3800
rect 20598 3760 20638 3800
rect 20638 3760 20663 3800
rect 20409 3737 20495 3760
rect 20577 3737 20663 3760
rect 24409 3800 24495 3823
rect 24577 3800 24663 3823
rect 24409 3760 24434 3800
rect 24434 3760 24474 3800
rect 24474 3760 24495 3800
rect 24577 3760 24598 3800
rect 24598 3760 24638 3800
rect 24638 3760 24663 3800
rect 24409 3737 24495 3760
rect 24577 3737 24663 3760
rect 28409 3800 28495 3823
rect 28577 3800 28663 3823
rect 28409 3760 28434 3800
rect 28434 3760 28474 3800
rect 28474 3760 28495 3800
rect 28577 3760 28598 3800
rect 28598 3760 28638 3800
rect 28638 3760 28663 3800
rect 28409 3737 28495 3760
rect 28577 3737 28663 3760
rect 32409 3800 32495 3823
rect 32577 3800 32663 3823
rect 32409 3760 32434 3800
rect 32434 3760 32474 3800
rect 32474 3760 32495 3800
rect 32577 3760 32598 3800
rect 32598 3760 32638 3800
rect 32638 3760 32663 3800
rect 32409 3737 32495 3760
rect 32577 3737 32663 3760
rect 36409 3800 36495 3823
rect 36577 3800 36663 3823
rect 36409 3760 36434 3800
rect 36434 3760 36474 3800
rect 36474 3760 36495 3800
rect 36577 3760 36598 3800
rect 36598 3760 36638 3800
rect 36638 3760 36663 3800
rect 36409 3737 36495 3760
rect 36577 3737 36663 3760
rect 40409 3800 40495 3823
rect 40577 3800 40663 3823
rect 40409 3760 40434 3800
rect 40434 3760 40474 3800
rect 40474 3760 40495 3800
rect 40577 3760 40598 3800
rect 40598 3760 40638 3800
rect 40638 3760 40663 3800
rect 40409 3737 40495 3760
rect 40577 3737 40663 3760
rect 44409 3800 44495 3823
rect 44577 3800 44663 3823
rect 44409 3760 44434 3800
rect 44434 3760 44474 3800
rect 44474 3760 44495 3800
rect 44577 3760 44598 3800
rect 44598 3760 44638 3800
rect 44638 3760 44663 3800
rect 44409 3737 44495 3760
rect 44577 3737 44663 3760
rect 48409 3800 48495 3823
rect 48577 3800 48663 3823
rect 48409 3760 48434 3800
rect 48434 3760 48474 3800
rect 48474 3760 48495 3800
rect 48577 3760 48598 3800
rect 48598 3760 48638 3800
rect 48638 3760 48663 3800
rect 48409 3737 48495 3760
rect 48577 3737 48663 3760
rect 52409 3800 52495 3823
rect 52577 3800 52663 3823
rect 52409 3760 52434 3800
rect 52434 3760 52474 3800
rect 52474 3760 52495 3800
rect 52577 3760 52598 3800
rect 52598 3760 52638 3800
rect 52638 3760 52663 3800
rect 52409 3737 52495 3760
rect 52577 3737 52663 3760
rect 56409 3800 56495 3823
rect 56577 3800 56663 3823
rect 56409 3760 56434 3800
rect 56434 3760 56474 3800
rect 56474 3760 56495 3800
rect 56577 3760 56598 3800
rect 56598 3760 56638 3800
rect 56638 3760 56663 3800
rect 56409 3737 56495 3760
rect 56577 3737 56663 3760
rect 60409 3800 60495 3823
rect 60577 3800 60663 3823
rect 60409 3760 60434 3800
rect 60434 3760 60474 3800
rect 60474 3760 60495 3800
rect 60577 3760 60598 3800
rect 60598 3760 60638 3800
rect 60638 3760 60663 3800
rect 60409 3737 60495 3760
rect 60577 3737 60663 3760
rect 64409 3800 64495 3823
rect 64577 3800 64663 3823
rect 64409 3760 64434 3800
rect 64434 3760 64474 3800
rect 64474 3760 64495 3800
rect 64577 3760 64598 3800
rect 64598 3760 64638 3800
rect 64638 3760 64663 3800
rect 64409 3737 64495 3760
rect 64577 3737 64663 3760
rect 68409 3800 68495 3823
rect 68577 3800 68663 3823
rect 68409 3760 68434 3800
rect 68434 3760 68474 3800
rect 68474 3760 68495 3800
rect 68577 3760 68598 3800
rect 68598 3760 68638 3800
rect 68638 3760 68663 3800
rect 68409 3737 68495 3760
rect 68577 3737 68663 3760
rect 72409 3800 72495 3823
rect 72577 3800 72663 3823
rect 72409 3760 72434 3800
rect 72434 3760 72474 3800
rect 72474 3760 72495 3800
rect 72577 3760 72598 3800
rect 72598 3760 72638 3800
rect 72638 3760 72663 3800
rect 72409 3737 72495 3760
rect 72577 3737 72663 3760
rect 76409 3800 76495 3823
rect 76577 3800 76663 3823
rect 76409 3760 76434 3800
rect 76434 3760 76474 3800
rect 76474 3760 76495 3800
rect 76577 3760 76598 3800
rect 76598 3760 76638 3800
rect 76638 3760 76663 3800
rect 76409 3737 76495 3760
rect 76577 3737 76663 3760
rect 80409 3800 80495 3823
rect 80577 3800 80663 3823
rect 80409 3760 80434 3800
rect 80434 3760 80474 3800
rect 80474 3760 80495 3800
rect 80577 3760 80598 3800
rect 80598 3760 80638 3800
rect 80638 3760 80663 3800
rect 80409 3737 80495 3760
rect 80577 3737 80663 3760
rect 84409 3800 84495 3823
rect 84577 3800 84663 3823
rect 84409 3760 84434 3800
rect 84434 3760 84474 3800
rect 84474 3760 84495 3800
rect 84577 3760 84598 3800
rect 84598 3760 84638 3800
rect 84638 3760 84663 3800
rect 84409 3737 84495 3760
rect 84577 3737 84663 3760
rect 88409 3800 88495 3823
rect 88577 3800 88663 3823
rect 88409 3760 88434 3800
rect 88434 3760 88474 3800
rect 88474 3760 88495 3800
rect 88577 3760 88598 3800
rect 88598 3760 88638 3800
rect 88638 3760 88663 3800
rect 88409 3737 88495 3760
rect 88577 3737 88663 3760
rect 92409 3800 92495 3823
rect 92577 3800 92663 3823
rect 92409 3760 92434 3800
rect 92434 3760 92474 3800
rect 92474 3760 92495 3800
rect 92577 3760 92598 3800
rect 92598 3760 92638 3800
rect 92638 3760 92663 3800
rect 92409 3737 92495 3760
rect 92577 3737 92663 3760
rect 96409 3800 96495 3823
rect 96577 3800 96663 3823
rect 96409 3760 96434 3800
rect 96434 3760 96474 3800
rect 96474 3760 96495 3800
rect 96577 3760 96598 3800
rect 96598 3760 96638 3800
rect 96638 3760 96663 3800
rect 96409 3737 96495 3760
rect 96577 3737 96663 3760
rect 3169 3044 3255 3067
rect 3337 3044 3423 3067
rect 3169 3004 3194 3044
rect 3194 3004 3234 3044
rect 3234 3004 3255 3044
rect 3337 3004 3358 3044
rect 3358 3004 3398 3044
rect 3398 3004 3423 3044
rect 3169 2981 3255 3004
rect 3337 2981 3423 3004
rect 7169 3044 7255 3067
rect 7337 3044 7423 3067
rect 7169 3004 7194 3044
rect 7194 3004 7234 3044
rect 7234 3004 7255 3044
rect 7337 3004 7358 3044
rect 7358 3004 7398 3044
rect 7398 3004 7423 3044
rect 7169 2981 7255 3004
rect 7337 2981 7423 3004
rect 11169 3044 11255 3067
rect 11337 3044 11423 3067
rect 11169 3004 11194 3044
rect 11194 3004 11234 3044
rect 11234 3004 11255 3044
rect 11337 3004 11358 3044
rect 11358 3004 11398 3044
rect 11398 3004 11423 3044
rect 11169 2981 11255 3004
rect 11337 2981 11423 3004
rect 15169 3044 15255 3067
rect 15337 3044 15423 3067
rect 15169 3004 15194 3044
rect 15194 3004 15234 3044
rect 15234 3004 15255 3044
rect 15337 3004 15358 3044
rect 15358 3004 15398 3044
rect 15398 3004 15423 3044
rect 15169 2981 15255 3004
rect 15337 2981 15423 3004
rect 19169 3044 19255 3067
rect 19337 3044 19423 3067
rect 19169 3004 19194 3044
rect 19194 3004 19234 3044
rect 19234 3004 19255 3044
rect 19337 3004 19358 3044
rect 19358 3004 19398 3044
rect 19398 3004 19423 3044
rect 19169 2981 19255 3004
rect 19337 2981 19423 3004
rect 23169 3044 23255 3067
rect 23337 3044 23423 3067
rect 23169 3004 23194 3044
rect 23194 3004 23234 3044
rect 23234 3004 23255 3044
rect 23337 3004 23358 3044
rect 23358 3004 23398 3044
rect 23398 3004 23423 3044
rect 23169 2981 23255 3004
rect 23337 2981 23423 3004
rect 27169 3044 27255 3067
rect 27337 3044 27423 3067
rect 27169 3004 27194 3044
rect 27194 3004 27234 3044
rect 27234 3004 27255 3044
rect 27337 3004 27358 3044
rect 27358 3004 27398 3044
rect 27398 3004 27423 3044
rect 27169 2981 27255 3004
rect 27337 2981 27423 3004
rect 31169 3044 31255 3067
rect 31337 3044 31423 3067
rect 31169 3004 31194 3044
rect 31194 3004 31234 3044
rect 31234 3004 31255 3044
rect 31337 3004 31358 3044
rect 31358 3004 31398 3044
rect 31398 3004 31423 3044
rect 31169 2981 31255 3004
rect 31337 2981 31423 3004
rect 35169 3044 35255 3067
rect 35337 3044 35423 3067
rect 35169 3004 35194 3044
rect 35194 3004 35234 3044
rect 35234 3004 35255 3044
rect 35337 3004 35358 3044
rect 35358 3004 35398 3044
rect 35398 3004 35423 3044
rect 35169 2981 35255 3004
rect 35337 2981 35423 3004
rect 39169 3044 39255 3067
rect 39337 3044 39423 3067
rect 39169 3004 39194 3044
rect 39194 3004 39234 3044
rect 39234 3004 39255 3044
rect 39337 3004 39358 3044
rect 39358 3004 39398 3044
rect 39398 3004 39423 3044
rect 39169 2981 39255 3004
rect 39337 2981 39423 3004
rect 43169 3044 43255 3067
rect 43337 3044 43423 3067
rect 43169 3004 43194 3044
rect 43194 3004 43234 3044
rect 43234 3004 43255 3044
rect 43337 3004 43358 3044
rect 43358 3004 43398 3044
rect 43398 3004 43423 3044
rect 43169 2981 43255 3004
rect 43337 2981 43423 3004
rect 47169 3044 47255 3067
rect 47337 3044 47423 3067
rect 47169 3004 47194 3044
rect 47194 3004 47234 3044
rect 47234 3004 47255 3044
rect 47337 3004 47358 3044
rect 47358 3004 47398 3044
rect 47398 3004 47423 3044
rect 47169 2981 47255 3004
rect 47337 2981 47423 3004
rect 51169 3044 51255 3067
rect 51337 3044 51423 3067
rect 51169 3004 51194 3044
rect 51194 3004 51234 3044
rect 51234 3004 51255 3044
rect 51337 3004 51358 3044
rect 51358 3004 51398 3044
rect 51398 3004 51423 3044
rect 51169 2981 51255 3004
rect 51337 2981 51423 3004
rect 55169 3044 55255 3067
rect 55337 3044 55423 3067
rect 55169 3004 55194 3044
rect 55194 3004 55234 3044
rect 55234 3004 55255 3044
rect 55337 3004 55358 3044
rect 55358 3004 55398 3044
rect 55398 3004 55423 3044
rect 55169 2981 55255 3004
rect 55337 2981 55423 3004
rect 59169 3044 59255 3067
rect 59337 3044 59423 3067
rect 59169 3004 59194 3044
rect 59194 3004 59234 3044
rect 59234 3004 59255 3044
rect 59337 3004 59358 3044
rect 59358 3004 59398 3044
rect 59398 3004 59423 3044
rect 59169 2981 59255 3004
rect 59337 2981 59423 3004
rect 63169 3044 63255 3067
rect 63337 3044 63423 3067
rect 63169 3004 63194 3044
rect 63194 3004 63234 3044
rect 63234 3004 63255 3044
rect 63337 3004 63358 3044
rect 63358 3004 63398 3044
rect 63398 3004 63423 3044
rect 63169 2981 63255 3004
rect 63337 2981 63423 3004
rect 67169 3044 67255 3067
rect 67337 3044 67423 3067
rect 67169 3004 67194 3044
rect 67194 3004 67234 3044
rect 67234 3004 67255 3044
rect 67337 3004 67358 3044
rect 67358 3004 67398 3044
rect 67398 3004 67423 3044
rect 67169 2981 67255 3004
rect 67337 2981 67423 3004
rect 71169 3044 71255 3067
rect 71337 3044 71423 3067
rect 71169 3004 71194 3044
rect 71194 3004 71234 3044
rect 71234 3004 71255 3044
rect 71337 3004 71358 3044
rect 71358 3004 71398 3044
rect 71398 3004 71423 3044
rect 71169 2981 71255 3004
rect 71337 2981 71423 3004
rect 75169 3044 75255 3067
rect 75337 3044 75423 3067
rect 75169 3004 75194 3044
rect 75194 3004 75234 3044
rect 75234 3004 75255 3044
rect 75337 3004 75358 3044
rect 75358 3004 75398 3044
rect 75398 3004 75423 3044
rect 75169 2981 75255 3004
rect 75337 2981 75423 3004
rect 79169 3044 79255 3067
rect 79337 3044 79423 3067
rect 79169 3004 79194 3044
rect 79194 3004 79234 3044
rect 79234 3004 79255 3044
rect 79337 3004 79358 3044
rect 79358 3004 79398 3044
rect 79398 3004 79423 3044
rect 79169 2981 79255 3004
rect 79337 2981 79423 3004
rect 83169 3044 83255 3067
rect 83337 3044 83423 3067
rect 83169 3004 83194 3044
rect 83194 3004 83234 3044
rect 83234 3004 83255 3044
rect 83337 3004 83358 3044
rect 83358 3004 83398 3044
rect 83398 3004 83423 3044
rect 83169 2981 83255 3004
rect 83337 2981 83423 3004
rect 87169 3044 87255 3067
rect 87337 3044 87423 3067
rect 87169 3004 87194 3044
rect 87194 3004 87234 3044
rect 87234 3004 87255 3044
rect 87337 3004 87358 3044
rect 87358 3004 87398 3044
rect 87398 3004 87423 3044
rect 87169 2981 87255 3004
rect 87337 2981 87423 3004
rect 91169 3044 91255 3067
rect 91337 3044 91423 3067
rect 91169 3004 91194 3044
rect 91194 3004 91234 3044
rect 91234 3004 91255 3044
rect 91337 3004 91358 3044
rect 91358 3004 91398 3044
rect 91398 3004 91423 3044
rect 91169 2981 91255 3004
rect 91337 2981 91423 3004
rect 95169 3044 95255 3067
rect 95337 3044 95423 3067
rect 95169 3004 95194 3044
rect 95194 3004 95234 3044
rect 95234 3004 95255 3044
rect 95337 3004 95358 3044
rect 95358 3004 95398 3044
rect 95398 3004 95423 3044
rect 95169 2981 95255 3004
rect 95337 2981 95423 3004
rect 99169 3044 99255 3067
rect 99337 3044 99423 3067
rect 99169 3004 99194 3044
rect 99194 3004 99234 3044
rect 99234 3004 99255 3044
rect 99337 3004 99358 3044
rect 99358 3004 99398 3044
rect 99398 3004 99423 3044
rect 99169 2981 99255 3004
rect 99337 2981 99423 3004
rect 4409 2288 4495 2311
rect 4577 2288 4663 2311
rect 4409 2248 4434 2288
rect 4434 2248 4474 2288
rect 4474 2248 4495 2288
rect 4577 2248 4598 2288
rect 4598 2248 4638 2288
rect 4638 2248 4663 2288
rect 4409 2225 4495 2248
rect 4577 2225 4663 2248
rect 8409 2288 8495 2311
rect 8577 2288 8663 2311
rect 8409 2248 8434 2288
rect 8434 2248 8474 2288
rect 8474 2248 8495 2288
rect 8577 2248 8598 2288
rect 8598 2248 8638 2288
rect 8638 2248 8663 2288
rect 8409 2225 8495 2248
rect 8577 2225 8663 2248
rect 12409 2288 12495 2311
rect 12577 2288 12663 2311
rect 12409 2248 12434 2288
rect 12434 2248 12474 2288
rect 12474 2248 12495 2288
rect 12577 2248 12598 2288
rect 12598 2248 12638 2288
rect 12638 2248 12663 2288
rect 12409 2225 12495 2248
rect 12577 2225 12663 2248
rect 16409 2288 16495 2311
rect 16577 2288 16663 2311
rect 16409 2248 16434 2288
rect 16434 2248 16474 2288
rect 16474 2248 16495 2288
rect 16577 2248 16598 2288
rect 16598 2248 16638 2288
rect 16638 2248 16663 2288
rect 16409 2225 16495 2248
rect 16577 2225 16663 2248
rect 20409 2288 20495 2311
rect 20577 2288 20663 2311
rect 20409 2248 20434 2288
rect 20434 2248 20474 2288
rect 20474 2248 20495 2288
rect 20577 2248 20598 2288
rect 20598 2248 20638 2288
rect 20638 2248 20663 2288
rect 20409 2225 20495 2248
rect 20577 2225 20663 2248
rect 24409 2288 24495 2311
rect 24577 2288 24663 2311
rect 24409 2248 24434 2288
rect 24434 2248 24474 2288
rect 24474 2248 24495 2288
rect 24577 2248 24598 2288
rect 24598 2248 24638 2288
rect 24638 2248 24663 2288
rect 24409 2225 24495 2248
rect 24577 2225 24663 2248
rect 28409 2288 28495 2311
rect 28577 2288 28663 2311
rect 28409 2248 28434 2288
rect 28434 2248 28474 2288
rect 28474 2248 28495 2288
rect 28577 2248 28598 2288
rect 28598 2248 28638 2288
rect 28638 2248 28663 2288
rect 28409 2225 28495 2248
rect 28577 2225 28663 2248
rect 32409 2288 32495 2311
rect 32577 2288 32663 2311
rect 32409 2248 32434 2288
rect 32434 2248 32474 2288
rect 32474 2248 32495 2288
rect 32577 2248 32598 2288
rect 32598 2248 32638 2288
rect 32638 2248 32663 2288
rect 32409 2225 32495 2248
rect 32577 2225 32663 2248
rect 36409 2288 36495 2311
rect 36577 2288 36663 2311
rect 36409 2248 36434 2288
rect 36434 2248 36474 2288
rect 36474 2248 36495 2288
rect 36577 2248 36598 2288
rect 36598 2248 36638 2288
rect 36638 2248 36663 2288
rect 36409 2225 36495 2248
rect 36577 2225 36663 2248
rect 40409 2288 40495 2311
rect 40577 2288 40663 2311
rect 40409 2248 40434 2288
rect 40434 2248 40474 2288
rect 40474 2248 40495 2288
rect 40577 2248 40598 2288
rect 40598 2248 40638 2288
rect 40638 2248 40663 2288
rect 40409 2225 40495 2248
rect 40577 2225 40663 2248
rect 44409 2288 44495 2311
rect 44577 2288 44663 2311
rect 44409 2248 44434 2288
rect 44434 2248 44474 2288
rect 44474 2248 44495 2288
rect 44577 2248 44598 2288
rect 44598 2248 44638 2288
rect 44638 2248 44663 2288
rect 44409 2225 44495 2248
rect 44577 2225 44663 2248
rect 48409 2288 48495 2311
rect 48577 2288 48663 2311
rect 48409 2248 48434 2288
rect 48434 2248 48474 2288
rect 48474 2248 48495 2288
rect 48577 2248 48598 2288
rect 48598 2248 48638 2288
rect 48638 2248 48663 2288
rect 48409 2225 48495 2248
rect 48577 2225 48663 2248
rect 52409 2288 52495 2311
rect 52577 2288 52663 2311
rect 52409 2248 52434 2288
rect 52434 2248 52474 2288
rect 52474 2248 52495 2288
rect 52577 2248 52598 2288
rect 52598 2248 52638 2288
rect 52638 2248 52663 2288
rect 52409 2225 52495 2248
rect 52577 2225 52663 2248
rect 56409 2288 56495 2311
rect 56577 2288 56663 2311
rect 56409 2248 56434 2288
rect 56434 2248 56474 2288
rect 56474 2248 56495 2288
rect 56577 2248 56598 2288
rect 56598 2248 56638 2288
rect 56638 2248 56663 2288
rect 56409 2225 56495 2248
rect 56577 2225 56663 2248
rect 60409 2288 60495 2311
rect 60577 2288 60663 2311
rect 60409 2248 60434 2288
rect 60434 2248 60474 2288
rect 60474 2248 60495 2288
rect 60577 2248 60598 2288
rect 60598 2248 60638 2288
rect 60638 2248 60663 2288
rect 60409 2225 60495 2248
rect 60577 2225 60663 2248
rect 64409 2288 64495 2311
rect 64577 2288 64663 2311
rect 64409 2248 64434 2288
rect 64434 2248 64474 2288
rect 64474 2248 64495 2288
rect 64577 2248 64598 2288
rect 64598 2248 64638 2288
rect 64638 2248 64663 2288
rect 64409 2225 64495 2248
rect 64577 2225 64663 2248
rect 68409 2288 68495 2311
rect 68577 2288 68663 2311
rect 68409 2248 68434 2288
rect 68434 2248 68474 2288
rect 68474 2248 68495 2288
rect 68577 2248 68598 2288
rect 68598 2248 68638 2288
rect 68638 2248 68663 2288
rect 68409 2225 68495 2248
rect 68577 2225 68663 2248
rect 72409 2288 72495 2311
rect 72577 2288 72663 2311
rect 72409 2248 72434 2288
rect 72434 2248 72474 2288
rect 72474 2248 72495 2288
rect 72577 2248 72598 2288
rect 72598 2248 72638 2288
rect 72638 2248 72663 2288
rect 72409 2225 72495 2248
rect 72577 2225 72663 2248
rect 76409 2288 76495 2311
rect 76577 2288 76663 2311
rect 76409 2248 76434 2288
rect 76434 2248 76474 2288
rect 76474 2248 76495 2288
rect 76577 2248 76598 2288
rect 76598 2248 76638 2288
rect 76638 2248 76663 2288
rect 76409 2225 76495 2248
rect 76577 2225 76663 2248
rect 80409 2288 80495 2311
rect 80577 2288 80663 2311
rect 80409 2248 80434 2288
rect 80434 2248 80474 2288
rect 80474 2248 80495 2288
rect 80577 2248 80598 2288
rect 80598 2248 80638 2288
rect 80638 2248 80663 2288
rect 80409 2225 80495 2248
rect 80577 2225 80663 2248
rect 84409 2288 84495 2311
rect 84577 2288 84663 2311
rect 84409 2248 84434 2288
rect 84434 2248 84474 2288
rect 84474 2248 84495 2288
rect 84577 2248 84598 2288
rect 84598 2248 84638 2288
rect 84638 2248 84663 2288
rect 84409 2225 84495 2248
rect 84577 2225 84663 2248
rect 88409 2288 88495 2311
rect 88577 2288 88663 2311
rect 88409 2248 88434 2288
rect 88434 2248 88474 2288
rect 88474 2248 88495 2288
rect 88577 2248 88598 2288
rect 88598 2248 88638 2288
rect 88638 2248 88663 2288
rect 88409 2225 88495 2248
rect 88577 2225 88663 2248
rect 92409 2288 92495 2311
rect 92577 2288 92663 2311
rect 92409 2248 92434 2288
rect 92434 2248 92474 2288
rect 92474 2248 92495 2288
rect 92577 2248 92598 2288
rect 92598 2248 92638 2288
rect 92638 2248 92663 2288
rect 92409 2225 92495 2248
rect 92577 2225 92663 2248
rect 96409 2288 96495 2311
rect 96577 2288 96663 2311
rect 96409 2248 96434 2288
rect 96434 2248 96474 2288
rect 96474 2248 96495 2288
rect 96577 2248 96598 2288
rect 96598 2248 96638 2288
rect 96638 2248 96663 2288
rect 96409 2225 96495 2248
rect 96577 2225 96663 2248
rect 3169 1532 3255 1555
rect 3337 1532 3423 1555
rect 3169 1492 3194 1532
rect 3194 1492 3234 1532
rect 3234 1492 3255 1532
rect 3337 1492 3358 1532
rect 3358 1492 3398 1532
rect 3398 1492 3423 1532
rect 3169 1469 3255 1492
rect 3337 1469 3423 1492
rect 7169 1532 7255 1555
rect 7337 1532 7423 1555
rect 7169 1492 7194 1532
rect 7194 1492 7234 1532
rect 7234 1492 7255 1532
rect 7337 1492 7358 1532
rect 7358 1492 7398 1532
rect 7398 1492 7423 1532
rect 7169 1469 7255 1492
rect 7337 1469 7423 1492
rect 11169 1532 11255 1555
rect 11337 1532 11423 1555
rect 11169 1492 11194 1532
rect 11194 1492 11234 1532
rect 11234 1492 11255 1532
rect 11337 1492 11358 1532
rect 11358 1492 11398 1532
rect 11398 1492 11423 1532
rect 11169 1469 11255 1492
rect 11337 1469 11423 1492
rect 15169 1532 15255 1555
rect 15337 1532 15423 1555
rect 15169 1492 15194 1532
rect 15194 1492 15234 1532
rect 15234 1492 15255 1532
rect 15337 1492 15358 1532
rect 15358 1492 15398 1532
rect 15398 1492 15423 1532
rect 15169 1469 15255 1492
rect 15337 1469 15423 1492
rect 19169 1532 19255 1555
rect 19337 1532 19423 1555
rect 19169 1492 19194 1532
rect 19194 1492 19234 1532
rect 19234 1492 19255 1532
rect 19337 1492 19358 1532
rect 19358 1492 19398 1532
rect 19398 1492 19423 1532
rect 19169 1469 19255 1492
rect 19337 1469 19423 1492
rect 23169 1532 23255 1555
rect 23337 1532 23423 1555
rect 23169 1492 23194 1532
rect 23194 1492 23234 1532
rect 23234 1492 23255 1532
rect 23337 1492 23358 1532
rect 23358 1492 23398 1532
rect 23398 1492 23423 1532
rect 23169 1469 23255 1492
rect 23337 1469 23423 1492
rect 27169 1532 27255 1555
rect 27337 1532 27423 1555
rect 27169 1492 27194 1532
rect 27194 1492 27234 1532
rect 27234 1492 27255 1532
rect 27337 1492 27358 1532
rect 27358 1492 27398 1532
rect 27398 1492 27423 1532
rect 27169 1469 27255 1492
rect 27337 1469 27423 1492
rect 31169 1532 31255 1555
rect 31337 1532 31423 1555
rect 31169 1492 31194 1532
rect 31194 1492 31234 1532
rect 31234 1492 31255 1532
rect 31337 1492 31358 1532
rect 31358 1492 31398 1532
rect 31398 1492 31423 1532
rect 31169 1469 31255 1492
rect 31337 1469 31423 1492
rect 35169 1532 35255 1555
rect 35337 1532 35423 1555
rect 35169 1492 35194 1532
rect 35194 1492 35234 1532
rect 35234 1492 35255 1532
rect 35337 1492 35358 1532
rect 35358 1492 35398 1532
rect 35398 1492 35423 1532
rect 35169 1469 35255 1492
rect 35337 1469 35423 1492
rect 39169 1532 39255 1555
rect 39337 1532 39423 1555
rect 39169 1492 39194 1532
rect 39194 1492 39234 1532
rect 39234 1492 39255 1532
rect 39337 1492 39358 1532
rect 39358 1492 39398 1532
rect 39398 1492 39423 1532
rect 39169 1469 39255 1492
rect 39337 1469 39423 1492
rect 43169 1532 43255 1555
rect 43337 1532 43423 1555
rect 43169 1492 43194 1532
rect 43194 1492 43234 1532
rect 43234 1492 43255 1532
rect 43337 1492 43358 1532
rect 43358 1492 43398 1532
rect 43398 1492 43423 1532
rect 43169 1469 43255 1492
rect 43337 1469 43423 1492
rect 47169 1532 47255 1555
rect 47337 1532 47423 1555
rect 47169 1492 47194 1532
rect 47194 1492 47234 1532
rect 47234 1492 47255 1532
rect 47337 1492 47358 1532
rect 47358 1492 47398 1532
rect 47398 1492 47423 1532
rect 47169 1469 47255 1492
rect 47337 1469 47423 1492
rect 51169 1532 51255 1555
rect 51337 1532 51423 1555
rect 51169 1492 51194 1532
rect 51194 1492 51234 1532
rect 51234 1492 51255 1532
rect 51337 1492 51358 1532
rect 51358 1492 51398 1532
rect 51398 1492 51423 1532
rect 51169 1469 51255 1492
rect 51337 1469 51423 1492
rect 55169 1532 55255 1555
rect 55337 1532 55423 1555
rect 55169 1492 55194 1532
rect 55194 1492 55234 1532
rect 55234 1492 55255 1532
rect 55337 1492 55358 1532
rect 55358 1492 55398 1532
rect 55398 1492 55423 1532
rect 55169 1469 55255 1492
rect 55337 1469 55423 1492
rect 59169 1532 59255 1555
rect 59337 1532 59423 1555
rect 59169 1492 59194 1532
rect 59194 1492 59234 1532
rect 59234 1492 59255 1532
rect 59337 1492 59358 1532
rect 59358 1492 59398 1532
rect 59398 1492 59423 1532
rect 59169 1469 59255 1492
rect 59337 1469 59423 1492
rect 63169 1532 63255 1555
rect 63337 1532 63423 1555
rect 63169 1492 63194 1532
rect 63194 1492 63234 1532
rect 63234 1492 63255 1532
rect 63337 1492 63358 1532
rect 63358 1492 63398 1532
rect 63398 1492 63423 1532
rect 63169 1469 63255 1492
rect 63337 1469 63423 1492
rect 67169 1532 67255 1555
rect 67337 1532 67423 1555
rect 67169 1492 67194 1532
rect 67194 1492 67234 1532
rect 67234 1492 67255 1532
rect 67337 1492 67358 1532
rect 67358 1492 67398 1532
rect 67398 1492 67423 1532
rect 67169 1469 67255 1492
rect 67337 1469 67423 1492
rect 71169 1532 71255 1555
rect 71337 1532 71423 1555
rect 71169 1492 71194 1532
rect 71194 1492 71234 1532
rect 71234 1492 71255 1532
rect 71337 1492 71358 1532
rect 71358 1492 71398 1532
rect 71398 1492 71423 1532
rect 71169 1469 71255 1492
rect 71337 1469 71423 1492
rect 75169 1532 75255 1555
rect 75337 1532 75423 1555
rect 75169 1492 75194 1532
rect 75194 1492 75234 1532
rect 75234 1492 75255 1532
rect 75337 1492 75358 1532
rect 75358 1492 75398 1532
rect 75398 1492 75423 1532
rect 75169 1469 75255 1492
rect 75337 1469 75423 1492
rect 79169 1532 79255 1555
rect 79337 1532 79423 1555
rect 79169 1492 79194 1532
rect 79194 1492 79234 1532
rect 79234 1492 79255 1532
rect 79337 1492 79358 1532
rect 79358 1492 79398 1532
rect 79398 1492 79423 1532
rect 79169 1469 79255 1492
rect 79337 1469 79423 1492
rect 83169 1532 83255 1555
rect 83337 1532 83423 1555
rect 83169 1492 83194 1532
rect 83194 1492 83234 1532
rect 83234 1492 83255 1532
rect 83337 1492 83358 1532
rect 83358 1492 83398 1532
rect 83398 1492 83423 1532
rect 83169 1469 83255 1492
rect 83337 1469 83423 1492
rect 87169 1532 87255 1555
rect 87337 1532 87423 1555
rect 87169 1492 87194 1532
rect 87194 1492 87234 1532
rect 87234 1492 87255 1532
rect 87337 1492 87358 1532
rect 87358 1492 87398 1532
rect 87398 1492 87423 1532
rect 87169 1469 87255 1492
rect 87337 1469 87423 1492
rect 91169 1532 91255 1555
rect 91337 1532 91423 1555
rect 91169 1492 91194 1532
rect 91194 1492 91234 1532
rect 91234 1492 91255 1532
rect 91337 1492 91358 1532
rect 91358 1492 91398 1532
rect 91398 1492 91423 1532
rect 91169 1469 91255 1492
rect 91337 1469 91423 1492
rect 95169 1532 95255 1555
rect 95337 1532 95423 1555
rect 95169 1492 95194 1532
rect 95194 1492 95234 1532
rect 95234 1492 95255 1532
rect 95337 1492 95358 1532
rect 95358 1492 95398 1532
rect 95398 1492 95423 1532
rect 95169 1469 95255 1492
rect 95337 1469 95423 1492
rect 99169 1532 99255 1555
rect 99337 1532 99423 1555
rect 99169 1492 99194 1532
rect 99194 1492 99234 1532
rect 99234 1492 99255 1532
rect 99337 1492 99358 1532
rect 99358 1492 99398 1532
rect 99398 1492 99423 1532
rect 99169 1469 99255 1492
rect 99337 1469 99423 1492
rect 4409 776 4495 799
rect 4577 776 4663 799
rect 4409 736 4434 776
rect 4434 736 4474 776
rect 4474 736 4495 776
rect 4577 736 4598 776
rect 4598 736 4638 776
rect 4638 736 4663 776
rect 4409 713 4495 736
rect 4577 713 4663 736
rect 8409 776 8495 799
rect 8577 776 8663 799
rect 8409 736 8434 776
rect 8434 736 8474 776
rect 8474 736 8495 776
rect 8577 736 8598 776
rect 8598 736 8638 776
rect 8638 736 8663 776
rect 8409 713 8495 736
rect 8577 713 8663 736
rect 12409 776 12495 799
rect 12577 776 12663 799
rect 12409 736 12434 776
rect 12434 736 12474 776
rect 12474 736 12495 776
rect 12577 736 12598 776
rect 12598 736 12638 776
rect 12638 736 12663 776
rect 12409 713 12495 736
rect 12577 713 12663 736
rect 16409 776 16495 799
rect 16577 776 16663 799
rect 16409 736 16434 776
rect 16434 736 16474 776
rect 16474 736 16495 776
rect 16577 736 16598 776
rect 16598 736 16638 776
rect 16638 736 16663 776
rect 16409 713 16495 736
rect 16577 713 16663 736
rect 20409 776 20495 799
rect 20577 776 20663 799
rect 20409 736 20434 776
rect 20434 736 20474 776
rect 20474 736 20495 776
rect 20577 736 20598 776
rect 20598 736 20638 776
rect 20638 736 20663 776
rect 20409 713 20495 736
rect 20577 713 20663 736
rect 24409 776 24495 799
rect 24577 776 24663 799
rect 24409 736 24434 776
rect 24434 736 24474 776
rect 24474 736 24495 776
rect 24577 736 24598 776
rect 24598 736 24638 776
rect 24638 736 24663 776
rect 24409 713 24495 736
rect 24577 713 24663 736
rect 28409 776 28495 799
rect 28577 776 28663 799
rect 28409 736 28434 776
rect 28434 736 28474 776
rect 28474 736 28495 776
rect 28577 736 28598 776
rect 28598 736 28638 776
rect 28638 736 28663 776
rect 28409 713 28495 736
rect 28577 713 28663 736
rect 32409 776 32495 799
rect 32577 776 32663 799
rect 32409 736 32434 776
rect 32434 736 32474 776
rect 32474 736 32495 776
rect 32577 736 32598 776
rect 32598 736 32638 776
rect 32638 736 32663 776
rect 32409 713 32495 736
rect 32577 713 32663 736
rect 36409 776 36495 799
rect 36577 776 36663 799
rect 36409 736 36434 776
rect 36434 736 36474 776
rect 36474 736 36495 776
rect 36577 736 36598 776
rect 36598 736 36638 776
rect 36638 736 36663 776
rect 36409 713 36495 736
rect 36577 713 36663 736
rect 40409 776 40495 799
rect 40577 776 40663 799
rect 40409 736 40434 776
rect 40434 736 40474 776
rect 40474 736 40495 776
rect 40577 736 40598 776
rect 40598 736 40638 776
rect 40638 736 40663 776
rect 40409 713 40495 736
rect 40577 713 40663 736
rect 44409 776 44495 799
rect 44577 776 44663 799
rect 44409 736 44434 776
rect 44434 736 44474 776
rect 44474 736 44495 776
rect 44577 736 44598 776
rect 44598 736 44638 776
rect 44638 736 44663 776
rect 44409 713 44495 736
rect 44577 713 44663 736
rect 48409 776 48495 799
rect 48577 776 48663 799
rect 48409 736 48434 776
rect 48434 736 48474 776
rect 48474 736 48495 776
rect 48577 736 48598 776
rect 48598 736 48638 776
rect 48638 736 48663 776
rect 48409 713 48495 736
rect 48577 713 48663 736
rect 52409 776 52495 799
rect 52577 776 52663 799
rect 52409 736 52434 776
rect 52434 736 52474 776
rect 52474 736 52495 776
rect 52577 736 52598 776
rect 52598 736 52638 776
rect 52638 736 52663 776
rect 52409 713 52495 736
rect 52577 713 52663 736
rect 56409 776 56495 799
rect 56577 776 56663 799
rect 56409 736 56434 776
rect 56434 736 56474 776
rect 56474 736 56495 776
rect 56577 736 56598 776
rect 56598 736 56638 776
rect 56638 736 56663 776
rect 56409 713 56495 736
rect 56577 713 56663 736
rect 60409 776 60495 799
rect 60577 776 60663 799
rect 60409 736 60434 776
rect 60434 736 60474 776
rect 60474 736 60495 776
rect 60577 736 60598 776
rect 60598 736 60638 776
rect 60638 736 60663 776
rect 60409 713 60495 736
rect 60577 713 60663 736
rect 64409 776 64495 799
rect 64577 776 64663 799
rect 64409 736 64434 776
rect 64434 736 64474 776
rect 64474 736 64495 776
rect 64577 736 64598 776
rect 64598 736 64638 776
rect 64638 736 64663 776
rect 64409 713 64495 736
rect 64577 713 64663 736
rect 68409 776 68495 799
rect 68577 776 68663 799
rect 68409 736 68434 776
rect 68434 736 68474 776
rect 68474 736 68495 776
rect 68577 736 68598 776
rect 68598 736 68638 776
rect 68638 736 68663 776
rect 68409 713 68495 736
rect 68577 713 68663 736
rect 72409 776 72495 799
rect 72577 776 72663 799
rect 72409 736 72434 776
rect 72434 736 72474 776
rect 72474 736 72495 776
rect 72577 736 72598 776
rect 72598 736 72638 776
rect 72638 736 72663 776
rect 72409 713 72495 736
rect 72577 713 72663 736
rect 76409 776 76495 799
rect 76577 776 76663 799
rect 76409 736 76434 776
rect 76434 736 76474 776
rect 76474 736 76495 776
rect 76577 736 76598 776
rect 76598 736 76638 776
rect 76638 736 76663 776
rect 76409 713 76495 736
rect 76577 713 76663 736
rect 80409 776 80495 799
rect 80577 776 80663 799
rect 80409 736 80434 776
rect 80434 736 80474 776
rect 80474 736 80495 776
rect 80577 736 80598 776
rect 80598 736 80638 776
rect 80638 736 80663 776
rect 80409 713 80495 736
rect 80577 713 80663 736
rect 84409 776 84495 799
rect 84577 776 84663 799
rect 84409 736 84434 776
rect 84434 736 84474 776
rect 84474 736 84495 776
rect 84577 736 84598 776
rect 84598 736 84638 776
rect 84638 736 84663 776
rect 84409 713 84495 736
rect 84577 713 84663 736
rect 88409 776 88495 799
rect 88577 776 88663 799
rect 88409 736 88434 776
rect 88434 736 88474 776
rect 88474 736 88495 776
rect 88577 736 88598 776
rect 88598 736 88638 776
rect 88638 736 88663 776
rect 88409 713 88495 736
rect 88577 713 88663 736
rect 92409 776 92495 799
rect 92577 776 92663 799
rect 92409 736 92434 776
rect 92434 736 92474 776
rect 92474 736 92495 776
rect 92577 736 92598 776
rect 92598 736 92638 776
rect 92638 736 92663 776
rect 92409 713 92495 736
rect 92577 713 92663 736
rect 96409 776 96495 799
rect 96577 776 96663 799
rect 96409 736 96434 776
rect 96434 736 96474 776
rect 96474 736 96495 776
rect 96577 736 96598 776
rect 96598 736 96638 776
rect 96638 736 96663 776
rect 96409 713 96495 736
rect 96577 713 96663 736
<< metal6 >>
rect 3076 37843 3516 38600
rect 3076 37757 3169 37843
rect 3255 37757 3337 37843
rect 3423 37757 3516 37843
rect 3076 36331 3516 37757
rect 3076 36245 3169 36331
rect 3255 36245 3337 36331
rect 3423 36245 3516 36331
rect 3076 35666 3516 36245
rect 3076 35286 3106 35666
rect 3486 35286 3516 35666
rect 3076 34819 3516 35286
rect 3076 34733 3169 34819
rect 3255 34733 3337 34819
rect 3423 34733 3516 34819
rect 3076 33307 3516 34733
rect 3076 33221 3169 33307
rect 3255 33221 3337 33307
rect 3423 33221 3516 33307
rect 3076 31795 3516 33221
rect 3076 31709 3169 31795
rect 3255 31709 3337 31795
rect 3423 31709 3516 31795
rect 3076 31666 3516 31709
rect 3076 31286 3106 31666
rect 3486 31286 3516 31666
rect 3076 30283 3516 31286
rect 3076 30197 3169 30283
rect 3255 30197 3337 30283
rect 3423 30197 3516 30283
rect 3076 28771 3516 30197
rect 3076 28685 3169 28771
rect 3255 28685 3337 28771
rect 3423 28685 3516 28771
rect 3076 27666 3516 28685
rect 3076 27286 3106 27666
rect 3486 27286 3516 27666
rect 3076 27259 3516 27286
rect 3076 27173 3169 27259
rect 3255 27173 3337 27259
rect 3423 27173 3516 27259
rect 3076 25747 3516 27173
rect 3076 25661 3169 25747
rect 3255 25661 3337 25747
rect 3423 25661 3516 25747
rect 3076 24235 3516 25661
rect 3076 24149 3169 24235
rect 3255 24149 3337 24235
rect 3423 24149 3516 24235
rect 3076 23666 3516 24149
rect 3076 23286 3106 23666
rect 3486 23286 3516 23666
rect 3076 22723 3516 23286
rect 3076 22637 3169 22723
rect 3255 22637 3337 22723
rect 3423 22637 3516 22723
rect 3076 21211 3516 22637
rect 3076 21125 3169 21211
rect 3255 21125 3337 21211
rect 3423 21125 3516 21211
rect 3076 19699 3516 21125
rect 3076 19666 3169 19699
rect 3255 19666 3337 19699
rect 3423 19666 3516 19699
rect 3076 19286 3106 19666
rect 3486 19286 3516 19666
rect 3076 18187 3516 19286
rect 3076 18101 3169 18187
rect 3255 18101 3337 18187
rect 3423 18101 3516 18187
rect 3076 16675 3516 18101
rect 3076 16589 3169 16675
rect 3255 16589 3337 16675
rect 3423 16589 3516 16675
rect 3076 15666 3516 16589
rect 3076 15286 3106 15666
rect 3486 15286 3516 15666
rect 3076 15163 3516 15286
rect 3076 15077 3169 15163
rect 3255 15077 3337 15163
rect 3423 15077 3516 15163
rect 3076 13651 3516 15077
rect 3076 13565 3169 13651
rect 3255 13565 3337 13651
rect 3423 13565 3516 13651
rect 3076 12139 3516 13565
rect 3076 12053 3169 12139
rect 3255 12053 3337 12139
rect 3423 12053 3516 12139
rect 3076 11666 3516 12053
rect 3076 11286 3106 11666
rect 3486 11286 3516 11666
rect 3076 10627 3516 11286
rect 3076 10541 3169 10627
rect 3255 10541 3337 10627
rect 3423 10541 3516 10627
rect 3076 9115 3516 10541
rect 3076 9029 3169 9115
rect 3255 9029 3337 9115
rect 3423 9029 3516 9115
rect 3076 7666 3516 9029
rect 3076 7286 3106 7666
rect 3486 7286 3516 7666
rect 3076 6091 3516 7286
rect 3076 6005 3169 6091
rect 3255 6005 3337 6091
rect 3423 6005 3516 6091
rect 3076 4579 3516 6005
rect 3076 4493 3169 4579
rect 3255 4493 3337 4579
rect 3423 4493 3516 4579
rect 3076 3666 3516 4493
rect 3076 3286 3106 3666
rect 3486 3286 3516 3666
rect 3076 3067 3516 3286
rect 3076 2981 3169 3067
rect 3255 2981 3337 3067
rect 3423 2981 3516 3067
rect 3076 1555 3516 2981
rect 3076 1469 3169 1555
rect 3255 1469 3337 1555
rect 3423 1469 3516 1555
rect 3076 712 3516 1469
rect 4316 38599 4756 38682
rect 4316 38513 4409 38599
rect 4495 38513 4577 38599
rect 4663 38513 4756 38599
rect 4316 37087 4756 38513
rect 4316 37001 4409 37087
rect 4495 37001 4577 37087
rect 4663 37001 4756 37087
rect 4316 36906 4756 37001
rect 4316 36526 4346 36906
rect 4726 36526 4756 36906
rect 4316 35575 4756 36526
rect 4316 35489 4409 35575
rect 4495 35489 4577 35575
rect 4663 35489 4756 35575
rect 4316 34063 4756 35489
rect 4316 33977 4409 34063
rect 4495 33977 4577 34063
rect 4663 33977 4756 34063
rect 4316 32906 4756 33977
rect 4316 32526 4346 32906
rect 4726 32526 4756 32906
rect 4316 32465 4409 32526
rect 4495 32465 4577 32526
rect 4663 32465 4756 32526
rect 4316 31039 4756 32465
rect 4316 30953 4409 31039
rect 4495 30953 4577 31039
rect 4663 30953 4756 31039
rect 4316 29527 4756 30953
rect 4316 29441 4409 29527
rect 4495 29441 4577 29527
rect 4663 29441 4756 29527
rect 4316 28906 4756 29441
rect 4316 28526 4346 28906
rect 4726 28526 4756 28906
rect 4316 28015 4756 28526
rect 4316 27929 4409 28015
rect 4495 27929 4577 28015
rect 4663 27929 4756 28015
rect 4316 26503 4756 27929
rect 4316 26417 4409 26503
rect 4495 26417 4577 26503
rect 4663 26417 4756 26503
rect 4316 24991 4756 26417
rect 4316 24906 4409 24991
rect 4495 24906 4577 24991
rect 4663 24906 4756 24991
rect 4316 24526 4346 24906
rect 4726 24526 4756 24906
rect 4316 23479 4756 24526
rect 4316 23393 4409 23479
rect 4495 23393 4577 23479
rect 4663 23393 4756 23479
rect 4316 21967 4756 23393
rect 4316 21881 4409 21967
rect 4495 21881 4577 21967
rect 4663 21881 4756 21967
rect 4316 20906 4756 21881
rect 4316 20526 4346 20906
rect 4726 20526 4756 20906
rect 4316 20455 4756 20526
rect 4316 20369 4409 20455
rect 4495 20369 4577 20455
rect 4663 20369 4756 20455
rect 4316 18943 4756 20369
rect 4316 18857 4409 18943
rect 4495 18857 4577 18943
rect 4663 18857 4756 18943
rect 4316 17431 4756 18857
rect 4316 17345 4409 17431
rect 4495 17345 4577 17431
rect 4663 17345 4756 17431
rect 4316 16906 4756 17345
rect 4316 16526 4346 16906
rect 4726 16526 4756 16906
rect 4316 15919 4756 16526
rect 4316 15833 4409 15919
rect 4495 15833 4577 15919
rect 4663 15833 4756 15919
rect 4316 14407 4756 15833
rect 4316 14321 4409 14407
rect 4495 14321 4577 14407
rect 4663 14321 4756 14407
rect 4316 12906 4756 14321
rect 4316 12526 4346 12906
rect 4726 12526 4756 12906
rect 4316 11383 4756 12526
rect 4316 11297 4409 11383
rect 4495 11297 4577 11383
rect 4663 11297 4756 11383
rect 4316 9871 4756 11297
rect 4316 9785 4409 9871
rect 4495 9785 4577 9871
rect 4663 9785 4756 9871
rect 4316 8906 4756 9785
rect 4316 8526 4346 8906
rect 4726 8526 4756 8906
rect 4316 8359 4756 8526
rect 4316 8273 4409 8359
rect 4495 8273 4577 8359
rect 4663 8273 4756 8359
rect 4316 6847 4756 8273
rect 4316 6761 4409 6847
rect 4495 6761 4577 6847
rect 4663 6761 4756 6847
rect 4316 5335 4756 6761
rect 4316 5249 4409 5335
rect 4495 5249 4577 5335
rect 4663 5249 4756 5335
rect 4316 4906 4756 5249
rect 4316 4526 4346 4906
rect 4726 4526 4756 4906
rect 4316 3823 4756 4526
rect 4316 3737 4409 3823
rect 4495 3737 4577 3823
rect 4663 3737 4756 3823
rect 4316 2311 4756 3737
rect 4316 2225 4409 2311
rect 4495 2225 4577 2311
rect 4663 2225 4756 2311
rect 4316 799 4756 2225
rect 4316 713 4409 799
rect 4495 713 4577 799
rect 4663 713 4756 799
rect 4316 630 4756 713
rect 7076 37843 7516 38600
rect 7076 37757 7169 37843
rect 7255 37757 7337 37843
rect 7423 37757 7516 37843
rect 7076 36331 7516 37757
rect 7076 36245 7169 36331
rect 7255 36245 7337 36331
rect 7423 36245 7516 36331
rect 7076 35666 7516 36245
rect 7076 35286 7106 35666
rect 7486 35286 7516 35666
rect 7076 34819 7516 35286
rect 7076 34733 7169 34819
rect 7255 34733 7337 34819
rect 7423 34733 7516 34819
rect 7076 33307 7516 34733
rect 7076 33221 7169 33307
rect 7255 33221 7337 33307
rect 7423 33221 7516 33307
rect 7076 31795 7516 33221
rect 7076 31709 7169 31795
rect 7255 31709 7337 31795
rect 7423 31709 7516 31795
rect 7076 31666 7516 31709
rect 7076 31286 7106 31666
rect 7486 31286 7516 31666
rect 7076 30283 7516 31286
rect 7076 30197 7169 30283
rect 7255 30197 7337 30283
rect 7423 30197 7516 30283
rect 7076 28771 7516 30197
rect 7076 28685 7169 28771
rect 7255 28685 7337 28771
rect 7423 28685 7516 28771
rect 7076 27666 7516 28685
rect 7076 27286 7106 27666
rect 7486 27286 7516 27666
rect 7076 27259 7516 27286
rect 7076 27173 7169 27259
rect 7255 27173 7337 27259
rect 7423 27173 7516 27259
rect 7076 25747 7516 27173
rect 7076 25661 7169 25747
rect 7255 25661 7337 25747
rect 7423 25661 7516 25747
rect 7076 24235 7516 25661
rect 7076 24149 7169 24235
rect 7255 24149 7337 24235
rect 7423 24149 7516 24235
rect 7076 23666 7516 24149
rect 7076 23286 7106 23666
rect 7486 23286 7516 23666
rect 7076 22723 7516 23286
rect 7076 22637 7169 22723
rect 7255 22637 7337 22723
rect 7423 22637 7516 22723
rect 7076 21211 7516 22637
rect 7076 21125 7169 21211
rect 7255 21125 7337 21211
rect 7423 21125 7516 21211
rect 7076 19699 7516 21125
rect 7076 19666 7169 19699
rect 7255 19666 7337 19699
rect 7423 19666 7516 19699
rect 7076 19286 7106 19666
rect 7486 19286 7516 19666
rect 7076 18187 7516 19286
rect 7076 18101 7169 18187
rect 7255 18101 7337 18187
rect 7423 18101 7516 18187
rect 7076 16675 7516 18101
rect 7076 16589 7169 16675
rect 7255 16589 7337 16675
rect 7423 16589 7516 16675
rect 7076 15666 7516 16589
rect 7076 15286 7106 15666
rect 7486 15286 7516 15666
rect 7076 15163 7516 15286
rect 7076 15077 7169 15163
rect 7255 15077 7337 15163
rect 7423 15077 7516 15163
rect 7076 13651 7516 15077
rect 7076 13565 7169 13651
rect 7255 13565 7337 13651
rect 7423 13565 7516 13651
rect 7076 12139 7516 13565
rect 7076 12053 7169 12139
rect 7255 12053 7337 12139
rect 7423 12053 7516 12139
rect 7076 11666 7516 12053
rect 7076 11286 7106 11666
rect 7486 11286 7516 11666
rect 7076 10627 7516 11286
rect 7076 10541 7169 10627
rect 7255 10541 7337 10627
rect 7423 10541 7516 10627
rect 7076 9115 7516 10541
rect 7076 9029 7169 9115
rect 7255 9029 7337 9115
rect 7423 9029 7516 9115
rect 7076 7666 7516 9029
rect 7076 7286 7106 7666
rect 7486 7286 7516 7666
rect 7076 6091 7516 7286
rect 7076 6005 7169 6091
rect 7255 6005 7337 6091
rect 7423 6005 7516 6091
rect 7076 4579 7516 6005
rect 7076 4493 7169 4579
rect 7255 4493 7337 4579
rect 7423 4493 7516 4579
rect 7076 3666 7516 4493
rect 7076 3286 7106 3666
rect 7486 3286 7516 3666
rect 7076 3067 7516 3286
rect 7076 2981 7169 3067
rect 7255 2981 7337 3067
rect 7423 2981 7516 3067
rect 7076 1555 7516 2981
rect 7076 1469 7169 1555
rect 7255 1469 7337 1555
rect 7423 1469 7516 1555
rect 7076 712 7516 1469
rect 8316 38599 8756 38682
rect 8316 38513 8409 38599
rect 8495 38513 8577 38599
rect 8663 38513 8756 38599
rect 8316 37087 8756 38513
rect 8316 37001 8409 37087
rect 8495 37001 8577 37087
rect 8663 37001 8756 37087
rect 8316 36906 8756 37001
rect 8316 36526 8346 36906
rect 8726 36526 8756 36906
rect 8316 35575 8756 36526
rect 8316 35489 8409 35575
rect 8495 35489 8577 35575
rect 8663 35489 8756 35575
rect 8316 34063 8756 35489
rect 8316 33977 8409 34063
rect 8495 33977 8577 34063
rect 8663 33977 8756 34063
rect 8316 32906 8756 33977
rect 8316 32526 8346 32906
rect 8726 32526 8756 32906
rect 8316 32465 8409 32526
rect 8495 32465 8577 32526
rect 8663 32465 8756 32526
rect 8316 31039 8756 32465
rect 8316 30953 8409 31039
rect 8495 30953 8577 31039
rect 8663 30953 8756 31039
rect 8316 29527 8756 30953
rect 8316 29441 8409 29527
rect 8495 29441 8577 29527
rect 8663 29441 8756 29527
rect 8316 28906 8756 29441
rect 8316 28526 8346 28906
rect 8726 28526 8756 28906
rect 8316 28015 8756 28526
rect 8316 27929 8409 28015
rect 8495 27929 8577 28015
rect 8663 27929 8756 28015
rect 8316 26503 8756 27929
rect 8316 26417 8409 26503
rect 8495 26417 8577 26503
rect 8663 26417 8756 26503
rect 8316 24991 8756 26417
rect 8316 24906 8409 24991
rect 8495 24906 8577 24991
rect 8663 24906 8756 24991
rect 8316 24526 8346 24906
rect 8726 24526 8756 24906
rect 8316 23479 8756 24526
rect 8316 23393 8409 23479
rect 8495 23393 8577 23479
rect 8663 23393 8756 23479
rect 8316 21967 8756 23393
rect 8316 21881 8409 21967
rect 8495 21881 8577 21967
rect 8663 21881 8756 21967
rect 8316 20906 8756 21881
rect 8316 20526 8346 20906
rect 8726 20526 8756 20906
rect 8316 20455 8756 20526
rect 8316 20369 8409 20455
rect 8495 20369 8577 20455
rect 8663 20369 8756 20455
rect 8316 18943 8756 20369
rect 8316 18857 8409 18943
rect 8495 18857 8577 18943
rect 8663 18857 8756 18943
rect 8316 17431 8756 18857
rect 8316 17345 8409 17431
rect 8495 17345 8577 17431
rect 8663 17345 8756 17431
rect 8316 16906 8756 17345
rect 8316 16526 8346 16906
rect 8726 16526 8756 16906
rect 8316 15919 8756 16526
rect 8316 15833 8409 15919
rect 8495 15833 8577 15919
rect 8663 15833 8756 15919
rect 8316 14407 8756 15833
rect 8316 14321 8409 14407
rect 8495 14321 8577 14407
rect 8663 14321 8756 14407
rect 8316 12906 8756 14321
rect 8316 12526 8346 12906
rect 8726 12526 8756 12906
rect 8316 11383 8756 12526
rect 8316 11297 8409 11383
rect 8495 11297 8577 11383
rect 8663 11297 8756 11383
rect 8316 9871 8756 11297
rect 8316 9785 8409 9871
rect 8495 9785 8577 9871
rect 8663 9785 8756 9871
rect 8316 8906 8756 9785
rect 8316 8526 8346 8906
rect 8726 8526 8756 8906
rect 8316 8359 8756 8526
rect 8316 8273 8409 8359
rect 8495 8273 8577 8359
rect 8663 8273 8756 8359
rect 8316 6847 8756 8273
rect 8316 6761 8409 6847
rect 8495 6761 8577 6847
rect 8663 6761 8756 6847
rect 8316 5335 8756 6761
rect 8316 5249 8409 5335
rect 8495 5249 8577 5335
rect 8663 5249 8756 5335
rect 8316 4906 8756 5249
rect 8316 4526 8346 4906
rect 8726 4526 8756 4906
rect 8316 3823 8756 4526
rect 8316 3737 8409 3823
rect 8495 3737 8577 3823
rect 8663 3737 8756 3823
rect 8316 2311 8756 3737
rect 8316 2225 8409 2311
rect 8495 2225 8577 2311
rect 8663 2225 8756 2311
rect 8316 799 8756 2225
rect 8316 713 8409 799
rect 8495 713 8577 799
rect 8663 713 8756 799
rect 8316 630 8756 713
rect 11076 37843 11516 38600
rect 11076 37757 11169 37843
rect 11255 37757 11337 37843
rect 11423 37757 11516 37843
rect 11076 36331 11516 37757
rect 11076 36245 11169 36331
rect 11255 36245 11337 36331
rect 11423 36245 11516 36331
rect 11076 35666 11516 36245
rect 11076 35286 11106 35666
rect 11486 35286 11516 35666
rect 11076 34819 11516 35286
rect 11076 34733 11169 34819
rect 11255 34733 11337 34819
rect 11423 34733 11516 34819
rect 11076 33307 11516 34733
rect 11076 33221 11169 33307
rect 11255 33221 11337 33307
rect 11423 33221 11516 33307
rect 11076 31795 11516 33221
rect 11076 31709 11169 31795
rect 11255 31709 11337 31795
rect 11423 31709 11516 31795
rect 11076 31666 11516 31709
rect 11076 31286 11106 31666
rect 11486 31286 11516 31666
rect 11076 30283 11516 31286
rect 11076 30197 11169 30283
rect 11255 30197 11337 30283
rect 11423 30197 11516 30283
rect 11076 28771 11516 30197
rect 11076 28685 11169 28771
rect 11255 28685 11337 28771
rect 11423 28685 11516 28771
rect 11076 27666 11516 28685
rect 11076 27286 11106 27666
rect 11486 27286 11516 27666
rect 11076 27259 11516 27286
rect 11076 27173 11169 27259
rect 11255 27173 11337 27259
rect 11423 27173 11516 27259
rect 11076 25747 11516 27173
rect 11076 25661 11169 25747
rect 11255 25661 11337 25747
rect 11423 25661 11516 25747
rect 11076 24235 11516 25661
rect 11076 24149 11169 24235
rect 11255 24149 11337 24235
rect 11423 24149 11516 24235
rect 11076 23666 11516 24149
rect 11076 23286 11106 23666
rect 11486 23286 11516 23666
rect 11076 22723 11516 23286
rect 11076 22637 11169 22723
rect 11255 22637 11337 22723
rect 11423 22637 11516 22723
rect 11076 21211 11516 22637
rect 11076 21125 11169 21211
rect 11255 21125 11337 21211
rect 11423 21125 11516 21211
rect 11076 19699 11516 21125
rect 11076 19666 11169 19699
rect 11255 19666 11337 19699
rect 11423 19666 11516 19699
rect 11076 19286 11106 19666
rect 11486 19286 11516 19666
rect 11076 18187 11516 19286
rect 11076 18101 11169 18187
rect 11255 18101 11337 18187
rect 11423 18101 11516 18187
rect 11076 16675 11516 18101
rect 11076 16589 11169 16675
rect 11255 16589 11337 16675
rect 11423 16589 11516 16675
rect 11076 15666 11516 16589
rect 11076 15286 11106 15666
rect 11486 15286 11516 15666
rect 11076 15163 11516 15286
rect 11076 15077 11169 15163
rect 11255 15077 11337 15163
rect 11423 15077 11516 15163
rect 11076 13651 11516 15077
rect 11076 13565 11169 13651
rect 11255 13565 11337 13651
rect 11423 13565 11516 13651
rect 11076 12139 11516 13565
rect 11076 12053 11169 12139
rect 11255 12053 11337 12139
rect 11423 12053 11516 12139
rect 11076 11666 11516 12053
rect 11076 11286 11106 11666
rect 11486 11286 11516 11666
rect 11076 10627 11516 11286
rect 11076 10541 11169 10627
rect 11255 10541 11337 10627
rect 11423 10541 11516 10627
rect 11076 9115 11516 10541
rect 11076 9029 11169 9115
rect 11255 9029 11337 9115
rect 11423 9029 11516 9115
rect 11076 7666 11516 9029
rect 11076 7286 11106 7666
rect 11486 7286 11516 7666
rect 11076 6091 11516 7286
rect 11076 6005 11169 6091
rect 11255 6005 11337 6091
rect 11423 6005 11516 6091
rect 11076 4579 11516 6005
rect 11076 4493 11169 4579
rect 11255 4493 11337 4579
rect 11423 4493 11516 4579
rect 11076 3666 11516 4493
rect 11076 3286 11106 3666
rect 11486 3286 11516 3666
rect 11076 3067 11516 3286
rect 11076 2981 11169 3067
rect 11255 2981 11337 3067
rect 11423 2981 11516 3067
rect 11076 1555 11516 2981
rect 11076 1469 11169 1555
rect 11255 1469 11337 1555
rect 11423 1469 11516 1555
rect 11076 712 11516 1469
rect 12316 38599 12756 38682
rect 12316 38513 12409 38599
rect 12495 38513 12577 38599
rect 12663 38513 12756 38599
rect 12316 37087 12756 38513
rect 12316 37001 12409 37087
rect 12495 37001 12577 37087
rect 12663 37001 12756 37087
rect 12316 36906 12756 37001
rect 12316 36526 12346 36906
rect 12726 36526 12756 36906
rect 12316 35575 12756 36526
rect 12316 35489 12409 35575
rect 12495 35489 12577 35575
rect 12663 35489 12756 35575
rect 12316 34063 12756 35489
rect 12316 33977 12409 34063
rect 12495 33977 12577 34063
rect 12663 33977 12756 34063
rect 12316 32906 12756 33977
rect 12316 32526 12346 32906
rect 12726 32526 12756 32906
rect 12316 32465 12409 32526
rect 12495 32465 12577 32526
rect 12663 32465 12756 32526
rect 12316 31039 12756 32465
rect 12316 30953 12409 31039
rect 12495 30953 12577 31039
rect 12663 30953 12756 31039
rect 12316 29527 12756 30953
rect 12316 29441 12409 29527
rect 12495 29441 12577 29527
rect 12663 29441 12756 29527
rect 12316 28906 12756 29441
rect 12316 28526 12346 28906
rect 12726 28526 12756 28906
rect 12316 28015 12756 28526
rect 12316 27929 12409 28015
rect 12495 27929 12577 28015
rect 12663 27929 12756 28015
rect 12316 26503 12756 27929
rect 12316 26417 12409 26503
rect 12495 26417 12577 26503
rect 12663 26417 12756 26503
rect 12316 24991 12756 26417
rect 12316 24906 12409 24991
rect 12495 24906 12577 24991
rect 12663 24906 12756 24991
rect 12316 24526 12346 24906
rect 12726 24526 12756 24906
rect 12316 23479 12756 24526
rect 12316 23393 12409 23479
rect 12495 23393 12577 23479
rect 12663 23393 12756 23479
rect 12316 21967 12756 23393
rect 12316 21881 12409 21967
rect 12495 21881 12577 21967
rect 12663 21881 12756 21967
rect 12316 20906 12756 21881
rect 12316 20526 12346 20906
rect 12726 20526 12756 20906
rect 12316 20455 12756 20526
rect 12316 20369 12409 20455
rect 12495 20369 12577 20455
rect 12663 20369 12756 20455
rect 12316 18943 12756 20369
rect 12316 18857 12409 18943
rect 12495 18857 12577 18943
rect 12663 18857 12756 18943
rect 12316 17431 12756 18857
rect 12316 17345 12409 17431
rect 12495 17345 12577 17431
rect 12663 17345 12756 17431
rect 12316 16906 12756 17345
rect 12316 16526 12346 16906
rect 12726 16526 12756 16906
rect 12316 15919 12756 16526
rect 12316 15833 12409 15919
rect 12495 15833 12577 15919
rect 12663 15833 12756 15919
rect 12316 14407 12756 15833
rect 12316 14321 12409 14407
rect 12495 14321 12577 14407
rect 12663 14321 12756 14407
rect 12316 12906 12756 14321
rect 12316 12526 12346 12906
rect 12726 12526 12756 12906
rect 12316 11383 12756 12526
rect 12316 11297 12409 11383
rect 12495 11297 12577 11383
rect 12663 11297 12756 11383
rect 12316 9871 12756 11297
rect 12316 9785 12409 9871
rect 12495 9785 12577 9871
rect 12663 9785 12756 9871
rect 12316 8906 12756 9785
rect 12316 8526 12346 8906
rect 12726 8526 12756 8906
rect 12316 8359 12756 8526
rect 12316 8273 12409 8359
rect 12495 8273 12577 8359
rect 12663 8273 12756 8359
rect 12316 6847 12756 8273
rect 12316 6761 12409 6847
rect 12495 6761 12577 6847
rect 12663 6761 12756 6847
rect 12316 5335 12756 6761
rect 12316 5249 12409 5335
rect 12495 5249 12577 5335
rect 12663 5249 12756 5335
rect 12316 4906 12756 5249
rect 12316 4526 12346 4906
rect 12726 4526 12756 4906
rect 12316 3823 12756 4526
rect 12316 3737 12409 3823
rect 12495 3737 12577 3823
rect 12663 3737 12756 3823
rect 12316 2311 12756 3737
rect 12316 2225 12409 2311
rect 12495 2225 12577 2311
rect 12663 2225 12756 2311
rect 12316 799 12756 2225
rect 12316 713 12409 799
rect 12495 713 12577 799
rect 12663 713 12756 799
rect 12316 630 12756 713
rect 15076 37843 15516 38600
rect 15076 37757 15169 37843
rect 15255 37757 15337 37843
rect 15423 37757 15516 37843
rect 15076 36331 15516 37757
rect 15076 36245 15169 36331
rect 15255 36245 15337 36331
rect 15423 36245 15516 36331
rect 15076 35666 15516 36245
rect 15076 35286 15106 35666
rect 15486 35286 15516 35666
rect 15076 34819 15516 35286
rect 15076 34733 15169 34819
rect 15255 34733 15337 34819
rect 15423 34733 15516 34819
rect 15076 33307 15516 34733
rect 15076 33221 15169 33307
rect 15255 33221 15337 33307
rect 15423 33221 15516 33307
rect 15076 31795 15516 33221
rect 15076 31709 15169 31795
rect 15255 31709 15337 31795
rect 15423 31709 15516 31795
rect 15076 31666 15516 31709
rect 15076 31286 15106 31666
rect 15486 31286 15516 31666
rect 15076 30283 15516 31286
rect 15076 30197 15169 30283
rect 15255 30197 15337 30283
rect 15423 30197 15516 30283
rect 15076 28771 15516 30197
rect 15076 28685 15169 28771
rect 15255 28685 15337 28771
rect 15423 28685 15516 28771
rect 15076 27666 15516 28685
rect 15076 27286 15106 27666
rect 15486 27286 15516 27666
rect 15076 27259 15516 27286
rect 15076 27173 15169 27259
rect 15255 27173 15337 27259
rect 15423 27173 15516 27259
rect 15076 25747 15516 27173
rect 15076 25661 15169 25747
rect 15255 25661 15337 25747
rect 15423 25661 15516 25747
rect 15076 24235 15516 25661
rect 15076 24149 15169 24235
rect 15255 24149 15337 24235
rect 15423 24149 15516 24235
rect 15076 23666 15516 24149
rect 15076 23286 15106 23666
rect 15486 23286 15516 23666
rect 15076 22723 15516 23286
rect 15076 22637 15169 22723
rect 15255 22637 15337 22723
rect 15423 22637 15516 22723
rect 15076 21211 15516 22637
rect 15076 21125 15169 21211
rect 15255 21125 15337 21211
rect 15423 21125 15516 21211
rect 15076 19699 15516 21125
rect 15076 19666 15169 19699
rect 15255 19666 15337 19699
rect 15423 19666 15516 19699
rect 15076 19286 15106 19666
rect 15486 19286 15516 19666
rect 15076 18187 15516 19286
rect 15076 18101 15169 18187
rect 15255 18101 15337 18187
rect 15423 18101 15516 18187
rect 15076 16675 15516 18101
rect 15076 16589 15169 16675
rect 15255 16589 15337 16675
rect 15423 16589 15516 16675
rect 15076 15666 15516 16589
rect 15076 15286 15106 15666
rect 15486 15286 15516 15666
rect 15076 15163 15516 15286
rect 15076 15077 15169 15163
rect 15255 15077 15337 15163
rect 15423 15077 15516 15163
rect 15076 13651 15516 15077
rect 15076 13565 15169 13651
rect 15255 13565 15337 13651
rect 15423 13565 15516 13651
rect 15076 12139 15516 13565
rect 15076 12053 15169 12139
rect 15255 12053 15337 12139
rect 15423 12053 15516 12139
rect 15076 11666 15516 12053
rect 15076 11286 15106 11666
rect 15486 11286 15516 11666
rect 15076 10627 15516 11286
rect 15076 10541 15169 10627
rect 15255 10541 15337 10627
rect 15423 10541 15516 10627
rect 15076 9115 15516 10541
rect 15076 9029 15169 9115
rect 15255 9029 15337 9115
rect 15423 9029 15516 9115
rect 15076 7666 15516 9029
rect 15076 7286 15106 7666
rect 15486 7286 15516 7666
rect 15076 6091 15516 7286
rect 15076 6005 15169 6091
rect 15255 6005 15337 6091
rect 15423 6005 15516 6091
rect 15076 4579 15516 6005
rect 15076 4493 15169 4579
rect 15255 4493 15337 4579
rect 15423 4493 15516 4579
rect 15076 3666 15516 4493
rect 15076 3286 15106 3666
rect 15486 3286 15516 3666
rect 15076 3067 15516 3286
rect 15076 2981 15169 3067
rect 15255 2981 15337 3067
rect 15423 2981 15516 3067
rect 15076 1555 15516 2981
rect 15076 1469 15169 1555
rect 15255 1469 15337 1555
rect 15423 1469 15516 1555
rect 15076 712 15516 1469
rect 16316 38599 16756 38682
rect 16316 38513 16409 38599
rect 16495 38513 16577 38599
rect 16663 38513 16756 38599
rect 16316 37087 16756 38513
rect 16316 37001 16409 37087
rect 16495 37001 16577 37087
rect 16663 37001 16756 37087
rect 16316 36906 16756 37001
rect 16316 36526 16346 36906
rect 16726 36526 16756 36906
rect 16316 35575 16756 36526
rect 16316 35489 16409 35575
rect 16495 35489 16577 35575
rect 16663 35489 16756 35575
rect 16316 34063 16756 35489
rect 16316 33977 16409 34063
rect 16495 33977 16577 34063
rect 16663 33977 16756 34063
rect 16316 32906 16756 33977
rect 16316 32526 16346 32906
rect 16726 32526 16756 32906
rect 16316 32465 16409 32526
rect 16495 32465 16577 32526
rect 16663 32465 16756 32526
rect 16316 31039 16756 32465
rect 16316 30953 16409 31039
rect 16495 30953 16577 31039
rect 16663 30953 16756 31039
rect 16316 29527 16756 30953
rect 16316 29441 16409 29527
rect 16495 29441 16577 29527
rect 16663 29441 16756 29527
rect 16316 28906 16756 29441
rect 16316 28526 16346 28906
rect 16726 28526 16756 28906
rect 16316 28015 16756 28526
rect 16316 27929 16409 28015
rect 16495 27929 16577 28015
rect 16663 27929 16756 28015
rect 16316 26503 16756 27929
rect 16316 26417 16409 26503
rect 16495 26417 16577 26503
rect 16663 26417 16756 26503
rect 16316 24991 16756 26417
rect 16316 24906 16409 24991
rect 16495 24906 16577 24991
rect 16663 24906 16756 24991
rect 16316 24526 16346 24906
rect 16726 24526 16756 24906
rect 16316 23479 16756 24526
rect 16316 23393 16409 23479
rect 16495 23393 16577 23479
rect 16663 23393 16756 23479
rect 16316 21967 16756 23393
rect 16316 21881 16409 21967
rect 16495 21881 16577 21967
rect 16663 21881 16756 21967
rect 16316 20906 16756 21881
rect 16316 20526 16346 20906
rect 16726 20526 16756 20906
rect 16316 20455 16756 20526
rect 16316 20369 16409 20455
rect 16495 20369 16577 20455
rect 16663 20369 16756 20455
rect 16316 18943 16756 20369
rect 16316 18857 16409 18943
rect 16495 18857 16577 18943
rect 16663 18857 16756 18943
rect 16316 17431 16756 18857
rect 16316 17345 16409 17431
rect 16495 17345 16577 17431
rect 16663 17345 16756 17431
rect 16316 16906 16756 17345
rect 16316 16526 16346 16906
rect 16726 16526 16756 16906
rect 16316 15919 16756 16526
rect 16316 15833 16409 15919
rect 16495 15833 16577 15919
rect 16663 15833 16756 15919
rect 16316 14407 16756 15833
rect 16316 14321 16409 14407
rect 16495 14321 16577 14407
rect 16663 14321 16756 14407
rect 16316 12906 16756 14321
rect 16316 12526 16346 12906
rect 16726 12526 16756 12906
rect 16316 11383 16756 12526
rect 16316 11297 16409 11383
rect 16495 11297 16577 11383
rect 16663 11297 16756 11383
rect 16316 9871 16756 11297
rect 16316 9785 16409 9871
rect 16495 9785 16577 9871
rect 16663 9785 16756 9871
rect 16316 8906 16756 9785
rect 16316 8526 16346 8906
rect 16726 8526 16756 8906
rect 16316 8359 16756 8526
rect 16316 8273 16409 8359
rect 16495 8273 16577 8359
rect 16663 8273 16756 8359
rect 16316 6847 16756 8273
rect 16316 6761 16409 6847
rect 16495 6761 16577 6847
rect 16663 6761 16756 6847
rect 16316 5335 16756 6761
rect 16316 5249 16409 5335
rect 16495 5249 16577 5335
rect 16663 5249 16756 5335
rect 16316 4906 16756 5249
rect 16316 4526 16346 4906
rect 16726 4526 16756 4906
rect 16316 3823 16756 4526
rect 16316 3737 16409 3823
rect 16495 3737 16577 3823
rect 16663 3737 16756 3823
rect 16316 2311 16756 3737
rect 16316 2225 16409 2311
rect 16495 2225 16577 2311
rect 16663 2225 16756 2311
rect 16316 799 16756 2225
rect 16316 713 16409 799
rect 16495 713 16577 799
rect 16663 713 16756 799
rect 16316 630 16756 713
rect 19076 37843 19516 38600
rect 19076 37757 19169 37843
rect 19255 37757 19337 37843
rect 19423 37757 19516 37843
rect 19076 36331 19516 37757
rect 19076 36245 19169 36331
rect 19255 36245 19337 36331
rect 19423 36245 19516 36331
rect 19076 35666 19516 36245
rect 19076 35286 19106 35666
rect 19486 35286 19516 35666
rect 19076 34819 19516 35286
rect 19076 34733 19169 34819
rect 19255 34733 19337 34819
rect 19423 34733 19516 34819
rect 19076 33307 19516 34733
rect 19076 33221 19169 33307
rect 19255 33221 19337 33307
rect 19423 33221 19516 33307
rect 19076 31795 19516 33221
rect 19076 31709 19169 31795
rect 19255 31709 19337 31795
rect 19423 31709 19516 31795
rect 19076 31666 19516 31709
rect 19076 31286 19106 31666
rect 19486 31286 19516 31666
rect 19076 30283 19516 31286
rect 19076 30197 19169 30283
rect 19255 30197 19337 30283
rect 19423 30197 19516 30283
rect 19076 28771 19516 30197
rect 19076 28685 19169 28771
rect 19255 28685 19337 28771
rect 19423 28685 19516 28771
rect 19076 27666 19516 28685
rect 19076 27286 19106 27666
rect 19486 27286 19516 27666
rect 19076 27259 19516 27286
rect 19076 27173 19169 27259
rect 19255 27173 19337 27259
rect 19423 27173 19516 27259
rect 19076 25747 19516 27173
rect 19076 25661 19169 25747
rect 19255 25661 19337 25747
rect 19423 25661 19516 25747
rect 19076 24235 19516 25661
rect 19076 24149 19169 24235
rect 19255 24149 19337 24235
rect 19423 24149 19516 24235
rect 19076 23666 19516 24149
rect 19076 23286 19106 23666
rect 19486 23286 19516 23666
rect 19076 22723 19516 23286
rect 19076 22637 19169 22723
rect 19255 22637 19337 22723
rect 19423 22637 19516 22723
rect 19076 21211 19516 22637
rect 19076 21125 19169 21211
rect 19255 21125 19337 21211
rect 19423 21125 19516 21211
rect 19076 19699 19516 21125
rect 19076 19666 19169 19699
rect 19255 19666 19337 19699
rect 19423 19666 19516 19699
rect 19076 19286 19106 19666
rect 19486 19286 19516 19666
rect 19076 18187 19516 19286
rect 19076 18101 19169 18187
rect 19255 18101 19337 18187
rect 19423 18101 19516 18187
rect 19076 16675 19516 18101
rect 19076 16589 19169 16675
rect 19255 16589 19337 16675
rect 19423 16589 19516 16675
rect 19076 15666 19516 16589
rect 19076 15286 19106 15666
rect 19486 15286 19516 15666
rect 19076 15163 19516 15286
rect 19076 15077 19169 15163
rect 19255 15077 19337 15163
rect 19423 15077 19516 15163
rect 19076 13651 19516 15077
rect 19076 13565 19169 13651
rect 19255 13565 19337 13651
rect 19423 13565 19516 13651
rect 19076 12139 19516 13565
rect 19076 12053 19169 12139
rect 19255 12053 19337 12139
rect 19423 12053 19516 12139
rect 19076 11666 19516 12053
rect 19076 11286 19106 11666
rect 19486 11286 19516 11666
rect 19076 10627 19516 11286
rect 19076 10541 19169 10627
rect 19255 10541 19337 10627
rect 19423 10541 19516 10627
rect 19076 9115 19516 10541
rect 19076 9029 19169 9115
rect 19255 9029 19337 9115
rect 19423 9029 19516 9115
rect 19076 7666 19516 9029
rect 19076 7286 19106 7666
rect 19486 7286 19516 7666
rect 19076 6091 19516 7286
rect 19076 6005 19169 6091
rect 19255 6005 19337 6091
rect 19423 6005 19516 6091
rect 19076 4579 19516 6005
rect 19076 4493 19169 4579
rect 19255 4493 19337 4579
rect 19423 4493 19516 4579
rect 19076 3666 19516 4493
rect 19076 3286 19106 3666
rect 19486 3286 19516 3666
rect 19076 3067 19516 3286
rect 19076 2981 19169 3067
rect 19255 2981 19337 3067
rect 19423 2981 19516 3067
rect 19076 1555 19516 2981
rect 19076 1469 19169 1555
rect 19255 1469 19337 1555
rect 19423 1469 19516 1555
rect 19076 712 19516 1469
rect 20316 38599 20756 38682
rect 20316 38513 20409 38599
rect 20495 38513 20577 38599
rect 20663 38513 20756 38599
rect 20316 37087 20756 38513
rect 20316 37001 20409 37087
rect 20495 37001 20577 37087
rect 20663 37001 20756 37087
rect 20316 36906 20756 37001
rect 20316 36526 20346 36906
rect 20726 36526 20756 36906
rect 20316 35575 20756 36526
rect 20316 35489 20409 35575
rect 20495 35489 20577 35575
rect 20663 35489 20756 35575
rect 20316 34063 20756 35489
rect 20316 33977 20409 34063
rect 20495 33977 20577 34063
rect 20663 33977 20756 34063
rect 20316 32906 20756 33977
rect 20316 32526 20346 32906
rect 20726 32526 20756 32906
rect 20316 32465 20409 32526
rect 20495 32465 20577 32526
rect 20663 32465 20756 32526
rect 20316 31039 20756 32465
rect 20316 30953 20409 31039
rect 20495 30953 20577 31039
rect 20663 30953 20756 31039
rect 20316 29527 20756 30953
rect 20316 29441 20409 29527
rect 20495 29441 20577 29527
rect 20663 29441 20756 29527
rect 20316 28906 20756 29441
rect 20316 28526 20346 28906
rect 20726 28526 20756 28906
rect 20316 28015 20756 28526
rect 20316 27929 20409 28015
rect 20495 27929 20577 28015
rect 20663 27929 20756 28015
rect 20316 26503 20756 27929
rect 20316 26417 20409 26503
rect 20495 26417 20577 26503
rect 20663 26417 20756 26503
rect 20316 24991 20756 26417
rect 20316 24906 20409 24991
rect 20495 24906 20577 24991
rect 20663 24906 20756 24991
rect 20316 24526 20346 24906
rect 20726 24526 20756 24906
rect 20316 23479 20756 24526
rect 20316 23393 20409 23479
rect 20495 23393 20577 23479
rect 20663 23393 20756 23479
rect 20316 21967 20756 23393
rect 20316 21881 20409 21967
rect 20495 21881 20577 21967
rect 20663 21881 20756 21967
rect 20316 20906 20756 21881
rect 20316 20526 20346 20906
rect 20726 20526 20756 20906
rect 20316 20455 20756 20526
rect 20316 20369 20409 20455
rect 20495 20369 20577 20455
rect 20663 20369 20756 20455
rect 20316 18943 20756 20369
rect 20316 18857 20409 18943
rect 20495 18857 20577 18943
rect 20663 18857 20756 18943
rect 20316 17431 20756 18857
rect 20316 17345 20409 17431
rect 20495 17345 20577 17431
rect 20663 17345 20756 17431
rect 20316 16906 20756 17345
rect 20316 16526 20346 16906
rect 20726 16526 20756 16906
rect 20316 15919 20756 16526
rect 20316 15833 20409 15919
rect 20495 15833 20577 15919
rect 20663 15833 20756 15919
rect 20316 14407 20756 15833
rect 20316 14321 20409 14407
rect 20495 14321 20577 14407
rect 20663 14321 20756 14407
rect 20316 12906 20756 14321
rect 20316 12526 20346 12906
rect 20726 12526 20756 12906
rect 20316 11383 20756 12526
rect 20316 11297 20409 11383
rect 20495 11297 20577 11383
rect 20663 11297 20756 11383
rect 20316 9871 20756 11297
rect 20316 9785 20409 9871
rect 20495 9785 20577 9871
rect 20663 9785 20756 9871
rect 20316 8906 20756 9785
rect 20316 8526 20346 8906
rect 20726 8526 20756 8906
rect 20316 8359 20756 8526
rect 20316 8273 20409 8359
rect 20495 8273 20577 8359
rect 20663 8273 20756 8359
rect 20316 6847 20756 8273
rect 20316 6761 20409 6847
rect 20495 6761 20577 6847
rect 20663 6761 20756 6847
rect 20316 5335 20756 6761
rect 20316 5249 20409 5335
rect 20495 5249 20577 5335
rect 20663 5249 20756 5335
rect 20316 4906 20756 5249
rect 20316 4526 20346 4906
rect 20726 4526 20756 4906
rect 20316 3823 20756 4526
rect 20316 3737 20409 3823
rect 20495 3737 20577 3823
rect 20663 3737 20756 3823
rect 20316 2311 20756 3737
rect 20316 2225 20409 2311
rect 20495 2225 20577 2311
rect 20663 2225 20756 2311
rect 20316 799 20756 2225
rect 20316 713 20409 799
rect 20495 713 20577 799
rect 20663 713 20756 799
rect 20316 630 20756 713
rect 23076 37843 23516 38600
rect 23076 37757 23169 37843
rect 23255 37757 23337 37843
rect 23423 37757 23516 37843
rect 23076 36331 23516 37757
rect 23076 36245 23169 36331
rect 23255 36245 23337 36331
rect 23423 36245 23516 36331
rect 23076 35666 23516 36245
rect 23076 35286 23106 35666
rect 23486 35286 23516 35666
rect 23076 34819 23516 35286
rect 23076 34733 23169 34819
rect 23255 34733 23337 34819
rect 23423 34733 23516 34819
rect 23076 33307 23516 34733
rect 23076 33221 23169 33307
rect 23255 33221 23337 33307
rect 23423 33221 23516 33307
rect 23076 31795 23516 33221
rect 23076 31709 23169 31795
rect 23255 31709 23337 31795
rect 23423 31709 23516 31795
rect 23076 31666 23516 31709
rect 23076 31286 23106 31666
rect 23486 31286 23516 31666
rect 23076 30283 23516 31286
rect 23076 30197 23169 30283
rect 23255 30197 23337 30283
rect 23423 30197 23516 30283
rect 23076 28771 23516 30197
rect 23076 28685 23169 28771
rect 23255 28685 23337 28771
rect 23423 28685 23516 28771
rect 23076 27666 23516 28685
rect 23076 27286 23106 27666
rect 23486 27286 23516 27666
rect 23076 27259 23516 27286
rect 23076 27173 23169 27259
rect 23255 27173 23337 27259
rect 23423 27173 23516 27259
rect 23076 25747 23516 27173
rect 23076 25661 23169 25747
rect 23255 25661 23337 25747
rect 23423 25661 23516 25747
rect 23076 24235 23516 25661
rect 23076 24149 23169 24235
rect 23255 24149 23337 24235
rect 23423 24149 23516 24235
rect 23076 23666 23516 24149
rect 23076 23286 23106 23666
rect 23486 23286 23516 23666
rect 23076 22723 23516 23286
rect 23076 22637 23169 22723
rect 23255 22637 23337 22723
rect 23423 22637 23516 22723
rect 23076 21211 23516 22637
rect 23076 21125 23169 21211
rect 23255 21125 23337 21211
rect 23423 21125 23516 21211
rect 23076 19699 23516 21125
rect 23076 19666 23169 19699
rect 23255 19666 23337 19699
rect 23423 19666 23516 19699
rect 23076 19286 23106 19666
rect 23486 19286 23516 19666
rect 23076 18187 23516 19286
rect 23076 18101 23169 18187
rect 23255 18101 23337 18187
rect 23423 18101 23516 18187
rect 23076 16675 23516 18101
rect 23076 16589 23169 16675
rect 23255 16589 23337 16675
rect 23423 16589 23516 16675
rect 23076 15666 23516 16589
rect 23076 15286 23106 15666
rect 23486 15286 23516 15666
rect 23076 15163 23516 15286
rect 23076 15077 23169 15163
rect 23255 15077 23337 15163
rect 23423 15077 23516 15163
rect 23076 13651 23516 15077
rect 23076 13565 23169 13651
rect 23255 13565 23337 13651
rect 23423 13565 23516 13651
rect 23076 12139 23516 13565
rect 23076 12053 23169 12139
rect 23255 12053 23337 12139
rect 23423 12053 23516 12139
rect 23076 11666 23516 12053
rect 23076 11286 23106 11666
rect 23486 11286 23516 11666
rect 23076 10627 23516 11286
rect 23076 10541 23169 10627
rect 23255 10541 23337 10627
rect 23423 10541 23516 10627
rect 23076 9115 23516 10541
rect 23076 9029 23169 9115
rect 23255 9029 23337 9115
rect 23423 9029 23516 9115
rect 23076 7666 23516 9029
rect 23076 7286 23106 7666
rect 23486 7286 23516 7666
rect 23076 6091 23516 7286
rect 23076 6005 23169 6091
rect 23255 6005 23337 6091
rect 23423 6005 23516 6091
rect 23076 4579 23516 6005
rect 23076 4493 23169 4579
rect 23255 4493 23337 4579
rect 23423 4493 23516 4579
rect 23076 3666 23516 4493
rect 23076 3286 23106 3666
rect 23486 3286 23516 3666
rect 23076 3067 23516 3286
rect 23076 2981 23169 3067
rect 23255 2981 23337 3067
rect 23423 2981 23516 3067
rect 23076 1555 23516 2981
rect 23076 1469 23169 1555
rect 23255 1469 23337 1555
rect 23423 1469 23516 1555
rect 23076 712 23516 1469
rect 24316 38599 24756 38682
rect 24316 38513 24409 38599
rect 24495 38513 24577 38599
rect 24663 38513 24756 38599
rect 24316 37087 24756 38513
rect 24316 37001 24409 37087
rect 24495 37001 24577 37087
rect 24663 37001 24756 37087
rect 24316 36906 24756 37001
rect 24316 36526 24346 36906
rect 24726 36526 24756 36906
rect 24316 35575 24756 36526
rect 24316 35489 24409 35575
rect 24495 35489 24577 35575
rect 24663 35489 24756 35575
rect 24316 34063 24756 35489
rect 24316 33977 24409 34063
rect 24495 33977 24577 34063
rect 24663 33977 24756 34063
rect 24316 32906 24756 33977
rect 24316 32526 24346 32906
rect 24726 32526 24756 32906
rect 24316 32465 24409 32526
rect 24495 32465 24577 32526
rect 24663 32465 24756 32526
rect 24316 31039 24756 32465
rect 24316 30953 24409 31039
rect 24495 30953 24577 31039
rect 24663 30953 24756 31039
rect 24316 29527 24756 30953
rect 24316 29441 24409 29527
rect 24495 29441 24577 29527
rect 24663 29441 24756 29527
rect 24316 28906 24756 29441
rect 24316 28526 24346 28906
rect 24726 28526 24756 28906
rect 24316 28015 24756 28526
rect 24316 27929 24409 28015
rect 24495 27929 24577 28015
rect 24663 27929 24756 28015
rect 24316 26503 24756 27929
rect 24316 26417 24409 26503
rect 24495 26417 24577 26503
rect 24663 26417 24756 26503
rect 24316 24991 24756 26417
rect 24316 24906 24409 24991
rect 24495 24906 24577 24991
rect 24663 24906 24756 24991
rect 24316 24526 24346 24906
rect 24726 24526 24756 24906
rect 24316 23479 24756 24526
rect 24316 23393 24409 23479
rect 24495 23393 24577 23479
rect 24663 23393 24756 23479
rect 24316 21967 24756 23393
rect 24316 21881 24409 21967
rect 24495 21881 24577 21967
rect 24663 21881 24756 21967
rect 24316 20906 24756 21881
rect 24316 20526 24346 20906
rect 24726 20526 24756 20906
rect 24316 20455 24756 20526
rect 24316 20369 24409 20455
rect 24495 20369 24577 20455
rect 24663 20369 24756 20455
rect 24316 18943 24756 20369
rect 24316 18857 24409 18943
rect 24495 18857 24577 18943
rect 24663 18857 24756 18943
rect 24316 17431 24756 18857
rect 24316 17345 24409 17431
rect 24495 17345 24577 17431
rect 24663 17345 24756 17431
rect 24316 16906 24756 17345
rect 24316 16526 24346 16906
rect 24726 16526 24756 16906
rect 24316 15919 24756 16526
rect 24316 15833 24409 15919
rect 24495 15833 24577 15919
rect 24663 15833 24756 15919
rect 24316 14407 24756 15833
rect 24316 14321 24409 14407
rect 24495 14321 24577 14407
rect 24663 14321 24756 14407
rect 24316 12906 24756 14321
rect 24316 12526 24346 12906
rect 24726 12526 24756 12906
rect 24316 11383 24756 12526
rect 24316 11297 24409 11383
rect 24495 11297 24577 11383
rect 24663 11297 24756 11383
rect 24316 9871 24756 11297
rect 24316 9785 24409 9871
rect 24495 9785 24577 9871
rect 24663 9785 24756 9871
rect 24316 8906 24756 9785
rect 24316 8526 24346 8906
rect 24726 8526 24756 8906
rect 24316 8359 24756 8526
rect 24316 8273 24409 8359
rect 24495 8273 24577 8359
rect 24663 8273 24756 8359
rect 24316 6847 24756 8273
rect 24316 6761 24409 6847
rect 24495 6761 24577 6847
rect 24663 6761 24756 6847
rect 24316 5335 24756 6761
rect 24316 5249 24409 5335
rect 24495 5249 24577 5335
rect 24663 5249 24756 5335
rect 24316 4906 24756 5249
rect 24316 4526 24346 4906
rect 24726 4526 24756 4906
rect 24316 3823 24756 4526
rect 24316 3737 24409 3823
rect 24495 3737 24577 3823
rect 24663 3737 24756 3823
rect 24316 2311 24756 3737
rect 24316 2225 24409 2311
rect 24495 2225 24577 2311
rect 24663 2225 24756 2311
rect 24316 799 24756 2225
rect 24316 713 24409 799
rect 24495 713 24577 799
rect 24663 713 24756 799
rect 24316 630 24756 713
rect 27076 37843 27516 38600
rect 27076 37757 27169 37843
rect 27255 37757 27337 37843
rect 27423 37757 27516 37843
rect 27076 36331 27516 37757
rect 27076 36245 27169 36331
rect 27255 36245 27337 36331
rect 27423 36245 27516 36331
rect 27076 35666 27516 36245
rect 27076 35286 27106 35666
rect 27486 35286 27516 35666
rect 27076 34819 27516 35286
rect 27076 34733 27169 34819
rect 27255 34733 27337 34819
rect 27423 34733 27516 34819
rect 27076 33307 27516 34733
rect 27076 33221 27169 33307
rect 27255 33221 27337 33307
rect 27423 33221 27516 33307
rect 27076 31795 27516 33221
rect 27076 31709 27169 31795
rect 27255 31709 27337 31795
rect 27423 31709 27516 31795
rect 27076 31666 27516 31709
rect 27076 31286 27106 31666
rect 27486 31286 27516 31666
rect 27076 30283 27516 31286
rect 27076 30197 27169 30283
rect 27255 30197 27337 30283
rect 27423 30197 27516 30283
rect 27076 28771 27516 30197
rect 27076 28685 27169 28771
rect 27255 28685 27337 28771
rect 27423 28685 27516 28771
rect 27076 27666 27516 28685
rect 27076 27286 27106 27666
rect 27486 27286 27516 27666
rect 27076 27259 27516 27286
rect 27076 27173 27169 27259
rect 27255 27173 27337 27259
rect 27423 27173 27516 27259
rect 27076 25747 27516 27173
rect 27076 25661 27169 25747
rect 27255 25661 27337 25747
rect 27423 25661 27516 25747
rect 27076 24235 27516 25661
rect 27076 24149 27169 24235
rect 27255 24149 27337 24235
rect 27423 24149 27516 24235
rect 27076 23666 27516 24149
rect 27076 23286 27106 23666
rect 27486 23286 27516 23666
rect 27076 22723 27516 23286
rect 27076 22637 27169 22723
rect 27255 22637 27337 22723
rect 27423 22637 27516 22723
rect 27076 21211 27516 22637
rect 27076 21125 27169 21211
rect 27255 21125 27337 21211
rect 27423 21125 27516 21211
rect 27076 19699 27516 21125
rect 27076 19666 27169 19699
rect 27255 19666 27337 19699
rect 27423 19666 27516 19699
rect 27076 19286 27106 19666
rect 27486 19286 27516 19666
rect 27076 18187 27516 19286
rect 27076 18101 27169 18187
rect 27255 18101 27337 18187
rect 27423 18101 27516 18187
rect 27076 16675 27516 18101
rect 27076 16589 27169 16675
rect 27255 16589 27337 16675
rect 27423 16589 27516 16675
rect 27076 15666 27516 16589
rect 27076 15286 27106 15666
rect 27486 15286 27516 15666
rect 27076 15163 27516 15286
rect 27076 15077 27169 15163
rect 27255 15077 27337 15163
rect 27423 15077 27516 15163
rect 27076 13651 27516 15077
rect 27076 13565 27169 13651
rect 27255 13565 27337 13651
rect 27423 13565 27516 13651
rect 27076 12139 27516 13565
rect 27076 12053 27169 12139
rect 27255 12053 27337 12139
rect 27423 12053 27516 12139
rect 27076 11666 27516 12053
rect 27076 11286 27106 11666
rect 27486 11286 27516 11666
rect 27076 10627 27516 11286
rect 27076 10541 27169 10627
rect 27255 10541 27337 10627
rect 27423 10541 27516 10627
rect 27076 9115 27516 10541
rect 27076 9029 27169 9115
rect 27255 9029 27337 9115
rect 27423 9029 27516 9115
rect 27076 7666 27516 9029
rect 27076 7286 27106 7666
rect 27486 7286 27516 7666
rect 27076 6091 27516 7286
rect 27076 6005 27169 6091
rect 27255 6005 27337 6091
rect 27423 6005 27516 6091
rect 27076 4579 27516 6005
rect 27076 4493 27169 4579
rect 27255 4493 27337 4579
rect 27423 4493 27516 4579
rect 27076 3666 27516 4493
rect 27076 3286 27106 3666
rect 27486 3286 27516 3666
rect 27076 3067 27516 3286
rect 27076 2981 27169 3067
rect 27255 2981 27337 3067
rect 27423 2981 27516 3067
rect 27076 1555 27516 2981
rect 27076 1469 27169 1555
rect 27255 1469 27337 1555
rect 27423 1469 27516 1555
rect 27076 712 27516 1469
rect 28316 38599 28756 38682
rect 28316 38513 28409 38599
rect 28495 38513 28577 38599
rect 28663 38513 28756 38599
rect 28316 37087 28756 38513
rect 28316 37001 28409 37087
rect 28495 37001 28577 37087
rect 28663 37001 28756 37087
rect 28316 36906 28756 37001
rect 28316 36526 28346 36906
rect 28726 36526 28756 36906
rect 28316 35575 28756 36526
rect 28316 35489 28409 35575
rect 28495 35489 28577 35575
rect 28663 35489 28756 35575
rect 28316 34063 28756 35489
rect 28316 33977 28409 34063
rect 28495 33977 28577 34063
rect 28663 33977 28756 34063
rect 28316 32906 28756 33977
rect 28316 32526 28346 32906
rect 28726 32526 28756 32906
rect 28316 32465 28409 32526
rect 28495 32465 28577 32526
rect 28663 32465 28756 32526
rect 28316 31039 28756 32465
rect 28316 30953 28409 31039
rect 28495 30953 28577 31039
rect 28663 30953 28756 31039
rect 28316 29527 28756 30953
rect 28316 29441 28409 29527
rect 28495 29441 28577 29527
rect 28663 29441 28756 29527
rect 28316 28906 28756 29441
rect 28316 28526 28346 28906
rect 28726 28526 28756 28906
rect 28316 28015 28756 28526
rect 28316 27929 28409 28015
rect 28495 27929 28577 28015
rect 28663 27929 28756 28015
rect 28316 26503 28756 27929
rect 28316 26417 28409 26503
rect 28495 26417 28577 26503
rect 28663 26417 28756 26503
rect 28316 24991 28756 26417
rect 28316 24906 28409 24991
rect 28495 24906 28577 24991
rect 28663 24906 28756 24991
rect 28316 24526 28346 24906
rect 28726 24526 28756 24906
rect 28316 23479 28756 24526
rect 28316 23393 28409 23479
rect 28495 23393 28577 23479
rect 28663 23393 28756 23479
rect 28316 21967 28756 23393
rect 28316 21881 28409 21967
rect 28495 21881 28577 21967
rect 28663 21881 28756 21967
rect 28316 20906 28756 21881
rect 28316 20526 28346 20906
rect 28726 20526 28756 20906
rect 28316 20455 28756 20526
rect 28316 20369 28409 20455
rect 28495 20369 28577 20455
rect 28663 20369 28756 20455
rect 28316 18943 28756 20369
rect 28316 18857 28409 18943
rect 28495 18857 28577 18943
rect 28663 18857 28756 18943
rect 28316 17431 28756 18857
rect 28316 17345 28409 17431
rect 28495 17345 28577 17431
rect 28663 17345 28756 17431
rect 28316 16906 28756 17345
rect 28316 16526 28346 16906
rect 28726 16526 28756 16906
rect 28316 15919 28756 16526
rect 28316 15833 28409 15919
rect 28495 15833 28577 15919
rect 28663 15833 28756 15919
rect 28316 14407 28756 15833
rect 28316 14321 28409 14407
rect 28495 14321 28577 14407
rect 28663 14321 28756 14407
rect 28316 12906 28756 14321
rect 28316 12526 28346 12906
rect 28726 12526 28756 12906
rect 28316 11383 28756 12526
rect 28316 11297 28409 11383
rect 28495 11297 28577 11383
rect 28663 11297 28756 11383
rect 28316 9871 28756 11297
rect 28316 9785 28409 9871
rect 28495 9785 28577 9871
rect 28663 9785 28756 9871
rect 28316 8906 28756 9785
rect 28316 8526 28346 8906
rect 28726 8526 28756 8906
rect 28316 8359 28756 8526
rect 28316 8273 28409 8359
rect 28495 8273 28577 8359
rect 28663 8273 28756 8359
rect 28316 6847 28756 8273
rect 28316 6761 28409 6847
rect 28495 6761 28577 6847
rect 28663 6761 28756 6847
rect 28316 5335 28756 6761
rect 28316 5249 28409 5335
rect 28495 5249 28577 5335
rect 28663 5249 28756 5335
rect 28316 4906 28756 5249
rect 28316 4526 28346 4906
rect 28726 4526 28756 4906
rect 28316 3823 28756 4526
rect 28316 3737 28409 3823
rect 28495 3737 28577 3823
rect 28663 3737 28756 3823
rect 28316 2311 28756 3737
rect 28316 2225 28409 2311
rect 28495 2225 28577 2311
rect 28663 2225 28756 2311
rect 28316 799 28756 2225
rect 28316 713 28409 799
rect 28495 713 28577 799
rect 28663 713 28756 799
rect 28316 630 28756 713
rect 31076 37843 31516 38600
rect 31076 37757 31169 37843
rect 31255 37757 31337 37843
rect 31423 37757 31516 37843
rect 31076 36331 31516 37757
rect 31076 36245 31169 36331
rect 31255 36245 31337 36331
rect 31423 36245 31516 36331
rect 31076 35666 31516 36245
rect 31076 35286 31106 35666
rect 31486 35286 31516 35666
rect 31076 34819 31516 35286
rect 31076 34733 31169 34819
rect 31255 34733 31337 34819
rect 31423 34733 31516 34819
rect 31076 33307 31516 34733
rect 31076 33221 31169 33307
rect 31255 33221 31337 33307
rect 31423 33221 31516 33307
rect 31076 31795 31516 33221
rect 31076 31709 31169 31795
rect 31255 31709 31337 31795
rect 31423 31709 31516 31795
rect 31076 31666 31516 31709
rect 31076 31286 31106 31666
rect 31486 31286 31516 31666
rect 31076 30283 31516 31286
rect 31076 30197 31169 30283
rect 31255 30197 31337 30283
rect 31423 30197 31516 30283
rect 31076 28771 31516 30197
rect 31076 28685 31169 28771
rect 31255 28685 31337 28771
rect 31423 28685 31516 28771
rect 31076 27666 31516 28685
rect 31076 27286 31106 27666
rect 31486 27286 31516 27666
rect 31076 27259 31516 27286
rect 31076 27173 31169 27259
rect 31255 27173 31337 27259
rect 31423 27173 31516 27259
rect 31076 25747 31516 27173
rect 31076 25661 31169 25747
rect 31255 25661 31337 25747
rect 31423 25661 31516 25747
rect 31076 24235 31516 25661
rect 31076 24149 31169 24235
rect 31255 24149 31337 24235
rect 31423 24149 31516 24235
rect 31076 23666 31516 24149
rect 31076 23286 31106 23666
rect 31486 23286 31516 23666
rect 31076 22723 31516 23286
rect 31076 22637 31169 22723
rect 31255 22637 31337 22723
rect 31423 22637 31516 22723
rect 31076 21211 31516 22637
rect 31076 21125 31169 21211
rect 31255 21125 31337 21211
rect 31423 21125 31516 21211
rect 31076 19699 31516 21125
rect 31076 19666 31169 19699
rect 31255 19666 31337 19699
rect 31423 19666 31516 19699
rect 31076 19286 31106 19666
rect 31486 19286 31516 19666
rect 31076 18187 31516 19286
rect 31076 18101 31169 18187
rect 31255 18101 31337 18187
rect 31423 18101 31516 18187
rect 31076 16675 31516 18101
rect 31076 16589 31169 16675
rect 31255 16589 31337 16675
rect 31423 16589 31516 16675
rect 31076 15666 31516 16589
rect 31076 15286 31106 15666
rect 31486 15286 31516 15666
rect 31076 15163 31516 15286
rect 31076 15077 31169 15163
rect 31255 15077 31337 15163
rect 31423 15077 31516 15163
rect 31076 13651 31516 15077
rect 31076 13565 31169 13651
rect 31255 13565 31337 13651
rect 31423 13565 31516 13651
rect 31076 12139 31516 13565
rect 31076 12053 31169 12139
rect 31255 12053 31337 12139
rect 31423 12053 31516 12139
rect 31076 11666 31516 12053
rect 31076 11286 31106 11666
rect 31486 11286 31516 11666
rect 31076 10627 31516 11286
rect 31076 10541 31169 10627
rect 31255 10541 31337 10627
rect 31423 10541 31516 10627
rect 31076 9115 31516 10541
rect 31076 9029 31169 9115
rect 31255 9029 31337 9115
rect 31423 9029 31516 9115
rect 31076 7666 31516 9029
rect 31076 7286 31106 7666
rect 31486 7286 31516 7666
rect 31076 6091 31516 7286
rect 31076 6005 31169 6091
rect 31255 6005 31337 6091
rect 31423 6005 31516 6091
rect 31076 4579 31516 6005
rect 31076 4493 31169 4579
rect 31255 4493 31337 4579
rect 31423 4493 31516 4579
rect 31076 3666 31516 4493
rect 31076 3286 31106 3666
rect 31486 3286 31516 3666
rect 31076 3067 31516 3286
rect 31076 2981 31169 3067
rect 31255 2981 31337 3067
rect 31423 2981 31516 3067
rect 31076 1555 31516 2981
rect 31076 1469 31169 1555
rect 31255 1469 31337 1555
rect 31423 1469 31516 1555
rect 31076 712 31516 1469
rect 32316 38599 32756 38682
rect 32316 38513 32409 38599
rect 32495 38513 32577 38599
rect 32663 38513 32756 38599
rect 32316 37087 32756 38513
rect 32316 37001 32409 37087
rect 32495 37001 32577 37087
rect 32663 37001 32756 37087
rect 32316 36906 32756 37001
rect 32316 36526 32346 36906
rect 32726 36526 32756 36906
rect 32316 35575 32756 36526
rect 32316 35489 32409 35575
rect 32495 35489 32577 35575
rect 32663 35489 32756 35575
rect 32316 34063 32756 35489
rect 32316 33977 32409 34063
rect 32495 33977 32577 34063
rect 32663 33977 32756 34063
rect 32316 32906 32756 33977
rect 32316 32526 32346 32906
rect 32726 32526 32756 32906
rect 32316 32465 32409 32526
rect 32495 32465 32577 32526
rect 32663 32465 32756 32526
rect 32316 31039 32756 32465
rect 32316 30953 32409 31039
rect 32495 30953 32577 31039
rect 32663 30953 32756 31039
rect 32316 29527 32756 30953
rect 32316 29441 32409 29527
rect 32495 29441 32577 29527
rect 32663 29441 32756 29527
rect 32316 28906 32756 29441
rect 32316 28526 32346 28906
rect 32726 28526 32756 28906
rect 32316 28015 32756 28526
rect 32316 27929 32409 28015
rect 32495 27929 32577 28015
rect 32663 27929 32756 28015
rect 32316 26503 32756 27929
rect 32316 26417 32409 26503
rect 32495 26417 32577 26503
rect 32663 26417 32756 26503
rect 32316 24991 32756 26417
rect 32316 24906 32409 24991
rect 32495 24906 32577 24991
rect 32663 24906 32756 24991
rect 32316 24526 32346 24906
rect 32726 24526 32756 24906
rect 32316 23479 32756 24526
rect 32316 23393 32409 23479
rect 32495 23393 32577 23479
rect 32663 23393 32756 23479
rect 32316 21967 32756 23393
rect 32316 21881 32409 21967
rect 32495 21881 32577 21967
rect 32663 21881 32756 21967
rect 32316 20906 32756 21881
rect 32316 20526 32346 20906
rect 32726 20526 32756 20906
rect 32316 20455 32756 20526
rect 32316 20369 32409 20455
rect 32495 20369 32577 20455
rect 32663 20369 32756 20455
rect 32316 18943 32756 20369
rect 32316 18857 32409 18943
rect 32495 18857 32577 18943
rect 32663 18857 32756 18943
rect 32316 17431 32756 18857
rect 32316 17345 32409 17431
rect 32495 17345 32577 17431
rect 32663 17345 32756 17431
rect 32316 16906 32756 17345
rect 32316 16526 32346 16906
rect 32726 16526 32756 16906
rect 32316 15919 32756 16526
rect 32316 15833 32409 15919
rect 32495 15833 32577 15919
rect 32663 15833 32756 15919
rect 32316 14407 32756 15833
rect 32316 14321 32409 14407
rect 32495 14321 32577 14407
rect 32663 14321 32756 14407
rect 32316 12906 32756 14321
rect 32316 12526 32346 12906
rect 32726 12526 32756 12906
rect 32316 11383 32756 12526
rect 32316 11297 32409 11383
rect 32495 11297 32577 11383
rect 32663 11297 32756 11383
rect 32316 9871 32756 11297
rect 32316 9785 32409 9871
rect 32495 9785 32577 9871
rect 32663 9785 32756 9871
rect 32316 8906 32756 9785
rect 32316 8526 32346 8906
rect 32726 8526 32756 8906
rect 32316 8359 32756 8526
rect 32316 8273 32409 8359
rect 32495 8273 32577 8359
rect 32663 8273 32756 8359
rect 32316 6847 32756 8273
rect 32316 6761 32409 6847
rect 32495 6761 32577 6847
rect 32663 6761 32756 6847
rect 32316 5335 32756 6761
rect 32316 5249 32409 5335
rect 32495 5249 32577 5335
rect 32663 5249 32756 5335
rect 32316 4906 32756 5249
rect 32316 4526 32346 4906
rect 32726 4526 32756 4906
rect 32316 3823 32756 4526
rect 32316 3737 32409 3823
rect 32495 3737 32577 3823
rect 32663 3737 32756 3823
rect 32316 2311 32756 3737
rect 32316 2225 32409 2311
rect 32495 2225 32577 2311
rect 32663 2225 32756 2311
rect 32316 799 32756 2225
rect 32316 713 32409 799
rect 32495 713 32577 799
rect 32663 713 32756 799
rect 32316 630 32756 713
rect 35076 37843 35516 38600
rect 35076 37757 35169 37843
rect 35255 37757 35337 37843
rect 35423 37757 35516 37843
rect 35076 36331 35516 37757
rect 35076 36245 35169 36331
rect 35255 36245 35337 36331
rect 35423 36245 35516 36331
rect 35076 35666 35516 36245
rect 35076 35286 35106 35666
rect 35486 35286 35516 35666
rect 35076 34819 35516 35286
rect 35076 34733 35169 34819
rect 35255 34733 35337 34819
rect 35423 34733 35516 34819
rect 35076 33307 35516 34733
rect 35076 33221 35169 33307
rect 35255 33221 35337 33307
rect 35423 33221 35516 33307
rect 35076 31795 35516 33221
rect 35076 31709 35169 31795
rect 35255 31709 35337 31795
rect 35423 31709 35516 31795
rect 35076 31666 35516 31709
rect 35076 31286 35106 31666
rect 35486 31286 35516 31666
rect 35076 30283 35516 31286
rect 35076 30197 35169 30283
rect 35255 30197 35337 30283
rect 35423 30197 35516 30283
rect 35076 28771 35516 30197
rect 35076 28685 35169 28771
rect 35255 28685 35337 28771
rect 35423 28685 35516 28771
rect 35076 27666 35516 28685
rect 35076 27286 35106 27666
rect 35486 27286 35516 27666
rect 35076 27259 35516 27286
rect 35076 27173 35169 27259
rect 35255 27173 35337 27259
rect 35423 27173 35516 27259
rect 35076 25747 35516 27173
rect 35076 25661 35169 25747
rect 35255 25661 35337 25747
rect 35423 25661 35516 25747
rect 35076 24235 35516 25661
rect 35076 24149 35169 24235
rect 35255 24149 35337 24235
rect 35423 24149 35516 24235
rect 35076 23666 35516 24149
rect 35076 23286 35106 23666
rect 35486 23286 35516 23666
rect 35076 22723 35516 23286
rect 35076 22637 35169 22723
rect 35255 22637 35337 22723
rect 35423 22637 35516 22723
rect 35076 21211 35516 22637
rect 35076 21125 35169 21211
rect 35255 21125 35337 21211
rect 35423 21125 35516 21211
rect 35076 19699 35516 21125
rect 35076 19666 35169 19699
rect 35255 19666 35337 19699
rect 35423 19666 35516 19699
rect 35076 19286 35106 19666
rect 35486 19286 35516 19666
rect 35076 18187 35516 19286
rect 35076 18101 35169 18187
rect 35255 18101 35337 18187
rect 35423 18101 35516 18187
rect 35076 16675 35516 18101
rect 35076 16589 35169 16675
rect 35255 16589 35337 16675
rect 35423 16589 35516 16675
rect 35076 15666 35516 16589
rect 35076 15286 35106 15666
rect 35486 15286 35516 15666
rect 35076 15163 35516 15286
rect 35076 15077 35169 15163
rect 35255 15077 35337 15163
rect 35423 15077 35516 15163
rect 35076 13651 35516 15077
rect 35076 13565 35169 13651
rect 35255 13565 35337 13651
rect 35423 13565 35516 13651
rect 35076 12139 35516 13565
rect 35076 12053 35169 12139
rect 35255 12053 35337 12139
rect 35423 12053 35516 12139
rect 35076 11666 35516 12053
rect 35076 11286 35106 11666
rect 35486 11286 35516 11666
rect 35076 10627 35516 11286
rect 35076 10541 35169 10627
rect 35255 10541 35337 10627
rect 35423 10541 35516 10627
rect 35076 9115 35516 10541
rect 35076 9029 35169 9115
rect 35255 9029 35337 9115
rect 35423 9029 35516 9115
rect 35076 7666 35516 9029
rect 35076 7286 35106 7666
rect 35486 7286 35516 7666
rect 35076 6091 35516 7286
rect 35076 6005 35169 6091
rect 35255 6005 35337 6091
rect 35423 6005 35516 6091
rect 35076 4579 35516 6005
rect 35076 4493 35169 4579
rect 35255 4493 35337 4579
rect 35423 4493 35516 4579
rect 35076 3666 35516 4493
rect 35076 3286 35106 3666
rect 35486 3286 35516 3666
rect 35076 3067 35516 3286
rect 35076 2981 35169 3067
rect 35255 2981 35337 3067
rect 35423 2981 35516 3067
rect 35076 1555 35516 2981
rect 35076 1469 35169 1555
rect 35255 1469 35337 1555
rect 35423 1469 35516 1555
rect 35076 712 35516 1469
rect 36316 38599 36756 38682
rect 36316 38513 36409 38599
rect 36495 38513 36577 38599
rect 36663 38513 36756 38599
rect 36316 37087 36756 38513
rect 36316 37001 36409 37087
rect 36495 37001 36577 37087
rect 36663 37001 36756 37087
rect 36316 36906 36756 37001
rect 36316 36526 36346 36906
rect 36726 36526 36756 36906
rect 36316 35575 36756 36526
rect 36316 35489 36409 35575
rect 36495 35489 36577 35575
rect 36663 35489 36756 35575
rect 36316 34063 36756 35489
rect 36316 33977 36409 34063
rect 36495 33977 36577 34063
rect 36663 33977 36756 34063
rect 36316 32906 36756 33977
rect 36316 32526 36346 32906
rect 36726 32526 36756 32906
rect 36316 32465 36409 32526
rect 36495 32465 36577 32526
rect 36663 32465 36756 32526
rect 36316 31039 36756 32465
rect 36316 30953 36409 31039
rect 36495 30953 36577 31039
rect 36663 30953 36756 31039
rect 36316 29527 36756 30953
rect 36316 29441 36409 29527
rect 36495 29441 36577 29527
rect 36663 29441 36756 29527
rect 36316 28906 36756 29441
rect 36316 28526 36346 28906
rect 36726 28526 36756 28906
rect 36316 28015 36756 28526
rect 36316 27929 36409 28015
rect 36495 27929 36577 28015
rect 36663 27929 36756 28015
rect 36316 26503 36756 27929
rect 36316 26417 36409 26503
rect 36495 26417 36577 26503
rect 36663 26417 36756 26503
rect 36316 24991 36756 26417
rect 36316 24906 36409 24991
rect 36495 24906 36577 24991
rect 36663 24906 36756 24991
rect 36316 24526 36346 24906
rect 36726 24526 36756 24906
rect 36316 23479 36756 24526
rect 36316 23393 36409 23479
rect 36495 23393 36577 23479
rect 36663 23393 36756 23479
rect 36316 21967 36756 23393
rect 36316 21881 36409 21967
rect 36495 21881 36577 21967
rect 36663 21881 36756 21967
rect 36316 20906 36756 21881
rect 36316 20526 36346 20906
rect 36726 20526 36756 20906
rect 36316 20455 36756 20526
rect 36316 20369 36409 20455
rect 36495 20369 36577 20455
rect 36663 20369 36756 20455
rect 36316 18943 36756 20369
rect 36316 18857 36409 18943
rect 36495 18857 36577 18943
rect 36663 18857 36756 18943
rect 36316 17431 36756 18857
rect 36316 17345 36409 17431
rect 36495 17345 36577 17431
rect 36663 17345 36756 17431
rect 36316 16906 36756 17345
rect 36316 16526 36346 16906
rect 36726 16526 36756 16906
rect 36316 15919 36756 16526
rect 36316 15833 36409 15919
rect 36495 15833 36577 15919
rect 36663 15833 36756 15919
rect 36316 14407 36756 15833
rect 36316 14321 36409 14407
rect 36495 14321 36577 14407
rect 36663 14321 36756 14407
rect 36316 12906 36756 14321
rect 36316 12526 36346 12906
rect 36726 12526 36756 12906
rect 36316 11383 36756 12526
rect 36316 11297 36409 11383
rect 36495 11297 36577 11383
rect 36663 11297 36756 11383
rect 36316 9871 36756 11297
rect 36316 9785 36409 9871
rect 36495 9785 36577 9871
rect 36663 9785 36756 9871
rect 36316 8906 36756 9785
rect 36316 8526 36346 8906
rect 36726 8526 36756 8906
rect 36316 8359 36756 8526
rect 36316 8273 36409 8359
rect 36495 8273 36577 8359
rect 36663 8273 36756 8359
rect 36316 6847 36756 8273
rect 36316 6761 36409 6847
rect 36495 6761 36577 6847
rect 36663 6761 36756 6847
rect 36316 5335 36756 6761
rect 36316 5249 36409 5335
rect 36495 5249 36577 5335
rect 36663 5249 36756 5335
rect 36316 4906 36756 5249
rect 36316 4526 36346 4906
rect 36726 4526 36756 4906
rect 36316 3823 36756 4526
rect 36316 3737 36409 3823
rect 36495 3737 36577 3823
rect 36663 3737 36756 3823
rect 36316 2311 36756 3737
rect 36316 2225 36409 2311
rect 36495 2225 36577 2311
rect 36663 2225 36756 2311
rect 36316 799 36756 2225
rect 36316 713 36409 799
rect 36495 713 36577 799
rect 36663 713 36756 799
rect 36316 630 36756 713
rect 39076 37843 39516 38600
rect 39076 37757 39169 37843
rect 39255 37757 39337 37843
rect 39423 37757 39516 37843
rect 39076 36331 39516 37757
rect 39076 36245 39169 36331
rect 39255 36245 39337 36331
rect 39423 36245 39516 36331
rect 39076 35666 39516 36245
rect 39076 35286 39106 35666
rect 39486 35286 39516 35666
rect 39076 34819 39516 35286
rect 39076 34733 39169 34819
rect 39255 34733 39337 34819
rect 39423 34733 39516 34819
rect 39076 33307 39516 34733
rect 39076 33221 39169 33307
rect 39255 33221 39337 33307
rect 39423 33221 39516 33307
rect 39076 31795 39516 33221
rect 39076 31709 39169 31795
rect 39255 31709 39337 31795
rect 39423 31709 39516 31795
rect 39076 31666 39516 31709
rect 39076 31286 39106 31666
rect 39486 31286 39516 31666
rect 39076 30283 39516 31286
rect 39076 30197 39169 30283
rect 39255 30197 39337 30283
rect 39423 30197 39516 30283
rect 39076 28771 39516 30197
rect 39076 28685 39169 28771
rect 39255 28685 39337 28771
rect 39423 28685 39516 28771
rect 39076 27666 39516 28685
rect 39076 27286 39106 27666
rect 39486 27286 39516 27666
rect 39076 27259 39516 27286
rect 39076 27173 39169 27259
rect 39255 27173 39337 27259
rect 39423 27173 39516 27259
rect 39076 25747 39516 27173
rect 39076 25661 39169 25747
rect 39255 25661 39337 25747
rect 39423 25661 39516 25747
rect 39076 24235 39516 25661
rect 39076 24149 39169 24235
rect 39255 24149 39337 24235
rect 39423 24149 39516 24235
rect 39076 23666 39516 24149
rect 39076 23286 39106 23666
rect 39486 23286 39516 23666
rect 39076 22723 39516 23286
rect 39076 22637 39169 22723
rect 39255 22637 39337 22723
rect 39423 22637 39516 22723
rect 39076 21211 39516 22637
rect 39076 21125 39169 21211
rect 39255 21125 39337 21211
rect 39423 21125 39516 21211
rect 39076 19699 39516 21125
rect 39076 19666 39169 19699
rect 39255 19666 39337 19699
rect 39423 19666 39516 19699
rect 39076 19286 39106 19666
rect 39486 19286 39516 19666
rect 39076 18187 39516 19286
rect 39076 18101 39169 18187
rect 39255 18101 39337 18187
rect 39423 18101 39516 18187
rect 39076 16675 39516 18101
rect 39076 16589 39169 16675
rect 39255 16589 39337 16675
rect 39423 16589 39516 16675
rect 39076 15666 39516 16589
rect 39076 15286 39106 15666
rect 39486 15286 39516 15666
rect 39076 15163 39516 15286
rect 39076 15077 39169 15163
rect 39255 15077 39337 15163
rect 39423 15077 39516 15163
rect 39076 13651 39516 15077
rect 39076 13565 39169 13651
rect 39255 13565 39337 13651
rect 39423 13565 39516 13651
rect 39076 12139 39516 13565
rect 39076 12053 39169 12139
rect 39255 12053 39337 12139
rect 39423 12053 39516 12139
rect 39076 11666 39516 12053
rect 39076 11286 39106 11666
rect 39486 11286 39516 11666
rect 39076 10627 39516 11286
rect 39076 10541 39169 10627
rect 39255 10541 39337 10627
rect 39423 10541 39516 10627
rect 39076 9115 39516 10541
rect 39076 9029 39169 9115
rect 39255 9029 39337 9115
rect 39423 9029 39516 9115
rect 39076 7666 39516 9029
rect 39076 7286 39106 7666
rect 39486 7286 39516 7666
rect 39076 6091 39516 7286
rect 39076 6005 39169 6091
rect 39255 6005 39337 6091
rect 39423 6005 39516 6091
rect 39076 4579 39516 6005
rect 39076 4493 39169 4579
rect 39255 4493 39337 4579
rect 39423 4493 39516 4579
rect 39076 3666 39516 4493
rect 39076 3286 39106 3666
rect 39486 3286 39516 3666
rect 39076 3067 39516 3286
rect 39076 2981 39169 3067
rect 39255 2981 39337 3067
rect 39423 2981 39516 3067
rect 39076 1555 39516 2981
rect 39076 1469 39169 1555
rect 39255 1469 39337 1555
rect 39423 1469 39516 1555
rect 39076 712 39516 1469
rect 40316 38599 40756 38682
rect 40316 38513 40409 38599
rect 40495 38513 40577 38599
rect 40663 38513 40756 38599
rect 40316 37087 40756 38513
rect 40316 37001 40409 37087
rect 40495 37001 40577 37087
rect 40663 37001 40756 37087
rect 40316 36906 40756 37001
rect 40316 36526 40346 36906
rect 40726 36526 40756 36906
rect 40316 35575 40756 36526
rect 40316 35489 40409 35575
rect 40495 35489 40577 35575
rect 40663 35489 40756 35575
rect 40316 34063 40756 35489
rect 40316 33977 40409 34063
rect 40495 33977 40577 34063
rect 40663 33977 40756 34063
rect 40316 32906 40756 33977
rect 40316 32526 40346 32906
rect 40726 32526 40756 32906
rect 40316 32465 40409 32526
rect 40495 32465 40577 32526
rect 40663 32465 40756 32526
rect 40316 31039 40756 32465
rect 40316 30953 40409 31039
rect 40495 30953 40577 31039
rect 40663 30953 40756 31039
rect 40316 29527 40756 30953
rect 40316 29441 40409 29527
rect 40495 29441 40577 29527
rect 40663 29441 40756 29527
rect 40316 28906 40756 29441
rect 40316 28526 40346 28906
rect 40726 28526 40756 28906
rect 40316 28015 40756 28526
rect 40316 27929 40409 28015
rect 40495 27929 40577 28015
rect 40663 27929 40756 28015
rect 40316 26503 40756 27929
rect 40316 26417 40409 26503
rect 40495 26417 40577 26503
rect 40663 26417 40756 26503
rect 40316 24991 40756 26417
rect 40316 24906 40409 24991
rect 40495 24906 40577 24991
rect 40663 24906 40756 24991
rect 40316 24526 40346 24906
rect 40726 24526 40756 24906
rect 40316 23479 40756 24526
rect 40316 23393 40409 23479
rect 40495 23393 40577 23479
rect 40663 23393 40756 23479
rect 40316 21967 40756 23393
rect 40316 21881 40409 21967
rect 40495 21881 40577 21967
rect 40663 21881 40756 21967
rect 40316 20906 40756 21881
rect 40316 20526 40346 20906
rect 40726 20526 40756 20906
rect 40316 20455 40756 20526
rect 40316 20369 40409 20455
rect 40495 20369 40577 20455
rect 40663 20369 40756 20455
rect 40316 18943 40756 20369
rect 40316 18857 40409 18943
rect 40495 18857 40577 18943
rect 40663 18857 40756 18943
rect 40316 17431 40756 18857
rect 40316 17345 40409 17431
rect 40495 17345 40577 17431
rect 40663 17345 40756 17431
rect 40316 16906 40756 17345
rect 40316 16526 40346 16906
rect 40726 16526 40756 16906
rect 40316 15919 40756 16526
rect 40316 15833 40409 15919
rect 40495 15833 40577 15919
rect 40663 15833 40756 15919
rect 40316 14407 40756 15833
rect 40316 14321 40409 14407
rect 40495 14321 40577 14407
rect 40663 14321 40756 14407
rect 40316 12906 40756 14321
rect 40316 12526 40346 12906
rect 40726 12526 40756 12906
rect 40316 11383 40756 12526
rect 40316 11297 40409 11383
rect 40495 11297 40577 11383
rect 40663 11297 40756 11383
rect 40316 9871 40756 11297
rect 40316 9785 40409 9871
rect 40495 9785 40577 9871
rect 40663 9785 40756 9871
rect 40316 8906 40756 9785
rect 40316 8526 40346 8906
rect 40726 8526 40756 8906
rect 40316 8359 40756 8526
rect 40316 8273 40409 8359
rect 40495 8273 40577 8359
rect 40663 8273 40756 8359
rect 40316 6847 40756 8273
rect 40316 6761 40409 6847
rect 40495 6761 40577 6847
rect 40663 6761 40756 6847
rect 40316 5335 40756 6761
rect 40316 5249 40409 5335
rect 40495 5249 40577 5335
rect 40663 5249 40756 5335
rect 40316 4906 40756 5249
rect 40316 4526 40346 4906
rect 40726 4526 40756 4906
rect 40316 3823 40756 4526
rect 40316 3737 40409 3823
rect 40495 3737 40577 3823
rect 40663 3737 40756 3823
rect 40316 2311 40756 3737
rect 40316 2225 40409 2311
rect 40495 2225 40577 2311
rect 40663 2225 40756 2311
rect 40316 799 40756 2225
rect 40316 713 40409 799
rect 40495 713 40577 799
rect 40663 713 40756 799
rect 40316 630 40756 713
rect 43076 37843 43516 38600
rect 43076 37757 43169 37843
rect 43255 37757 43337 37843
rect 43423 37757 43516 37843
rect 43076 36331 43516 37757
rect 43076 36245 43169 36331
rect 43255 36245 43337 36331
rect 43423 36245 43516 36331
rect 43076 35666 43516 36245
rect 43076 35286 43106 35666
rect 43486 35286 43516 35666
rect 43076 34819 43516 35286
rect 43076 34733 43169 34819
rect 43255 34733 43337 34819
rect 43423 34733 43516 34819
rect 43076 33307 43516 34733
rect 43076 33221 43169 33307
rect 43255 33221 43337 33307
rect 43423 33221 43516 33307
rect 43076 31795 43516 33221
rect 43076 31709 43169 31795
rect 43255 31709 43337 31795
rect 43423 31709 43516 31795
rect 43076 31666 43516 31709
rect 43076 31286 43106 31666
rect 43486 31286 43516 31666
rect 43076 30283 43516 31286
rect 43076 30197 43169 30283
rect 43255 30197 43337 30283
rect 43423 30197 43516 30283
rect 43076 28771 43516 30197
rect 43076 28685 43169 28771
rect 43255 28685 43337 28771
rect 43423 28685 43516 28771
rect 43076 27666 43516 28685
rect 43076 27286 43106 27666
rect 43486 27286 43516 27666
rect 43076 27259 43516 27286
rect 43076 27173 43169 27259
rect 43255 27173 43337 27259
rect 43423 27173 43516 27259
rect 43076 25747 43516 27173
rect 43076 25661 43169 25747
rect 43255 25661 43337 25747
rect 43423 25661 43516 25747
rect 43076 24235 43516 25661
rect 43076 24149 43169 24235
rect 43255 24149 43337 24235
rect 43423 24149 43516 24235
rect 43076 23666 43516 24149
rect 43076 23286 43106 23666
rect 43486 23286 43516 23666
rect 43076 22723 43516 23286
rect 43076 22637 43169 22723
rect 43255 22637 43337 22723
rect 43423 22637 43516 22723
rect 43076 21211 43516 22637
rect 43076 21125 43169 21211
rect 43255 21125 43337 21211
rect 43423 21125 43516 21211
rect 43076 19699 43516 21125
rect 43076 19666 43169 19699
rect 43255 19666 43337 19699
rect 43423 19666 43516 19699
rect 43076 19286 43106 19666
rect 43486 19286 43516 19666
rect 43076 18187 43516 19286
rect 43076 18101 43169 18187
rect 43255 18101 43337 18187
rect 43423 18101 43516 18187
rect 43076 16675 43516 18101
rect 43076 16589 43169 16675
rect 43255 16589 43337 16675
rect 43423 16589 43516 16675
rect 43076 15666 43516 16589
rect 43076 15286 43106 15666
rect 43486 15286 43516 15666
rect 43076 15163 43516 15286
rect 43076 15077 43169 15163
rect 43255 15077 43337 15163
rect 43423 15077 43516 15163
rect 43076 13651 43516 15077
rect 43076 13565 43169 13651
rect 43255 13565 43337 13651
rect 43423 13565 43516 13651
rect 43076 12139 43516 13565
rect 43076 12053 43169 12139
rect 43255 12053 43337 12139
rect 43423 12053 43516 12139
rect 43076 11666 43516 12053
rect 43076 11286 43106 11666
rect 43486 11286 43516 11666
rect 43076 10627 43516 11286
rect 43076 10541 43169 10627
rect 43255 10541 43337 10627
rect 43423 10541 43516 10627
rect 43076 9115 43516 10541
rect 43076 9029 43169 9115
rect 43255 9029 43337 9115
rect 43423 9029 43516 9115
rect 43076 7666 43516 9029
rect 43076 7286 43106 7666
rect 43486 7286 43516 7666
rect 43076 6091 43516 7286
rect 43076 6005 43169 6091
rect 43255 6005 43337 6091
rect 43423 6005 43516 6091
rect 43076 4579 43516 6005
rect 43076 4493 43169 4579
rect 43255 4493 43337 4579
rect 43423 4493 43516 4579
rect 43076 3666 43516 4493
rect 43076 3286 43106 3666
rect 43486 3286 43516 3666
rect 43076 3067 43516 3286
rect 43076 2981 43169 3067
rect 43255 2981 43337 3067
rect 43423 2981 43516 3067
rect 43076 1555 43516 2981
rect 43076 1469 43169 1555
rect 43255 1469 43337 1555
rect 43423 1469 43516 1555
rect 43076 712 43516 1469
rect 44316 38599 44756 38682
rect 44316 38513 44409 38599
rect 44495 38513 44577 38599
rect 44663 38513 44756 38599
rect 44316 37087 44756 38513
rect 44316 37001 44409 37087
rect 44495 37001 44577 37087
rect 44663 37001 44756 37087
rect 44316 36906 44756 37001
rect 44316 36526 44346 36906
rect 44726 36526 44756 36906
rect 44316 35575 44756 36526
rect 44316 35489 44409 35575
rect 44495 35489 44577 35575
rect 44663 35489 44756 35575
rect 44316 34063 44756 35489
rect 44316 33977 44409 34063
rect 44495 33977 44577 34063
rect 44663 33977 44756 34063
rect 44316 32906 44756 33977
rect 44316 32526 44346 32906
rect 44726 32526 44756 32906
rect 44316 32465 44409 32526
rect 44495 32465 44577 32526
rect 44663 32465 44756 32526
rect 44316 31039 44756 32465
rect 44316 30953 44409 31039
rect 44495 30953 44577 31039
rect 44663 30953 44756 31039
rect 44316 29527 44756 30953
rect 44316 29441 44409 29527
rect 44495 29441 44577 29527
rect 44663 29441 44756 29527
rect 44316 28906 44756 29441
rect 44316 28526 44346 28906
rect 44726 28526 44756 28906
rect 44316 28015 44756 28526
rect 44316 27929 44409 28015
rect 44495 27929 44577 28015
rect 44663 27929 44756 28015
rect 44316 26503 44756 27929
rect 44316 26417 44409 26503
rect 44495 26417 44577 26503
rect 44663 26417 44756 26503
rect 44316 24991 44756 26417
rect 44316 24906 44409 24991
rect 44495 24906 44577 24991
rect 44663 24906 44756 24991
rect 44316 24526 44346 24906
rect 44726 24526 44756 24906
rect 44316 23479 44756 24526
rect 44316 23393 44409 23479
rect 44495 23393 44577 23479
rect 44663 23393 44756 23479
rect 44316 21967 44756 23393
rect 44316 21881 44409 21967
rect 44495 21881 44577 21967
rect 44663 21881 44756 21967
rect 44316 20906 44756 21881
rect 44316 20526 44346 20906
rect 44726 20526 44756 20906
rect 44316 20455 44756 20526
rect 44316 20369 44409 20455
rect 44495 20369 44577 20455
rect 44663 20369 44756 20455
rect 44316 18943 44756 20369
rect 44316 18857 44409 18943
rect 44495 18857 44577 18943
rect 44663 18857 44756 18943
rect 44316 17431 44756 18857
rect 44316 17345 44409 17431
rect 44495 17345 44577 17431
rect 44663 17345 44756 17431
rect 44316 16906 44756 17345
rect 44316 16526 44346 16906
rect 44726 16526 44756 16906
rect 44316 15919 44756 16526
rect 44316 15833 44409 15919
rect 44495 15833 44577 15919
rect 44663 15833 44756 15919
rect 44316 14407 44756 15833
rect 44316 14321 44409 14407
rect 44495 14321 44577 14407
rect 44663 14321 44756 14407
rect 44316 12906 44756 14321
rect 44316 12526 44346 12906
rect 44726 12526 44756 12906
rect 44316 11383 44756 12526
rect 44316 11297 44409 11383
rect 44495 11297 44577 11383
rect 44663 11297 44756 11383
rect 44316 9871 44756 11297
rect 44316 9785 44409 9871
rect 44495 9785 44577 9871
rect 44663 9785 44756 9871
rect 44316 8906 44756 9785
rect 44316 8526 44346 8906
rect 44726 8526 44756 8906
rect 44316 8359 44756 8526
rect 44316 8273 44409 8359
rect 44495 8273 44577 8359
rect 44663 8273 44756 8359
rect 44316 6847 44756 8273
rect 44316 6761 44409 6847
rect 44495 6761 44577 6847
rect 44663 6761 44756 6847
rect 44316 5335 44756 6761
rect 44316 5249 44409 5335
rect 44495 5249 44577 5335
rect 44663 5249 44756 5335
rect 44316 4906 44756 5249
rect 44316 4526 44346 4906
rect 44726 4526 44756 4906
rect 44316 3823 44756 4526
rect 44316 3737 44409 3823
rect 44495 3737 44577 3823
rect 44663 3737 44756 3823
rect 44316 2311 44756 3737
rect 44316 2225 44409 2311
rect 44495 2225 44577 2311
rect 44663 2225 44756 2311
rect 44316 799 44756 2225
rect 44316 713 44409 799
rect 44495 713 44577 799
rect 44663 713 44756 799
rect 44316 630 44756 713
rect 47076 37843 47516 38600
rect 47076 37757 47169 37843
rect 47255 37757 47337 37843
rect 47423 37757 47516 37843
rect 47076 36331 47516 37757
rect 47076 36245 47169 36331
rect 47255 36245 47337 36331
rect 47423 36245 47516 36331
rect 47076 35666 47516 36245
rect 47076 35286 47106 35666
rect 47486 35286 47516 35666
rect 47076 34819 47516 35286
rect 47076 34733 47169 34819
rect 47255 34733 47337 34819
rect 47423 34733 47516 34819
rect 47076 33307 47516 34733
rect 47076 33221 47169 33307
rect 47255 33221 47337 33307
rect 47423 33221 47516 33307
rect 47076 31795 47516 33221
rect 47076 31709 47169 31795
rect 47255 31709 47337 31795
rect 47423 31709 47516 31795
rect 47076 31666 47516 31709
rect 47076 31286 47106 31666
rect 47486 31286 47516 31666
rect 47076 30283 47516 31286
rect 47076 30197 47169 30283
rect 47255 30197 47337 30283
rect 47423 30197 47516 30283
rect 47076 28771 47516 30197
rect 47076 28685 47169 28771
rect 47255 28685 47337 28771
rect 47423 28685 47516 28771
rect 47076 27666 47516 28685
rect 47076 27286 47106 27666
rect 47486 27286 47516 27666
rect 47076 27259 47516 27286
rect 47076 27173 47169 27259
rect 47255 27173 47337 27259
rect 47423 27173 47516 27259
rect 47076 25747 47516 27173
rect 47076 25661 47169 25747
rect 47255 25661 47337 25747
rect 47423 25661 47516 25747
rect 47076 24235 47516 25661
rect 47076 24149 47169 24235
rect 47255 24149 47337 24235
rect 47423 24149 47516 24235
rect 47076 23666 47516 24149
rect 47076 23286 47106 23666
rect 47486 23286 47516 23666
rect 47076 22723 47516 23286
rect 47076 22637 47169 22723
rect 47255 22637 47337 22723
rect 47423 22637 47516 22723
rect 47076 21211 47516 22637
rect 47076 21125 47169 21211
rect 47255 21125 47337 21211
rect 47423 21125 47516 21211
rect 47076 19699 47516 21125
rect 47076 19666 47169 19699
rect 47255 19666 47337 19699
rect 47423 19666 47516 19699
rect 47076 19286 47106 19666
rect 47486 19286 47516 19666
rect 47076 18187 47516 19286
rect 47076 18101 47169 18187
rect 47255 18101 47337 18187
rect 47423 18101 47516 18187
rect 47076 16675 47516 18101
rect 47076 16589 47169 16675
rect 47255 16589 47337 16675
rect 47423 16589 47516 16675
rect 47076 15666 47516 16589
rect 47076 15286 47106 15666
rect 47486 15286 47516 15666
rect 47076 15163 47516 15286
rect 47076 15077 47169 15163
rect 47255 15077 47337 15163
rect 47423 15077 47516 15163
rect 47076 13651 47516 15077
rect 47076 13565 47169 13651
rect 47255 13565 47337 13651
rect 47423 13565 47516 13651
rect 47076 12139 47516 13565
rect 47076 12053 47169 12139
rect 47255 12053 47337 12139
rect 47423 12053 47516 12139
rect 47076 11666 47516 12053
rect 47076 11286 47106 11666
rect 47486 11286 47516 11666
rect 47076 10627 47516 11286
rect 47076 10541 47169 10627
rect 47255 10541 47337 10627
rect 47423 10541 47516 10627
rect 47076 9115 47516 10541
rect 47076 9029 47169 9115
rect 47255 9029 47337 9115
rect 47423 9029 47516 9115
rect 47076 7666 47516 9029
rect 47076 7286 47106 7666
rect 47486 7286 47516 7666
rect 47076 6091 47516 7286
rect 47076 6005 47169 6091
rect 47255 6005 47337 6091
rect 47423 6005 47516 6091
rect 47076 4579 47516 6005
rect 47076 4493 47169 4579
rect 47255 4493 47337 4579
rect 47423 4493 47516 4579
rect 47076 3666 47516 4493
rect 47076 3286 47106 3666
rect 47486 3286 47516 3666
rect 47076 3067 47516 3286
rect 47076 2981 47169 3067
rect 47255 2981 47337 3067
rect 47423 2981 47516 3067
rect 47076 1555 47516 2981
rect 47076 1469 47169 1555
rect 47255 1469 47337 1555
rect 47423 1469 47516 1555
rect 47076 712 47516 1469
rect 48316 38599 48756 38682
rect 48316 38513 48409 38599
rect 48495 38513 48577 38599
rect 48663 38513 48756 38599
rect 48316 37087 48756 38513
rect 48316 37001 48409 37087
rect 48495 37001 48577 37087
rect 48663 37001 48756 37087
rect 48316 36906 48756 37001
rect 48316 36526 48346 36906
rect 48726 36526 48756 36906
rect 48316 35575 48756 36526
rect 48316 35489 48409 35575
rect 48495 35489 48577 35575
rect 48663 35489 48756 35575
rect 48316 34063 48756 35489
rect 48316 33977 48409 34063
rect 48495 33977 48577 34063
rect 48663 33977 48756 34063
rect 48316 32906 48756 33977
rect 48316 32526 48346 32906
rect 48726 32526 48756 32906
rect 48316 32465 48409 32526
rect 48495 32465 48577 32526
rect 48663 32465 48756 32526
rect 48316 31039 48756 32465
rect 48316 30953 48409 31039
rect 48495 30953 48577 31039
rect 48663 30953 48756 31039
rect 48316 29527 48756 30953
rect 48316 29441 48409 29527
rect 48495 29441 48577 29527
rect 48663 29441 48756 29527
rect 48316 28906 48756 29441
rect 48316 28526 48346 28906
rect 48726 28526 48756 28906
rect 48316 28015 48756 28526
rect 48316 27929 48409 28015
rect 48495 27929 48577 28015
rect 48663 27929 48756 28015
rect 48316 26503 48756 27929
rect 48316 26417 48409 26503
rect 48495 26417 48577 26503
rect 48663 26417 48756 26503
rect 48316 24991 48756 26417
rect 48316 24906 48409 24991
rect 48495 24906 48577 24991
rect 48663 24906 48756 24991
rect 48316 24526 48346 24906
rect 48726 24526 48756 24906
rect 48316 23479 48756 24526
rect 48316 23393 48409 23479
rect 48495 23393 48577 23479
rect 48663 23393 48756 23479
rect 48316 21967 48756 23393
rect 48316 21881 48409 21967
rect 48495 21881 48577 21967
rect 48663 21881 48756 21967
rect 48316 20906 48756 21881
rect 48316 20526 48346 20906
rect 48726 20526 48756 20906
rect 48316 20455 48756 20526
rect 48316 20369 48409 20455
rect 48495 20369 48577 20455
rect 48663 20369 48756 20455
rect 48316 18943 48756 20369
rect 48316 18857 48409 18943
rect 48495 18857 48577 18943
rect 48663 18857 48756 18943
rect 48316 17431 48756 18857
rect 48316 17345 48409 17431
rect 48495 17345 48577 17431
rect 48663 17345 48756 17431
rect 48316 16906 48756 17345
rect 48316 16526 48346 16906
rect 48726 16526 48756 16906
rect 48316 15919 48756 16526
rect 48316 15833 48409 15919
rect 48495 15833 48577 15919
rect 48663 15833 48756 15919
rect 48316 14407 48756 15833
rect 48316 14321 48409 14407
rect 48495 14321 48577 14407
rect 48663 14321 48756 14407
rect 48316 12906 48756 14321
rect 48316 12526 48346 12906
rect 48726 12526 48756 12906
rect 48316 11383 48756 12526
rect 48316 11297 48409 11383
rect 48495 11297 48577 11383
rect 48663 11297 48756 11383
rect 48316 9871 48756 11297
rect 48316 9785 48409 9871
rect 48495 9785 48577 9871
rect 48663 9785 48756 9871
rect 48316 8906 48756 9785
rect 48316 8526 48346 8906
rect 48726 8526 48756 8906
rect 48316 8359 48756 8526
rect 48316 8273 48409 8359
rect 48495 8273 48577 8359
rect 48663 8273 48756 8359
rect 48316 6847 48756 8273
rect 48316 6761 48409 6847
rect 48495 6761 48577 6847
rect 48663 6761 48756 6847
rect 48316 5335 48756 6761
rect 48316 5249 48409 5335
rect 48495 5249 48577 5335
rect 48663 5249 48756 5335
rect 48316 4906 48756 5249
rect 48316 4526 48346 4906
rect 48726 4526 48756 4906
rect 48316 3823 48756 4526
rect 48316 3737 48409 3823
rect 48495 3737 48577 3823
rect 48663 3737 48756 3823
rect 48316 2311 48756 3737
rect 48316 2225 48409 2311
rect 48495 2225 48577 2311
rect 48663 2225 48756 2311
rect 48316 799 48756 2225
rect 48316 713 48409 799
rect 48495 713 48577 799
rect 48663 713 48756 799
rect 48316 630 48756 713
rect 51076 37843 51516 38600
rect 51076 37757 51169 37843
rect 51255 37757 51337 37843
rect 51423 37757 51516 37843
rect 51076 36331 51516 37757
rect 51076 36245 51169 36331
rect 51255 36245 51337 36331
rect 51423 36245 51516 36331
rect 51076 35666 51516 36245
rect 51076 35286 51106 35666
rect 51486 35286 51516 35666
rect 51076 34819 51516 35286
rect 51076 34733 51169 34819
rect 51255 34733 51337 34819
rect 51423 34733 51516 34819
rect 51076 33307 51516 34733
rect 51076 33221 51169 33307
rect 51255 33221 51337 33307
rect 51423 33221 51516 33307
rect 51076 31795 51516 33221
rect 51076 31709 51169 31795
rect 51255 31709 51337 31795
rect 51423 31709 51516 31795
rect 51076 31666 51516 31709
rect 51076 31286 51106 31666
rect 51486 31286 51516 31666
rect 51076 30283 51516 31286
rect 51076 30197 51169 30283
rect 51255 30197 51337 30283
rect 51423 30197 51516 30283
rect 51076 28771 51516 30197
rect 51076 28685 51169 28771
rect 51255 28685 51337 28771
rect 51423 28685 51516 28771
rect 51076 27666 51516 28685
rect 51076 27286 51106 27666
rect 51486 27286 51516 27666
rect 51076 27259 51516 27286
rect 51076 27173 51169 27259
rect 51255 27173 51337 27259
rect 51423 27173 51516 27259
rect 51076 25747 51516 27173
rect 51076 25661 51169 25747
rect 51255 25661 51337 25747
rect 51423 25661 51516 25747
rect 51076 24235 51516 25661
rect 51076 24149 51169 24235
rect 51255 24149 51337 24235
rect 51423 24149 51516 24235
rect 51076 23666 51516 24149
rect 51076 23286 51106 23666
rect 51486 23286 51516 23666
rect 51076 22723 51516 23286
rect 51076 22637 51169 22723
rect 51255 22637 51337 22723
rect 51423 22637 51516 22723
rect 51076 21211 51516 22637
rect 51076 21125 51169 21211
rect 51255 21125 51337 21211
rect 51423 21125 51516 21211
rect 51076 19699 51516 21125
rect 51076 19666 51169 19699
rect 51255 19666 51337 19699
rect 51423 19666 51516 19699
rect 51076 19286 51106 19666
rect 51486 19286 51516 19666
rect 51076 18187 51516 19286
rect 51076 18101 51169 18187
rect 51255 18101 51337 18187
rect 51423 18101 51516 18187
rect 51076 16675 51516 18101
rect 51076 16589 51169 16675
rect 51255 16589 51337 16675
rect 51423 16589 51516 16675
rect 51076 15666 51516 16589
rect 51076 15286 51106 15666
rect 51486 15286 51516 15666
rect 51076 15163 51516 15286
rect 51076 15077 51169 15163
rect 51255 15077 51337 15163
rect 51423 15077 51516 15163
rect 51076 13651 51516 15077
rect 51076 13565 51169 13651
rect 51255 13565 51337 13651
rect 51423 13565 51516 13651
rect 51076 12139 51516 13565
rect 51076 12053 51169 12139
rect 51255 12053 51337 12139
rect 51423 12053 51516 12139
rect 51076 11666 51516 12053
rect 51076 11286 51106 11666
rect 51486 11286 51516 11666
rect 51076 10627 51516 11286
rect 51076 10541 51169 10627
rect 51255 10541 51337 10627
rect 51423 10541 51516 10627
rect 51076 9115 51516 10541
rect 51076 9029 51169 9115
rect 51255 9029 51337 9115
rect 51423 9029 51516 9115
rect 51076 7666 51516 9029
rect 51076 7286 51106 7666
rect 51486 7286 51516 7666
rect 51076 6091 51516 7286
rect 51076 6005 51169 6091
rect 51255 6005 51337 6091
rect 51423 6005 51516 6091
rect 51076 4579 51516 6005
rect 51076 4493 51169 4579
rect 51255 4493 51337 4579
rect 51423 4493 51516 4579
rect 51076 3666 51516 4493
rect 51076 3286 51106 3666
rect 51486 3286 51516 3666
rect 51076 3067 51516 3286
rect 51076 2981 51169 3067
rect 51255 2981 51337 3067
rect 51423 2981 51516 3067
rect 51076 1555 51516 2981
rect 51076 1469 51169 1555
rect 51255 1469 51337 1555
rect 51423 1469 51516 1555
rect 51076 712 51516 1469
rect 52316 38599 52756 38682
rect 52316 38513 52409 38599
rect 52495 38513 52577 38599
rect 52663 38513 52756 38599
rect 52316 37087 52756 38513
rect 52316 37001 52409 37087
rect 52495 37001 52577 37087
rect 52663 37001 52756 37087
rect 52316 36906 52756 37001
rect 52316 36526 52346 36906
rect 52726 36526 52756 36906
rect 52316 35575 52756 36526
rect 52316 35489 52409 35575
rect 52495 35489 52577 35575
rect 52663 35489 52756 35575
rect 52316 34063 52756 35489
rect 52316 33977 52409 34063
rect 52495 33977 52577 34063
rect 52663 33977 52756 34063
rect 52316 32906 52756 33977
rect 52316 32526 52346 32906
rect 52726 32526 52756 32906
rect 52316 32465 52409 32526
rect 52495 32465 52577 32526
rect 52663 32465 52756 32526
rect 52316 31039 52756 32465
rect 52316 30953 52409 31039
rect 52495 30953 52577 31039
rect 52663 30953 52756 31039
rect 52316 29527 52756 30953
rect 52316 29441 52409 29527
rect 52495 29441 52577 29527
rect 52663 29441 52756 29527
rect 52316 28906 52756 29441
rect 52316 28526 52346 28906
rect 52726 28526 52756 28906
rect 52316 28015 52756 28526
rect 52316 27929 52409 28015
rect 52495 27929 52577 28015
rect 52663 27929 52756 28015
rect 52316 26503 52756 27929
rect 52316 26417 52409 26503
rect 52495 26417 52577 26503
rect 52663 26417 52756 26503
rect 52316 24991 52756 26417
rect 52316 24906 52409 24991
rect 52495 24906 52577 24991
rect 52663 24906 52756 24991
rect 52316 24526 52346 24906
rect 52726 24526 52756 24906
rect 52316 23479 52756 24526
rect 52316 23393 52409 23479
rect 52495 23393 52577 23479
rect 52663 23393 52756 23479
rect 52316 21967 52756 23393
rect 52316 21881 52409 21967
rect 52495 21881 52577 21967
rect 52663 21881 52756 21967
rect 52316 20906 52756 21881
rect 52316 20526 52346 20906
rect 52726 20526 52756 20906
rect 52316 20455 52756 20526
rect 52316 20369 52409 20455
rect 52495 20369 52577 20455
rect 52663 20369 52756 20455
rect 52316 18943 52756 20369
rect 52316 18857 52409 18943
rect 52495 18857 52577 18943
rect 52663 18857 52756 18943
rect 52316 17431 52756 18857
rect 52316 17345 52409 17431
rect 52495 17345 52577 17431
rect 52663 17345 52756 17431
rect 52316 16906 52756 17345
rect 52316 16526 52346 16906
rect 52726 16526 52756 16906
rect 52316 15919 52756 16526
rect 52316 15833 52409 15919
rect 52495 15833 52577 15919
rect 52663 15833 52756 15919
rect 52316 14407 52756 15833
rect 52316 14321 52409 14407
rect 52495 14321 52577 14407
rect 52663 14321 52756 14407
rect 52316 12906 52756 14321
rect 52316 12526 52346 12906
rect 52726 12526 52756 12906
rect 52316 11383 52756 12526
rect 52316 11297 52409 11383
rect 52495 11297 52577 11383
rect 52663 11297 52756 11383
rect 52316 9871 52756 11297
rect 52316 9785 52409 9871
rect 52495 9785 52577 9871
rect 52663 9785 52756 9871
rect 52316 8906 52756 9785
rect 52316 8526 52346 8906
rect 52726 8526 52756 8906
rect 52316 8359 52756 8526
rect 52316 8273 52409 8359
rect 52495 8273 52577 8359
rect 52663 8273 52756 8359
rect 52316 6847 52756 8273
rect 52316 6761 52409 6847
rect 52495 6761 52577 6847
rect 52663 6761 52756 6847
rect 52316 5335 52756 6761
rect 52316 5249 52409 5335
rect 52495 5249 52577 5335
rect 52663 5249 52756 5335
rect 52316 4906 52756 5249
rect 52316 4526 52346 4906
rect 52726 4526 52756 4906
rect 52316 3823 52756 4526
rect 52316 3737 52409 3823
rect 52495 3737 52577 3823
rect 52663 3737 52756 3823
rect 52316 2311 52756 3737
rect 52316 2225 52409 2311
rect 52495 2225 52577 2311
rect 52663 2225 52756 2311
rect 52316 799 52756 2225
rect 52316 713 52409 799
rect 52495 713 52577 799
rect 52663 713 52756 799
rect 52316 630 52756 713
rect 55076 37843 55516 38600
rect 55076 37757 55169 37843
rect 55255 37757 55337 37843
rect 55423 37757 55516 37843
rect 55076 36331 55516 37757
rect 55076 36245 55169 36331
rect 55255 36245 55337 36331
rect 55423 36245 55516 36331
rect 55076 35666 55516 36245
rect 55076 35286 55106 35666
rect 55486 35286 55516 35666
rect 55076 34819 55516 35286
rect 55076 34733 55169 34819
rect 55255 34733 55337 34819
rect 55423 34733 55516 34819
rect 55076 33307 55516 34733
rect 55076 33221 55169 33307
rect 55255 33221 55337 33307
rect 55423 33221 55516 33307
rect 55076 31795 55516 33221
rect 55076 31709 55169 31795
rect 55255 31709 55337 31795
rect 55423 31709 55516 31795
rect 55076 31666 55516 31709
rect 55076 31286 55106 31666
rect 55486 31286 55516 31666
rect 55076 30283 55516 31286
rect 55076 30197 55169 30283
rect 55255 30197 55337 30283
rect 55423 30197 55516 30283
rect 55076 28771 55516 30197
rect 55076 28685 55169 28771
rect 55255 28685 55337 28771
rect 55423 28685 55516 28771
rect 55076 27666 55516 28685
rect 55076 27286 55106 27666
rect 55486 27286 55516 27666
rect 55076 27259 55516 27286
rect 55076 27173 55169 27259
rect 55255 27173 55337 27259
rect 55423 27173 55516 27259
rect 55076 25747 55516 27173
rect 55076 25661 55169 25747
rect 55255 25661 55337 25747
rect 55423 25661 55516 25747
rect 55076 24235 55516 25661
rect 55076 24149 55169 24235
rect 55255 24149 55337 24235
rect 55423 24149 55516 24235
rect 55076 23666 55516 24149
rect 55076 23286 55106 23666
rect 55486 23286 55516 23666
rect 55076 22723 55516 23286
rect 55076 22637 55169 22723
rect 55255 22637 55337 22723
rect 55423 22637 55516 22723
rect 55076 21211 55516 22637
rect 55076 21125 55169 21211
rect 55255 21125 55337 21211
rect 55423 21125 55516 21211
rect 55076 19699 55516 21125
rect 55076 19666 55169 19699
rect 55255 19666 55337 19699
rect 55423 19666 55516 19699
rect 55076 19286 55106 19666
rect 55486 19286 55516 19666
rect 55076 18187 55516 19286
rect 55076 18101 55169 18187
rect 55255 18101 55337 18187
rect 55423 18101 55516 18187
rect 55076 16675 55516 18101
rect 55076 16589 55169 16675
rect 55255 16589 55337 16675
rect 55423 16589 55516 16675
rect 55076 15666 55516 16589
rect 55076 15286 55106 15666
rect 55486 15286 55516 15666
rect 55076 15163 55516 15286
rect 55076 15077 55169 15163
rect 55255 15077 55337 15163
rect 55423 15077 55516 15163
rect 55076 13651 55516 15077
rect 55076 13565 55169 13651
rect 55255 13565 55337 13651
rect 55423 13565 55516 13651
rect 55076 12139 55516 13565
rect 55076 12053 55169 12139
rect 55255 12053 55337 12139
rect 55423 12053 55516 12139
rect 55076 11666 55516 12053
rect 55076 11286 55106 11666
rect 55486 11286 55516 11666
rect 55076 10627 55516 11286
rect 55076 10541 55169 10627
rect 55255 10541 55337 10627
rect 55423 10541 55516 10627
rect 55076 9115 55516 10541
rect 55076 9029 55169 9115
rect 55255 9029 55337 9115
rect 55423 9029 55516 9115
rect 55076 7666 55516 9029
rect 55076 7286 55106 7666
rect 55486 7286 55516 7666
rect 55076 6091 55516 7286
rect 55076 6005 55169 6091
rect 55255 6005 55337 6091
rect 55423 6005 55516 6091
rect 55076 4579 55516 6005
rect 55076 4493 55169 4579
rect 55255 4493 55337 4579
rect 55423 4493 55516 4579
rect 55076 3666 55516 4493
rect 55076 3286 55106 3666
rect 55486 3286 55516 3666
rect 55076 3067 55516 3286
rect 55076 2981 55169 3067
rect 55255 2981 55337 3067
rect 55423 2981 55516 3067
rect 55076 1555 55516 2981
rect 55076 1469 55169 1555
rect 55255 1469 55337 1555
rect 55423 1469 55516 1555
rect 55076 712 55516 1469
rect 56316 38599 56756 38682
rect 56316 38513 56409 38599
rect 56495 38513 56577 38599
rect 56663 38513 56756 38599
rect 56316 37087 56756 38513
rect 56316 37001 56409 37087
rect 56495 37001 56577 37087
rect 56663 37001 56756 37087
rect 56316 36906 56756 37001
rect 56316 36526 56346 36906
rect 56726 36526 56756 36906
rect 56316 35575 56756 36526
rect 56316 35489 56409 35575
rect 56495 35489 56577 35575
rect 56663 35489 56756 35575
rect 56316 34063 56756 35489
rect 56316 33977 56409 34063
rect 56495 33977 56577 34063
rect 56663 33977 56756 34063
rect 56316 32906 56756 33977
rect 56316 32526 56346 32906
rect 56726 32526 56756 32906
rect 56316 32465 56409 32526
rect 56495 32465 56577 32526
rect 56663 32465 56756 32526
rect 56316 31039 56756 32465
rect 56316 30953 56409 31039
rect 56495 30953 56577 31039
rect 56663 30953 56756 31039
rect 56316 29527 56756 30953
rect 56316 29441 56409 29527
rect 56495 29441 56577 29527
rect 56663 29441 56756 29527
rect 56316 28906 56756 29441
rect 56316 28526 56346 28906
rect 56726 28526 56756 28906
rect 56316 28015 56756 28526
rect 56316 27929 56409 28015
rect 56495 27929 56577 28015
rect 56663 27929 56756 28015
rect 56316 26503 56756 27929
rect 56316 26417 56409 26503
rect 56495 26417 56577 26503
rect 56663 26417 56756 26503
rect 56316 24991 56756 26417
rect 56316 24906 56409 24991
rect 56495 24906 56577 24991
rect 56663 24906 56756 24991
rect 56316 24526 56346 24906
rect 56726 24526 56756 24906
rect 56316 23479 56756 24526
rect 56316 23393 56409 23479
rect 56495 23393 56577 23479
rect 56663 23393 56756 23479
rect 56316 21967 56756 23393
rect 56316 21881 56409 21967
rect 56495 21881 56577 21967
rect 56663 21881 56756 21967
rect 56316 20906 56756 21881
rect 56316 20526 56346 20906
rect 56726 20526 56756 20906
rect 56316 20455 56756 20526
rect 56316 20369 56409 20455
rect 56495 20369 56577 20455
rect 56663 20369 56756 20455
rect 56316 18943 56756 20369
rect 56316 18857 56409 18943
rect 56495 18857 56577 18943
rect 56663 18857 56756 18943
rect 56316 17431 56756 18857
rect 56316 17345 56409 17431
rect 56495 17345 56577 17431
rect 56663 17345 56756 17431
rect 56316 16906 56756 17345
rect 56316 16526 56346 16906
rect 56726 16526 56756 16906
rect 56316 15919 56756 16526
rect 56316 15833 56409 15919
rect 56495 15833 56577 15919
rect 56663 15833 56756 15919
rect 56316 14407 56756 15833
rect 56316 14321 56409 14407
rect 56495 14321 56577 14407
rect 56663 14321 56756 14407
rect 56316 12906 56756 14321
rect 56316 12526 56346 12906
rect 56726 12526 56756 12906
rect 56316 11383 56756 12526
rect 56316 11297 56409 11383
rect 56495 11297 56577 11383
rect 56663 11297 56756 11383
rect 56316 9871 56756 11297
rect 56316 9785 56409 9871
rect 56495 9785 56577 9871
rect 56663 9785 56756 9871
rect 56316 8906 56756 9785
rect 56316 8526 56346 8906
rect 56726 8526 56756 8906
rect 56316 8359 56756 8526
rect 56316 8273 56409 8359
rect 56495 8273 56577 8359
rect 56663 8273 56756 8359
rect 56316 6847 56756 8273
rect 56316 6761 56409 6847
rect 56495 6761 56577 6847
rect 56663 6761 56756 6847
rect 56316 5335 56756 6761
rect 56316 5249 56409 5335
rect 56495 5249 56577 5335
rect 56663 5249 56756 5335
rect 56316 4906 56756 5249
rect 56316 4526 56346 4906
rect 56726 4526 56756 4906
rect 56316 3823 56756 4526
rect 56316 3737 56409 3823
rect 56495 3737 56577 3823
rect 56663 3737 56756 3823
rect 56316 2311 56756 3737
rect 56316 2225 56409 2311
rect 56495 2225 56577 2311
rect 56663 2225 56756 2311
rect 56316 799 56756 2225
rect 56316 713 56409 799
rect 56495 713 56577 799
rect 56663 713 56756 799
rect 56316 630 56756 713
rect 59076 37843 59516 38600
rect 59076 37757 59169 37843
rect 59255 37757 59337 37843
rect 59423 37757 59516 37843
rect 59076 36331 59516 37757
rect 59076 36245 59169 36331
rect 59255 36245 59337 36331
rect 59423 36245 59516 36331
rect 59076 35666 59516 36245
rect 59076 35286 59106 35666
rect 59486 35286 59516 35666
rect 59076 34819 59516 35286
rect 59076 34733 59169 34819
rect 59255 34733 59337 34819
rect 59423 34733 59516 34819
rect 59076 33307 59516 34733
rect 59076 33221 59169 33307
rect 59255 33221 59337 33307
rect 59423 33221 59516 33307
rect 59076 31795 59516 33221
rect 59076 31709 59169 31795
rect 59255 31709 59337 31795
rect 59423 31709 59516 31795
rect 59076 31666 59516 31709
rect 59076 31286 59106 31666
rect 59486 31286 59516 31666
rect 59076 30283 59516 31286
rect 59076 30197 59169 30283
rect 59255 30197 59337 30283
rect 59423 30197 59516 30283
rect 59076 28771 59516 30197
rect 59076 28685 59169 28771
rect 59255 28685 59337 28771
rect 59423 28685 59516 28771
rect 59076 27666 59516 28685
rect 59076 27286 59106 27666
rect 59486 27286 59516 27666
rect 59076 27259 59516 27286
rect 59076 27173 59169 27259
rect 59255 27173 59337 27259
rect 59423 27173 59516 27259
rect 59076 25747 59516 27173
rect 59076 25661 59169 25747
rect 59255 25661 59337 25747
rect 59423 25661 59516 25747
rect 59076 24235 59516 25661
rect 59076 24149 59169 24235
rect 59255 24149 59337 24235
rect 59423 24149 59516 24235
rect 59076 23666 59516 24149
rect 59076 23286 59106 23666
rect 59486 23286 59516 23666
rect 59076 22723 59516 23286
rect 59076 22637 59169 22723
rect 59255 22637 59337 22723
rect 59423 22637 59516 22723
rect 59076 21211 59516 22637
rect 59076 21125 59169 21211
rect 59255 21125 59337 21211
rect 59423 21125 59516 21211
rect 59076 19699 59516 21125
rect 59076 19666 59169 19699
rect 59255 19666 59337 19699
rect 59423 19666 59516 19699
rect 59076 19286 59106 19666
rect 59486 19286 59516 19666
rect 59076 18187 59516 19286
rect 59076 18101 59169 18187
rect 59255 18101 59337 18187
rect 59423 18101 59516 18187
rect 59076 16675 59516 18101
rect 59076 16589 59169 16675
rect 59255 16589 59337 16675
rect 59423 16589 59516 16675
rect 59076 15666 59516 16589
rect 59076 15286 59106 15666
rect 59486 15286 59516 15666
rect 59076 15163 59516 15286
rect 59076 15077 59169 15163
rect 59255 15077 59337 15163
rect 59423 15077 59516 15163
rect 59076 13651 59516 15077
rect 59076 13565 59169 13651
rect 59255 13565 59337 13651
rect 59423 13565 59516 13651
rect 59076 12139 59516 13565
rect 59076 12053 59169 12139
rect 59255 12053 59337 12139
rect 59423 12053 59516 12139
rect 59076 11666 59516 12053
rect 59076 11286 59106 11666
rect 59486 11286 59516 11666
rect 59076 10627 59516 11286
rect 59076 10541 59169 10627
rect 59255 10541 59337 10627
rect 59423 10541 59516 10627
rect 59076 9115 59516 10541
rect 59076 9029 59169 9115
rect 59255 9029 59337 9115
rect 59423 9029 59516 9115
rect 59076 7666 59516 9029
rect 59076 7286 59106 7666
rect 59486 7286 59516 7666
rect 59076 6091 59516 7286
rect 59076 6005 59169 6091
rect 59255 6005 59337 6091
rect 59423 6005 59516 6091
rect 59076 4579 59516 6005
rect 59076 4493 59169 4579
rect 59255 4493 59337 4579
rect 59423 4493 59516 4579
rect 59076 3666 59516 4493
rect 59076 3286 59106 3666
rect 59486 3286 59516 3666
rect 59076 3067 59516 3286
rect 59076 2981 59169 3067
rect 59255 2981 59337 3067
rect 59423 2981 59516 3067
rect 59076 1555 59516 2981
rect 59076 1469 59169 1555
rect 59255 1469 59337 1555
rect 59423 1469 59516 1555
rect 59076 712 59516 1469
rect 60316 38599 60756 38682
rect 60316 38513 60409 38599
rect 60495 38513 60577 38599
rect 60663 38513 60756 38599
rect 60316 37087 60756 38513
rect 60316 37001 60409 37087
rect 60495 37001 60577 37087
rect 60663 37001 60756 37087
rect 60316 36906 60756 37001
rect 60316 36526 60346 36906
rect 60726 36526 60756 36906
rect 60316 35575 60756 36526
rect 60316 35489 60409 35575
rect 60495 35489 60577 35575
rect 60663 35489 60756 35575
rect 60316 34063 60756 35489
rect 60316 33977 60409 34063
rect 60495 33977 60577 34063
rect 60663 33977 60756 34063
rect 60316 32906 60756 33977
rect 60316 32526 60346 32906
rect 60726 32526 60756 32906
rect 60316 32465 60409 32526
rect 60495 32465 60577 32526
rect 60663 32465 60756 32526
rect 60316 31039 60756 32465
rect 60316 30953 60409 31039
rect 60495 30953 60577 31039
rect 60663 30953 60756 31039
rect 60316 29527 60756 30953
rect 60316 29441 60409 29527
rect 60495 29441 60577 29527
rect 60663 29441 60756 29527
rect 60316 28906 60756 29441
rect 60316 28526 60346 28906
rect 60726 28526 60756 28906
rect 60316 28015 60756 28526
rect 60316 27929 60409 28015
rect 60495 27929 60577 28015
rect 60663 27929 60756 28015
rect 60316 26503 60756 27929
rect 60316 26417 60409 26503
rect 60495 26417 60577 26503
rect 60663 26417 60756 26503
rect 60316 24991 60756 26417
rect 60316 24906 60409 24991
rect 60495 24906 60577 24991
rect 60663 24906 60756 24991
rect 60316 24526 60346 24906
rect 60726 24526 60756 24906
rect 60316 23479 60756 24526
rect 60316 23393 60409 23479
rect 60495 23393 60577 23479
rect 60663 23393 60756 23479
rect 60316 21967 60756 23393
rect 60316 21881 60409 21967
rect 60495 21881 60577 21967
rect 60663 21881 60756 21967
rect 60316 20906 60756 21881
rect 60316 20526 60346 20906
rect 60726 20526 60756 20906
rect 60316 20455 60756 20526
rect 60316 20369 60409 20455
rect 60495 20369 60577 20455
rect 60663 20369 60756 20455
rect 60316 18943 60756 20369
rect 60316 18857 60409 18943
rect 60495 18857 60577 18943
rect 60663 18857 60756 18943
rect 60316 17431 60756 18857
rect 60316 17345 60409 17431
rect 60495 17345 60577 17431
rect 60663 17345 60756 17431
rect 60316 16906 60756 17345
rect 60316 16526 60346 16906
rect 60726 16526 60756 16906
rect 60316 15919 60756 16526
rect 60316 15833 60409 15919
rect 60495 15833 60577 15919
rect 60663 15833 60756 15919
rect 60316 14407 60756 15833
rect 60316 14321 60409 14407
rect 60495 14321 60577 14407
rect 60663 14321 60756 14407
rect 60316 12906 60756 14321
rect 60316 12526 60346 12906
rect 60726 12526 60756 12906
rect 60316 11383 60756 12526
rect 60316 11297 60409 11383
rect 60495 11297 60577 11383
rect 60663 11297 60756 11383
rect 60316 9871 60756 11297
rect 60316 9785 60409 9871
rect 60495 9785 60577 9871
rect 60663 9785 60756 9871
rect 60316 8906 60756 9785
rect 60316 8526 60346 8906
rect 60726 8526 60756 8906
rect 60316 8359 60756 8526
rect 60316 8273 60409 8359
rect 60495 8273 60577 8359
rect 60663 8273 60756 8359
rect 60316 6847 60756 8273
rect 60316 6761 60409 6847
rect 60495 6761 60577 6847
rect 60663 6761 60756 6847
rect 60316 5335 60756 6761
rect 60316 5249 60409 5335
rect 60495 5249 60577 5335
rect 60663 5249 60756 5335
rect 60316 4906 60756 5249
rect 60316 4526 60346 4906
rect 60726 4526 60756 4906
rect 60316 3823 60756 4526
rect 60316 3737 60409 3823
rect 60495 3737 60577 3823
rect 60663 3737 60756 3823
rect 60316 2311 60756 3737
rect 60316 2225 60409 2311
rect 60495 2225 60577 2311
rect 60663 2225 60756 2311
rect 60316 799 60756 2225
rect 60316 713 60409 799
rect 60495 713 60577 799
rect 60663 713 60756 799
rect 60316 630 60756 713
rect 63076 37843 63516 38600
rect 63076 37757 63169 37843
rect 63255 37757 63337 37843
rect 63423 37757 63516 37843
rect 63076 36331 63516 37757
rect 63076 36245 63169 36331
rect 63255 36245 63337 36331
rect 63423 36245 63516 36331
rect 63076 35666 63516 36245
rect 63076 35286 63106 35666
rect 63486 35286 63516 35666
rect 63076 34819 63516 35286
rect 63076 34733 63169 34819
rect 63255 34733 63337 34819
rect 63423 34733 63516 34819
rect 63076 33307 63516 34733
rect 63076 33221 63169 33307
rect 63255 33221 63337 33307
rect 63423 33221 63516 33307
rect 63076 31795 63516 33221
rect 63076 31709 63169 31795
rect 63255 31709 63337 31795
rect 63423 31709 63516 31795
rect 63076 31666 63516 31709
rect 63076 31286 63106 31666
rect 63486 31286 63516 31666
rect 63076 30283 63516 31286
rect 63076 30197 63169 30283
rect 63255 30197 63337 30283
rect 63423 30197 63516 30283
rect 63076 28771 63516 30197
rect 63076 28685 63169 28771
rect 63255 28685 63337 28771
rect 63423 28685 63516 28771
rect 63076 27666 63516 28685
rect 63076 27286 63106 27666
rect 63486 27286 63516 27666
rect 63076 27259 63516 27286
rect 63076 27173 63169 27259
rect 63255 27173 63337 27259
rect 63423 27173 63516 27259
rect 63076 25747 63516 27173
rect 63076 25661 63169 25747
rect 63255 25661 63337 25747
rect 63423 25661 63516 25747
rect 63076 24235 63516 25661
rect 63076 24149 63169 24235
rect 63255 24149 63337 24235
rect 63423 24149 63516 24235
rect 63076 23666 63516 24149
rect 63076 23286 63106 23666
rect 63486 23286 63516 23666
rect 63076 22723 63516 23286
rect 63076 22637 63169 22723
rect 63255 22637 63337 22723
rect 63423 22637 63516 22723
rect 63076 21211 63516 22637
rect 63076 21125 63169 21211
rect 63255 21125 63337 21211
rect 63423 21125 63516 21211
rect 63076 19699 63516 21125
rect 63076 19666 63169 19699
rect 63255 19666 63337 19699
rect 63423 19666 63516 19699
rect 63076 19286 63106 19666
rect 63486 19286 63516 19666
rect 63076 18187 63516 19286
rect 63076 18101 63169 18187
rect 63255 18101 63337 18187
rect 63423 18101 63516 18187
rect 63076 16675 63516 18101
rect 63076 16589 63169 16675
rect 63255 16589 63337 16675
rect 63423 16589 63516 16675
rect 63076 15666 63516 16589
rect 63076 15286 63106 15666
rect 63486 15286 63516 15666
rect 63076 15163 63516 15286
rect 63076 15077 63169 15163
rect 63255 15077 63337 15163
rect 63423 15077 63516 15163
rect 63076 13651 63516 15077
rect 63076 13565 63169 13651
rect 63255 13565 63337 13651
rect 63423 13565 63516 13651
rect 63076 12139 63516 13565
rect 63076 12053 63169 12139
rect 63255 12053 63337 12139
rect 63423 12053 63516 12139
rect 63076 11666 63516 12053
rect 63076 11286 63106 11666
rect 63486 11286 63516 11666
rect 63076 10627 63516 11286
rect 63076 10541 63169 10627
rect 63255 10541 63337 10627
rect 63423 10541 63516 10627
rect 63076 9115 63516 10541
rect 63076 9029 63169 9115
rect 63255 9029 63337 9115
rect 63423 9029 63516 9115
rect 63076 7666 63516 9029
rect 63076 7286 63106 7666
rect 63486 7286 63516 7666
rect 63076 6091 63516 7286
rect 63076 6005 63169 6091
rect 63255 6005 63337 6091
rect 63423 6005 63516 6091
rect 63076 4579 63516 6005
rect 63076 4493 63169 4579
rect 63255 4493 63337 4579
rect 63423 4493 63516 4579
rect 63076 3666 63516 4493
rect 63076 3286 63106 3666
rect 63486 3286 63516 3666
rect 63076 3067 63516 3286
rect 63076 2981 63169 3067
rect 63255 2981 63337 3067
rect 63423 2981 63516 3067
rect 63076 1555 63516 2981
rect 63076 1469 63169 1555
rect 63255 1469 63337 1555
rect 63423 1469 63516 1555
rect 63076 712 63516 1469
rect 64316 38599 64756 38682
rect 64316 38513 64409 38599
rect 64495 38513 64577 38599
rect 64663 38513 64756 38599
rect 64316 37087 64756 38513
rect 64316 37001 64409 37087
rect 64495 37001 64577 37087
rect 64663 37001 64756 37087
rect 64316 36906 64756 37001
rect 64316 36526 64346 36906
rect 64726 36526 64756 36906
rect 64316 35575 64756 36526
rect 64316 35489 64409 35575
rect 64495 35489 64577 35575
rect 64663 35489 64756 35575
rect 64316 34063 64756 35489
rect 64316 33977 64409 34063
rect 64495 33977 64577 34063
rect 64663 33977 64756 34063
rect 64316 32906 64756 33977
rect 64316 32526 64346 32906
rect 64726 32526 64756 32906
rect 64316 32465 64409 32526
rect 64495 32465 64577 32526
rect 64663 32465 64756 32526
rect 64316 31039 64756 32465
rect 64316 30953 64409 31039
rect 64495 30953 64577 31039
rect 64663 30953 64756 31039
rect 64316 29527 64756 30953
rect 64316 29441 64409 29527
rect 64495 29441 64577 29527
rect 64663 29441 64756 29527
rect 64316 28906 64756 29441
rect 64316 28526 64346 28906
rect 64726 28526 64756 28906
rect 64316 28015 64756 28526
rect 64316 27929 64409 28015
rect 64495 27929 64577 28015
rect 64663 27929 64756 28015
rect 64316 26503 64756 27929
rect 64316 26417 64409 26503
rect 64495 26417 64577 26503
rect 64663 26417 64756 26503
rect 64316 24991 64756 26417
rect 64316 24906 64409 24991
rect 64495 24906 64577 24991
rect 64663 24906 64756 24991
rect 64316 24526 64346 24906
rect 64726 24526 64756 24906
rect 64316 23479 64756 24526
rect 64316 23393 64409 23479
rect 64495 23393 64577 23479
rect 64663 23393 64756 23479
rect 64316 21967 64756 23393
rect 64316 21881 64409 21967
rect 64495 21881 64577 21967
rect 64663 21881 64756 21967
rect 64316 20906 64756 21881
rect 64316 20526 64346 20906
rect 64726 20526 64756 20906
rect 64316 20455 64756 20526
rect 64316 20369 64409 20455
rect 64495 20369 64577 20455
rect 64663 20369 64756 20455
rect 64316 18943 64756 20369
rect 64316 18857 64409 18943
rect 64495 18857 64577 18943
rect 64663 18857 64756 18943
rect 64316 17431 64756 18857
rect 64316 17345 64409 17431
rect 64495 17345 64577 17431
rect 64663 17345 64756 17431
rect 64316 16906 64756 17345
rect 64316 16526 64346 16906
rect 64726 16526 64756 16906
rect 64316 15919 64756 16526
rect 64316 15833 64409 15919
rect 64495 15833 64577 15919
rect 64663 15833 64756 15919
rect 64316 14407 64756 15833
rect 64316 14321 64409 14407
rect 64495 14321 64577 14407
rect 64663 14321 64756 14407
rect 64316 12906 64756 14321
rect 64316 12526 64346 12906
rect 64726 12526 64756 12906
rect 64316 11383 64756 12526
rect 64316 11297 64409 11383
rect 64495 11297 64577 11383
rect 64663 11297 64756 11383
rect 64316 9871 64756 11297
rect 64316 9785 64409 9871
rect 64495 9785 64577 9871
rect 64663 9785 64756 9871
rect 64316 8906 64756 9785
rect 64316 8526 64346 8906
rect 64726 8526 64756 8906
rect 64316 8359 64756 8526
rect 64316 8273 64409 8359
rect 64495 8273 64577 8359
rect 64663 8273 64756 8359
rect 64316 6847 64756 8273
rect 64316 6761 64409 6847
rect 64495 6761 64577 6847
rect 64663 6761 64756 6847
rect 64316 5335 64756 6761
rect 64316 5249 64409 5335
rect 64495 5249 64577 5335
rect 64663 5249 64756 5335
rect 64316 4906 64756 5249
rect 64316 4526 64346 4906
rect 64726 4526 64756 4906
rect 64316 3823 64756 4526
rect 64316 3737 64409 3823
rect 64495 3737 64577 3823
rect 64663 3737 64756 3823
rect 64316 2311 64756 3737
rect 64316 2225 64409 2311
rect 64495 2225 64577 2311
rect 64663 2225 64756 2311
rect 64316 799 64756 2225
rect 64316 713 64409 799
rect 64495 713 64577 799
rect 64663 713 64756 799
rect 64316 630 64756 713
rect 67076 37843 67516 38600
rect 67076 37757 67169 37843
rect 67255 37757 67337 37843
rect 67423 37757 67516 37843
rect 67076 36331 67516 37757
rect 67076 36245 67169 36331
rect 67255 36245 67337 36331
rect 67423 36245 67516 36331
rect 67076 35666 67516 36245
rect 67076 35286 67106 35666
rect 67486 35286 67516 35666
rect 67076 34819 67516 35286
rect 67076 34733 67169 34819
rect 67255 34733 67337 34819
rect 67423 34733 67516 34819
rect 67076 33307 67516 34733
rect 67076 33221 67169 33307
rect 67255 33221 67337 33307
rect 67423 33221 67516 33307
rect 67076 31795 67516 33221
rect 67076 31709 67169 31795
rect 67255 31709 67337 31795
rect 67423 31709 67516 31795
rect 67076 31666 67516 31709
rect 67076 31286 67106 31666
rect 67486 31286 67516 31666
rect 67076 30283 67516 31286
rect 67076 30197 67169 30283
rect 67255 30197 67337 30283
rect 67423 30197 67516 30283
rect 67076 28771 67516 30197
rect 67076 28685 67169 28771
rect 67255 28685 67337 28771
rect 67423 28685 67516 28771
rect 67076 27666 67516 28685
rect 67076 27286 67106 27666
rect 67486 27286 67516 27666
rect 67076 27259 67516 27286
rect 67076 27173 67169 27259
rect 67255 27173 67337 27259
rect 67423 27173 67516 27259
rect 67076 25747 67516 27173
rect 67076 25661 67169 25747
rect 67255 25661 67337 25747
rect 67423 25661 67516 25747
rect 67076 24235 67516 25661
rect 67076 24149 67169 24235
rect 67255 24149 67337 24235
rect 67423 24149 67516 24235
rect 67076 23666 67516 24149
rect 67076 23286 67106 23666
rect 67486 23286 67516 23666
rect 67076 22723 67516 23286
rect 67076 22637 67169 22723
rect 67255 22637 67337 22723
rect 67423 22637 67516 22723
rect 67076 21211 67516 22637
rect 67076 21125 67169 21211
rect 67255 21125 67337 21211
rect 67423 21125 67516 21211
rect 67076 19699 67516 21125
rect 67076 19666 67169 19699
rect 67255 19666 67337 19699
rect 67423 19666 67516 19699
rect 67076 19286 67106 19666
rect 67486 19286 67516 19666
rect 67076 18187 67516 19286
rect 67076 18101 67169 18187
rect 67255 18101 67337 18187
rect 67423 18101 67516 18187
rect 67076 16675 67516 18101
rect 67076 16589 67169 16675
rect 67255 16589 67337 16675
rect 67423 16589 67516 16675
rect 67076 15666 67516 16589
rect 67076 15286 67106 15666
rect 67486 15286 67516 15666
rect 67076 15163 67516 15286
rect 67076 15077 67169 15163
rect 67255 15077 67337 15163
rect 67423 15077 67516 15163
rect 67076 13651 67516 15077
rect 67076 13565 67169 13651
rect 67255 13565 67337 13651
rect 67423 13565 67516 13651
rect 67076 12139 67516 13565
rect 67076 12053 67169 12139
rect 67255 12053 67337 12139
rect 67423 12053 67516 12139
rect 67076 11666 67516 12053
rect 67076 11286 67106 11666
rect 67486 11286 67516 11666
rect 67076 10627 67516 11286
rect 67076 10541 67169 10627
rect 67255 10541 67337 10627
rect 67423 10541 67516 10627
rect 67076 9115 67516 10541
rect 67076 9029 67169 9115
rect 67255 9029 67337 9115
rect 67423 9029 67516 9115
rect 67076 7666 67516 9029
rect 67076 7286 67106 7666
rect 67486 7286 67516 7666
rect 67076 6091 67516 7286
rect 67076 6005 67169 6091
rect 67255 6005 67337 6091
rect 67423 6005 67516 6091
rect 67076 4579 67516 6005
rect 67076 4493 67169 4579
rect 67255 4493 67337 4579
rect 67423 4493 67516 4579
rect 67076 3666 67516 4493
rect 67076 3286 67106 3666
rect 67486 3286 67516 3666
rect 67076 3067 67516 3286
rect 67076 2981 67169 3067
rect 67255 2981 67337 3067
rect 67423 2981 67516 3067
rect 67076 1555 67516 2981
rect 67076 1469 67169 1555
rect 67255 1469 67337 1555
rect 67423 1469 67516 1555
rect 67076 712 67516 1469
rect 68316 38599 68756 38682
rect 68316 38513 68409 38599
rect 68495 38513 68577 38599
rect 68663 38513 68756 38599
rect 68316 37087 68756 38513
rect 68316 37001 68409 37087
rect 68495 37001 68577 37087
rect 68663 37001 68756 37087
rect 68316 36906 68756 37001
rect 68316 36526 68346 36906
rect 68726 36526 68756 36906
rect 68316 35575 68756 36526
rect 68316 35489 68409 35575
rect 68495 35489 68577 35575
rect 68663 35489 68756 35575
rect 68316 34063 68756 35489
rect 68316 33977 68409 34063
rect 68495 33977 68577 34063
rect 68663 33977 68756 34063
rect 68316 32906 68756 33977
rect 68316 32526 68346 32906
rect 68726 32526 68756 32906
rect 68316 32465 68409 32526
rect 68495 32465 68577 32526
rect 68663 32465 68756 32526
rect 68316 31039 68756 32465
rect 68316 30953 68409 31039
rect 68495 30953 68577 31039
rect 68663 30953 68756 31039
rect 68316 29527 68756 30953
rect 68316 29441 68409 29527
rect 68495 29441 68577 29527
rect 68663 29441 68756 29527
rect 68316 28906 68756 29441
rect 68316 28526 68346 28906
rect 68726 28526 68756 28906
rect 68316 28015 68756 28526
rect 68316 27929 68409 28015
rect 68495 27929 68577 28015
rect 68663 27929 68756 28015
rect 68316 26503 68756 27929
rect 68316 26417 68409 26503
rect 68495 26417 68577 26503
rect 68663 26417 68756 26503
rect 68316 24991 68756 26417
rect 68316 24906 68409 24991
rect 68495 24906 68577 24991
rect 68663 24906 68756 24991
rect 68316 24526 68346 24906
rect 68726 24526 68756 24906
rect 68316 23479 68756 24526
rect 68316 23393 68409 23479
rect 68495 23393 68577 23479
rect 68663 23393 68756 23479
rect 68316 21967 68756 23393
rect 68316 21881 68409 21967
rect 68495 21881 68577 21967
rect 68663 21881 68756 21967
rect 68316 20906 68756 21881
rect 68316 20526 68346 20906
rect 68726 20526 68756 20906
rect 68316 20455 68756 20526
rect 68316 20369 68409 20455
rect 68495 20369 68577 20455
rect 68663 20369 68756 20455
rect 68316 18943 68756 20369
rect 68316 18857 68409 18943
rect 68495 18857 68577 18943
rect 68663 18857 68756 18943
rect 68316 17431 68756 18857
rect 68316 17345 68409 17431
rect 68495 17345 68577 17431
rect 68663 17345 68756 17431
rect 68316 16906 68756 17345
rect 68316 16526 68346 16906
rect 68726 16526 68756 16906
rect 68316 15919 68756 16526
rect 68316 15833 68409 15919
rect 68495 15833 68577 15919
rect 68663 15833 68756 15919
rect 68316 14407 68756 15833
rect 68316 14321 68409 14407
rect 68495 14321 68577 14407
rect 68663 14321 68756 14407
rect 68316 12906 68756 14321
rect 68316 12526 68346 12906
rect 68726 12526 68756 12906
rect 68316 11383 68756 12526
rect 68316 11297 68409 11383
rect 68495 11297 68577 11383
rect 68663 11297 68756 11383
rect 68316 9871 68756 11297
rect 68316 9785 68409 9871
rect 68495 9785 68577 9871
rect 68663 9785 68756 9871
rect 68316 8906 68756 9785
rect 68316 8526 68346 8906
rect 68726 8526 68756 8906
rect 68316 8359 68756 8526
rect 68316 8273 68409 8359
rect 68495 8273 68577 8359
rect 68663 8273 68756 8359
rect 68316 6847 68756 8273
rect 68316 6761 68409 6847
rect 68495 6761 68577 6847
rect 68663 6761 68756 6847
rect 68316 5335 68756 6761
rect 68316 5249 68409 5335
rect 68495 5249 68577 5335
rect 68663 5249 68756 5335
rect 68316 4906 68756 5249
rect 68316 4526 68346 4906
rect 68726 4526 68756 4906
rect 68316 3823 68756 4526
rect 68316 3737 68409 3823
rect 68495 3737 68577 3823
rect 68663 3737 68756 3823
rect 68316 2311 68756 3737
rect 68316 2225 68409 2311
rect 68495 2225 68577 2311
rect 68663 2225 68756 2311
rect 68316 799 68756 2225
rect 68316 713 68409 799
rect 68495 713 68577 799
rect 68663 713 68756 799
rect 68316 630 68756 713
rect 71076 37843 71516 38600
rect 71076 37757 71169 37843
rect 71255 37757 71337 37843
rect 71423 37757 71516 37843
rect 71076 36331 71516 37757
rect 71076 36245 71169 36331
rect 71255 36245 71337 36331
rect 71423 36245 71516 36331
rect 71076 35666 71516 36245
rect 71076 35286 71106 35666
rect 71486 35286 71516 35666
rect 71076 34819 71516 35286
rect 71076 34733 71169 34819
rect 71255 34733 71337 34819
rect 71423 34733 71516 34819
rect 71076 31666 71516 34733
rect 71076 31286 71106 31666
rect 71486 31286 71516 31666
rect 71076 27666 71516 31286
rect 71076 27286 71106 27666
rect 71486 27286 71516 27666
rect 71076 24235 71516 27286
rect 71076 24149 71169 24235
rect 71255 24149 71337 24235
rect 71423 24149 71516 24235
rect 71076 23666 71516 24149
rect 71076 23286 71106 23666
rect 71486 23286 71516 23666
rect 71076 22723 71516 23286
rect 71076 22637 71169 22723
rect 71255 22637 71337 22723
rect 71423 22637 71516 22723
rect 71076 21211 71516 22637
rect 71076 21125 71169 21211
rect 71255 21125 71337 21211
rect 71423 21125 71516 21211
rect 71076 19699 71516 21125
rect 71076 19666 71169 19699
rect 71255 19666 71337 19699
rect 71423 19666 71516 19699
rect 71076 19286 71106 19666
rect 71486 19286 71516 19666
rect 71076 18187 71516 19286
rect 71076 18101 71169 18187
rect 71255 18101 71337 18187
rect 71423 18101 71516 18187
rect 71076 16675 71516 18101
rect 71076 16589 71169 16675
rect 71255 16589 71337 16675
rect 71423 16589 71516 16675
rect 71076 15666 71516 16589
rect 71076 15286 71106 15666
rect 71486 15286 71516 15666
rect 71076 11666 71516 15286
rect 71076 11286 71106 11666
rect 71486 11286 71516 11666
rect 71076 7666 71516 11286
rect 71076 7286 71106 7666
rect 71486 7286 71516 7666
rect 71076 4579 71516 7286
rect 71076 4493 71169 4579
rect 71255 4493 71337 4579
rect 71423 4493 71516 4579
rect 71076 3666 71516 4493
rect 71076 3286 71106 3666
rect 71486 3286 71516 3666
rect 71076 3067 71516 3286
rect 71076 2981 71169 3067
rect 71255 2981 71337 3067
rect 71423 2981 71516 3067
rect 71076 1555 71516 2981
rect 71076 1469 71169 1555
rect 71255 1469 71337 1555
rect 71423 1469 71516 1555
rect 71076 712 71516 1469
rect 72316 38599 72756 38682
rect 72316 38513 72409 38599
rect 72495 38513 72577 38599
rect 72663 38513 72756 38599
rect 72316 37087 72756 38513
rect 72316 37001 72409 37087
rect 72495 37001 72577 37087
rect 72663 37001 72756 37087
rect 72316 36906 72756 37001
rect 72316 36526 72346 36906
rect 72726 36526 72756 36906
rect 72316 35575 72756 36526
rect 72316 35489 72409 35575
rect 72495 35489 72577 35575
rect 72663 35489 72756 35575
rect 72316 32906 72756 35489
rect 75076 37843 75516 38600
rect 75076 37757 75169 37843
rect 75255 37757 75337 37843
rect 75423 37757 75516 37843
rect 75076 36331 75516 37757
rect 75076 36245 75169 36331
rect 75255 36245 75337 36331
rect 75423 36245 75516 36331
rect 75076 35666 75516 36245
rect 75076 35286 75106 35666
rect 75486 35286 75516 35666
rect 75076 34819 75516 35286
rect 75076 34733 75169 34819
rect 75255 34733 75337 34819
rect 75423 34733 75516 34819
rect 72316 32526 72346 32906
rect 72726 32526 72756 32906
rect 72316 31856 72756 32526
rect 72316 31770 72409 31856
rect 72495 31770 72577 31856
rect 72663 31770 72756 31856
rect 72316 31688 72756 31770
rect 72316 31602 72409 31688
rect 72495 31602 72577 31688
rect 72663 31602 72756 31688
rect 72316 31520 72756 31602
rect 72316 31434 72409 31520
rect 72495 31434 72577 31520
rect 72663 31434 72756 31520
rect 72316 31352 72756 31434
rect 72316 31266 72409 31352
rect 72495 31266 72577 31352
rect 72663 31266 72756 31352
rect 72316 31184 72756 31266
rect 72316 31098 72409 31184
rect 72495 31098 72577 31184
rect 72663 31098 72756 31184
rect 72316 31016 72756 31098
rect 72316 30930 72409 31016
rect 72495 30930 72577 31016
rect 72663 30930 72756 31016
rect 72316 30848 72756 30930
rect 72316 30762 72409 30848
rect 72495 30762 72577 30848
rect 72663 30762 72756 30848
rect 72316 30680 72756 30762
rect 72316 30594 72409 30680
rect 72495 30594 72577 30680
rect 72663 30594 72756 30680
rect 72316 30512 72756 30594
rect 72316 30426 72409 30512
rect 72495 30426 72577 30512
rect 72663 30426 72756 30512
rect 72316 30344 72756 30426
rect 72316 30258 72409 30344
rect 72495 30258 72577 30344
rect 72663 30258 72756 30344
rect 72316 30176 72756 30258
rect 72316 30090 72409 30176
rect 72495 30090 72577 30176
rect 72663 30090 72756 30176
rect 72316 30008 72756 30090
rect 72316 29922 72409 30008
rect 72495 29922 72577 30008
rect 72663 29922 72756 30008
rect 72316 29840 72756 29922
rect 72316 29754 72409 29840
rect 72495 29754 72577 29840
rect 72663 29754 72756 29840
rect 72316 28906 72756 29754
rect 72316 28526 72346 28906
rect 72726 28526 72756 28906
rect 72316 24906 72756 28526
rect 73124 32887 73452 33008
rect 73124 32801 73245 32887
rect 73331 32801 73452 32887
rect 73124 26587 73452 32801
rect 73124 26501 73245 26587
rect 73331 26501 73452 26587
rect 73124 26380 73452 26501
rect 75076 31666 75516 34733
rect 75076 31286 75106 31666
rect 75486 31286 75516 31666
rect 75076 28980 75516 31286
rect 75076 28894 75169 28980
rect 75255 28894 75337 28980
rect 75423 28894 75516 28980
rect 75076 28812 75516 28894
rect 75076 28726 75169 28812
rect 75255 28726 75337 28812
rect 75423 28726 75516 28812
rect 75076 28644 75516 28726
rect 75076 28558 75169 28644
rect 75255 28558 75337 28644
rect 75423 28558 75516 28644
rect 75076 28476 75516 28558
rect 75076 28390 75169 28476
rect 75255 28390 75337 28476
rect 75423 28390 75516 28476
rect 75076 28308 75516 28390
rect 75076 28222 75169 28308
rect 75255 28222 75337 28308
rect 75423 28222 75516 28308
rect 75076 28140 75516 28222
rect 75076 28054 75169 28140
rect 75255 28054 75337 28140
rect 75423 28054 75516 28140
rect 75076 27972 75516 28054
rect 75076 27886 75169 27972
rect 75255 27886 75337 27972
rect 75423 27886 75516 27972
rect 75076 27804 75516 27886
rect 75076 27718 75169 27804
rect 75255 27718 75337 27804
rect 75423 27718 75516 27804
rect 75076 27666 75516 27718
rect 75076 27286 75106 27666
rect 75486 27286 75516 27666
rect 75076 27214 75169 27286
rect 75255 27214 75337 27286
rect 75423 27214 75516 27286
rect 75076 27132 75516 27214
rect 75076 27046 75169 27132
rect 75255 27046 75337 27132
rect 75423 27046 75516 27132
rect 75076 26964 75516 27046
rect 75076 26878 75169 26964
rect 75255 26878 75337 26964
rect 75423 26878 75516 26964
rect 72316 24526 72346 24906
rect 72726 24526 72756 24906
rect 72316 23479 72756 24526
rect 72316 23393 72409 23479
rect 72495 23393 72577 23479
rect 72663 23393 72756 23479
rect 72316 21967 72756 23393
rect 72316 21881 72409 21967
rect 72495 21881 72577 21967
rect 72663 21881 72756 21967
rect 72316 20906 72756 21881
rect 72316 20526 72346 20906
rect 72726 20526 72756 20906
rect 72316 20455 72756 20526
rect 72316 20369 72409 20455
rect 72495 20369 72577 20455
rect 72663 20369 72756 20455
rect 72316 18943 72756 20369
rect 72316 18857 72409 18943
rect 72495 18857 72577 18943
rect 72663 18857 72756 18943
rect 72316 17431 72756 18857
rect 72316 17345 72409 17431
rect 72495 17345 72577 17431
rect 72663 17345 72756 17431
rect 72316 16906 72756 17345
rect 72316 16526 72346 16906
rect 72726 16526 72756 16906
rect 72316 15919 72756 16526
rect 72316 15833 72409 15919
rect 72495 15833 72577 15919
rect 72663 15833 72756 15919
rect 72316 13122 72756 15833
rect 72316 13036 72409 13122
rect 72495 13036 72577 13122
rect 72663 13036 72756 13122
rect 72316 12954 72756 13036
rect 72316 12906 72409 12954
rect 72495 12906 72577 12954
rect 72663 12906 72756 12954
rect 72316 12526 72346 12906
rect 72726 12526 72756 12906
rect 72316 12450 72756 12526
rect 72316 12364 72409 12450
rect 72495 12364 72577 12450
rect 72663 12364 72756 12450
rect 72316 12282 72756 12364
rect 72316 12196 72409 12282
rect 72495 12196 72577 12282
rect 72663 12196 72756 12282
rect 72316 12114 72756 12196
rect 72316 12028 72409 12114
rect 72495 12028 72577 12114
rect 72663 12028 72756 12114
rect 72316 11946 72756 12028
rect 72316 11860 72409 11946
rect 72495 11860 72577 11946
rect 72663 11860 72756 11946
rect 72316 11778 72756 11860
rect 72316 11692 72409 11778
rect 72495 11692 72577 11778
rect 72663 11692 72756 11778
rect 72316 11610 72756 11692
rect 72316 11524 72409 11610
rect 72495 11524 72577 11610
rect 72663 11524 72756 11610
rect 72316 11442 72756 11524
rect 72316 11356 72409 11442
rect 72495 11356 72577 11442
rect 72663 11356 72756 11442
rect 72316 11274 72756 11356
rect 72316 11188 72409 11274
rect 72495 11188 72577 11274
rect 72663 11188 72756 11274
rect 72316 11106 72756 11188
rect 72316 11020 72409 11106
rect 72495 11020 72577 11106
rect 72663 11020 72756 11106
rect 72316 8906 72756 11020
rect 72316 8526 72346 8906
rect 72726 8526 72756 8906
rect 72316 5335 72756 8526
rect 72316 5249 72409 5335
rect 72495 5249 72577 5335
rect 72663 5249 72756 5335
rect 72316 4906 72756 5249
rect 72316 4526 72346 4906
rect 72726 4526 72756 4906
rect 72316 3823 72756 4526
rect 72316 3737 72409 3823
rect 72495 3737 72577 3823
rect 72663 3737 72756 3823
rect 72316 2311 72756 3737
rect 72316 2225 72409 2311
rect 72495 2225 72577 2311
rect 72663 2225 72756 2311
rect 72316 799 72756 2225
rect 72316 713 72409 799
rect 72495 713 72577 799
rect 72663 713 72756 799
rect 72316 630 72756 713
rect 75076 24235 75516 26878
rect 75076 24149 75169 24235
rect 75255 24149 75337 24235
rect 75423 24149 75516 24235
rect 75076 23666 75516 24149
rect 75076 23286 75106 23666
rect 75486 23286 75516 23666
rect 75076 22723 75516 23286
rect 75076 22637 75169 22723
rect 75255 22637 75337 22723
rect 75423 22637 75516 22723
rect 75076 21211 75516 22637
rect 75076 21125 75169 21211
rect 75255 21125 75337 21211
rect 75423 21125 75516 21211
rect 75076 19699 75516 21125
rect 75076 19666 75169 19699
rect 75255 19666 75337 19699
rect 75423 19666 75516 19699
rect 75076 19286 75106 19666
rect 75486 19286 75516 19666
rect 75076 18187 75516 19286
rect 75076 18101 75169 18187
rect 75255 18101 75337 18187
rect 75423 18101 75516 18187
rect 75076 16675 75516 18101
rect 75076 16589 75169 16675
rect 75255 16589 75337 16675
rect 75423 16589 75516 16675
rect 75076 15666 75516 16589
rect 75076 15286 75106 15666
rect 75486 15286 75516 15666
rect 75076 11666 75516 15286
rect 75076 11286 75106 11666
rect 75486 11286 75516 11666
rect 75076 10246 75516 11286
rect 75076 10160 75169 10246
rect 75255 10160 75337 10246
rect 75423 10160 75516 10246
rect 75076 10078 75516 10160
rect 75076 9992 75169 10078
rect 75255 9992 75337 10078
rect 75423 9992 75516 10078
rect 75076 9910 75516 9992
rect 75076 9824 75169 9910
rect 75255 9824 75337 9910
rect 75423 9824 75516 9910
rect 75076 9742 75516 9824
rect 75076 9656 75169 9742
rect 75255 9656 75337 9742
rect 75423 9656 75516 9742
rect 75076 9574 75516 9656
rect 75076 9488 75169 9574
rect 75255 9488 75337 9574
rect 75423 9488 75516 9574
rect 75076 9406 75516 9488
rect 75076 9320 75169 9406
rect 75255 9320 75337 9406
rect 75423 9320 75516 9406
rect 75076 9238 75516 9320
rect 75076 9152 75169 9238
rect 75255 9152 75337 9238
rect 75423 9152 75516 9238
rect 75076 9070 75516 9152
rect 75076 8984 75169 9070
rect 75255 8984 75337 9070
rect 75423 8984 75516 9070
rect 75076 8902 75516 8984
rect 75076 8816 75169 8902
rect 75255 8816 75337 8902
rect 75423 8816 75516 8902
rect 75076 8734 75516 8816
rect 75076 8648 75169 8734
rect 75255 8648 75337 8734
rect 75423 8648 75516 8734
rect 75076 8566 75516 8648
rect 75076 8480 75169 8566
rect 75255 8480 75337 8566
rect 75423 8480 75516 8566
rect 75076 8398 75516 8480
rect 75076 8312 75169 8398
rect 75255 8312 75337 8398
rect 75423 8312 75516 8398
rect 75076 8230 75516 8312
rect 75076 8144 75169 8230
rect 75255 8144 75337 8230
rect 75423 8144 75516 8230
rect 75076 7666 75516 8144
rect 75076 7286 75106 7666
rect 75486 7286 75516 7666
rect 75076 4579 75516 7286
rect 75076 4493 75169 4579
rect 75255 4493 75337 4579
rect 75423 4493 75516 4579
rect 75076 3666 75516 4493
rect 75076 3286 75106 3666
rect 75486 3286 75516 3666
rect 75076 3067 75516 3286
rect 75076 2981 75169 3067
rect 75255 2981 75337 3067
rect 75423 2981 75516 3067
rect 75076 1555 75516 2981
rect 75076 1469 75169 1555
rect 75255 1469 75337 1555
rect 75423 1469 75516 1555
rect 75076 712 75516 1469
rect 76316 38599 76756 38682
rect 76316 38513 76409 38599
rect 76495 38513 76577 38599
rect 76663 38513 76756 38599
rect 76316 37087 76756 38513
rect 76316 37001 76409 37087
rect 76495 37001 76577 37087
rect 76663 37001 76756 37087
rect 76316 36906 76756 37001
rect 76316 36526 76346 36906
rect 76726 36526 76756 36906
rect 76316 35575 76756 36526
rect 76316 35489 76409 35575
rect 76495 35489 76577 35575
rect 76663 35489 76756 35575
rect 76316 32906 76756 35489
rect 76316 32526 76346 32906
rect 76726 32526 76756 32906
rect 76316 31856 76756 32526
rect 76316 31770 76409 31856
rect 76495 31770 76577 31856
rect 76663 31770 76756 31856
rect 76316 31688 76756 31770
rect 76316 31602 76409 31688
rect 76495 31602 76577 31688
rect 76663 31602 76756 31688
rect 76316 31520 76756 31602
rect 76316 31434 76409 31520
rect 76495 31434 76577 31520
rect 76663 31434 76756 31520
rect 76316 31352 76756 31434
rect 76316 31266 76409 31352
rect 76495 31266 76577 31352
rect 76663 31266 76756 31352
rect 76316 31184 76756 31266
rect 76316 31098 76409 31184
rect 76495 31098 76577 31184
rect 76663 31098 76756 31184
rect 76316 31016 76756 31098
rect 76316 30930 76409 31016
rect 76495 30930 76577 31016
rect 76663 30930 76756 31016
rect 76316 30848 76756 30930
rect 76316 30762 76409 30848
rect 76495 30762 76577 30848
rect 76663 30762 76756 30848
rect 76316 30680 76756 30762
rect 76316 30594 76409 30680
rect 76495 30594 76577 30680
rect 76663 30594 76756 30680
rect 76316 30512 76756 30594
rect 76316 30426 76409 30512
rect 76495 30426 76577 30512
rect 76663 30426 76756 30512
rect 76316 30344 76756 30426
rect 76316 30258 76409 30344
rect 76495 30258 76577 30344
rect 76663 30258 76756 30344
rect 76316 30176 76756 30258
rect 76316 30090 76409 30176
rect 76495 30090 76577 30176
rect 76663 30090 76756 30176
rect 76316 30008 76756 30090
rect 76316 29922 76409 30008
rect 76495 29922 76577 30008
rect 76663 29922 76756 30008
rect 76316 29840 76756 29922
rect 76316 29754 76409 29840
rect 76495 29754 76577 29840
rect 76663 29754 76756 29840
rect 76316 28906 76756 29754
rect 76316 28526 76346 28906
rect 76726 28526 76756 28906
rect 76316 24906 76756 28526
rect 76316 24526 76346 24906
rect 76726 24526 76756 24906
rect 76316 23479 76756 24526
rect 76316 23393 76409 23479
rect 76495 23393 76577 23479
rect 76663 23393 76756 23479
rect 76316 21967 76756 23393
rect 76316 21881 76409 21967
rect 76495 21881 76577 21967
rect 76663 21881 76756 21967
rect 76316 20906 76756 21881
rect 76316 20526 76346 20906
rect 76726 20526 76756 20906
rect 76316 20455 76756 20526
rect 76316 20369 76409 20455
rect 76495 20369 76577 20455
rect 76663 20369 76756 20455
rect 76316 18943 76756 20369
rect 76316 18857 76409 18943
rect 76495 18857 76577 18943
rect 76663 18857 76756 18943
rect 76316 17431 76756 18857
rect 76316 17345 76409 17431
rect 76495 17345 76577 17431
rect 76663 17345 76756 17431
rect 76316 16906 76756 17345
rect 76316 16526 76346 16906
rect 76726 16526 76756 16906
rect 76316 15919 76756 16526
rect 76316 15833 76409 15919
rect 76495 15833 76577 15919
rect 76663 15833 76756 15919
rect 76316 13122 76756 15833
rect 76316 13036 76409 13122
rect 76495 13036 76577 13122
rect 76663 13036 76756 13122
rect 76316 12954 76756 13036
rect 76316 12906 76409 12954
rect 76495 12906 76577 12954
rect 76663 12906 76756 12954
rect 76316 12526 76346 12906
rect 76726 12526 76756 12906
rect 76316 12450 76756 12526
rect 76316 12364 76409 12450
rect 76495 12364 76577 12450
rect 76663 12364 76756 12450
rect 76316 12282 76756 12364
rect 76316 12196 76409 12282
rect 76495 12196 76577 12282
rect 76663 12196 76756 12282
rect 76316 12114 76756 12196
rect 76316 12028 76409 12114
rect 76495 12028 76577 12114
rect 76663 12028 76756 12114
rect 76316 11946 76756 12028
rect 76316 11860 76409 11946
rect 76495 11860 76577 11946
rect 76663 11860 76756 11946
rect 76316 11778 76756 11860
rect 76316 11692 76409 11778
rect 76495 11692 76577 11778
rect 76663 11692 76756 11778
rect 76316 11610 76756 11692
rect 76316 11524 76409 11610
rect 76495 11524 76577 11610
rect 76663 11524 76756 11610
rect 76316 11442 76756 11524
rect 76316 11356 76409 11442
rect 76495 11356 76577 11442
rect 76663 11356 76756 11442
rect 76316 11274 76756 11356
rect 76316 11188 76409 11274
rect 76495 11188 76577 11274
rect 76663 11188 76756 11274
rect 76316 11106 76756 11188
rect 76316 11020 76409 11106
rect 76495 11020 76577 11106
rect 76663 11020 76756 11106
rect 76316 8906 76756 11020
rect 76316 8526 76346 8906
rect 76726 8526 76756 8906
rect 76316 5335 76756 8526
rect 76316 5249 76409 5335
rect 76495 5249 76577 5335
rect 76663 5249 76756 5335
rect 76316 4906 76756 5249
rect 76316 4526 76346 4906
rect 76726 4526 76756 4906
rect 76316 3823 76756 4526
rect 76316 3737 76409 3823
rect 76495 3737 76577 3823
rect 76663 3737 76756 3823
rect 76316 2311 76756 3737
rect 76316 2225 76409 2311
rect 76495 2225 76577 2311
rect 76663 2225 76756 2311
rect 76316 799 76756 2225
rect 76316 713 76409 799
rect 76495 713 76577 799
rect 76663 713 76756 799
rect 76316 630 76756 713
rect 79076 37843 79516 38600
rect 79076 37757 79169 37843
rect 79255 37757 79337 37843
rect 79423 37757 79516 37843
rect 79076 36331 79516 37757
rect 79076 36245 79169 36331
rect 79255 36245 79337 36331
rect 79423 36245 79516 36331
rect 79076 35666 79516 36245
rect 79076 35286 79106 35666
rect 79486 35286 79516 35666
rect 79076 34819 79516 35286
rect 79076 34733 79169 34819
rect 79255 34733 79337 34819
rect 79423 34733 79516 34819
rect 79076 31666 79516 34733
rect 79076 31286 79106 31666
rect 79486 31286 79516 31666
rect 79076 28980 79516 31286
rect 79076 28894 79169 28980
rect 79255 28894 79337 28980
rect 79423 28894 79516 28980
rect 79076 28812 79516 28894
rect 79076 28726 79169 28812
rect 79255 28726 79337 28812
rect 79423 28726 79516 28812
rect 79076 28644 79516 28726
rect 79076 28558 79169 28644
rect 79255 28558 79337 28644
rect 79423 28558 79516 28644
rect 79076 28476 79516 28558
rect 79076 28390 79169 28476
rect 79255 28390 79337 28476
rect 79423 28390 79516 28476
rect 79076 28308 79516 28390
rect 79076 28222 79169 28308
rect 79255 28222 79337 28308
rect 79423 28222 79516 28308
rect 79076 28140 79516 28222
rect 79076 28054 79169 28140
rect 79255 28054 79337 28140
rect 79423 28054 79516 28140
rect 79076 27972 79516 28054
rect 79076 27886 79169 27972
rect 79255 27886 79337 27972
rect 79423 27886 79516 27972
rect 79076 27804 79516 27886
rect 79076 27718 79169 27804
rect 79255 27718 79337 27804
rect 79423 27718 79516 27804
rect 79076 27666 79516 27718
rect 79076 27286 79106 27666
rect 79486 27286 79516 27666
rect 79076 27214 79169 27286
rect 79255 27214 79337 27286
rect 79423 27214 79516 27286
rect 79076 27132 79516 27214
rect 79076 27046 79169 27132
rect 79255 27046 79337 27132
rect 79423 27046 79516 27132
rect 79076 26964 79516 27046
rect 79076 26878 79169 26964
rect 79255 26878 79337 26964
rect 79423 26878 79516 26964
rect 79076 24235 79516 26878
rect 79076 24149 79169 24235
rect 79255 24149 79337 24235
rect 79423 24149 79516 24235
rect 79076 23666 79516 24149
rect 79076 23286 79106 23666
rect 79486 23286 79516 23666
rect 79076 22723 79516 23286
rect 79076 22637 79169 22723
rect 79255 22637 79337 22723
rect 79423 22637 79516 22723
rect 79076 21211 79516 22637
rect 79076 21125 79169 21211
rect 79255 21125 79337 21211
rect 79423 21125 79516 21211
rect 79076 19699 79516 21125
rect 79076 19666 79169 19699
rect 79255 19666 79337 19699
rect 79423 19666 79516 19699
rect 79076 19286 79106 19666
rect 79486 19286 79516 19666
rect 79076 18187 79516 19286
rect 79076 18101 79169 18187
rect 79255 18101 79337 18187
rect 79423 18101 79516 18187
rect 79076 16675 79516 18101
rect 79076 16589 79169 16675
rect 79255 16589 79337 16675
rect 79423 16589 79516 16675
rect 79076 15666 79516 16589
rect 79076 15286 79106 15666
rect 79486 15286 79516 15666
rect 79076 11666 79516 15286
rect 79076 11286 79106 11666
rect 79486 11286 79516 11666
rect 79076 10246 79516 11286
rect 79076 10160 79169 10246
rect 79255 10160 79337 10246
rect 79423 10160 79516 10246
rect 79076 10078 79516 10160
rect 79076 9992 79169 10078
rect 79255 9992 79337 10078
rect 79423 9992 79516 10078
rect 79076 9910 79516 9992
rect 79076 9824 79169 9910
rect 79255 9824 79337 9910
rect 79423 9824 79516 9910
rect 79076 9742 79516 9824
rect 79076 9656 79169 9742
rect 79255 9656 79337 9742
rect 79423 9656 79516 9742
rect 79076 9574 79516 9656
rect 79076 9488 79169 9574
rect 79255 9488 79337 9574
rect 79423 9488 79516 9574
rect 79076 9406 79516 9488
rect 79076 9320 79169 9406
rect 79255 9320 79337 9406
rect 79423 9320 79516 9406
rect 79076 9238 79516 9320
rect 79076 9152 79169 9238
rect 79255 9152 79337 9238
rect 79423 9152 79516 9238
rect 79076 9070 79516 9152
rect 79076 8984 79169 9070
rect 79255 8984 79337 9070
rect 79423 8984 79516 9070
rect 79076 8902 79516 8984
rect 79076 8816 79169 8902
rect 79255 8816 79337 8902
rect 79423 8816 79516 8902
rect 79076 8734 79516 8816
rect 79076 8648 79169 8734
rect 79255 8648 79337 8734
rect 79423 8648 79516 8734
rect 79076 8566 79516 8648
rect 79076 8480 79169 8566
rect 79255 8480 79337 8566
rect 79423 8480 79516 8566
rect 79076 8398 79516 8480
rect 79076 8312 79169 8398
rect 79255 8312 79337 8398
rect 79423 8312 79516 8398
rect 79076 8230 79516 8312
rect 79076 8144 79169 8230
rect 79255 8144 79337 8230
rect 79423 8144 79516 8230
rect 79076 7666 79516 8144
rect 79076 7286 79106 7666
rect 79486 7286 79516 7666
rect 79076 4579 79516 7286
rect 79076 4493 79169 4579
rect 79255 4493 79337 4579
rect 79423 4493 79516 4579
rect 79076 3666 79516 4493
rect 79076 3286 79106 3666
rect 79486 3286 79516 3666
rect 79076 3067 79516 3286
rect 79076 2981 79169 3067
rect 79255 2981 79337 3067
rect 79423 2981 79516 3067
rect 79076 1555 79516 2981
rect 79076 1469 79169 1555
rect 79255 1469 79337 1555
rect 79423 1469 79516 1555
rect 79076 712 79516 1469
rect 80316 38599 80756 38682
rect 80316 38513 80409 38599
rect 80495 38513 80577 38599
rect 80663 38513 80756 38599
rect 80316 37087 80756 38513
rect 80316 37001 80409 37087
rect 80495 37001 80577 37087
rect 80663 37001 80756 37087
rect 80316 36906 80756 37001
rect 80316 36526 80346 36906
rect 80726 36526 80756 36906
rect 80316 35575 80756 36526
rect 80316 35489 80409 35575
rect 80495 35489 80577 35575
rect 80663 35489 80756 35575
rect 80316 32906 80756 35489
rect 80316 32526 80346 32906
rect 80726 32526 80756 32906
rect 80316 31856 80756 32526
rect 80316 31770 80409 31856
rect 80495 31770 80577 31856
rect 80663 31770 80756 31856
rect 80316 31688 80756 31770
rect 80316 31602 80409 31688
rect 80495 31602 80577 31688
rect 80663 31602 80756 31688
rect 80316 31520 80756 31602
rect 80316 31434 80409 31520
rect 80495 31434 80577 31520
rect 80663 31434 80756 31520
rect 80316 31352 80756 31434
rect 80316 31266 80409 31352
rect 80495 31266 80577 31352
rect 80663 31266 80756 31352
rect 80316 31184 80756 31266
rect 80316 31098 80409 31184
rect 80495 31098 80577 31184
rect 80663 31098 80756 31184
rect 80316 31016 80756 31098
rect 80316 30930 80409 31016
rect 80495 30930 80577 31016
rect 80663 30930 80756 31016
rect 80316 30848 80756 30930
rect 80316 30762 80409 30848
rect 80495 30762 80577 30848
rect 80663 30762 80756 30848
rect 80316 30680 80756 30762
rect 80316 30594 80409 30680
rect 80495 30594 80577 30680
rect 80663 30594 80756 30680
rect 80316 30512 80756 30594
rect 80316 30426 80409 30512
rect 80495 30426 80577 30512
rect 80663 30426 80756 30512
rect 80316 30344 80756 30426
rect 80316 30258 80409 30344
rect 80495 30258 80577 30344
rect 80663 30258 80756 30344
rect 80316 30176 80756 30258
rect 80316 30090 80409 30176
rect 80495 30090 80577 30176
rect 80663 30090 80756 30176
rect 80316 30008 80756 30090
rect 80316 29922 80409 30008
rect 80495 29922 80577 30008
rect 80663 29922 80756 30008
rect 80316 29840 80756 29922
rect 80316 29754 80409 29840
rect 80495 29754 80577 29840
rect 80663 29754 80756 29840
rect 80316 28906 80756 29754
rect 80316 28526 80346 28906
rect 80726 28526 80756 28906
rect 80316 24906 80756 28526
rect 80316 24526 80346 24906
rect 80726 24526 80756 24906
rect 80316 23479 80756 24526
rect 80316 23393 80409 23479
rect 80495 23393 80577 23479
rect 80663 23393 80756 23479
rect 80316 21967 80756 23393
rect 80316 21881 80409 21967
rect 80495 21881 80577 21967
rect 80663 21881 80756 21967
rect 80316 20906 80756 21881
rect 80316 20526 80346 20906
rect 80726 20526 80756 20906
rect 80316 20455 80756 20526
rect 80316 20369 80409 20455
rect 80495 20369 80577 20455
rect 80663 20369 80756 20455
rect 80316 18943 80756 20369
rect 80316 18857 80409 18943
rect 80495 18857 80577 18943
rect 80663 18857 80756 18943
rect 80316 17431 80756 18857
rect 80316 17345 80409 17431
rect 80495 17345 80577 17431
rect 80663 17345 80756 17431
rect 80316 16906 80756 17345
rect 80316 16526 80346 16906
rect 80726 16526 80756 16906
rect 80316 15919 80756 16526
rect 80316 15833 80409 15919
rect 80495 15833 80577 15919
rect 80663 15833 80756 15919
rect 80316 13122 80756 15833
rect 80316 13036 80409 13122
rect 80495 13036 80577 13122
rect 80663 13036 80756 13122
rect 80316 12954 80756 13036
rect 80316 12906 80409 12954
rect 80495 12906 80577 12954
rect 80663 12906 80756 12954
rect 80316 12526 80346 12906
rect 80726 12526 80756 12906
rect 80316 12450 80756 12526
rect 80316 12364 80409 12450
rect 80495 12364 80577 12450
rect 80663 12364 80756 12450
rect 80316 12282 80756 12364
rect 80316 12196 80409 12282
rect 80495 12196 80577 12282
rect 80663 12196 80756 12282
rect 80316 12114 80756 12196
rect 80316 12028 80409 12114
rect 80495 12028 80577 12114
rect 80663 12028 80756 12114
rect 80316 11946 80756 12028
rect 80316 11860 80409 11946
rect 80495 11860 80577 11946
rect 80663 11860 80756 11946
rect 80316 11778 80756 11860
rect 80316 11692 80409 11778
rect 80495 11692 80577 11778
rect 80663 11692 80756 11778
rect 80316 11610 80756 11692
rect 80316 11524 80409 11610
rect 80495 11524 80577 11610
rect 80663 11524 80756 11610
rect 80316 11442 80756 11524
rect 80316 11356 80409 11442
rect 80495 11356 80577 11442
rect 80663 11356 80756 11442
rect 80316 11274 80756 11356
rect 80316 11188 80409 11274
rect 80495 11188 80577 11274
rect 80663 11188 80756 11274
rect 80316 11106 80756 11188
rect 80316 11020 80409 11106
rect 80495 11020 80577 11106
rect 80663 11020 80756 11106
rect 80316 8906 80756 11020
rect 80316 8526 80346 8906
rect 80726 8526 80756 8906
rect 80316 5335 80756 8526
rect 80316 5249 80409 5335
rect 80495 5249 80577 5335
rect 80663 5249 80756 5335
rect 80316 4906 80756 5249
rect 80316 4526 80346 4906
rect 80726 4526 80756 4906
rect 80316 3823 80756 4526
rect 80316 3737 80409 3823
rect 80495 3737 80577 3823
rect 80663 3737 80756 3823
rect 80316 2311 80756 3737
rect 80316 2225 80409 2311
rect 80495 2225 80577 2311
rect 80663 2225 80756 2311
rect 80316 799 80756 2225
rect 80316 713 80409 799
rect 80495 713 80577 799
rect 80663 713 80756 799
rect 80316 630 80756 713
rect 83076 37843 83516 38600
rect 83076 37757 83169 37843
rect 83255 37757 83337 37843
rect 83423 37757 83516 37843
rect 83076 36331 83516 37757
rect 83076 36245 83169 36331
rect 83255 36245 83337 36331
rect 83423 36245 83516 36331
rect 83076 35666 83516 36245
rect 83076 35286 83106 35666
rect 83486 35286 83516 35666
rect 83076 34819 83516 35286
rect 83076 34733 83169 34819
rect 83255 34733 83337 34819
rect 83423 34733 83516 34819
rect 83076 31666 83516 34733
rect 83076 31286 83106 31666
rect 83486 31286 83516 31666
rect 83076 28980 83516 31286
rect 83076 28894 83169 28980
rect 83255 28894 83337 28980
rect 83423 28894 83516 28980
rect 83076 28812 83516 28894
rect 83076 28726 83169 28812
rect 83255 28726 83337 28812
rect 83423 28726 83516 28812
rect 83076 28644 83516 28726
rect 83076 28558 83169 28644
rect 83255 28558 83337 28644
rect 83423 28558 83516 28644
rect 83076 28476 83516 28558
rect 83076 28390 83169 28476
rect 83255 28390 83337 28476
rect 83423 28390 83516 28476
rect 83076 28308 83516 28390
rect 83076 28222 83169 28308
rect 83255 28222 83337 28308
rect 83423 28222 83516 28308
rect 83076 28140 83516 28222
rect 83076 28054 83169 28140
rect 83255 28054 83337 28140
rect 83423 28054 83516 28140
rect 83076 27972 83516 28054
rect 83076 27886 83169 27972
rect 83255 27886 83337 27972
rect 83423 27886 83516 27972
rect 83076 27804 83516 27886
rect 83076 27718 83169 27804
rect 83255 27718 83337 27804
rect 83423 27718 83516 27804
rect 83076 27666 83516 27718
rect 83076 27286 83106 27666
rect 83486 27286 83516 27666
rect 83076 27214 83169 27286
rect 83255 27214 83337 27286
rect 83423 27214 83516 27286
rect 83076 27132 83516 27214
rect 83076 27046 83169 27132
rect 83255 27046 83337 27132
rect 83423 27046 83516 27132
rect 83076 26964 83516 27046
rect 83076 26878 83169 26964
rect 83255 26878 83337 26964
rect 83423 26878 83516 26964
rect 83076 24235 83516 26878
rect 83076 24149 83169 24235
rect 83255 24149 83337 24235
rect 83423 24149 83516 24235
rect 83076 23666 83516 24149
rect 83076 23286 83106 23666
rect 83486 23286 83516 23666
rect 83076 22723 83516 23286
rect 83076 22637 83169 22723
rect 83255 22637 83337 22723
rect 83423 22637 83516 22723
rect 83076 21211 83516 22637
rect 83076 21125 83169 21211
rect 83255 21125 83337 21211
rect 83423 21125 83516 21211
rect 83076 19699 83516 21125
rect 83076 19666 83169 19699
rect 83255 19666 83337 19699
rect 83423 19666 83516 19699
rect 83076 19286 83106 19666
rect 83486 19286 83516 19666
rect 83076 18187 83516 19286
rect 83076 18101 83169 18187
rect 83255 18101 83337 18187
rect 83423 18101 83516 18187
rect 83076 16675 83516 18101
rect 83076 16589 83169 16675
rect 83255 16589 83337 16675
rect 83423 16589 83516 16675
rect 83076 15666 83516 16589
rect 83076 15286 83106 15666
rect 83486 15286 83516 15666
rect 83076 11666 83516 15286
rect 83076 11286 83106 11666
rect 83486 11286 83516 11666
rect 83076 10246 83516 11286
rect 83076 10160 83169 10246
rect 83255 10160 83337 10246
rect 83423 10160 83516 10246
rect 83076 10078 83516 10160
rect 83076 9992 83169 10078
rect 83255 9992 83337 10078
rect 83423 9992 83516 10078
rect 83076 9910 83516 9992
rect 83076 9824 83169 9910
rect 83255 9824 83337 9910
rect 83423 9824 83516 9910
rect 83076 9742 83516 9824
rect 83076 9656 83169 9742
rect 83255 9656 83337 9742
rect 83423 9656 83516 9742
rect 83076 9574 83516 9656
rect 83076 9488 83169 9574
rect 83255 9488 83337 9574
rect 83423 9488 83516 9574
rect 83076 9406 83516 9488
rect 83076 9320 83169 9406
rect 83255 9320 83337 9406
rect 83423 9320 83516 9406
rect 83076 9238 83516 9320
rect 83076 9152 83169 9238
rect 83255 9152 83337 9238
rect 83423 9152 83516 9238
rect 83076 9070 83516 9152
rect 83076 8984 83169 9070
rect 83255 8984 83337 9070
rect 83423 8984 83516 9070
rect 83076 8902 83516 8984
rect 83076 8816 83169 8902
rect 83255 8816 83337 8902
rect 83423 8816 83516 8902
rect 83076 8734 83516 8816
rect 83076 8648 83169 8734
rect 83255 8648 83337 8734
rect 83423 8648 83516 8734
rect 83076 8566 83516 8648
rect 83076 8480 83169 8566
rect 83255 8480 83337 8566
rect 83423 8480 83516 8566
rect 83076 8398 83516 8480
rect 83076 8312 83169 8398
rect 83255 8312 83337 8398
rect 83423 8312 83516 8398
rect 83076 8230 83516 8312
rect 83076 8144 83169 8230
rect 83255 8144 83337 8230
rect 83423 8144 83516 8230
rect 83076 7666 83516 8144
rect 83076 7286 83106 7666
rect 83486 7286 83516 7666
rect 83076 4579 83516 7286
rect 83076 4493 83169 4579
rect 83255 4493 83337 4579
rect 83423 4493 83516 4579
rect 83076 3666 83516 4493
rect 83076 3286 83106 3666
rect 83486 3286 83516 3666
rect 83076 3067 83516 3286
rect 83076 2981 83169 3067
rect 83255 2981 83337 3067
rect 83423 2981 83516 3067
rect 83076 1555 83516 2981
rect 83076 1469 83169 1555
rect 83255 1469 83337 1555
rect 83423 1469 83516 1555
rect 83076 712 83516 1469
rect 84316 38599 84756 38682
rect 84316 38513 84409 38599
rect 84495 38513 84577 38599
rect 84663 38513 84756 38599
rect 84316 37087 84756 38513
rect 84316 37001 84409 37087
rect 84495 37001 84577 37087
rect 84663 37001 84756 37087
rect 84316 36906 84756 37001
rect 84316 36526 84346 36906
rect 84726 36526 84756 36906
rect 84316 35575 84756 36526
rect 84316 35489 84409 35575
rect 84495 35489 84577 35575
rect 84663 35489 84756 35575
rect 84316 32906 84756 35489
rect 87076 37843 87516 38600
rect 87076 37757 87169 37843
rect 87255 37757 87337 37843
rect 87423 37757 87516 37843
rect 87076 36331 87516 37757
rect 87076 36245 87169 36331
rect 87255 36245 87337 36331
rect 87423 36245 87516 36331
rect 87076 35666 87516 36245
rect 87076 35286 87106 35666
rect 87486 35286 87516 35666
rect 87076 34819 87516 35286
rect 87076 34733 87169 34819
rect 87255 34733 87337 34819
rect 87423 34733 87516 34819
rect 84316 32526 84346 32906
rect 84726 32526 84756 32906
rect 84316 31856 84756 32526
rect 84316 31770 84409 31856
rect 84495 31770 84577 31856
rect 84663 31770 84756 31856
rect 84316 31688 84756 31770
rect 84316 31602 84409 31688
rect 84495 31602 84577 31688
rect 84663 31602 84756 31688
rect 84316 31520 84756 31602
rect 84316 31434 84409 31520
rect 84495 31434 84577 31520
rect 84663 31434 84756 31520
rect 84316 31352 84756 31434
rect 84316 31266 84409 31352
rect 84495 31266 84577 31352
rect 84663 31266 84756 31352
rect 84316 31184 84756 31266
rect 84316 31098 84409 31184
rect 84495 31098 84577 31184
rect 84663 31098 84756 31184
rect 84316 31016 84756 31098
rect 84316 30930 84409 31016
rect 84495 30930 84577 31016
rect 84663 30930 84756 31016
rect 84316 30848 84756 30930
rect 84316 30762 84409 30848
rect 84495 30762 84577 30848
rect 84663 30762 84756 30848
rect 84316 30680 84756 30762
rect 84316 30594 84409 30680
rect 84495 30594 84577 30680
rect 84663 30594 84756 30680
rect 84316 30512 84756 30594
rect 84316 30426 84409 30512
rect 84495 30426 84577 30512
rect 84663 30426 84756 30512
rect 84316 30344 84756 30426
rect 84316 30258 84409 30344
rect 84495 30258 84577 30344
rect 84663 30258 84756 30344
rect 84316 30176 84756 30258
rect 84316 30090 84409 30176
rect 84495 30090 84577 30176
rect 84663 30090 84756 30176
rect 84316 30008 84756 30090
rect 84316 29922 84409 30008
rect 84495 29922 84577 30008
rect 84663 29922 84756 30008
rect 84316 29840 84756 29922
rect 84316 29754 84409 29840
rect 84495 29754 84577 29840
rect 84663 29754 84756 29840
rect 84316 28906 84756 29754
rect 84316 28526 84346 28906
rect 84726 28526 84756 28906
rect 84316 24906 84756 28526
rect 86348 33475 86676 33596
rect 86348 33389 86469 33475
rect 86555 33389 86676 33475
rect 86348 25411 86676 33389
rect 86348 25325 86469 25411
rect 86555 25325 86676 25411
rect 86348 25204 86676 25325
rect 87076 31666 87516 34733
rect 87076 31286 87106 31666
rect 87486 31286 87516 31666
rect 87076 28980 87516 31286
rect 87076 28894 87169 28980
rect 87255 28894 87337 28980
rect 87423 28894 87516 28980
rect 87076 28812 87516 28894
rect 87076 28726 87169 28812
rect 87255 28726 87337 28812
rect 87423 28726 87516 28812
rect 87076 28644 87516 28726
rect 87076 28558 87169 28644
rect 87255 28558 87337 28644
rect 87423 28558 87516 28644
rect 87076 28476 87516 28558
rect 87076 28390 87169 28476
rect 87255 28390 87337 28476
rect 87423 28390 87516 28476
rect 87076 28308 87516 28390
rect 87076 28222 87169 28308
rect 87255 28222 87337 28308
rect 87423 28222 87516 28308
rect 87076 28140 87516 28222
rect 87076 28054 87169 28140
rect 87255 28054 87337 28140
rect 87423 28054 87516 28140
rect 87076 27972 87516 28054
rect 87076 27886 87169 27972
rect 87255 27886 87337 27972
rect 87423 27886 87516 27972
rect 87076 27804 87516 27886
rect 87076 27718 87169 27804
rect 87255 27718 87337 27804
rect 87423 27718 87516 27804
rect 87076 27666 87516 27718
rect 87076 27286 87106 27666
rect 87486 27286 87516 27666
rect 87076 27214 87169 27286
rect 87255 27214 87337 27286
rect 87423 27214 87516 27286
rect 87076 27132 87516 27214
rect 87076 27046 87169 27132
rect 87255 27046 87337 27132
rect 87423 27046 87516 27132
rect 87076 26964 87516 27046
rect 87076 26878 87169 26964
rect 87255 26878 87337 26964
rect 87423 26878 87516 26964
rect 84316 24526 84346 24906
rect 84726 24526 84756 24906
rect 84316 23479 84756 24526
rect 84316 23393 84409 23479
rect 84495 23393 84577 23479
rect 84663 23393 84756 23479
rect 84316 21967 84756 23393
rect 84316 21881 84409 21967
rect 84495 21881 84577 21967
rect 84663 21881 84756 21967
rect 84316 20906 84756 21881
rect 84316 20526 84346 20906
rect 84726 20526 84756 20906
rect 84316 20455 84756 20526
rect 84316 20369 84409 20455
rect 84495 20369 84577 20455
rect 84663 20369 84756 20455
rect 84316 18943 84756 20369
rect 84316 18857 84409 18943
rect 84495 18857 84577 18943
rect 84663 18857 84756 18943
rect 84316 17431 84756 18857
rect 84316 17345 84409 17431
rect 84495 17345 84577 17431
rect 84663 17345 84756 17431
rect 84316 16906 84756 17345
rect 84316 16526 84346 16906
rect 84726 16526 84756 16906
rect 87076 24235 87516 26878
rect 87076 24149 87169 24235
rect 87255 24149 87337 24235
rect 87423 24149 87516 24235
rect 87076 23666 87516 24149
rect 87076 23286 87106 23666
rect 87486 23286 87516 23666
rect 87076 22723 87516 23286
rect 87076 22637 87169 22723
rect 87255 22637 87337 22723
rect 87423 22637 87516 22723
rect 87076 21211 87516 22637
rect 87076 21125 87169 21211
rect 87255 21125 87337 21211
rect 87423 21125 87516 21211
rect 87076 19699 87516 21125
rect 87076 19666 87169 19699
rect 87255 19666 87337 19699
rect 87423 19666 87516 19699
rect 87076 19286 87106 19666
rect 87486 19286 87516 19666
rect 87076 18187 87516 19286
rect 87076 18101 87169 18187
rect 87255 18101 87337 18187
rect 87423 18101 87516 18187
rect 87076 16675 87516 18101
rect 87076 16589 87169 16675
rect 87255 16589 87337 16675
rect 87423 16589 87516 16675
rect 84316 15919 84756 16526
rect 84316 15833 84409 15919
rect 84495 15833 84577 15919
rect 84663 15833 84756 15919
rect 84316 13122 84756 15833
rect 84316 13036 84409 13122
rect 84495 13036 84577 13122
rect 84663 13036 84756 13122
rect 84316 12954 84756 13036
rect 84316 12906 84409 12954
rect 84495 12906 84577 12954
rect 84663 12906 84756 12954
rect 84316 12526 84346 12906
rect 84726 12526 84756 12906
rect 84316 12450 84756 12526
rect 84316 12364 84409 12450
rect 84495 12364 84577 12450
rect 84663 12364 84756 12450
rect 84316 12282 84756 12364
rect 84316 12196 84409 12282
rect 84495 12196 84577 12282
rect 84663 12196 84756 12282
rect 84316 12114 84756 12196
rect 84316 12028 84409 12114
rect 84495 12028 84577 12114
rect 84663 12028 84756 12114
rect 84316 11946 84756 12028
rect 84316 11860 84409 11946
rect 84495 11860 84577 11946
rect 84663 11860 84756 11946
rect 84316 11778 84756 11860
rect 84316 11692 84409 11778
rect 84495 11692 84577 11778
rect 84663 11692 84756 11778
rect 84316 11610 84756 11692
rect 84316 11524 84409 11610
rect 84495 11524 84577 11610
rect 84663 11524 84756 11610
rect 84316 11442 84756 11524
rect 84316 11356 84409 11442
rect 84495 11356 84577 11442
rect 84663 11356 84756 11442
rect 84316 11274 84756 11356
rect 84316 11188 84409 11274
rect 84495 11188 84577 11274
rect 84663 11188 84756 11274
rect 84316 11106 84756 11188
rect 84316 11020 84409 11106
rect 84495 11020 84577 11106
rect 84663 11020 84756 11106
rect 84316 8906 84756 11020
rect 84316 8526 84346 8906
rect 84726 8526 84756 8906
rect 84316 5335 84756 8526
rect 86348 16423 86676 16544
rect 86348 16337 86469 16423
rect 86555 16337 86676 16423
rect 86348 7519 86676 16337
rect 86348 7433 86469 7519
rect 86555 7433 86676 7519
rect 86348 7312 86676 7433
rect 87076 15666 87516 16589
rect 87076 15286 87106 15666
rect 87486 15286 87516 15666
rect 87076 11666 87516 15286
rect 87076 11286 87106 11666
rect 87486 11286 87516 11666
rect 87076 10246 87516 11286
rect 87076 10160 87169 10246
rect 87255 10160 87337 10246
rect 87423 10160 87516 10246
rect 87076 10078 87516 10160
rect 87076 9992 87169 10078
rect 87255 9992 87337 10078
rect 87423 9992 87516 10078
rect 87076 9910 87516 9992
rect 87076 9824 87169 9910
rect 87255 9824 87337 9910
rect 87423 9824 87516 9910
rect 87076 9742 87516 9824
rect 87076 9656 87169 9742
rect 87255 9656 87337 9742
rect 87423 9656 87516 9742
rect 87076 9574 87516 9656
rect 87076 9488 87169 9574
rect 87255 9488 87337 9574
rect 87423 9488 87516 9574
rect 87076 9406 87516 9488
rect 87076 9320 87169 9406
rect 87255 9320 87337 9406
rect 87423 9320 87516 9406
rect 87076 9238 87516 9320
rect 87076 9152 87169 9238
rect 87255 9152 87337 9238
rect 87423 9152 87516 9238
rect 87076 9070 87516 9152
rect 87076 8984 87169 9070
rect 87255 8984 87337 9070
rect 87423 8984 87516 9070
rect 87076 8902 87516 8984
rect 87076 8816 87169 8902
rect 87255 8816 87337 8902
rect 87423 8816 87516 8902
rect 87076 8734 87516 8816
rect 87076 8648 87169 8734
rect 87255 8648 87337 8734
rect 87423 8648 87516 8734
rect 87076 8566 87516 8648
rect 87076 8480 87169 8566
rect 87255 8480 87337 8566
rect 87423 8480 87516 8566
rect 87076 8398 87516 8480
rect 87076 8312 87169 8398
rect 87255 8312 87337 8398
rect 87423 8312 87516 8398
rect 87076 8230 87516 8312
rect 87076 8144 87169 8230
rect 87255 8144 87337 8230
rect 87423 8144 87516 8230
rect 87076 7666 87516 8144
rect 84316 5249 84409 5335
rect 84495 5249 84577 5335
rect 84663 5249 84756 5335
rect 84316 4906 84756 5249
rect 84316 4526 84346 4906
rect 84726 4526 84756 4906
rect 84316 3823 84756 4526
rect 84316 3737 84409 3823
rect 84495 3737 84577 3823
rect 84663 3737 84756 3823
rect 84316 2311 84756 3737
rect 84316 2225 84409 2311
rect 84495 2225 84577 2311
rect 84663 2225 84756 2311
rect 84316 799 84756 2225
rect 84316 713 84409 799
rect 84495 713 84577 799
rect 84663 713 84756 799
rect 84316 630 84756 713
rect 87076 7286 87106 7666
rect 87486 7286 87516 7666
rect 87076 4579 87516 7286
rect 87076 4493 87169 4579
rect 87255 4493 87337 4579
rect 87423 4493 87516 4579
rect 87076 3666 87516 4493
rect 87076 3286 87106 3666
rect 87486 3286 87516 3666
rect 87076 3067 87516 3286
rect 87076 2981 87169 3067
rect 87255 2981 87337 3067
rect 87423 2981 87516 3067
rect 87076 1555 87516 2981
rect 87076 1469 87169 1555
rect 87255 1469 87337 1555
rect 87423 1469 87516 1555
rect 87076 712 87516 1469
rect 88316 38599 88756 38682
rect 88316 38513 88409 38599
rect 88495 38513 88577 38599
rect 88663 38513 88756 38599
rect 88316 37087 88756 38513
rect 88316 37001 88409 37087
rect 88495 37001 88577 37087
rect 88663 37001 88756 37087
rect 88316 36906 88756 37001
rect 88316 36526 88346 36906
rect 88726 36526 88756 36906
rect 88316 35575 88756 36526
rect 88316 35489 88409 35575
rect 88495 35489 88577 35575
rect 88663 35489 88756 35575
rect 88316 32906 88756 35489
rect 88316 32526 88346 32906
rect 88726 32526 88756 32906
rect 88316 31856 88756 32526
rect 88316 31770 88409 31856
rect 88495 31770 88577 31856
rect 88663 31770 88756 31856
rect 88316 31688 88756 31770
rect 88316 31602 88409 31688
rect 88495 31602 88577 31688
rect 88663 31602 88756 31688
rect 88316 31520 88756 31602
rect 88316 31434 88409 31520
rect 88495 31434 88577 31520
rect 88663 31434 88756 31520
rect 88316 31352 88756 31434
rect 88316 31266 88409 31352
rect 88495 31266 88577 31352
rect 88663 31266 88756 31352
rect 88316 31184 88756 31266
rect 88316 31098 88409 31184
rect 88495 31098 88577 31184
rect 88663 31098 88756 31184
rect 88316 31016 88756 31098
rect 88316 30930 88409 31016
rect 88495 30930 88577 31016
rect 88663 30930 88756 31016
rect 88316 30848 88756 30930
rect 88316 30762 88409 30848
rect 88495 30762 88577 30848
rect 88663 30762 88756 30848
rect 88316 30680 88756 30762
rect 88316 30594 88409 30680
rect 88495 30594 88577 30680
rect 88663 30594 88756 30680
rect 88316 30512 88756 30594
rect 88316 30426 88409 30512
rect 88495 30426 88577 30512
rect 88663 30426 88756 30512
rect 88316 30344 88756 30426
rect 88316 30258 88409 30344
rect 88495 30258 88577 30344
rect 88663 30258 88756 30344
rect 88316 30176 88756 30258
rect 88316 30090 88409 30176
rect 88495 30090 88577 30176
rect 88663 30090 88756 30176
rect 88316 30008 88756 30090
rect 88316 29922 88409 30008
rect 88495 29922 88577 30008
rect 88663 29922 88756 30008
rect 88316 29840 88756 29922
rect 88316 29754 88409 29840
rect 88495 29754 88577 29840
rect 88663 29754 88756 29840
rect 88316 28906 88756 29754
rect 88316 28526 88346 28906
rect 88726 28526 88756 28906
rect 88316 24906 88756 28526
rect 88316 24526 88346 24906
rect 88726 24526 88756 24906
rect 88316 23479 88756 24526
rect 88316 23393 88409 23479
rect 88495 23393 88577 23479
rect 88663 23393 88756 23479
rect 88316 21967 88756 23393
rect 88316 21881 88409 21967
rect 88495 21881 88577 21967
rect 88663 21881 88756 21967
rect 88316 20906 88756 21881
rect 88316 20526 88346 20906
rect 88726 20526 88756 20906
rect 88316 20455 88756 20526
rect 88316 20369 88409 20455
rect 88495 20369 88577 20455
rect 88663 20369 88756 20455
rect 88316 18943 88756 20369
rect 88316 18857 88409 18943
rect 88495 18857 88577 18943
rect 88663 18857 88756 18943
rect 88316 17431 88756 18857
rect 88316 17345 88409 17431
rect 88495 17345 88577 17431
rect 88663 17345 88756 17431
rect 88316 16906 88756 17345
rect 88316 16526 88346 16906
rect 88726 16526 88756 16906
rect 88316 15919 88756 16526
rect 88316 15833 88409 15919
rect 88495 15833 88577 15919
rect 88663 15833 88756 15919
rect 88316 13122 88756 15833
rect 88316 13036 88409 13122
rect 88495 13036 88577 13122
rect 88663 13036 88756 13122
rect 88316 12954 88756 13036
rect 88316 12906 88409 12954
rect 88495 12906 88577 12954
rect 88663 12906 88756 12954
rect 88316 12526 88346 12906
rect 88726 12526 88756 12906
rect 88316 12450 88756 12526
rect 88316 12364 88409 12450
rect 88495 12364 88577 12450
rect 88663 12364 88756 12450
rect 88316 12282 88756 12364
rect 88316 12196 88409 12282
rect 88495 12196 88577 12282
rect 88663 12196 88756 12282
rect 88316 12114 88756 12196
rect 88316 12028 88409 12114
rect 88495 12028 88577 12114
rect 88663 12028 88756 12114
rect 88316 11946 88756 12028
rect 88316 11860 88409 11946
rect 88495 11860 88577 11946
rect 88663 11860 88756 11946
rect 88316 11778 88756 11860
rect 88316 11692 88409 11778
rect 88495 11692 88577 11778
rect 88663 11692 88756 11778
rect 88316 11610 88756 11692
rect 88316 11524 88409 11610
rect 88495 11524 88577 11610
rect 88663 11524 88756 11610
rect 88316 11442 88756 11524
rect 88316 11356 88409 11442
rect 88495 11356 88577 11442
rect 88663 11356 88756 11442
rect 88316 11274 88756 11356
rect 88316 11188 88409 11274
rect 88495 11188 88577 11274
rect 88663 11188 88756 11274
rect 88316 11106 88756 11188
rect 88316 11020 88409 11106
rect 88495 11020 88577 11106
rect 88663 11020 88756 11106
rect 88316 8906 88756 11020
rect 88316 8526 88346 8906
rect 88726 8526 88756 8906
rect 88316 5335 88756 8526
rect 88316 5249 88409 5335
rect 88495 5249 88577 5335
rect 88663 5249 88756 5335
rect 88316 4906 88756 5249
rect 88316 4526 88346 4906
rect 88726 4526 88756 4906
rect 88316 3823 88756 4526
rect 88316 3737 88409 3823
rect 88495 3737 88577 3823
rect 88663 3737 88756 3823
rect 88316 2311 88756 3737
rect 88316 2225 88409 2311
rect 88495 2225 88577 2311
rect 88663 2225 88756 2311
rect 88316 799 88756 2225
rect 88316 713 88409 799
rect 88495 713 88577 799
rect 88663 713 88756 799
rect 88316 630 88756 713
rect 91076 37843 91516 38600
rect 91076 37757 91169 37843
rect 91255 37757 91337 37843
rect 91423 37757 91516 37843
rect 91076 36331 91516 37757
rect 91076 36245 91169 36331
rect 91255 36245 91337 36331
rect 91423 36245 91516 36331
rect 91076 35666 91516 36245
rect 91076 35286 91106 35666
rect 91486 35286 91516 35666
rect 91076 34819 91516 35286
rect 91076 34733 91169 34819
rect 91255 34733 91337 34819
rect 91423 34733 91516 34819
rect 91076 31666 91516 34733
rect 91076 31286 91106 31666
rect 91486 31286 91516 31666
rect 91076 28980 91516 31286
rect 91076 28894 91169 28980
rect 91255 28894 91337 28980
rect 91423 28894 91516 28980
rect 91076 28812 91516 28894
rect 91076 28726 91169 28812
rect 91255 28726 91337 28812
rect 91423 28726 91516 28812
rect 91076 28644 91516 28726
rect 91076 28558 91169 28644
rect 91255 28558 91337 28644
rect 91423 28558 91516 28644
rect 91076 28476 91516 28558
rect 91076 28390 91169 28476
rect 91255 28390 91337 28476
rect 91423 28390 91516 28476
rect 91076 28308 91516 28390
rect 91076 28222 91169 28308
rect 91255 28222 91337 28308
rect 91423 28222 91516 28308
rect 91076 28140 91516 28222
rect 91076 28054 91169 28140
rect 91255 28054 91337 28140
rect 91423 28054 91516 28140
rect 91076 27972 91516 28054
rect 91076 27886 91169 27972
rect 91255 27886 91337 27972
rect 91423 27886 91516 27972
rect 91076 27804 91516 27886
rect 91076 27718 91169 27804
rect 91255 27718 91337 27804
rect 91423 27718 91516 27804
rect 91076 27666 91516 27718
rect 91076 27286 91106 27666
rect 91486 27286 91516 27666
rect 91076 27214 91169 27286
rect 91255 27214 91337 27286
rect 91423 27214 91516 27286
rect 91076 27132 91516 27214
rect 91076 27046 91169 27132
rect 91255 27046 91337 27132
rect 91423 27046 91516 27132
rect 91076 26964 91516 27046
rect 91076 26878 91169 26964
rect 91255 26878 91337 26964
rect 91423 26878 91516 26964
rect 91076 24235 91516 26878
rect 91076 24149 91169 24235
rect 91255 24149 91337 24235
rect 91423 24149 91516 24235
rect 91076 23666 91516 24149
rect 91076 23286 91106 23666
rect 91486 23286 91516 23666
rect 91076 22723 91516 23286
rect 91076 22637 91169 22723
rect 91255 22637 91337 22723
rect 91423 22637 91516 22723
rect 91076 21211 91516 22637
rect 91076 21125 91169 21211
rect 91255 21125 91337 21211
rect 91423 21125 91516 21211
rect 91076 19699 91516 21125
rect 91076 19666 91169 19699
rect 91255 19666 91337 19699
rect 91423 19666 91516 19699
rect 91076 19286 91106 19666
rect 91486 19286 91516 19666
rect 91076 18187 91516 19286
rect 91076 18101 91169 18187
rect 91255 18101 91337 18187
rect 91423 18101 91516 18187
rect 91076 16675 91516 18101
rect 91076 16589 91169 16675
rect 91255 16589 91337 16675
rect 91423 16589 91516 16675
rect 91076 15666 91516 16589
rect 91076 15286 91106 15666
rect 91486 15286 91516 15666
rect 91076 11666 91516 15286
rect 91076 11286 91106 11666
rect 91486 11286 91516 11666
rect 91076 10246 91516 11286
rect 91076 10160 91169 10246
rect 91255 10160 91337 10246
rect 91423 10160 91516 10246
rect 91076 10078 91516 10160
rect 91076 9992 91169 10078
rect 91255 9992 91337 10078
rect 91423 9992 91516 10078
rect 91076 9910 91516 9992
rect 91076 9824 91169 9910
rect 91255 9824 91337 9910
rect 91423 9824 91516 9910
rect 91076 9742 91516 9824
rect 91076 9656 91169 9742
rect 91255 9656 91337 9742
rect 91423 9656 91516 9742
rect 91076 9574 91516 9656
rect 91076 9488 91169 9574
rect 91255 9488 91337 9574
rect 91423 9488 91516 9574
rect 91076 9406 91516 9488
rect 91076 9320 91169 9406
rect 91255 9320 91337 9406
rect 91423 9320 91516 9406
rect 91076 9238 91516 9320
rect 91076 9152 91169 9238
rect 91255 9152 91337 9238
rect 91423 9152 91516 9238
rect 91076 9070 91516 9152
rect 91076 8984 91169 9070
rect 91255 8984 91337 9070
rect 91423 8984 91516 9070
rect 91076 8902 91516 8984
rect 91076 8816 91169 8902
rect 91255 8816 91337 8902
rect 91423 8816 91516 8902
rect 91076 8734 91516 8816
rect 91076 8648 91169 8734
rect 91255 8648 91337 8734
rect 91423 8648 91516 8734
rect 91076 8566 91516 8648
rect 91076 8480 91169 8566
rect 91255 8480 91337 8566
rect 91423 8480 91516 8566
rect 91076 8398 91516 8480
rect 91076 8312 91169 8398
rect 91255 8312 91337 8398
rect 91423 8312 91516 8398
rect 91076 8230 91516 8312
rect 91076 8144 91169 8230
rect 91255 8144 91337 8230
rect 91423 8144 91516 8230
rect 91076 7666 91516 8144
rect 91076 7286 91106 7666
rect 91486 7286 91516 7666
rect 91076 4579 91516 7286
rect 91076 4493 91169 4579
rect 91255 4493 91337 4579
rect 91423 4493 91516 4579
rect 91076 3666 91516 4493
rect 91076 3286 91106 3666
rect 91486 3286 91516 3666
rect 91076 3067 91516 3286
rect 91076 2981 91169 3067
rect 91255 2981 91337 3067
rect 91423 2981 91516 3067
rect 91076 1555 91516 2981
rect 91076 1469 91169 1555
rect 91255 1469 91337 1555
rect 91423 1469 91516 1555
rect 91076 712 91516 1469
rect 92316 38599 92756 38682
rect 92316 38513 92409 38599
rect 92495 38513 92577 38599
rect 92663 38513 92756 38599
rect 92316 37087 92756 38513
rect 92316 37001 92409 37087
rect 92495 37001 92577 37087
rect 92663 37001 92756 37087
rect 92316 36906 92756 37001
rect 92316 36526 92346 36906
rect 92726 36526 92756 36906
rect 92316 35575 92756 36526
rect 92316 35489 92409 35575
rect 92495 35489 92577 35575
rect 92663 35489 92756 35575
rect 92316 32906 92756 35489
rect 92316 32526 92346 32906
rect 92726 32526 92756 32906
rect 92316 31856 92756 32526
rect 92316 31770 92409 31856
rect 92495 31770 92577 31856
rect 92663 31770 92756 31856
rect 92316 31688 92756 31770
rect 92316 31602 92409 31688
rect 92495 31602 92577 31688
rect 92663 31602 92756 31688
rect 92316 31520 92756 31602
rect 92316 31434 92409 31520
rect 92495 31434 92577 31520
rect 92663 31434 92756 31520
rect 92316 31352 92756 31434
rect 92316 31266 92409 31352
rect 92495 31266 92577 31352
rect 92663 31266 92756 31352
rect 92316 31184 92756 31266
rect 92316 31098 92409 31184
rect 92495 31098 92577 31184
rect 92663 31098 92756 31184
rect 92316 31016 92756 31098
rect 92316 30930 92409 31016
rect 92495 30930 92577 31016
rect 92663 30930 92756 31016
rect 92316 30848 92756 30930
rect 92316 30762 92409 30848
rect 92495 30762 92577 30848
rect 92663 30762 92756 30848
rect 92316 30680 92756 30762
rect 92316 30594 92409 30680
rect 92495 30594 92577 30680
rect 92663 30594 92756 30680
rect 92316 30512 92756 30594
rect 92316 30426 92409 30512
rect 92495 30426 92577 30512
rect 92663 30426 92756 30512
rect 92316 30344 92756 30426
rect 92316 30258 92409 30344
rect 92495 30258 92577 30344
rect 92663 30258 92756 30344
rect 92316 30176 92756 30258
rect 92316 30090 92409 30176
rect 92495 30090 92577 30176
rect 92663 30090 92756 30176
rect 92316 30008 92756 30090
rect 92316 29922 92409 30008
rect 92495 29922 92577 30008
rect 92663 29922 92756 30008
rect 92316 29840 92756 29922
rect 92316 29754 92409 29840
rect 92495 29754 92577 29840
rect 92663 29754 92756 29840
rect 92316 28906 92756 29754
rect 92316 28526 92346 28906
rect 92726 28526 92756 28906
rect 92316 24906 92756 28526
rect 92316 24526 92346 24906
rect 92726 24526 92756 24906
rect 92316 23479 92756 24526
rect 92316 23393 92409 23479
rect 92495 23393 92577 23479
rect 92663 23393 92756 23479
rect 92316 21967 92756 23393
rect 92316 21881 92409 21967
rect 92495 21881 92577 21967
rect 92663 21881 92756 21967
rect 92316 20906 92756 21881
rect 92316 20526 92346 20906
rect 92726 20526 92756 20906
rect 92316 20455 92756 20526
rect 92316 20369 92409 20455
rect 92495 20369 92577 20455
rect 92663 20369 92756 20455
rect 92316 18943 92756 20369
rect 92316 18857 92409 18943
rect 92495 18857 92577 18943
rect 92663 18857 92756 18943
rect 92316 17431 92756 18857
rect 92316 17345 92409 17431
rect 92495 17345 92577 17431
rect 92663 17345 92756 17431
rect 92316 16906 92756 17345
rect 92316 16526 92346 16906
rect 92726 16526 92756 16906
rect 92316 15919 92756 16526
rect 92316 15833 92409 15919
rect 92495 15833 92577 15919
rect 92663 15833 92756 15919
rect 92316 13122 92756 15833
rect 92316 13036 92409 13122
rect 92495 13036 92577 13122
rect 92663 13036 92756 13122
rect 92316 12954 92756 13036
rect 92316 12906 92409 12954
rect 92495 12906 92577 12954
rect 92663 12906 92756 12954
rect 92316 12526 92346 12906
rect 92726 12526 92756 12906
rect 92316 12450 92756 12526
rect 92316 12364 92409 12450
rect 92495 12364 92577 12450
rect 92663 12364 92756 12450
rect 92316 12282 92756 12364
rect 92316 12196 92409 12282
rect 92495 12196 92577 12282
rect 92663 12196 92756 12282
rect 92316 12114 92756 12196
rect 92316 12028 92409 12114
rect 92495 12028 92577 12114
rect 92663 12028 92756 12114
rect 92316 11946 92756 12028
rect 92316 11860 92409 11946
rect 92495 11860 92577 11946
rect 92663 11860 92756 11946
rect 92316 11778 92756 11860
rect 92316 11692 92409 11778
rect 92495 11692 92577 11778
rect 92663 11692 92756 11778
rect 92316 11610 92756 11692
rect 92316 11524 92409 11610
rect 92495 11524 92577 11610
rect 92663 11524 92756 11610
rect 92316 11442 92756 11524
rect 92316 11356 92409 11442
rect 92495 11356 92577 11442
rect 92663 11356 92756 11442
rect 92316 11274 92756 11356
rect 92316 11188 92409 11274
rect 92495 11188 92577 11274
rect 92663 11188 92756 11274
rect 92316 11106 92756 11188
rect 92316 11020 92409 11106
rect 92495 11020 92577 11106
rect 92663 11020 92756 11106
rect 92316 8906 92756 11020
rect 92316 8526 92346 8906
rect 92726 8526 92756 8906
rect 92316 5335 92756 8526
rect 92316 5249 92409 5335
rect 92495 5249 92577 5335
rect 92663 5249 92756 5335
rect 92316 4906 92756 5249
rect 92316 4526 92346 4906
rect 92726 4526 92756 4906
rect 92316 3823 92756 4526
rect 92316 3737 92409 3823
rect 92495 3737 92577 3823
rect 92663 3737 92756 3823
rect 92316 2311 92756 3737
rect 92316 2225 92409 2311
rect 92495 2225 92577 2311
rect 92663 2225 92756 2311
rect 92316 799 92756 2225
rect 92316 713 92409 799
rect 92495 713 92577 799
rect 92663 713 92756 799
rect 92316 630 92756 713
rect 95076 37843 95516 38600
rect 95076 37757 95169 37843
rect 95255 37757 95337 37843
rect 95423 37757 95516 37843
rect 95076 36331 95516 37757
rect 95076 36245 95169 36331
rect 95255 36245 95337 36331
rect 95423 36245 95516 36331
rect 95076 35666 95516 36245
rect 95076 35286 95106 35666
rect 95486 35286 95516 35666
rect 95076 34819 95516 35286
rect 95076 34733 95169 34819
rect 95255 34733 95337 34819
rect 95423 34733 95516 34819
rect 95076 31666 95516 34733
rect 95076 31286 95106 31666
rect 95486 31286 95516 31666
rect 95076 28980 95516 31286
rect 95076 28894 95169 28980
rect 95255 28894 95337 28980
rect 95423 28894 95516 28980
rect 95076 28812 95516 28894
rect 95076 28726 95169 28812
rect 95255 28726 95337 28812
rect 95423 28726 95516 28812
rect 95076 28644 95516 28726
rect 95076 28558 95169 28644
rect 95255 28558 95337 28644
rect 95423 28558 95516 28644
rect 95076 28476 95516 28558
rect 95076 28390 95169 28476
rect 95255 28390 95337 28476
rect 95423 28390 95516 28476
rect 95076 28308 95516 28390
rect 95076 28222 95169 28308
rect 95255 28222 95337 28308
rect 95423 28222 95516 28308
rect 95076 28140 95516 28222
rect 95076 28054 95169 28140
rect 95255 28054 95337 28140
rect 95423 28054 95516 28140
rect 95076 27972 95516 28054
rect 95076 27886 95169 27972
rect 95255 27886 95337 27972
rect 95423 27886 95516 27972
rect 95076 27804 95516 27886
rect 95076 27718 95169 27804
rect 95255 27718 95337 27804
rect 95423 27718 95516 27804
rect 95076 27666 95516 27718
rect 95076 27286 95106 27666
rect 95486 27286 95516 27666
rect 95076 27214 95169 27286
rect 95255 27214 95337 27286
rect 95423 27214 95516 27286
rect 95076 27132 95516 27214
rect 95076 27046 95169 27132
rect 95255 27046 95337 27132
rect 95423 27046 95516 27132
rect 95076 26964 95516 27046
rect 95076 26878 95169 26964
rect 95255 26878 95337 26964
rect 95423 26878 95516 26964
rect 95076 24235 95516 26878
rect 95076 24149 95169 24235
rect 95255 24149 95337 24235
rect 95423 24149 95516 24235
rect 95076 23666 95516 24149
rect 95076 23286 95106 23666
rect 95486 23286 95516 23666
rect 95076 22723 95516 23286
rect 95076 22637 95169 22723
rect 95255 22637 95337 22723
rect 95423 22637 95516 22723
rect 95076 21211 95516 22637
rect 95076 21125 95169 21211
rect 95255 21125 95337 21211
rect 95423 21125 95516 21211
rect 95076 19699 95516 21125
rect 95076 19666 95169 19699
rect 95255 19666 95337 19699
rect 95423 19666 95516 19699
rect 95076 19286 95106 19666
rect 95486 19286 95516 19666
rect 95076 18187 95516 19286
rect 95076 18101 95169 18187
rect 95255 18101 95337 18187
rect 95423 18101 95516 18187
rect 95076 16675 95516 18101
rect 95076 16589 95169 16675
rect 95255 16589 95337 16675
rect 95423 16589 95516 16675
rect 95076 15666 95516 16589
rect 95076 15286 95106 15666
rect 95486 15286 95516 15666
rect 95076 11666 95516 15286
rect 95076 11286 95106 11666
rect 95486 11286 95516 11666
rect 95076 10246 95516 11286
rect 95076 10160 95169 10246
rect 95255 10160 95337 10246
rect 95423 10160 95516 10246
rect 95076 10078 95516 10160
rect 95076 9992 95169 10078
rect 95255 9992 95337 10078
rect 95423 9992 95516 10078
rect 95076 9910 95516 9992
rect 95076 9824 95169 9910
rect 95255 9824 95337 9910
rect 95423 9824 95516 9910
rect 95076 9742 95516 9824
rect 95076 9656 95169 9742
rect 95255 9656 95337 9742
rect 95423 9656 95516 9742
rect 95076 9574 95516 9656
rect 95076 9488 95169 9574
rect 95255 9488 95337 9574
rect 95423 9488 95516 9574
rect 95076 9406 95516 9488
rect 95076 9320 95169 9406
rect 95255 9320 95337 9406
rect 95423 9320 95516 9406
rect 95076 9238 95516 9320
rect 95076 9152 95169 9238
rect 95255 9152 95337 9238
rect 95423 9152 95516 9238
rect 95076 9070 95516 9152
rect 95076 8984 95169 9070
rect 95255 8984 95337 9070
rect 95423 8984 95516 9070
rect 95076 8902 95516 8984
rect 95076 8816 95169 8902
rect 95255 8816 95337 8902
rect 95423 8816 95516 8902
rect 95076 8734 95516 8816
rect 95076 8648 95169 8734
rect 95255 8648 95337 8734
rect 95423 8648 95516 8734
rect 95076 8566 95516 8648
rect 95076 8480 95169 8566
rect 95255 8480 95337 8566
rect 95423 8480 95516 8566
rect 95076 8398 95516 8480
rect 95076 8312 95169 8398
rect 95255 8312 95337 8398
rect 95423 8312 95516 8398
rect 95076 8230 95516 8312
rect 95076 8144 95169 8230
rect 95255 8144 95337 8230
rect 95423 8144 95516 8230
rect 95076 7666 95516 8144
rect 95076 7286 95106 7666
rect 95486 7286 95516 7666
rect 95076 4579 95516 7286
rect 95076 4493 95169 4579
rect 95255 4493 95337 4579
rect 95423 4493 95516 4579
rect 95076 3666 95516 4493
rect 95076 3286 95106 3666
rect 95486 3286 95516 3666
rect 95076 3067 95516 3286
rect 95076 2981 95169 3067
rect 95255 2981 95337 3067
rect 95423 2981 95516 3067
rect 95076 1555 95516 2981
rect 95076 1469 95169 1555
rect 95255 1469 95337 1555
rect 95423 1469 95516 1555
rect 95076 712 95516 1469
rect 96316 38599 96756 38682
rect 96316 38513 96409 38599
rect 96495 38513 96577 38599
rect 96663 38513 96756 38599
rect 96316 37087 96756 38513
rect 96316 37001 96409 37087
rect 96495 37001 96577 37087
rect 96663 37001 96756 37087
rect 96316 36906 96756 37001
rect 96316 36526 96346 36906
rect 96726 36526 96756 36906
rect 96316 35575 96756 36526
rect 96316 35489 96409 35575
rect 96495 35489 96577 35575
rect 96663 35489 96756 35575
rect 96316 32906 96756 35489
rect 96316 32526 96346 32906
rect 96726 32526 96756 32906
rect 96316 31856 96756 32526
rect 96316 31770 96409 31856
rect 96495 31770 96577 31856
rect 96663 31770 96756 31856
rect 96316 31688 96756 31770
rect 96316 31602 96409 31688
rect 96495 31602 96577 31688
rect 96663 31602 96756 31688
rect 96316 31520 96756 31602
rect 96316 31434 96409 31520
rect 96495 31434 96577 31520
rect 96663 31434 96756 31520
rect 96316 31352 96756 31434
rect 96316 31266 96409 31352
rect 96495 31266 96577 31352
rect 96663 31266 96756 31352
rect 96316 31184 96756 31266
rect 96316 31098 96409 31184
rect 96495 31098 96577 31184
rect 96663 31098 96756 31184
rect 96316 31016 96756 31098
rect 96316 30930 96409 31016
rect 96495 30930 96577 31016
rect 96663 30930 96756 31016
rect 96316 30848 96756 30930
rect 96316 30762 96409 30848
rect 96495 30762 96577 30848
rect 96663 30762 96756 30848
rect 96316 30680 96756 30762
rect 96316 30594 96409 30680
rect 96495 30594 96577 30680
rect 96663 30594 96756 30680
rect 96316 30512 96756 30594
rect 96316 30426 96409 30512
rect 96495 30426 96577 30512
rect 96663 30426 96756 30512
rect 96316 30344 96756 30426
rect 96316 30258 96409 30344
rect 96495 30258 96577 30344
rect 96663 30258 96756 30344
rect 96316 30176 96756 30258
rect 96316 30090 96409 30176
rect 96495 30090 96577 30176
rect 96663 30090 96756 30176
rect 96316 30008 96756 30090
rect 96316 29922 96409 30008
rect 96495 29922 96577 30008
rect 96663 29922 96756 30008
rect 96316 29840 96756 29922
rect 96316 29754 96409 29840
rect 96495 29754 96577 29840
rect 96663 29754 96756 29840
rect 96316 28906 96756 29754
rect 96316 28526 96346 28906
rect 96726 28526 96756 28906
rect 96316 24906 96756 28526
rect 96316 24526 96346 24906
rect 96726 24526 96756 24906
rect 96316 23479 96756 24526
rect 96316 23393 96409 23479
rect 96495 23393 96577 23479
rect 96663 23393 96756 23479
rect 96316 21967 96756 23393
rect 96316 21881 96409 21967
rect 96495 21881 96577 21967
rect 96663 21881 96756 21967
rect 96316 20906 96756 21881
rect 96316 20526 96346 20906
rect 96726 20526 96756 20906
rect 96316 20455 96756 20526
rect 96316 20369 96409 20455
rect 96495 20369 96577 20455
rect 96663 20369 96756 20455
rect 96316 18943 96756 20369
rect 96316 18857 96409 18943
rect 96495 18857 96577 18943
rect 96663 18857 96756 18943
rect 96316 17431 96756 18857
rect 96316 17345 96409 17431
rect 96495 17345 96577 17431
rect 96663 17345 96756 17431
rect 96316 16906 96756 17345
rect 96316 16526 96346 16906
rect 96726 16526 96756 16906
rect 96316 15919 96756 16526
rect 96316 15833 96409 15919
rect 96495 15833 96577 15919
rect 96663 15833 96756 15919
rect 96316 13122 96756 15833
rect 96316 13036 96409 13122
rect 96495 13036 96577 13122
rect 96663 13036 96756 13122
rect 96316 12954 96756 13036
rect 96316 12906 96409 12954
rect 96495 12906 96577 12954
rect 96663 12906 96756 12954
rect 96316 12526 96346 12906
rect 96726 12526 96756 12906
rect 96316 12450 96756 12526
rect 96316 12364 96409 12450
rect 96495 12364 96577 12450
rect 96663 12364 96756 12450
rect 96316 12282 96756 12364
rect 96316 12196 96409 12282
rect 96495 12196 96577 12282
rect 96663 12196 96756 12282
rect 96316 12114 96756 12196
rect 96316 12028 96409 12114
rect 96495 12028 96577 12114
rect 96663 12028 96756 12114
rect 96316 11946 96756 12028
rect 96316 11860 96409 11946
rect 96495 11860 96577 11946
rect 96663 11860 96756 11946
rect 96316 11778 96756 11860
rect 96316 11692 96409 11778
rect 96495 11692 96577 11778
rect 96663 11692 96756 11778
rect 96316 11610 96756 11692
rect 96316 11524 96409 11610
rect 96495 11524 96577 11610
rect 96663 11524 96756 11610
rect 96316 11442 96756 11524
rect 96316 11356 96409 11442
rect 96495 11356 96577 11442
rect 96663 11356 96756 11442
rect 96316 11274 96756 11356
rect 96316 11188 96409 11274
rect 96495 11188 96577 11274
rect 96663 11188 96756 11274
rect 96316 11106 96756 11188
rect 96316 11020 96409 11106
rect 96495 11020 96577 11106
rect 96663 11020 96756 11106
rect 96316 8906 96756 11020
rect 96316 8526 96346 8906
rect 96726 8526 96756 8906
rect 96316 5335 96756 8526
rect 96316 5249 96409 5335
rect 96495 5249 96577 5335
rect 96663 5249 96756 5335
rect 96316 4906 96756 5249
rect 96316 4526 96346 4906
rect 96726 4526 96756 4906
rect 96316 3823 96756 4526
rect 96316 3737 96409 3823
rect 96495 3737 96577 3823
rect 96663 3737 96756 3823
rect 96316 2311 96756 3737
rect 96316 2225 96409 2311
rect 96495 2225 96577 2311
rect 96663 2225 96756 2311
rect 96316 799 96756 2225
rect 96316 713 96409 799
rect 96495 713 96577 799
rect 96663 713 96756 799
rect 96316 630 96756 713
rect 99076 37843 99516 38600
rect 99076 37757 99169 37843
rect 99255 37757 99337 37843
rect 99423 37757 99516 37843
rect 99076 36331 99516 37757
rect 99076 36245 99169 36331
rect 99255 36245 99337 36331
rect 99423 36245 99516 36331
rect 99076 35666 99516 36245
rect 99076 35286 99106 35666
rect 99486 35286 99516 35666
rect 99076 34819 99516 35286
rect 99076 34733 99169 34819
rect 99255 34733 99337 34819
rect 99423 34733 99516 34819
rect 99076 31666 99516 34733
rect 99076 31286 99106 31666
rect 99486 31286 99516 31666
rect 99076 27666 99516 31286
rect 99076 27286 99106 27666
rect 99486 27286 99516 27666
rect 99076 24235 99516 27286
rect 99076 24149 99169 24235
rect 99255 24149 99337 24235
rect 99423 24149 99516 24235
rect 99076 23666 99516 24149
rect 99076 23286 99106 23666
rect 99486 23286 99516 23666
rect 99076 22723 99516 23286
rect 99076 22637 99169 22723
rect 99255 22637 99337 22723
rect 99423 22637 99516 22723
rect 99076 21211 99516 22637
rect 99076 21125 99169 21211
rect 99255 21125 99337 21211
rect 99423 21125 99516 21211
rect 99076 19699 99516 21125
rect 99076 19666 99169 19699
rect 99255 19666 99337 19699
rect 99423 19666 99516 19699
rect 99076 19286 99106 19666
rect 99486 19286 99516 19666
rect 99076 18187 99516 19286
rect 99076 18101 99169 18187
rect 99255 18101 99337 18187
rect 99423 18101 99516 18187
rect 99076 16675 99516 18101
rect 99076 16589 99169 16675
rect 99255 16589 99337 16675
rect 99423 16589 99516 16675
rect 99076 15666 99516 16589
rect 99076 15286 99106 15666
rect 99486 15286 99516 15666
rect 99076 11666 99516 15286
rect 99076 11286 99106 11666
rect 99486 11286 99516 11666
rect 99076 7666 99516 11286
rect 99076 7286 99106 7666
rect 99486 7286 99516 7666
rect 99076 4579 99516 7286
rect 99076 4493 99169 4579
rect 99255 4493 99337 4579
rect 99423 4493 99516 4579
rect 99076 3666 99516 4493
rect 99076 3286 99106 3666
rect 99486 3286 99516 3666
rect 99076 3067 99516 3286
rect 99076 2981 99169 3067
rect 99255 2981 99337 3067
rect 99423 2981 99516 3067
rect 99076 1555 99516 2981
rect 99076 1469 99169 1555
rect 99255 1469 99337 1555
rect 99423 1469 99516 1555
rect 99076 712 99516 1469
<< via6 >>
rect 3106 35286 3486 35666
rect 3106 31286 3486 31666
rect 3106 27286 3486 27666
rect 3106 23286 3486 23666
rect 3106 19613 3169 19666
rect 3169 19613 3255 19666
rect 3255 19613 3337 19666
rect 3337 19613 3423 19666
rect 3423 19613 3486 19666
rect 3106 19286 3486 19613
rect 3106 15286 3486 15666
rect 3106 11286 3486 11666
rect 3106 7603 3486 7666
rect 3106 7517 3169 7603
rect 3169 7517 3255 7603
rect 3255 7517 3337 7603
rect 3337 7517 3423 7603
rect 3423 7517 3486 7603
rect 3106 7286 3486 7517
rect 3106 3286 3486 3666
rect 4346 36526 4726 36906
rect 4346 32551 4726 32906
rect 4346 32526 4409 32551
rect 4409 32526 4495 32551
rect 4495 32526 4577 32551
rect 4577 32526 4663 32551
rect 4663 32526 4726 32551
rect 4346 28526 4726 28906
rect 4346 24905 4409 24906
rect 4409 24905 4495 24906
rect 4495 24905 4577 24906
rect 4577 24905 4663 24906
rect 4663 24905 4726 24906
rect 4346 24526 4726 24905
rect 4346 20526 4726 20906
rect 4346 16526 4726 16906
rect 4346 12895 4726 12906
rect 4346 12809 4409 12895
rect 4409 12809 4495 12895
rect 4495 12809 4577 12895
rect 4577 12809 4663 12895
rect 4663 12809 4726 12895
rect 4346 12526 4726 12809
rect 4346 8526 4726 8906
rect 4346 4526 4726 4906
rect 7106 35286 7486 35666
rect 7106 31286 7486 31666
rect 7106 27286 7486 27666
rect 7106 23286 7486 23666
rect 7106 19613 7169 19666
rect 7169 19613 7255 19666
rect 7255 19613 7337 19666
rect 7337 19613 7423 19666
rect 7423 19613 7486 19666
rect 7106 19286 7486 19613
rect 7106 15286 7486 15666
rect 7106 11286 7486 11666
rect 7106 7603 7486 7666
rect 7106 7517 7169 7603
rect 7169 7517 7255 7603
rect 7255 7517 7337 7603
rect 7337 7517 7423 7603
rect 7423 7517 7486 7603
rect 7106 7286 7486 7517
rect 7106 3286 7486 3666
rect 8346 36526 8726 36906
rect 8346 32551 8726 32906
rect 8346 32526 8409 32551
rect 8409 32526 8495 32551
rect 8495 32526 8577 32551
rect 8577 32526 8663 32551
rect 8663 32526 8726 32551
rect 8346 28526 8726 28906
rect 8346 24905 8409 24906
rect 8409 24905 8495 24906
rect 8495 24905 8577 24906
rect 8577 24905 8663 24906
rect 8663 24905 8726 24906
rect 8346 24526 8726 24905
rect 8346 20526 8726 20906
rect 8346 16526 8726 16906
rect 8346 12895 8726 12906
rect 8346 12809 8409 12895
rect 8409 12809 8495 12895
rect 8495 12809 8577 12895
rect 8577 12809 8663 12895
rect 8663 12809 8726 12895
rect 8346 12526 8726 12809
rect 8346 8526 8726 8906
rect 8346 4526 8726 4906
rect 11106 35286 11486 35666
rect 11106 31286 11486 31666
rect 11106 27286 11486 27666
rect 11106 23286 11486 23666
rect 11106 19613 11169 19666
rect 11169 19613 11255 19666
rect 11255 19613 11337 19666
rect 11337 19613 11423 19666
rect 11423 19613 11486 19666
rect 11106 19286 11486 19613
rect 11106 15286 11486 15666
rect 11106 11286 11486 11666
rect 11106 7603 11486 7666
rect 11106 7517 11169 7603
rect 11169 7517 11255 7603
rect 11255 7517 11337 7603
rect 11337 7517 11423 7603
rect 11423 7517 11486 7603
rect 11106 7286 11486 7517
rect 11106 3286 11486 3666
rect 12346 36526 12726 36906
rect 12346 32551 12726 32906
rect 12346 32526 12409 32551
rect 12409 32526 12495 32551
rect 12495 32526 12577 32551
rect 12577 32526 12663 32551
rect 12663 32526 12726 32551
rect 12346 28526 12726 28906
rect 12346 24905 12409 24906
rect 12409 24905 12495 24906
rect 12495 24905 12577 24906
rect 12577 24905 12663 24906
rect 12663 24905 12726 24906
rect 12346 24526 12726 24905
rect 12346 20526 12726 20906
rect 12346 16526 12726 16906
rect 12346 12895 12726 12906
rect 12346 12809 12409 12895
rect 12409 12809 12495 12895
rect 12495 12809 12577 12895
rect 12577 12809 12663 12895
rect 12663 12809 12726 12895
rect 12346 12526 12726 12809
rect 12346 8526 12726 8906
rect 12346 4526 12726 4906
rect 15106 35286 15486 35666
rect 15106 31286 15486 31666
rect 15106 27286 15486 27666
rect 15106 23286 15486 23666
rect 15106 19613 15169 19666
rect 15169 19613 15255 19666
rect 15255 19613 15337 19666
rect 15337 19613 15423 19666
rect 15423 19613 15486 19666
rect 15106 19286 15486 19613
rect 15106 15286 15486 15666
rect 15106 11286 15486 11666
rect 15106 7603 15486 7666
rect 15106 7517 15169 7603
rect 15169 7517 15255 7603
rect 15255 7517 15337 7603
rect 15337 7517 15423 7603
rect 15423 7517 15486 7603
rect 15106 7286 15486 7517
rect 15106 3286 15486 3666
rect 16346 36526 16726 36906
rect 16346 32551 16726 32906
rect 16346 32526 16409 32551
rect 16409 32526 16495 32551
rect 16495 32526 16577 32551
rect 16577 32526 16663 32551
rect 16663 32526 16726 32551
rect 16346 28526 16726 28906
rect 16346 24905 16409 24906
rect 16409 24905 16495 24906
rect 16495 24905 16577 24906
rect 16577 24905 16663 24906
rect 16663 24905 16726 24906
rect 16346 24526 16726 24905
rect 16346 20526 16726 20906
rect 16346 16526 16726 16906
rect 16346 12895 16726 12906
rect 16346 12809 16409 12895
rect 16409 12809 16495 12895
rect 16495 12809 16577 12895
rect 16577 12809 16663 12895
rect 16663 12809 16726 12895
rect 16346 12526 16726 12809
rect 16346 8526 16726 8906
rect 16346 4526 16726 4906
rect 19106 35286 19486 35666
rect 19106 31286 19486 31666
rect 19106 27286 19486 27666
rect 19106 23286 19486 23666
rect 19106 19613 19169 19666
rect 19169 19613 19255 19666
rect 19255 19613 19337 19666
rect 19337 19613 19423 19666
rect 19423 19613 19486 19666
rect 19106 19286 19486 19613
rect 19106 15286 19486 15666
rect 19106 11286 19486 11666
rect 19106 7603 19486 7666
rect 19106 7517 19169 7603
rect 19169 7517 19255 7603
rect 19255 7517 19337 7603
rect 19337 7517 19423 7603
rect 19423 7517 19486 7603
rect 19106 7286 19486 7517
rect 19106 3286 19486 3666
rect 20346 36526 20726 36906
rect 20346 32551 20726 32906
rect 20346 32526 20409 32551
rect 20409 32526 20495 32551
rect 20495 32526 20577 32551
rect 20577 32526 20663 32551
rect 20663 32526 20726 32551
rect 20346 28526 20726 28906
rect 20346 24905 20409 24906
rect 20409 24905 20495 24906
rect 20495 24905 20577 24906
rect 20577 24905 20663 24906
rect 20663 24905 20726 24906
rect 20346 24526 20726 24905
rect 20346 20526 20726 20906
rect 20346 16526 20726 16906
rect 20346 12895 20726 12906
rect 20346 12809 20409 12895
rect 20409 12809 20495 12895
rect 20495 12809 20577 12895
rect 20577 12809 20663 12895
rect 20663 12809 20726 12895
rect 20346 12526 20726 12809
rect 20346 8526 20726 8906
rect 20346 4526 20726 4906
rect 23106 35286 23486 35666
rect 23106 31286 23486 31666
rect 23106 27286 23486 27666
rect 23106 23286 23486 23666
rect 23106 19613 23169 19666
rect 23169 19613 23255 19666
rect 23255 19613 23337 19666
rect 23337 19613 23423 19666
rect 23423 19613 23486 19666
rect 23106 19286 23486 19613
rect 23106 15286 23486 15666
rect 23106 11286 23486 11666
rect 23106 7603 23486 7666
rect 23106 7517 23169 7603
rect 23169 7517 23255 7603
rect 23255 7517 23337 7603
rect 23337 7517 23423 7603
rect 23423 7517 23486 7603
rect 23106 7286 23486 7517
rect 23106 3286 23486 3666
rect 24346 36526 24726 36906
rect 24346 32551 24726 32906
rect 24346 32526 24409 32551
rect 24409 32526 24495 32551
rect 24495 32526 24577 32551
rect 24577 32526 24663 32551
rect 24663 32526 24726 32551
rect 24346 28526 24726 28906
rect 24346 24905 24409 24906
rect 24409 24905 24495 24906
rect 24495 24905 24577 24906
rect 24577 24905 24663 24906
rect 24663 24905 24726 24906
rect 24346 24526 24726 24905
rect 24346 20526 24726 20906
rect 24346 16526 24726 16906
rect 24346 12895 24726 12906
rect 24346 12809 24409 12895
rect 24409 12809 24495 12895
rect 24495 12809 24577 12895
rect 24577 12809 24663 12895
rect 24663 12809 24726 12895
rect 24346 12526 24726 12809
rect 24346 8526 24726 8906
rect 24346 4526 24726 4906
rect 27106 35286 27486 35666
rect 27106 31286 27486 31666
rect 27106 27286 27486 27666
rect 27106 23286 27486 23666
rect 27106 19613 27169 19666
rect 27169 19613 27255 19666
rect 27255 19613 27337 19666
rect 27337 19613 27423 19666
rect 27423 19613 27486 19666
rect 27106 19286 27486 19613
rect 27106 15286 27486 15666
rect 27106 11286 27486 11666
rect 27106 7603 27486 7666
rect 27106 7517 27169 7603
rect 27169 7517 27255 7603
rect 27255 7517 27337 7603
rect 27337 7517 27423 7603
rect 27423 7517 27486 7603
rect 27106 7286 27486 7517
rect 27106 3286 27486 3666
rect 28346 36526 28726 36906
rect 28346 32551 28726 32906
rect 28346 32526 28409 32551
rect 28409 32526 28495 32551
rect 28495 32526 28577 32551
rect 28577 32526 28663 32551
rect 28663 32526 28726 32551
rect 28346 28526 28726 28906
rect 28346 24905 28409 24906
rect 28409 24905 28495 24906
rect 28495 24905 28577 24906
rect 28577 24905 28663 24906
rect 28663 24905 28726 24906
rect 28346 24526 28726 24905
rect 28346 20526 28726 20906
rect 28346 16526 28726 16906
rect 28346 12895 28726 12906
rect 28346 12809 28409 12895
rect 28409 12809 28495 12895
rect 28495 12809 28577 12895
rect 28577 12809 28663 12895
rect 28663 12809 28726 12895
rect 28346 12526 28726 12809
rect 28346 8526 28726 8906
rect 28346 4526 28726 4906
rect 31106 35286 31486 35666
rect 31106 31286 31486 31666
rect 31106 27286 31486 27666
rect 31106 23286 31486 23666
rect 31106 19613 31169 19666
rect 31169 19613 31255 19666
rect 31255 19613 31337 19666
rect 31337 19613 31423 19666
rect 31423 19613 31486 19666
rect 31106 19286 31486 19613
rect 31106 15286 31486 15666
rect 31106 11286 31486 11666
rect 31106 7603 31486 7666
rect 31106 7517 31169 7603
rect 31169 7517 31255 7603
rect 31255 7517 31337 7603
rect 31337 7517 31423 7603
rect 31423 7517 31486 7603
rect 31106 7286 31486 7517
rect 31106 3286 31486 3666
rect 32346 36526 32726 36906
rect 32346 32551 32726 32906
rect 32346 32526 32409 32551
rect 32409 32526 32495 32551
rect 32495 32526 32577 32551
rect 32577 32526 32663 32551
rect 32663 32526 32726 32551
rect 32346 28526 32726 28906
rect 32346 24905 32409 24906
rect 32409 24905 32495 24906
rect 32495 24905 32577 24906
rect 32577 24905 32663 24906
rect 32663 24905 32726 24906
rect 32346 24526 32726 24905
rect 32346 20526 32726 20906
rect 32346 16526 32726 16906
rect 32346 12895 32726 12906
rect 32346 12809 32409 12895
rect 32409 12809 32495 12895
rect 32495 12809 32577 12895
rect 32577 12809 32663 12895
rect 32663 12809 32726 12895
rect 32346 12526 32726 12809
rect 32346 8526 32726 8906
rect 32346 4526 32726 4906
rect 35106 35286 35486 35666
rect 35106 31286 35486 31666
rect 35106 27286 35486 27666
rect 35106 23286 35486 23666
rect 35106 19613 35169 19666
rect 35169 19613 35255 19666
rect 35255 19613 35337 19666
rect 35337 19613 35423 19666
rect 35423 19613 35486 19666
rect 35106 19286 35486 19613
rect 35106 15286 35486 15666
rect 35106 11286 35486 11666
rect 35106 7603 35486 7666
rect 35106 7517 35169 7603
rect 35169 7517 35255 7603
rect 35255 7517 35337 7603
rect 35337 7517 35423 7603
rect 35423 7517 35486 7603
rect 35106 7286 35486 7517
rect 35106 3286 35486 3666
rect 36346 36526 36726 36906
rect 36346 32551 36726 32906
rect 36346 32526 36409 32551
rect 36409 32526 36495 32551
rect 36495 32526 36577 32551
rect 36577 32526 36663 32551
rect 36663 32526 36726 32551
rect 36346 28526 36726 28906
rect 36346 24905 36409 24906
rect 36409 24905 36495 24906
rect 36495 24905 36577 24906
rect 36577 24905 36663 24906
rect 36663 24905 36726 24906
rect 36346 24526 36726 24905
rect 36346 20526 36726 20906
rect 36346 16526 36726 16906
rect 36346 12895 36726 12906
rect 36346 12809 36409 12895
rect 36409 12809 36495 12895
rect 36495 12809 36577 12895
rect 36577 12809 36663 12895
rect 36663 12809 36726 12895
rect 36346 12526 36726 12809
rect 36346 8526 36726 8906
rect 36346 4526 36726 4906
rect 39106 35286 39486 35666
rect 39106 31286 39486 31666
rect 39106 27286 39486 27666
rect 39106 23286 39486 23666
rect 39106 19613 39169 19666
rect 39169 19613 39255 19666
rect 39255 19613 39337 19666
rect 39337 19613 39423 19666
rect 39423 19613 39486 19666
rect 39106 19286 39486 19613
rect 39106 15286 39486 15666
rect 39106 11286 39486 11666
rect 39106 7603 39486 7666
rect 39106 7517 39169 7603
rect 39169 7517 39255 7603
rect 39255 7517 39337 7603
rect 39337 7517 39423 7603
rect 39423 7517 39486 7603
rect 39106 7286 39486 7517
rect 39106 3286 39486 3666
rect 40346 36526 40726 36906
rect 40346 32551 40726 32906
rect 40346 32526 40409 32551
rect 40409 32526 40495 32551
rect 40495 32526 40577 32551
rect 40577 32526 40663 32551
rect 40663 32526 40726 32551
rect 40346 28526 40726 28906
rect 40346 24905 40409 24906
rect 40409 24905 40495 24906
rect 40495 24905 40577 24906
rect 40577 24905 40663 24906
rect 40663 24905 40726 24906
rect 40346 24526 40726 24905
rect 40346 20526 40726 20906
rect 40346 16526 40726 16906
rect 40346 12895 40726 12906
rect 40346 12809 40409 12895
rect 40409 12809 40495 12895
rect 40495 12809 40577 12895
rect 40577 12809 40663 12895
rect 40663 12809 40726 12895
rect 40346 12526 40726 12809
rect 40346 8526 40726 8906
rect 40346 4526 40726 4906
rect 43106 35286 43486 35666
rect 43106 31286 43486 31666
rect 43106 27286 43486 27666
rect 43106 23286 43486 23666
rect 43106 19613 43169 19666
rect 43169 19613 43255 19666
rect 43255 19613 43337 19666
rect 43337 19613 43423 19666
rect 43423 19613 43486 19666
rect 43106 19286 43486 19613
rect 43106 15286 43486 15666
rect 43106 11286 43486 11666
rect 43106 7603 43486 7666
rect 43106 7517 43169 7603
rect 43169 7517 43255 7603
rect 43255 7517 43337 7603
rect 43337 7517 43423 7603
rect 43423 7517 43486 7603
rect 43106 7286 43486 7517
rect 43106 3286 43486 3666
rect 44346 36526 44726 36906
rect 44346 32551 44726 32906
rect 44346 32526 44409 32551
rect 44409 32526 44495 32551
rect 44495 32526 44577 32551
rect 44577 32526 44663 32551
rect 44663 32526 44726 32551
rect 44346 28526 44726 28906
rect 44346 24905 44409 24906
rect 44409 24905 44495 24906
rect 44495 24905 44577 24906
rect 44577 24905 44663 24906
rect 44663 24905 44726 24906
rect 44346 24526 44726 24905
rect 44346 20526 44726 20906
rect 44346 16526 44726 16906
rect 44346 12895 44726 12906
rect 44346 12809 44409 12895
rect 44409 12809 44495 12895
rect 44495 12809 44577 12895
rect 44577 12809 44663 12895
rect 44663 12809 44726 12895
rect 44346 12526 44726 12809
rect 44346 8526 44726 8906
rect 44346 4526 44726 4906
rect 47106 35286 47486 35666
rect 47106 31286 47486 31666
rect 47106 27286 47486 27666
rect 47106 23286 47486 23666
rect 47106 19613 47169 19666
rect 47169 19613 47255 19666
rect 47255 19613 47337 19666
rect 47337 19613 47423 19666
rect 47423 19613 47486 19666
rect 47106 19286 47486 19613
rect 47106 15286 47486 15666
rect 47106 11286 47486 11666
rect 47106 7603 47486 7666
rect 47106 7517 47169 7603
rect 47169 7517 47255 7603
rect 47255 7517 47337 7603
rect 47337 7517 47423 7603
rect 47423 7517 47486 7603
rect 47106 7286 47486 7517
rect 47106 3286 47486 3666
rect 48346 36526 48726 36906
rect 48346 32551 48726 32906
rect 48346 32526 48409 32551
rect 48409 32526 48495 32551
rect 48495 32526 48577 32551
rect 48577 32526 48663 32551
rect 48663 32526 48726 32551
rect 48346 28526 48726 28906
rect 48346 24905 48409 24906
rect 48409 24905 48495 24906
rect 48495 24905 48577 24906
rect 48577 24905 48663 24906
rect 48663 24905 48726 24906
rect 48346 24526 48726 24905
rect 48346 20526 48726 20906
rect 48346 16526 48726 16906
rect 48346 12895 48726 12906
rect 48346 12809 48409 12895
rect 48409 12809 48495 12895
rect 48495 12809 48577 12895
rect 48577 12809 48663 12895
rect 48663 12809 48726 12895
rect 48346 12526 48726 12809
rect 48346 8526 48726 8906
rect 48346 4526 48726 4906
rect 51106 35286 51486 35666
rect 51106 31286 51486 31666
rect 51106 27286 51486 27666
rect 51106 23286 51486 23666
rect 51106 19613 51169 19666
rect 51169 19613 51255 19666
rect 51255 19613 51337 19666
rect 51337 19613 51423 19666
rect 51423 19613 51486 19666
rect 51106 19286 51486 19613
rect 51106 15286 51486 15666
rect 51106 11286 51486 11666
rect 51106 7603 51486 7666
rect 51106 7517 51169 7603
rect 51169 7517 51255 7603
rect 51255 7517 51337 7603
rect 51337 7517 51423 7603
rect 51423 7517 51486 7603
rect 51106 7286 51486 7517
rect 51106 3286 51486 3666
rect 52346 36526 52726 36906
rect 52346 32551 52726 32906
rect 52346 32526 52409 32551
rect 52409 32526 52495 32551
rect 52495 32526 52577 32551
rect 52577 32526 52663 32551
rect 52663 32526 52726 32551
rect 52346 28526 52726 28906
rect 52346 24905 52409 24906
rect 52409 24905 52495 24906
rect 52495 24905 52577 24906
rect 52577 24905 52663 24906
rect 52663 24905 52726 24906
rect 52346 24526 52726 24905
rect 52346 20526 52726 20906
rect 52346 16526 52726 16906
rect 52346 12895 52726 12906
rect 52346 12809 52409 12895
rect 52409 12809 52495 12895
rect 52495 12809 52577 12895
rect 52577 12809 52663 12895
rect 52663 12809 52726 12895
rect 52346 12526 52726 12809
rect 52346 8526 52726 8906
rect 52346 4526 52726 4906
rect 55106 35286 55486 35666
rect 55106 31286 55486 31666
rect 55106 27286 55486 27666
rect 55106 23286 55486 23666
rect 55106 19613 55169 19666
rect 55169 19613 55255 19666
rect 55255 19613 55337 19666
rect 55337 19613 55423 19666
rect 55423 19613 55486 19666
rect 55106 19286 55486 19613
rect 55106 15286 55486 15666
rect 55106 11286 55486 11666
rect 55106 7603 55486 7666
rect 55106 7517 55169 7603
rect 55169 7517 55255 7603
rect 55255 7517 55337 7603
rect 55337 7517 55423 7603
rect 55423 7517 55486 7603
rect 55106 7286 55486 7517
rect 55106 3286 55486 3666
rect 56346 36526 56726 36906
rect 56346 32551 56726 32906
rect 56346 32526 56409 32551
rect 56409 32526 56495 32551
rect 56495 32526 56577 32551
rect 56577 32526 56663 32551
rect 56663 32526 56726 32551
rect 56346 28526 56726 28906
rect 56346 24905 56409 24906
rect 56409 24905 56495 24906
rect 56495 24905 56577 24906
rect 56577 24905 56663 24906
rect 56663 24905 56726 24906
rect 56346 24526 56726 24905
rect 56346 20526 56726 20906
rect 56346 16526 56726 16906
rect 56346 12895 56726 12906
rect 56346 12809 56409 12895
rect 56409 12809 56495 12895
rect 56495 12809 56577 12895
rect 56577 12809 56663 12895
rect 56663 12809 56726 12895
rect 56346 12526 56726 12809
rect 56346 8526 56726 8906
rect 56346 4526 56726 4906
rect 59106 35286 59486 35666
rect 59106 31286 59486 31666
rect 59106 27286 59486 27666
rect 59106 23286 59486 23666
rect 59106 19613 59169 19666
rect 59169 19613 59255 19666
rect 59255 19613 59337 19666
rect 59337 19613 59423 19666
rect 59423 19613 59486 19666
rect 59106 19286 59486 19613
rect 59106 15286 59486 15666
rect 59106 11286 59486 11666
rect 59106 7603 59486 7666
rect 59106 7517 59169 7603
rect 59169 7517 59255 7603
rect 59255 7517 59337 7603
rect 59337 7517 59423 7603
rect 59423 7517 59486 7603
rect 59106 7286 59486 7517
rect 59106 3286 59486 3666
rect 60346 36526 60726 36906
rect 60346 32551 60726 32906
rect 60346 32526 60409 32551
rect 60409 32526 60495 32551
rect 60495 32526 60577 32551
rect 60577 32526 60663 32551
rect 60663 32526 60726 32551
rect 60346 28526 60726 28906
rect 60346 24905 60409 24906
rect 60409 24905 60495 24906
rect 60495 24905 60577 24906
rect 60577 24905 60663 24906
rect 60663 24905 60726 24906
rect 60346 24526 60726 24905
rect 60346 20526 60726 20906
rect 60346 16526 60726 16906
rect 60346 12895 60726 12906
rect 60346 12809 60409 12895
rect 60409 12809 60495 12895
rect 60495 12809 60577 12895
rect 60577 12809 60663 12895
rect 60663 12809 60726 12895
rect 60346 12526 60726 12809
rect 60346 8526 60726 8906
rect 60346 4526 60726 4906
rect 63106 35286 63486 35666
rect 63106 31286 63486 31666
rect 63106 27286 63486 27666
rect 63106 23286 63486 23666
rect 63106 19613 63169 19666
rect 63169 19613 63255 19666
rect 63255 19613 63337 19666
rect 63337 19613 63423 19666
rect 63423 19613 63486 19666
rect 63106 19286 63486 19613
rect 63106 15286 63486 15666
rect 63106 11286 63486 11666
rect 63106 7603 63486 7666
rect 63106 7517 63169 7603
rect 63169 7517 63255 7603
rect 63255 7517 63337 7603
rect 63337 7517 63423 7603
rect 63423 7517 63486 7603
rect 63106 7286 63486 7517
rect 63106 3286 63486 3666
rect 64346 36526 64726 36906
rect 64346 32551 64726 32906
rect 64346 32526 64409 32551
rect 64409 32526 64495 32551
rect 64495 32526 64577 32551
rect 64577 32526 64663 32551
rect 64663 32526 64726 32551
rect 64346 28526 64726 28906
rect 64346 24905 64409 24906
rect 64409 24905 64495 24906
rect 64495 24905 64577 24906
rect 64577 24905 64663 24906
rect 64663 24905 64726 24906
rect 64346 24526 64726 24905
rect 64346 20526 64726 20906
rect 64346 16526 64726 16906
rect 64346 12895 64726 12906
rect 64346 12809 64409 12895
rect 64409 12809 64495 12895
rect 64495 12809 64577 12895
rect 64577 12809 64663 12895
rect 64663 12809 64726 12895
rect 64346 12526 64726 12809
rect 64346 8526 64726 8906
rect 64346 4526 64726 4906
rect 67106 35286 67486 35666
rect 67106 31286 67486 31666
rect 67106 27286 67486 27666
rect 67106 23286 67486 23666
rect 67106 19613 67169 19666
rect 67169 19613 67255 19666
rect 67255 19613 67337 19666
rect 67337 19613 67423 19666
rect 67423 19613 67486 19666
rect 67106 19286 67486 19613
rect 67106 15286 67486 15666
rect 67106 11286 67486 11666
rect 67106 7603 67486 7666
rect 67106 7517 67169 7603
rect 67169 7517 67255 7603
rect 67255 7517 67337 7603
rect 67337 7517 67423 7603
rect 67423 7517 67486 7603
rect 67106 7286 67486 7517
rect 67106 3286 67486 3666
rect 68346 36526 68726 36906
rect 68346 32551 68726 32906
rect 68346 32526 68409 32551
rect 68409 32526 68495 32551
rect 68495 32526 68577 32551
rect 68577 32526 68663 32551
rect 68663 32526 68726 32551
rect 68346 28526 68726 28906
rect 68346 24905 68409 24906
rect 68409 24905 68495 24906
rect 68495 24905 68577 24906
rect 68577 24905 68663 24906
rect 68663 24905 68726 24906
rect 68346 24526 68726 24905
rect 68346 20526 68726 20906
rect 68346 16526 68726 16906
rect 68346 12895 68726 12906
rect 68346 12809 68409 12895
rect 68409 12809 68495 12895
rect 68495 12809 68577 12895
rect 68577 12809 68663 12895
rect 68663 12809 68726 12895
rect 68346 12526 68726 12809
rect 68346 8526 68726 8906
rect 68346 4526 68726 4906
rect 71106 35286 71486 35666
rect 71106 31286 71486 31666
rect 71106 27286 71486 27666
rect 71106 23286 71486 23666
rect 71106 19613 71169 19666
rect 71169 19613 71255 19666
rect 71255 19613 71337 19666
rect 71337 19613 71423 19666
rect 71423 19613 71486 19666
rect 71106 19286 71486 19613
rect 71106 15286 71486 15666
rect 71106 11286 71486 11666
rect 71106 7286 71486 7666
rect 71106 3286 71486 3666
rect 72346 36526 72726 36906
rect 75106 35286 75486 35666
rect 72346 32526 72726 32906
rect 72346 28526 72726 28906
rect 75106 31286 75486 31666
rect 75106 27636 75486 27666
rect 75106 27550 75169 27636
rect 75169 27550 75255 27636
rect 75255 27550 75337 27636
rect 75337 27550 75423 27636
rect 75423 27550 75486 27636
rect 75106 27468 75486 27550
rect 75106 27382 75169 27468
rect 75169 27382 75255 27468
rect 75255 27382 75337 27468
rect 75337 27382 75423 27468
rect 75423 27382 75486 27468
rect 75106 27300 75486 27382
rect 75106 27286 75169 27300
rect 75169 27286 75255 27300
rect 75255 27286 75337 27300
rect 75337 27286 75423 27300
rect 75423 27286 75486 27300
rect 72346 24526 72726 24906
rect 72346 20526 72726 20906
rect 72346 16526 72726 16906
rect 72346 12868 72409 12906
rect 72409 12868 72495 12906
rect 72495 12868 72577 12906
rect 72577 12868 72663 12906
rect 72663 12868 72726 12906
rect 72346 12786 72726 12868
rect 72346 12700 72409 12786
rect 72409 12700 72495 12786
rect 72495 12700 72577 12786
rect 72577 12700 72663 12786
rect 72663 12700 72726 12786
rect 72346 12618 72726 12700
rect 72346 12532 72409 12618
rect 72409 12532 72495 12618
rect 72495 12532 72577 12618
rect 72577 12532 72663 12618
rect 72663 12532 72726 12618
rect 72346 12526 72726 12532
rect 72346 8526 72726 8906
rect 72346 4526 72726 4906
rect 75106 23286 75486 23666
rect 75106 19613 75169 19666
rect 75169 19613 75255 19666
rect 75255 19613 75337 19666
rect 75337 19613 75423 19666
rect 75423 19613 75486 19666
rect 75106 19286 75486 19613
rect 75106 15286 75486 15666
rect 75106 11286 75486 11666
rect 75106 7286 75486 7666
rect 75106 3286 75486 3666
rect 76346 36526 76726 36906
rect 76346 32526 76726 32906
rect 76346 28526 76726 28906
rect 76346 24526 76726 24906
rect 76346 20526 76726 20906
rect 76346 16526 76726 16906
rect 76346 12868 76409 12906
rect 76409 12868 76495 12906
rect 76495 12868 76577 12906
rect 76577 12868 76663 12906
rect 76663 12868 76726 12906
rect 76346 12786 76726 12868
rect 76346 12700 76409 12786
rect 76409 12700 76495 12786
rect 76495 12700 76577 12786
rect 76577 12700 76663 12786
rect 76663 12700 76726 12786
rect 76346 12618 76726 12700
rect 76346 12532 76409 12618
rect 76409 12532 76495 12618
rect 76495 12532 76577 12618
rect 76577 12532 76663 12618
rect 76663 12532 76726 12618
rect 76346 12526 76726 12532
rect 76346 8526 76726 8906
rect 76346 4526 76726 4906
rect 79106 35286 79486 35666
rect 79106 31286 79486 31666
rect 79106 27636 79486 27666
rect 79106 27550 79169 27636
rect 79169 27550 79255 27636
rect 79255 27550 79337 27636
rect 79337 27550 79423 27636
rect 79423 27550 79486 27636
rect 79106 27468 79486 27550
rect 79106 27382 79169 27468
rect 79169 27382 79255 27468
rect 79255 27382 79337 27468
rect 79337 27382 79423 27468
rect 79423 27382 79486 27468
rect 79106 27300 79486 27382
rect 79106 27286 79169 27300
rect 79169 27286 79255 27300
rect 79255 27286 79337 27300
rect 79337 27286 79423 27300
rect 79423 27286 79486 27300
rect 79106 23286 79486 23666
rect 79106 19613 79169 19666
rect 79169 19613 79255 19666
rect 79255 19613 79337 19666
rect 79337 19613 79423 19666
rect 79423 19613 79486 19666
rect 79106 19286 79486 19613
rect 79106 15286 79486 15666
rect 79106 11286 79486 11666
rect 79106 7286 79486 7666
rect 79106 3286 79486 3666
rect 80346 36526 80726 36906
rect 80346 32526 80726 32906
rect 80346 28526 80726 28906
rect 80346 24526 80726 24906
rect 80346 20526 80726 20906
rect 80346 16526 80726 16906
rect 80346 12868 80409 12906
rect 80409 12868 80495 12906
rect 80495 12868 80577 12906
rect 80577 12868 80663 12906
rect 80663 12868 80726 12906
rect 80346 12786 80726 12868
rect 80346 12700 80409 12786
rect 80409 12700 80495 12786
rect 80495 12700 80577 12786
rect 80577 12700 80663 12786
rect 80663 12700 80726 12786
rect 80346 12618 80726 12700
rect 80346 12532 80409 12618
rect 80409 12532 80495 12618
rect 80495 12532 80577 12618
rect 80577 12532 80663 12618
rect 80663 12532 80726 12618
rect 80346 12526 80726 12532
rect 80346 8526 80726 8906
rect 80346 4526 80726 4906
rect 83106 35286 83486 35666
rect 83106 31286 83486 31666
rect 83106 27636 83486 27666
rect 83106 27550 83169 27636
rect 83169 27550 83255 27636
rect 83255 27550 83337 27636
rect 83337 27550 83423 27636
rect 83423 27550 83486 27636
rect 83106 27468 83486 27550
rect 83106 27382 83169 27468
rect 83169 27382 83255 27468
rect 83255 27382 83337 27468
rect 83337 27382 83423 27468
rect 83423 27382 83486 27468
rect 83106 27300 83486 27382
rect 83106 27286 83169 27300
rect 83169 27286 83255 27300
rect 83255 27286 83337 27300
rect 83337 27286 83423 27300
rect 83423 27286 83486 27300
rect 83106 23286 83486 23666
rect 83106 19613 83169 19666
rect 83169 19613 83255 19666
rect 83255 19613 83337 19666
rect 83337 19613 83423 19666
rect 83423 19613 83486 19666
rect 83106 19286 83486 19613
rect 83106 15286 83486 15666
rect 83106 11286 83486 11666
rect 83106 7286 83486 7666
rect 83106 3286 83486 3666
rect 84346 36526 84726 36906
rect 87106 35286 87486 35666
rect 84346 32526 84726 32906
rect 84346 28526 84726 28906
rect 87106 31286 87486 31666
rect 87106 27636 87486 27666
rect 87106 27550 87169 27636
rect 87169 27550 87255 27636
rect 87255 27550 87337 27636
rect 87337 27550 87423 27636
rect 87423 27550 87486 27636
rect 87106 27468 87486 27550
rect 87106 27382 87169 27468
rect 87169 27382 87255 27468
rect 87255 27382 87337 27468
rect 87337 27382 87423 27468
rect 87423 27382 87486 27468
rect 87106 27300 87486 27382
rect 87106 27286 87169 27300
rect 87169 27286 87255 27300
rect 87255 27286 87337 27300
rect 87337 27286 87423 27300
rect 87423 27286 87486 27300
rect 84346 24526 84726 24906
rect 84346 20526 84726 20906
rect 84346 16526 84726 16906
rect 87106 23286 87486 23666
rect 87106 19613 87169 19666
rect 87169 19613 87255 19666
rect 87255 19613 87337 19666
rect 87337 19613 87423 19666
rect 87423 19613 87486 19666
rect 87106 19286 87486 19613
rect 84346 12868 84409 12906
rect 84409 12868 84495 12906
rect 84495 12868 84577 12906
rect 84577 12868 84663 12906
rect 84663 12868 84726 12906
rect 84346 12786 84726 12868
rect 84346 12700 84409 12786
rect 84409 12700 84495 12786
rect 84495 12700 84577 12786
rect 84577 12700 84663 12786
rect 84663 12700 84726 12786
rect 84346 12618 84726 12700
rect 84346 12532 84409 12618
rect 84409 12532 84495 12618
rect 84495 12532 84577 12618
rect 84577 12532 84663 12618
rect 84663 12532 84726 12618
rect 84346 12526 84726 12532
rect 84346 8526 84726 8906
rect 87106 15286 87486 15666
rect 87106 11286 87486 11666
rect 84346 4526 84726 4906
rect 87106 7286 87486 7666
rect 87106 3286 87486 3666
rect 88346 36526 88726 36906
rect 88346 32526 88726 32906
rect 88346 28526 88726 28906
rect 88346 24526 88726 24906
rect 88346 20526 88726 20906
rect 88346 16526 88726 16906
rect 88346 12868 88409 12906
rect 88409 12868 88495 12906
rect 88495 12868 88577 12906
rect 88577 12868 88663 12906
rect 88663 12868 88726 12906
rect 88346 12786 88726 12868
rect 88346 12700 88409 12786
rect 88409 12700 88495 12786
rect 88495 12700 88577 12786
rect 88577 12700 88663 12786
rect 88663 12700 88726 12786
rect 88346 12618 88726 12700
rect 88346 12532 88409 12618
rect 88409 12532 88495 12618
rect 88495 12532 88577 12618
rect 88577 12532 88663 12618
rect 88663 12532 88726 12618
rect 88346 12526 88726 12532
rect 88346 8526 88726 8906
rect 88346 4526 88726 4906
rect 91106 35286 91486 35666
rect 91106 31286 91486 31666
rect 91106 27636 91486 27666
rect 91106 27550 91169 27636
rect 91169 27550 91255 27636
rect 91255 27550 91337 27636
rect 91337 27550 91423 27636
rect 91423 27550 91486 27636
rect 91106 27468 91486 27550
rect 91106 27382 91169 27468
rect 91169 27382 91255 27468
rect 91255 27382 91337 27468
rect 91337 27382 91423 27468
rect 91423 27382 91486 27468
rect 91106 27300 91486 27382
rect 91106 27286 91169 27300
rect 91169 27286 91255 27300
rect 91255 27286 91337 27300
rect 91337 27286 91423 27300
rect 91423 27286 91486 27300
rect 91106 23286 91486 23666
rect 91106 19613 91169 19666
rect 91169 19613 91255 19666
rect 91255 19613 91337 19666
rect 91337 19613 91423 19666
rect 91423 19613 91486 19666
rect 91106 19286 91486 19613
rect 91106 15286 91486 15666
rect 91106 11286 91486 11666
rect 91106 7286 91486 7666
rect 91106 3286 91486 3666
rect 92346 36526 92726 36906
rect 92346 32526 92726 32906
rect 92346 28526 92726 28906
rect 92346 24526 92726 24906
rect 92346 20526 92726 20906
rect 92346 16526 92726 16906
rect 92346 12868 92409 12906
rect 92409 12868 92495 12906
rect 92495 12868 92577 12906
rect 92577 12868 92663 12906
rect 92663 12868 92726 12906
rect 92346 12786 92726 12868
rect 92346 12700 92409 12786
rect 92409 12700 92495 12786
rect 92495 12700 92577 12786
rect 92577 12700 92663 12786
rect 92663 12700 92726 12786
rect 92346 12618 92726 12700
rect 92346 12532 92409 12618
rect 92409 12532 92495 12618
rect 92495 12532 92577 12618
rect 92577 12532 92663 12618
rect 92663 12532 92726 12618
rect 92346 12526 92726 12532
rect 92346 8526 92726 8906
rect 92346 4526 92726 4906
rect 95106 35286 95486 35666
rect 95106 31286 95486 31666
rect 95106 27636 95486 27666
rect 95106 27550 95169 27636
rect 95169 27550 95255 27636
rect 95255 27550 95337 27636
rect 95337 27550 95423 27636
rect 95423 27550 95486 27636
rect 95106 27468 95486 27550
rect 95106 27382 95169 27468
rect 95169 27382 95255 27468
rect 95255 27382 95337 27468
rect 95337 27382 95423 27468
rect 95423 27382 95486 27468
rect 95106 27300 95486 27382
rect 95106 27286 95169 27300
rect 95169 27286 95255 27300
rect 95255 27286 95337 27300
rect 95337 27286 95423 27300
rect 95423 27286 95486 27300
rect 95106 23286 95486 23666
rect 95106 19613 95169 19666
rect 95169 19613 95255 19666
rect 95255 19613 95337 19666
rect 95337 19613 95423 19666
rect 95423 19613 95486 19666
rect 95106 19286 95486 19613
rect 95106 15286 95486 15666
rect 95106 11286 95486 11666
rect 95106 7286 95486 7666
rect 95106 3286 95486 3666
rect 96346 36526 96726 36906
rect 96346 32526 96726 32906
rect 96346 28526 96726 28906
rect 96346 24526 96726 24906
rect 96346 20526 96726 20906
rect 96346 16526 96726 16906
rect 96346 12868 96409 12906
rect 96409 12868 96495 12906
rect 96495 12868 96577 12906
rect 96577 12868 96663 12906
rect 96663 12868 96726 12906
rect 96346 12786 96726 12868
rect 96346 12700 96409 12786
rect 96409 12700 96495 12786
rect 96495 12700 96577 12786
rect 96577 12700 96663 12786
rect 96663 12700 96726 12786
rect 96346 12618 96726 12700
rect 96346 12532 96409 12618
rect 96409 12532 96495 12618
rect 96495 12532 96577 12618
rect 96577 12532 96663 12618
rect 96663 12532 96726 12618
rect 96346 12526 96726 12532
rect 96346 8526 96726 8906
rect 96346 4526 96726 4906
rect 99106 35286 99486 35666
rect 99106 31286 99486 31666
rect 99106 27286 99486 27666
rect 99106 23286 99486 23666
rect 99106 19613 99169 19666
rect 99169 19613 99255 19666
rect 99255 19613 99337 19666
rect 99337 19613 99423 19666
rect 99423 19613 99486 19666
rect 99106 19286 99486 19613
rect 99106 15286 99486 15666
rect 99106 11286 99486 11666
rect 99106 7286 99486 7666
rect 99106 3286 99486 3666
<< metal7 >>
rect 532 36906 99404 36936
rect 532 36526 4346 36906
rect 4726 36526 8346 36906
rect 8726 36526 12346 36906
rect 12726 36526 16346 36906
rect 16726 36526 20346 36906
rect 20726 36526 24346 36906
rect 24726 36526 28346 36906
rect 28726 36526 32346 36906
rect 32726 36526 36346 36906
rect 36726 36526 40346 36906
rect 40726 36526 44346 36906
rect 44726 36526 48346 36906
rect 48726 36526 52346 36906
rect 52726 36526 56346 36906
rect 56726 36526 60346 36906
rect 60726 36526 64346 36906
rect 64726 36526 68346 36906
rect 68726 36526 72346 36906
rect 72726 36526 76346 36906
rect 76726 36526 80346 36906
rect 80726 36526 84346 36906
rect 84726 36526 88346 36906
rect 88726 36526 92346 36906
rect 92726 36526 96346 36906
rect 96726 36526 99404 36906
rect 532 36496 99404 36526
rect 532 35666 99516 35696
rect 532 35286 3106 35666
rect 3486 35286 7106 35666
rect 7486 35286 11106 35666
rect 11486 35286 15106 35666
rect 15486 35286 19106 35666
rect 19486 35286 23106 35666
rect 23486 35286 27106 35666
rect 27486 35286 31106 35666
rect 31486 35286 35106 35666
rect 35486 35286 39106 35666
rect 39486 35286 43106 35666
rect 43486 35286 47106 35666
rect 47486 35286 51106 35666
rect 51486 35286 55106 35666
rect 55486 35286 59106 35666
rect 59486 35286 63106 35666
rect 63486 35286 67106 35666
rect 67486 35286 71106 35666
rect 71486 35286 75106 35666
rect 75486 35286 79106 35666
rect 79486 35286 83106 35666
rect 83486 35286 87106 35666
rect 87486 35286 91106 35666
rect 91486 35286 95106 35666
rect 95486 35286 99106 35666
rect 99486 35286 99516 35666
rect 532 35256 99516 35286
rect 532 32906 99404 32936
rect 532 32526 4346 32906
rect 4726 32526 8346 32906
rect 8726 32526 12346 32906
rect 12726 32526 16346 32906
rect 16726 32526 20346 32906
rect 20726 32526 24346 32906
rect 24726 32526 28346 32906
rect 28726 32526 32346 32906
rect 32726 32526 36346 32906
rect 36726 32526 40346 32906
rect 40726 32526 44346 32906
rect 44726 32526 48346 32906
rect 48726 32526 52346 32906
rect 52726 32526 56346 32906
rect 56726 32526 60346 32906
rect 60726 32526 64346 32906
rect 64726 32526 68346 32906
rect 68726 32526 72346 32906
rect 72726 32526 76346 32906
rect 76726 32526 80346 32906
rect 80726 32526 84346 32906
rect 84726 32526 88346 32906
rect 88726 32526 92346 32906
rect 92726 32526 96346 32906
rect 96726 32526 99404 32906
rect 532 32496 99404 32526
rect 532 31666 99516 31696
rect 532 31286 3106 31666
rect 3486 31286 7106 31666
rect 7486 31286 11106 31666
rect 11486 31286 15106 31666
rect 15486 31286 19106 31666
rect 19486 31286 23106 31666
rect 23486 31286 27106 31666
rect 27486 31286 31106 31666
rect 31486 31286 35106 31666
rect 35486 31286 39106 31666
rect 39486 31286 43106 31666
rect 43486 31286 47106 31666
rect 47486 31286 51106 31666
rect 51486 31286 55106 31666
rect 55486 31286 59106 31666
rect 59486 31286 63106 31666
rect 63486 31286 67106 31666
rect 67486 31286 71106 31666
rect 71486 31286 75106 31666
rect 75486 31286 79106 31666
rect 79486 31286 83106 31666
rect 83486 31286 87106 31666
rect 87486 31286 91106 31666
rect 91486 31286 95106 31666
rect 95486 31286 99106 31666
rect 99486 31286 99516 31666
rect 532 31256 99516 31286
rect 532 28906 99404 28936
rect 532 28526 4346 28906
rect 4726 28526 8346 28906
rect 8726 28526 12346 28906
rect 12726 28526 16346 28906
rect 16726 28526 20346 28906
rect 20726 28526 24346 28906
rect 24726 28526 28346 28906
rect 28726 28526 32346 28906
rect 32726 28526 36346 28906
rect 36726 28526 40346 28906
rect 40726 28526 44346 28906
rect 44726 28526 48346 28906
rect 48726 28526 52346 28906
rect 52726 28526 56346 28906
rect 56726 28526 60346 28906
rect 60726 28526 64346 28906
rect 64726 28526 68346 28906
rect 68726 28526 72346 28906
rect 72726 28526 76346 28906
rect 76726 28526 80346 28906
rect 80726 28526 84346 28906
rect 84726 28526 88346 28906
rect 88726 28526 92346 28906
rect 92726 28526 96346 28906
rect 96726 28526 99404 28906
rect 532 28496 99404 28526
rect 532 27666 99516 27696
rect 532 27286 3106 27666
rect 3486 27286 7106 27666
rect 7486 27286 11106 27666
rect 11486 27286 15106 27666
rect 15486 27286 19106 27666
rect 19486 27286 23106 27666
rect 23486 27286 27106 27666
rect 27486 27286 31106 27666
rect 31486 27286 35106 27666
rect 35486 27286 39106 27666
rect 39486 27286 43106 27666
rect 43486 27286 47106 27666
rect 47486 27286 51106 27666
rect 51486 27286 55106 27666
rect 55486 27286 59106 27666
rect 59486 27286 63106 27666
rect 63486 27286 67106 27666
rect 67486 27286 71106 27666
rect 71486 27286 75106 27666
rect 75486 27286 79106 27666
rect 79486 27286 83106 27666
rect 83486 27286 87106 27666
rect 87486 27286 91106 27666
rect 91486 27286 95106 27666
rect 95486 27286 99106 27666
rect 99486 27286 99516 27666
rect 532 27256 99516 27286
rect 532 24906 99404 24936
rect 532 24526 4346 24906
rect 4726 24526 8346 24906
rect 8726 24526 12346 24906
rect 12726 24526 16346 24906
rect 16726 24526 20346 24906
rect 20726 24526 24346 24906
rect 24726 24526 28346 24906
rect 28726 24526 32346 24906
rect 32726 24526 36346 24906
rect 36726 24526 40346 24906
rect 40726 24526 44346 24906
rect 44726 24526 48346 24906
rect 48726 24526 52346 24906
rect 52726 24526 56346 24906
rect 56726 24526 60346 24906
rect 60726 24526 64346 24906
rect 64726 24526 68346 24906
rect 68726 24526 72346 24906
rect 72726 24526 76346 24906
rect 76726 24526 80346 24906
rect 80726 24526 84346 24906
rect 84726 24526 88346 24906
rect 88726 24526 92346 24906
rect 92726 24526 96346 24906
rect 96726 24526 99404 24906
rect 532 24496 99404 24526
rect 532 23666 99516 23696
rect 532 23286 3106 23666
rect 3486 23286 7106 23666
rect 7486 23286 11106 23666
rect 11486 23286 15106 23666
rect 15486 23286 19106 23666
rect 19486 23286 23106 23666
rect 23486 23286 27106 23666
rect 27486 23286 31106 23666
rect 31486 23286 35106 23666
rect 35486 23286 39106 23666
rect 39486 23286 43106 23666
rect 43486 23286 47106 23666
rect 47486 23286 51106 23666
rect 51486 23286 55106 23666
rect 55486 23286 59106 23666
rect 59486 23286 63106 23666
rect 63486 23286 67106 23666
rect 67486 23286 71106 23666
rect 71486 23286 75106 23666
rect 75486 23286 79106 23666
rect 79486 23286 83106 23666
rect 83486 23286 87106 23666
rect 87486 23286 91106 23666
rect 91486 23286 95106 23666
rect 95486 23286 99106 23666
rect 99486 23286 99516 23666
rect 532 23256 99516 23286
rect 532 20906 99404 20936
rect 532 20526 4346 20906
rect 4726 20526 8346 20906
rect 8726 20526 12346 20906
rect 12726 20526 16346 20906
rect 16726 20526 20346 20906
rect 20726 20526 24346 20906
rect 24726 20526 28346 20906
rect 28726 20526 32346 20906
rect 32726 20526 36346 20906
rect 36726 20526 40346 20906
rect 40726 20526 44346 20906
rect 44726 20526 48346 20906
rect 48726 20526 52346 20906
rect 52726 20526 56346 20906
rect 56726 20526 60346 20906
rect 60726 20526 64346 20906
rect 64726 20526 68346 20906
rect 68726 20526 72346 20906
rect 72726 20526 76346 20906
rect 76726 20526 80346 20906
rect 80726 20526 84346 20906
rect 84726 20526 88346 20906
rect 88726 20526 92346 20906
rect 92726 20526 96346 20906
rect 96726 20526 99404 20906
rect 532 20496 99404 20526
rect 532 19666 99516 19696
rect 532 19286 3106 19666
rect 3486 19286 7106 19666
rect 7486 19286 11106 19666
rect 11486 19286 15106 19666
rect 15486 19286 19106 19666
rect 19486 19286 23106 19666
rect 23486 19286 27106 19666
rect 27486 19286 31106 19666
rect 31486 19286 35106 19666
rect 35486 19286 39106 19666
rect 39486 19286 43106 19666
rect 43486 19286 47106 19666
rect 47486 19286 51106 19666
rect 51486 19286 55106 19666
rect 55486 19286 59106 19666
rect 59486 19286 63106 19666
rect 63486 19286 67106 19666
rect 67486 19286 71106 19666
rect 71486 19286 75106 19666
rect 75486 19286 79106 19666
rect 79486 19286 83106 19666
rect 83486 19286 87106 19666
rect 87486 19286 91106 19666
rect 91486 19286 95106 19666
rect 95486 19286 99106 19666
rect 99486 19286 99516 19666
rect 532 19256 99516 19286
rect 532 16906 99404 16936
rect 532 16526 4346 16906
rect 4726 16526 8346 16906
rect 8726 16526 12346 16906
rect 12726 16526 16346 16906
rect 16726 16526 20346 16906
rect 20726 16526 24346 16906
rect 24726 16526 28346 16906
rect 28726 16526 32346 16906
rect 32726 16526 36346 16906
rect 36726 16526 40346 16906
rect 40726 16526 44346 16906
rect 44726 16526 48346 16906
rect 48726 16526 52346 16906
rect 52726 16526 56346 16906
rect 56726 16526 60346 16906
rect 60726 16526 64346 16906
rect 64726 16526 68346 16906
rect 68726 16526 72346 16906
rect 72726 16526 76346 16906
rect 76726 16526 80346 16906
rect 80726 16526 84346 16906
rect 84726 16526 88346 16906
rect 88726 16526 92346 16906
rect 92726 16526 96346 16906
rect 96726 16526 99404 16906
rect 532 16496 99404 16526
rect 532 15666 99516 15696
rect 532 15286 3106 15666
rect 3486 15286 7106 15666
rect 7486 15286 11106 15666
rect 11486 15286 15106 15666
rect 15486 15286 19106 15666
rect 19486 15286 23106 15666
rect 23486 15286 27106 15666
rect 27486 15286 31106 15666
rect 31486 15286 35106 15666
rect 35486 15286 39106 15666
rect 39486 15286 43106 15666
rect 43486 15286 47106 15666
rect 47486 15286 51106 15666
rect 51486 15286 55106 15666
rect 55486 15286 59106 15666
rect 59486 15286 63106 15666
rect 63486 15286 67106 15666
rect 67486 15286 71106 15666
rect 71486 15286 75106 15666
rect 75486 15286 79106 15666
rect 79486 15286 83106 15666
rect 83486 15286 87106 15666
rect 87486 15286 91106 15666
rect 91486 15286 95106 15666
rect 95486 15286 99106 15666
rect 99486 15286 99516 15666
rect 532 15256 99516 15286
rect 532 12906 99404 12936
rect 532 12526 4346 12906
rect 4726 12526 8346 12906
rect 8726 12526 12346 12906
rect 12726 12526 16346 12906
rect 16726 12526 20346 12906
rect 20726 12526 24346 12906
rect 24726 12526 28346 12906
rect 28726 12526 32346 12906
rect 32726 12526 36346 12906
rect 36726 12526 40346 12906
rect 40726 12526 44346 12906
rect 44726 12526 48346 12906
rect 48726 12526 52346 12906
rect 52726 12526 56346 12906
rect 56726 12526 60346 12906
rect 60726 12526 64346 12906
rect 64726 12526 68346 12906
rect 68726 12526 72346 12906
rect 72726 12526 76346 12906
rect 76726 12526 80346 12906
rect 80726 12526 84346 12906
rect 84726 12526 88346 12906
rect 88726 12526 92346 12906
rect 92726 12526 96346 12906
rect 96726 12526 99404 12906
rect 532 12496 99404 12526
rect 532 11666 99516 11696
rect 532 11286 3106 11666
rect 3486 11286 7106 11666
rect 7486 11286 11106 11666
rect 11486 11286 15106 11666
rect 15486 11286 19106 11666
rect 19486 11286 23106 11666
rect 23486 11286 27106 11666
rect 27486 11286 31106 11666
rect 31486 11286 35106 11666
rect 35486 11286 39106 11666
rect 39486 11286 43106 11666
rect 43486 11286 47106 11666
rect 47486 11286 51106 11666
rect 51486 11286 55106 11666
rect 55486 11286 59106 11666
rect 59486 11286 63106 11666
rect 63486 11286 67106 11666
rect 67486 11286 71106 11666
rect 71486 11286 75106 11666
rect 75486 11286 79106 11666
rect 79486 11286 83106 11666
rect 83486 11286 87106 11666
rect 87486 11286 91106 11666
rect 91486 11286 95106 11666
rect 95486 11286 99106 11666
rect 99486 11286 99516 11666
rect 532 11256 99516 11286
rect 532 8906 99404 8936
rect 532 8526 4346 8906
rect 4726 8526 8346 8906
rect 8726 8526 12346 8906
rect 12726 8526 16346 8906
rect 16726 8526 20346 8906
rect 20726 8526 24346 8906
rect 24726 8526 28346 8906
rect 28726 8526 32346 8906
rect 32726 8526 36346 8906
rect 36726 8526 40346 8906
rect 40726 8526 44346 8906
rect 44726 8526 48346 8906
rect 48726 8526 52346 8906
rect 52726 8526 56346 8906
rect 56726 8526 60346 8906
rect 60726 8526 64346 8906
rect 64726 8526 68346 8906
rect 68726 8526 72346 8906
rect 72726 8526 76346 8906
rect 76726 8526 80346 8906
rect 80726 8526 84346 8906
rect 84726 8526 88346 8906
rect 88726 8526 92346 8906
rect 92726 8526 96346 8906
rect 96726 8526 99404 8906
rect 532 8496 99404 8526
rect 532 7666 99516 7696
rect 532 7286 3106 7666
rect 3486 7286 7106 7666
rect 7486 7286 11106 7666
rect 11486 7286 15106 7666
rect 15486 7286 19106 7666
rect 19486 7286 23106 7666
rect 23486 7286 27106 7666
rect 27486 7286 31106 7666
rect 31486 7286 35106 7666
rect 35486 7286 39106 7666
rect 39486 7286 43106 7666
rect 43486 7286 47106 7666
rect 47486 7286 51106 7666
rect 51486 7286 55106 7666
rect 55486 7286 59106 7666
rect 59486 7286 63106 7666
rect 63486 7286 67106 7666
rect 67486 7286 71106 7666
rect 71486 7286 75106 7666
rect 75486 7286 79106 7666
rect 79486 7286 83106 7666
rect 83486 7286 87106 7666
rect 87486 7286 91106 7666
rect 91486 7286 95106 7666
rect 95486 7286 99106 7666
rect 99486 7286 99516 7666
rect 532 7256 99516 7286
rect 532 4906 99404 4936
rect 532 4526 4346 4906
rect 4726 4526 8346 4906
rect 8726 4526 12346 4906
rect 12726 4526 16346 4906
rect 16726 4526 20346 4906
rect 20726 4526 24346 4906
rect 24726 4526 28346 4906
rect 28726 4526 32346 4906
rect 32726 4526 36346 4906
rect 36726 4526 40346 4906
rect 40726 4526 44346 4906
rect 44726 4526 48346 4906
rect 48726 4526 52346 4906
rect 52726 4526 56346 4906
rect 56726 4526 60346 4906
rect 60726 4526 64346 4906
rect 64726 4526 68346 4906
rect 68726 4526 72346 4906
rect 72726 4526 76346 4906
rect 76726 4526 80346 4906
rect 80726 4526 84346 4906
rect 84726 4526 88346 4906
rect 88726 4526 92346 4906
rect 92726 4526 96346 4906
rect 96726 4526 99404 4906
rect 532 4496 99404 4526
rect 532 3666 99516 3696
rect 532 3286 3106 3666
rect 3486 3286 7106 3666
rect 7486 3286 11106 3666
rect 11486 3286 15106 3666
rect 15486 3286 19106 3666
rect 19486 3286 23106 3666
rect 23486 3286 27106 3666
rect 27486 3286 31106 3666
rect 31486 3286 35106 3666
rect 35486 3286 39106 3666
rect 39486 3286 43106 3666
rect 43486 3286 47106 3666
rect 47486 3286 51106 3666
rect 51486 3286 55106 3666
rect 55486 3286 59106 3666
rect 59486 3286 63106 3666
rect 63486 3286 67106 3666
rect 67486 3286 71106 3666
rect 71486 3286 75106 3666
rect 75486 3286 79106 3666
rect 79486 3286 83106 3666
rect 83486 3286 87106 3666
rect 87486 3286 91106 3666
rect 91486 3286 95106 3666
rect 95486 3286 99106 3666
rect 99486 3286 99516 3666
rect 532 3256 99516 3286
use sg13g2_buf_1  _08_
timestamp 1676381911
transform -1 0 1536 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _09_
timestamp 1676381911
transform -1 0 1536 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _10_
timestamp 1676381911
transform -1 0 1920 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _11_
timestamp 1676381911
transform -1 0 1344 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _12_
timestamp 1676381911
transform -1 0 1728 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _13_
timestamp 1676381911
transform -1 0 2304 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _14_
timestamp 1676381911
transform -1 0 1152 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _15_
timestamp 1676381911
transform -1 0 1536 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _16_
timestamp 1676381911
transform -1 0 1920 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _17_
timestamp 1676381911
transform -1 0 1632 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _18_
timestamp 1676381911
transform -1 0 2016 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _19_
timestamp 1676381911
transform -1 0 1824 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _20_
timestamp 1676381911
transform -1 0 1440 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _21_
timestamp 1676381911
transform -1 0 1824 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _22_
timestamp 1676381911
transform -1 0 1344 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _23_
timestamp 1676381911
transform -1 0 1728 0 1 9828
box -48 -56 432 834
use dac128module  dacH
timestamp 0
transform 1 0 72000 0 1 26748
box 0 0 1 1
use dac128module  dacL
timestamp 0
transform 1 0 72000 0 1 8014
box 0 0 1 1
use sg13g2_buf_1  digitalenH.g\[0\].u.buff
timestamp 1676381911
transform 1 0 71136 0 -1 27972
box -48 -56 432 834
use sg13g2_inv_1  digitalenH.g\[0\].u.inv
timestamp 1676382929
transform 1 0 71232 0 -1 26460
box -48 -56 336 834
use sg13g2_buf_1  digitalenH.g\[1\].u.buff
timestamp 1676381911
transform -1 0 98688 0 1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalenH.g\[1\].u.inv
timestamp 1676382929
transform -1 0 98976 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalenH.g\[2\].u.buff
timestamp 1676381911
transform -1 0 98784 0 1 32508
box -48 -56 432 834
use sg13g2_inv_1  digitalenH.g\[2\].u.inv
timestamp 1676382929
transform 1 0 98784 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalenH.g\[3\].u.buff
timestamp 1676381911
transform 1 0 71136 0 -1 32508
box -48 -56 432 834
use sg13g2_inv_1  digitalenH.g\[3\].u.inv
timestamp 1676382929
transform 1 0 71424 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalenL.g\[0\].u.buff
timestamp 1676381911
transform 1 0 71136 0 -1 8316
box -48 -56 432 834
use sg13g2_inv_1  digitalenL.g\[0\].u.inv
timestamp 1676382929
transform 1 0 71232 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalenL.g\[1\].u.buff
timestamp 1676381911
transform -1 0 98784 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalenL.g\[1\].u.inv
timestamp 1676382929
transform -1 0 98592 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalenL.g\[2\].u.buff
timestamp 1676381911
transform -1 0 98880 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalenL.g\[2\].u.inv
timestamp 1676382929
transform -1 0 98496 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalenL.g\[3\].u.buff
timestamp 1676381911
transform 1 0 71040 0 1 12852
box -48 -56 432 834
use sg13g2_inv_1  digitalenL.g\[3\].u.inv
timestamp 1676382929
transform 1 0 71040 0 -1 12852
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[0\].u.buff
timestamp 1676381911
transform 1 0 71040 0 1 26460
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[0\].u.inv
timestamp 1676382929
transform 1 0 70848 0 -1 26460
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[1\].u.buff
timestamp 1676381911
transform 1 0 70272 0 1 26460
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[1\].u.inv
timestamp 1676382929
transform 1 0 72576 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[2\].u.buff
timestamp 1676381911
transform 1 0 70656 0 1 26460
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[2\].u.inv
timestamp 1676382929
transform 1 0 70848 0 -1 27972
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[3\].u.buff
timestamp 1676381911
transform 1 0 73248 0 1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[3\].u.inv
timestamp 1676382929
transform 1 0 73152 0 -1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[4\].u.buff
timestamp 1676381911
transform 1 0 73824 0 1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[4\].u.inv
timestamp 1676382929
transform -1 0 73728 0 -1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[5\].u.buff
timestamp 1676381911
transform 1 0 69696 0 1 26460
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[5\].u.inv
timestamp 1676382929
transform -1 0 76128 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[6\].u.buff
timestamp 1676381911
transform 1 0 74592 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[6\].u.inv
timestamp 1676382929
transform -1 0 76416 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[7\].u.buff
timestamp 1676381911
transform 1 0 75168 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[7\].u.inv
timestamp 1676382929
transform -1 0 75840 0 -1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[8\].u.buff
timestamp 1676381911
transform 1 0 75456 0 1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[8\].u.inv
timestamp 1676382929
transform -1 0 76704 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[9\].u.buff
timestamp 1676381911
transform 1 0 75936 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[9\].u.inv
timestamp 1676382929
transform 1 0 76704 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[10\].u.buff
timestamp 1676381911
transform 1 0 76320 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[10\].u.inv
timestamp 1676382929
transform 1 0 76992 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[11\].u.buff
timestamp 1676381911
transform 1 0 76800 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[11\].u.inv
timestamp 1676382929
transform -1 0 78720 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[12\].u.buff
timestamp 1676381911
transform 1 0 77184 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[12\].u.inv
timestamp 1676382929
transform -1 0 78144 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[13\].u.buff
timestamp 1676381911
transform -1 0 78336 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[13\].u.inv
timestamp 1676382929
transform -1 0 78432 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[14\].u.buff
timestamp 1676381911
transform -1 0 78720 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[14\].u.inv
timestamp 1676382929
transform -1 0 79968 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[15\].u.buff
timestamp 1676381911
transform -1 0 79104 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[15\].u.inv
timestamp 1676382929
transform -1 0 79008 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[16\].u.buff
timestamp 1676381911
transform -1 0 79488 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[16\].u.inv
timestamp 1676382929
transform 1 0 79008 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[17\].u.buff
timestamp 1676381911
transform -1 0 79872 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[17\].u.inv
timestamp 1676382929
transform 1 0 79392 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[18\].u.buff
timestamp 1676381911
transform -1 0 80256 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[18\].u.inv
timestamp 1676382929
transform 1 0 79968 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[19\].u.buff
timestamp 1676381911
transform -1 0 80448 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[19\].u.inv
timestamp 1676382929
transform -1 0 80544 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[20\].u.buff
timestamp 1676381911
transform -1 0 81504 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[20\].u.inv
timestamp 1676382929
transform 1 0 80640 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[21\].u.buff
timestamp 1676381911
transform -1 0 81888 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[21\].u.inv
timestamp 1676382929
transform 1 0 81024 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[22\].u.buff
timestamp 1676381911
transform -1 0 82272 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[22\].u.inv
timestamp 1676382929
transform 1 0 81408 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[23\].u.buff
timestamp 1676381911
transform 1 0 81600 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[23\].u.inv
timestamp 1676382929
transform 1 0 81888 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[24\].u.buff
timestamp 1676381911
transform -1 0 82656 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[24\].u.inv
timestamp 1676382929
transform 1 0 82176 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[25\].u.buff
timestamp 1676381911
transform 1 0 82368 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[25\].u.inv
timestamp 1676382929
transform 1 0 82560 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[26\].u.buff
timestamp 1676381911
transform 1 0 82848 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[26\].u.inv
timestamp 1676382929
transform -1 0 83328 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[27\].u.buff
timestamp 1676381911
transform 1 0 83232 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[27\].u.inv
timestamp 1676382929
transform -1 0 84192 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[28\].u.buff
timestamp 1676381911
transform 1 0 83616 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[28\].u.inv
timestamp 1676382929
transform -1 0 84480 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[29\].u.buff
timestamp 1676381911
transform -1 0 84768 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[29\].u.inv
timestamp 1676382929
transform -1 0 84768 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[30\].u.buff
timestamp 1676381911
transform -1 0 85152 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[30\].u.inv
timestamp 1676382929
transform -1 0 85056 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[31\].u.buff
timestamp 1676381911
transform 1 0 84864 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[31\].u.inv
timestamp 1676382929
transform 1 0 85056 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[32\].u.buff
timestamp 1676381911
transform 1 0 85248 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[32\].u.inv
timestamp 1676382929
transform 1 0 85440 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[33\].u.buff
timestamp 1676381911
transform 1 0 85632 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[33\].u.inv
timestamp 1676382929
transform 1 0 85824 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[34\].u.buff
timestamp 1676381911
transform 1 0 86016 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[34\].u.inv
timestamp 1676382929
transform -1 0 86592 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[35\].u.buff
timestamp 1676381911
transform 1 0 86400 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[35\].u.inv
timestamp 1676382929
transform -1 0 87744 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[36\].u.buff
timestamp 1676381911
transform 1 0 86880 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[36\].u.inv
timestamp 1676382929
transform -1 0 87936 0 -1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[37\].u.buff
timestamp 1676381911
transform 1 0 87264 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[37\].u.inv
timestamp 1676382929
transform -1 0 88032 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[38\].u.buff
timestamp 1676381911
transform 1 0 87648 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[38\].u.inv
timestamp 1676382929
transform -1 0 88320 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[39\].u.buff
timestamp 1676381911
transform 1 0 88032 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[39\].u.inv
timestamp 1676382929
transform -1 0 88608 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[40\].u.buff
timestamp 1676381911
transform 1 0 88416 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[40\].u.inv
timestamp 1676382929
transform 1 0 88608 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[41\].u.buff
timestamp 1676381911
transform 1 0 88800 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[41\].u.inv
timestamp 1676382929
transform 1 0 88992 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[42\].u.buff
timestamp 1676381911
transform 1 0 89184 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[42\].u.inv
timestamp 1676382929
transform -1 0 90144 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[43\].u.buff
timestamp 1676381911
transform 1 0 89664 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[43\].u.inv
timestamp 1676382929
transform -1 0 90432 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[44\].u.buff
timestamp 1676381911
transform 1 0 90048 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[44\].u.inv
timestamp 1676382929
transform -1 0 90720 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[45\].u.buff
timestamp 1676381911
transform 1 0 90432 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[45\].u.inv
timestamp 1676382929
transform -1 0 91008 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[46\].u.buff
timestamp 1676381911
transform 1 0 90912 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[46\].u.inv
timestamp 1676382929
transform -1 0 91392 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[47\].u.buff
timestamp 1676381911
transform 1 0 91200 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[47\].u.inv
timestamp 1676382929
transform 1 0 91392 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[48\].u.buff
timestamp 1676381911
transform 1 0 91584 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[48\].u.inv
timestamp 1676382929
transform 1 0 91872 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[49\].u.buff
timestamp 1676381911
transform -1 0 92448 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[49\].u.inv
timestamp 1676382929
transform 1 0 92256 0 1 23436
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[50\].u.buff
timestamp 1676381911
transform -1 0 93216 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[50\].u.inv
timestamp 1676382929
transform -1 0 93024 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[51\].u.buff
timestamp 1676381911
transform -1 0 93600 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[51\].u.inv
timestamp 1676382929
transform 1 0 93024 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[52\].u.buff
timestamp 1676381911
transform 1 0 93312 0 1 23436
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[52\].u.inv
timestamp 1676382929
transform -1 0 93792 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[53\].u.buff
timestamp 1676381911
transform 1 0 93696 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[53\].u.inv
timestamp 1676382929
transform 1 0 93888 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[54\].u.buff
timestamp 1676381911
transform 1 0 94080 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[54\].u.inv
timestamp 1676382929
transform 1 0 94176 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[55\].u.buff
timestamp 1676381911
transform 1 0 94464 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[55\].u.inv
timestamp 1676382929
transform -1 0 95040 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[56\].u.buff
timestamp 1676381911
transform 1 0 94848 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[56\].u.inv
timestamp 1676382929
transform -1 0 95424 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[57\].u.buff
timestamp 1676381911
transform 1 0 95328 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[57\].u.inv
timestamp 1676382929
transform -1 0 96288 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[58\].u.buff
timestamp 1676381911
transform -1 0 96480 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[58\].u.inv
timestamp 1676382929
transform -1 0 96576 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[59\].u.buff
timestamp 1676381911
transform -1 0 96864 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[59\].u.inv
timestamp 1676382929
transform -1 0 97632 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[60\].u.buff
timestamp 1676381911
transform -1 0 97248 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[60\].u.inv
timestamp 1676382929
transform 1 0 96672 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[61\].u.buff
timestamp 1676381911
transform -1 0 97632 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[61\].u.inv
timestamp 1676382929
transform 1 0 97056 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[62\].u.buff
timestamp 1676381911
transform -1 0 98016 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[62\].u.inv
timestamp 1676382929
transform -1 0 97920 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[63\].u.buff
timestamp 1676381911
transform -1 0 98400 0 -1 24948
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[63\].u.inv
timestamp 1676382929
transform 1 0 97920 0 1 24948
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[64\].u.buff
timestamp 1676381911
transform -1 0 98496 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[64\].u.inv
timestamp 1676382929
transform 1 0 99072 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[65\].u.buff
timestamp 1676381911
transform -1 0 98112 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[65\].u.inv
timestamp 1676382929
transform -1 0 98208 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[66\].u.buff
timestamp 1676381911
transform -1 0 97728 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[66\].u.inv
timestamp 1676382929
transform -1 0 97920 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[67\].u.buff
timestamp 1676381911
transform -1 0 97344 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[67\].u.inv
timestamp 1676382929
transform -1 0 97632 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[68\].u.buff
timestamp 1676381911
transform -1 0 96960 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[68\].u.inv
timestamp 1676382929
transform -1 0 97344 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[69\].u.buff
timestamp 1676381911
transform -1 0 96576 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[69\].u.inv
timestamp 1676382929
transform -1 0 96480 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[70\].u.buff
timestamp 1676381911
transform -1 0 96192 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[70\].u.inv
timestamp 1676382929
transform -1 0 96192 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[71\].u.buff
timestamp 1676381911
transform -1 0 95424 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[71\].u.inv
timestamp 1676382929
transform 1 0 95616 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[72\].u.buff
timestamp 1676381911
transform 1 0 94560 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[72\].u.inv
timestamp 1676382929
transform -1 0 95616 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[73\].u.buff
timestamp 1676381911
transform 1 0 94176 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[73\].u.inv
timestamp 1676382929
transform -1 0 95328 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[74\].u.buff
timestamp 1676381911
transform -1 0 94176 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[74\].u.inv
timestamp 1676382929
transform -1 0 94752 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[75\].u.buff
timestamp 1676381911
transform 1 0 93312 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[75\].u.inv
timestamp 1676382929
transform 1 0 94752 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[76\].u.buff
timestamp 1676381911
transform -1 0 93696 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[76\].u.inv
timestamp 1676382929
transform -1 0 94464 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[77\].u.buff
timestamp 1676381911
transform -1 0 93312 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[77\].u.inv
timestamp 1676382929
transform -1 0 93792 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[78\].u.buff
timestamp 1676381911
transform 1 0 92160 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[78\].u.inv
timestamp 1676382929
transform -1 0 93504 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[79\].u.buff
timestamp 1676381911
transform 1 0 91776 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[79\].u.inv
timestamp 1676382929
transform 1 0 92928 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[80\].u.buff
timestamp 1676381911
transform 1 0 91392 0 1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[80\].u.inv
timestamp 1676382929
transform -1 0 92928 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[81\].u.buff
timestamp 1676381911
transform -1 0 91776 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[81\].u.inv
timestamp 1676382929
transform -1 0 92160 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[82\].u.buff
timestamp 1676381911
transform -1 0 91392 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[82\].u.inv
timestamp 1676382929
transform -1 0 91872 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[83\].u.buff
timestamp 1676381911
transform -1 0 91008 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[83\].u.inv
timestamp 1676382929
transform -1 0 91584 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[84\].u.buff
timestamp 1676381911
transform -1 0 90624 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[84\].u.inv
timestamp 1676382929
transform -1 0 91296 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[85\].u.buff
timestamp 1676381911
transform -1 0 90240 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[85\].u.inv
timestamp 1676382929
transform -1 0 90432 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[86\].u.buff
timestamp 1676381911
transform 1 0 88896 0 1 32508
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[86\].u.inv
timestamp 1676382929
transform 1 0 89856 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[87\].u.buff
timestamp 1676381911
transform -1 0 89472 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[87\].u.inv
timestamp 1676382929
transform -1 0 89856 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[88\].u.buff
timestamp 1676381911
transform -1 0 89088 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[88\].u.inv
timestamp 1676382929
transform -1 0 89568 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[89\].u.buff
timestamp 1676381911
transform -1 0 88704 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[89\].u.inv
timestamp 1676382929
transform -1 0 88800 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[90\].u.buff
timestamp 1676381911
transform -1 0 88320 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[90\].u.inv
timestamp 1676382929
transform 1 0 88224 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[91\].u.buff
timestamp 1676381911
transform -1 0 87936 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[91\].u.inv
timestamp 1676382929
transform -1 0 87744 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[92\].u.buff
timestamp 1676381911
transform -1 0 87552 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[92\].u.inv
timestamp 1676382929
transform -1 0 87456 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[93\].u.buff
timestamp 1676381911
transform -1 0 86784 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[93\].u.inv
timestamp 1676382929
transform -1 0 87168 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[94\].u.buff
timestamp 1676381911
transform -1 0 86400 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[94\].u.inv
timestamp 1676382929
transform 1 0 86592 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[95\].u.buff
timestamp 1676381911
transform -1 0 86016 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[95\].u.inv
timestamp 1676382929
transform -1 0 86112 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[96\].u.buff
timestamp 1676381911
transform -1 0 85632 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[96\].u.inv
timestamp 1676382929
transform -1 0 85824 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[97\].u.buff
timestamp 1676381911
transform -1 0 85248 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[97\].u.inv
timestamp 1676382929
transform -1 0 85536 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[98\].u.buff
timestamp 1676381911
transform -1 0 84864 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[98\].u.inv
timestamp 1676382929
transform 1 0 84960 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[99\].u.buff
timestamp 1676381911
transform -1 0 84480 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[99\].u.inv
timestamp 1676382929
transform -1 0 84576 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[100\].u.buff
timestamp 1676381911
transform -1 0 84096 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[100\].u.inv
timestamp 1676382929
transform -1 0 84288 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[101\].u.buff
timestamp 1676381911
transform -1 0 83712 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[101\].u.inv
timestamp 1676382929
transform -1 0 84000 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[102\].u.buff
timestamp 1676381911
transform -1 0 83328 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[102\].u.inv
timestamp 1676382929
transform 1 0 83424 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[103\].u.buff
timestamp 1676381911
transform -1 0 82944 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[103\].u.inv
timestamp 1676382929
transform -1 0 83040 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[104\].u.buff
timestamp 1676381911
transform -1 0 82176 0 1 32508
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[104\].u.inv
timestamp 1676382929
transform -1 0 82752 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[105\].u.buff
timestamp 1676381911
transform -1 0 82176 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[105\].u.inv
timestamp 1676382929
transform 1 0 82176 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[106\].u.buff
timestamp 1676381911
transform -1 0 81792 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[106\].u.inv
timestamp 1676382929
transform -1 0 81792 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[107\].u.buff
timestamp 1676381911
transform 1 0 80544 0 1 32508
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[107\].u.inv
timestamp 1676382929
transform -1 0 81504 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[108\].u.buff
timestamp 1676381911
transform -1 0 81024 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[108\].u.inv
timestamp 1676382929
transform -1 0 81216 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[109\].u.buff
timestamp 1676381911
transform 1 0 79680 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[109\].u.inv
timestamp 1676382929
transform 1 0 80160 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[110\].u.buff
timestamp 1676381911
transform 1 0 79296 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[110\].u.inv
timestamp 1676382929
transform -1 0 80160 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[111\].u.buff
timestamp 1676381911
transform 1 0 78912 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[111\].u.inv
timestamp 1676382929
transform -1 0 79872 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[112\].u.buff
timestamp 1676381911
transform 1 0 78528 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[112\].u.inv
timestamp 1676382929
transform -1 0 79584 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[113\].u.buff
timestamp 1676381911
transform 1 0 78144 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[113\].u.inv
timestamp 1676382929
transform 1 0 79008 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[114\].u.buff
timestamp 1676381911
transform 1 0 77760 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[114\].u.inv
timestamp 1676382929
transform -1 0 78528 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[115\].u.buff
timestamp 1676381911
transform 1 0 77376 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[115\].u.inv
timestamp 1676382929
transform -1 0 78240 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[116\].u.buff
timestamp 1676381911
transform 1 0 76896 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[116\].u.inv
timestamp 1676382929
transform -1 0 77952 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[117\].u.buff
timestamp 1676381911
transform 1 0 76512 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[117\].u.inv
timestamp 1676382929
transform 1 0 77376 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[118\].u.buff
timestamp 1676381911
transform 1 0 76128 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[118\].u.inv
timestamp 1676382929
transform -1 0 76992 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[119\].u.buff
timestamp 1676381911
transform 1 0 75744 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[119\].u.inv
timestamp 1676382929
transform -1 0 76704 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[120\].u.buff
timestamp 1676381911
transform 1 0 75264 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[120\].u.inv
timestamp 1676382929
transform -1 0 76416 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[121\].u.buff
timestamp 1676381911
transform 1 0 74784 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[121\].u.inv
timestamp 1676382929
transform -1 0 75552 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[122\].u.buff
timestamp 1676381911
transform 1 0 74400 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[122\].u.inv
timestamp 1676382929
transform -1 0 75264 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[123\].u.buff
timestamp 1676381911
transform 1 0 74016 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[123\].u.inv
timestamp 1676382929
transform -1 0 74112 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[124\].u.buff
timestamp 1676381911
transform 1 0 73536 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[124\].u.inv
timestamp 1676382929
transform 1 0 73536 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[125\].u.buff
timestamp 1676381911
transform 1 0 73152 0 -1 34020
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[125\].u.inv
timestamp 1676382929
transform 1 0 72960 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[126\].u.buff
timestamp 1676381911
transform 1 0 72576 0 1 32508
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[126\].u.inv
timestamp 1676382929
transform 1 0 72288 0 1 32508
box -48 -56 336 834
use sg13g2_buf_1  digitalH.g\[127\].u.buff
timestamp 1676381911
transform 1 0 70560 0 1 30996
box -48 -56 432 834
use sg13g2_inv_1  digitalH.g\[127\].u.inv
timestamp 1676382929
transform 1 0 70944 0 1 30996
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[0\].u.buff
timestamp 1676381911
transform 1 0 70752 0 -1 8316
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[0\].u.inv
timestamp 1676382929
transform 1 0 72000 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[1\].u.buff
timestamp 1676381911
transform 1 0 72288 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[1\].u.inv
timestamp 1676382929
transform -1 0 73536 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[2\].u.buff
timestamp 1676381911
transform 1 0 72864 0 1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[2\].u.inv
timestamp 1676382929
transform 1 0 73536 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[3\].u.buff
timestamp 1676381911
transform 1 0 73440 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[3\].u.inv
timestamp 1676382929
transform 1 0 73152 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[4\].u.buff
timestamp 1676381911
transform 1 0 73920 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[4\].u.inv
timestamp 1676382929
transform -1 0 75072 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[5\].u.buff
timestamp 1676381911
transform 1 0 74304 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[5\].u.inv
timestamp 1676382929
transform -1 0 75360 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[6\].u.buff
timestamp 1676381911
transform 1 0 74784 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[6\].u.inv
timestamp 1676382929
transform -1 0 76128 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[7\].u.buff
timestamp 1676381911
transform 1 0 75168 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[7\].u.inv
timestamp 1676382929
transform -1 0 76416 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[8\].u.buff
timestamp 1676381911
transform 1 0 75552 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[8\].u.inv
timestamp 1676382929
transform -1 0 76704 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[9\].u.buff
timestamp 1676381911
transform 1 0 75936 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[9\].u.inv
timestamp 1676382929
transform -1 0 76992 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[10\].u.buff
timestamp 1676381911
transform 1 0 76416 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[10\].u.inv
timestamp 1676382929
transform 1 0 77472 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[11\].u.buff
timestamp 1676381911
transform 1 0 76800 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[11\].u.inv
timestamp 1676382929
transform -1 0 78048 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[12\].u.buff
timestamp 1676381911
transform 1 0 77184 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[12\].u.inv
timestamp 1676382929
transform -1 0 78336 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[13\].u.buff
timestamp 1676381911
transform 1 0 77568 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[13\].u.inv
timestamp 1676382929
transform -1 0 78624 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[14\].u.buff
timestamp 1676381911
transform 1 0 78048 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[14\].u.inv
timestamp 1676382929
transform 1 0 79104 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[15\].u.buff
timestamp 1676381911
transform 1 0 78432 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[15\].u.inv
timestamp 1676382929
transform -1 0 79680 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[16\].u.buff
timestamp 1676381911
transform 1 0 78816 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[16\].u.inv
timestamp 1676382929
transform -1 0 80736 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[17\].u.buff
timestamp 1676381911
transform 1 0 79200 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[17\].u.inv
timestamp 1676382929
transform 1 0 80736 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[18\].u.buff
timestamp 1676381911
transform 1 0 79680 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[18\].u.inv
timestamp 1676382929
transform -1 0 81312 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[19\].u.buff
timestamp 1676381911
transform 1 0 80064 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[19\].u.inv
timestamp 1676382929
transform -1 0 81120 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[20\].u.buff
timestamp 1676381911
transform 1 0 80448 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[20\].u.inv
timestamp 1676382929
transform -1 0 82176 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[21\].u.buff
timestamp 1676381911
transform 1 0 80832 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[21\].u.inv
timestamp 1676382929
transform 1 0 82176 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[22\].u.buff
timestamp 1676381911
transform 1 0 81216 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[22\].u.inv
timestamp 1676382929
transform -1 0 82752 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[23\].u.buff
timestamp 1676381911
transform 1 0 81600 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[23\].u.inv
timestamp 1676382929
transform -1 0 83040 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[24\].u.buff
timestamp 1676381911
transform 1 0 81984 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[24\].u.inv
timestamp 1676382929
transform -1 0 83808 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[25\].u.buff
timestamp 1676381911
transform 1 0 82464 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[25\].u.inv
timestamp 1676382929
transform 1 0 83808 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[26\].u.buff
timestamp 1676381911
transform 1 0 82848 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[26\].u.inv
timestamp 1676382929
transform -1 0 83520 0 -1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[27\].u.buff
timestamp 1676381911
transform 1 0 83232 0 1 5292
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[27\].u.inv
timestamp 1676382929
transform -1 0 84384 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[28\].u.buff
timestamp 1676381911
transform 1 0 83616 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[28\].u.inv
timestamp 1676382929
transform -1 0 84672 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[29\].u.buff
timestamp 1676381911
transform 1 0 84000 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[29\].u.inv
timestamp 1676382929
transform 1 0 85152 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[30\].u.buff
timestamp 1676381911
transform 1 0 84384 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[30\].u.inv
timestamp 1676382929
transform -1 0 85728 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[31\].u.buff
timestamp 1676381911
transform 1 0 84768 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[31\].u.inv
timestamp 1676382929
transform -1 0 86016 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[32\].u.buff
timestamp 1676381911
transform 1 0 85248 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[32\].u.inv
timestamp 1676382929
transform -1 0 87072 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[33\].u.buff
timestamp 1676381911
transform 1 0 85632 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[33\].u.inv
timestamp 1676382929
transform 1 0 87072 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[34\].u.buff
timestamp 1676381911
transform 1 0 86016 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[34\].u.inv
timestamp 1676382929
transform -1 0 87648 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[35\].u.buff
timestamp 1676381911
transform 1 0 86400 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[35\].u.inv
timestamp 1676382929
transform -1 0 87936 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[36\].u.buff
timestamp 1676381911
transform 1 0 86784 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[36\].u.inv
timestamp 1676382929
transform -1 0 88608 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[37\].u.buff
timestamp 1676381911
transform 1 0 87264 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[37\].u.inv
timestamp 1676382929
transform 1 0 88608 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[38\].u.buff
timestamp 1676381911
transform -1 0 88032 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[38\].u.inv
timestamp 1676382929
transform -1 0 89184 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[39\].u.buff
timestamp 1676381911
transform 1 0 88032 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[39\].u.inv
timestamp 1676382929
transform -1 0 89856 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[40\].u.buff
timestamp 1676381911
transform 1 0 88416 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[40\].u.inv
timestamp 1676382929
transform 1 0 89856 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[41\].u.buff
timestamp 1676381911
transform 1 0 88800 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[41\].u.inv
timestamp 1676382929
transform -1 0 90432 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[42\].u.buff
timestamp 1676381911
transform 1 0 89184 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[42\].u.inv
timestamp 1676382929
transform -1 0 90720 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[43\].u.buff
timestamp 1676381911
transform 1 0 89664 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[43\].u.inv
timestamp 1676382929
transform -1 0 91392 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[44\].u.buff
timestamp 1676381911
transform 1 0 90048 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[44\].u.inv
timestamp 1676382929
transform 1 0 91392 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[45\].u.buff
timestamp 1676381911
transform 1 0 90432 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[45\].u.inv
timestamp 1676382929
transform -1 0 91968 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[46\].u.buff
timestamp 1676381911
transform 1 0 90816 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[46\].u.inv
timestamp 1676382929
transform 1 0 91008 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[47\].u.buff
timestamp 1676381911
transform 1 0 91200 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[47\].u.inv
timestamp 1676382929
transform -1 0 93120 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[48\].u.buff
timestamp 1676381911
transform 1 0 91680 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[48\].u.inv
timestamp 1676382929
transform 1 0 93120 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[49\].u.buff
timestamp 1676381911
transform 1 0 92064 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[49\].u.inv
timestamp 1676382929
transform -1 0 93696 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[50\].u.buff
timestamp 1676381911
transform 1 0 92448 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[50\].u.inv
timestamp 1676382929
transform -1 0 93984 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[51\].u.buff
timestamp 1676381911
transform 1 0 92832 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[51\].u.inv
timestamp 1676382929
transform -1 0 94656 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[52\].u.buff
timestamp 1676381911
transform 1 0 93312 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[52\].u.inv
timestamp 1676382929
transform 1 0 94656 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[53\].u.buff
timestamp 1676381911
transform -1 0 94080 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[53\].u.inv
timestamp 1676382929
transform 1 0 93888 0 1 5292
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[54\].u.buff
timestamp 1676381911
transform 1 0 94080 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[54\].u.inv
timestamp 1676382929
transform -1 0 95808 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[55\].u.buff
timestamp 1676381911
transform 1 0 94464 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[55\].u.inv
timestamp 1676382929
transform 1 0 95808 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[56\].u.buff
timestamp 1676381911
transform 1 0 94848 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[56\].u.inv
timestamp 1676382929
transform -1 0 96384 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[57\].u.buff
timestamp 1676381911
transform 1 0 95328 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[57\].u.inv
timestamp 1676382929
transform -1 0 96672 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[58\].u.buff
timestamp 1676381911
transform 1 0 95712 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[58\].u.inv
timestamp 1676382929
transform -1 0 97440 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[59\].u.buff
timestamp 1676381911
transform 1 0 96096 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[59\].u.inv
timestamp 1676382929
transform 1 0 97440 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[60\].u.buff
timestamp 1676381911
transform 1 0 96480 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[60\].u.inv
timestamp 1676382929
transform -1 0 98016 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[61\].u.buff
timestamp 1676381911
transform -1 0 97344 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[61\].u.inv
timestamp 1676382929
transform -1 0 98304 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[62\].u.buff
timestamp 1676381911
transform -1 0 97824 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[62\].u.inv
timestamp 1676382929
transform -1 0 99072 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[63\].u.buff
timestamp 1676381911
transform -1 0 98208 0 -1 6804
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[63\].u.inv
timestamp 1676382929
transform 1 0 99072 0 1 6804
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[64\].u.buff
timestamp 1676381911
transform -1 0 98496 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[64\].u.inv
timestamp 1676382929
transform 1 0 98496 0 -1 15876
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[65\].u.buff
timestamp 1676381911
transform -1 0 98112 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[65\].u.inv
timestamp 1676382929
transform 1 0 97344 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[66\].u.buff
timestamp 1676381911
transform -1 0 97728 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[66\].u.inv
timestamp 1676382929
transform 1 0 97632 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[67\].u.buff
timestamp 1676381911
transform -1 0 96960 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[67\].u.inv
timestamp 1676382929
transform -1 0 97248 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[68\].u.buff
timestamp 1676381911
transform -1 0 96960 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[68\].u.inv
timestamp 1676382929
transform -1 0 96480 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[69\].u.buff
timestamp 1676381911
transform -1 0 96576 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[69\].u.inv
timestamp 1676382929
transform -1 0 96096 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[70\].u.buff
timestamp 1676381911
transform -1 0 96192 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[70\].u.inv
timestamp 1676382929
transform -1 0 95616 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[71\].u.buff
timestamp 1676381911
transform 1 0 94944 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[71\].u.inv
timestamp 1676382929
transform 1 0 94944 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[72\].u.buff
timestamp 1676381911
transform 1 0 94560 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[72\].u.inv
timestamp 1676382929
transform 1 0 94560 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[73\].u.buff
timestamp 1676381911
transform 1 0 94176 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[73\].u.inv
timestamp 1676382929
transform 1 0 94176 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[74\].u.buff
timestamp 1676381911
transform 1 0 93696 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[74\].u.inv
timestamp 1676382929
transform -1 0 94080 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[75\].u.buff
timestamp 1676381911
transform 1 0 93312 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[75\].u.inv
timestamp 1676382929
transform 1 0 93312 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[76\].u.buff
timestamp 1676381911
transform 1 0 92928 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[76\].u.inv
timestamp 1676382929
transform 1 0 92640 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[77\].u.buff
timestamp 1676381911
transform 1 0 92640 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[77\].u.inv
timestamp 1676382929
transform 1 0 92352 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[78\].u.buff
timestamp 1676381911
transform -1 0 92640 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[78\].u.inv
timestamp 1676382929
transform 1 0 92064 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[79\].u.buff
timestamp 1676381911
transform 1 0 91872 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[79\].u.inv
timestamp 1676382929
transform 1 0 91680 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[80\].u.buff
timestamp 1676381911
transform 1 0 91392 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[80\].u.inv
timestamp 1676382929
transform -1 0 91680 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[81\].u.buff
timestamp 1676381911
transform 1 0 91008 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[81\].u.inv
timestamp 1676382929
transform 1 0 90912 0 1 15876
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[82\].u.buff
timestamp 1676381911
transform 1 0 90432 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[82\].u.inv
timestamp 1676382929
transform 1 0 90528 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[83\].u.buff
timestamp 1676381911
transform -1 0 91200 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[83\].u.inv
timestamp 1676382929
transform 1 0 90144 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[84\].u.buff
timestamp 1676381911
transform 1 0 89760 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[84\].u.inv
timestamp 1676382929
transform -1 0 90144 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[85\].u.buff
timestamp 1676381911
transform 1 0 89376 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[85\].u.inv
timestamp 1676382929
transform -1 0 89760 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[86\].u.buff
timestamp 1676381911
transform 1 0 88992 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[86\].u.inv
timestamp 1676382929
transform 1 0 88896 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[87\].u.buff
timestamp 1676381911
transform 1 0 88608 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[87\].u.inv
timestamp 1676382929
transform 1 0 88512 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[88\].u.buff
timestamp 1676381911
transform 1 0 88224 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[88\].u.inv
timestamp 1676382929
transform 1 0 88128 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[89\].u.buff
timestamp 1676381911
transform 1 0 87840 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[89\].u.inv
timestamp 1676382929
transform -1 0 88032 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[90\].u.buff
timestamp 1676381911
transform 1 0 87360 0 1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[90\].u.inv
timestamp 1676382929
transform 1 0 87360 0 -1 15876
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[91\].u.buff
timestamp 1676381911
transform 1 0 86976 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[91\].u.inv
timestamp 1676382929
transform 1 0 86976 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[92\].u.buff
timestamp 1676381911
transform 1 0 86496 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[92\].u.inv
timestamp 1676382929
transform -1 0 86880 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[93\].u.buff
timestamp 1676381911
transform 1 0 86112 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[93\].u.inv
timestamp 1676382929
transform -1 0 86496 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[94\].u.buff
timestamp 1676381911
transform 1 0 85728 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[94\].u.inv
timestamp 1676382929
transform 1 0 85728 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[95\].u.buff
timestamp 1676381911
transform 1 0 85344 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[95\].u.inv
timestamp 1676382929
transform 1 0 85344 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[96\].u.buff
timestamp 1676381911
transform 1 0 84960 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[96\].u.inv
timestamp 1676382929
transform 1 0 84960 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[97\].u.buff
timestamp 1676381911
transform 1 0 84480 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[97\].u.inv
timestamp 1676382929
transform 1 0 84480 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[98\].u.buff
timestamp 1676381911
transform 1 0 84096 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[98\].u.inv
timestamp 1676382929
transform 1 0 83808 0 -1 15876
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[99\].u.buff
timestamp 1676381911
transform 1 0 83712 0 1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[99\].u.inv
timestamp 1676382929
transform 1 0 83712 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[100\].u.buff
timestamp 1676381911
transform 1 0 83328 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[100\].u.inv
timestamp 1676382929
transform 1 0 83328 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[101\].u.buff
timestamp 1676381911
transform 1 0 82944 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[101\].u.inv
timestamp 1676382929
transform 1 0 82944 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[102\].u.buff
timestamp 1676381911
transform 1 0 82464 0 1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[102\].u.inv
timestamp 1676382929
transform 1 0 82560 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[103\].u.buff
timestamp 1676381911
transform 1 0 82176 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[103\].u.inv
timestamp 1676382929
transform 1 0 81888 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[104\].u.buff
timestamp 1676381911
transform -1 0 82272 0 1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[104\].u.inv
timestamp 1676382929
transform 1 0 81696 0 -1 15876
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[105\].u.buff
timestamp 1676381911
transform 1 0 81120 0 1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[105\].u.inv
timestamp 1676382929
transform 1 0 81312 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[106\].u.buff
timestamp 1676381911
transform 1 0 81024 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[106\].u.inv
timestamp 1676382929
transform 1 0 80928 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[107\].u.buff
timestamp 1676381911
transform 1 0 80640 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[107\].u.inv
timestamp 1676382929
transform -1 0 80928 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[108\].u.buff
timestamp 1676381911
transform 1 0 80160 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[108\].u.inv
timestamp 1676382929
transform 1 0 80064 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[109\].u.buff
timestamp 1676381911
transform 1 0 79680 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[109\].u.inv
timestamp 1676382929
transform 1 0 80352 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[110\].u.buff
timestamp 1676381911
transform 1 0 79296 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[110\].u.inv
timestamp 1676382929
transform 1 0 79296 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[111\].u.buff
timestamp 1676381911
transform 1 0 78816 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[111\].u.inv
timestamp 1676382929
transform 1 0 79584 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[112\].u.buff
timestamp 1676381911
transform -1 0 79296 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[112\].u.inv
timestamp 1676382929
transform -1 0 78816 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[113\].u.buff
timestamp 1676381911
transform 1 0 78048 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[113\].u.inv
timestamp 1676382929
transform 1 0 78048 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[114\].u.buff
timestamp 1676381911
transform 1 0 77664 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[114\].u.inv
timestamp 1676382929
transform 1 0 77760 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[115\].u.buff
timestamp 1676381911
transform 1 0 77280 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[115\].u.inv
timestamp 1676382929
transform 1 0 77280 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[116\].u.buff
timestamp 1676381911
transform 1 0 76896 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[116\].u.inv
timestamp 1676382929
transform 1 0 76896 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[117\].u.buff
timestamp 1676381911
transform 1 0 76512 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[117\].u.inv
timestamp 1676382929
transform 1 0 76512 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[118\].u.buff
timestamp 1676381911
transform 1 0 76128 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[118\].u.inv
timestamp 1676382929
transform 1 0 76032 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[119\].u.buff
timestamp 1676381911
transform 1 0 75744 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[119\].u.inv
timestamp 1676382929
transform 1 0 75744 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[120\].u.buff
timestamp 1676381911
transform 1 0 75264 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[120\].u.inv
timestamp 1676382929
transform 1 0 75264 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[121\].u.buff
timestamp 1676381911
transform 1 0 74784 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[121\].u.inv
timestamp 1676382929
transform 1 0 74784 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[122\].u.buff
timestamp 1676381911
transform 1 0 74400 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[122\].u.inv
timestamp 1676382929
transform 1 0 74112 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[123\].u.buff
timestamp 1676381911
transform 1 0 73632 0 -1 15876
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[123\].u.inv
timestamp 1676382929
transform 1 0 72672 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[124\].u.buff
timestamp 1676381911
transform 1 0 73440 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[124\].u.inv
timestamp 1676382929
transform 1 0 73824 0 1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[125\].u.buff
timestamp 1676381911
transform 1 0 72960 0 1 14364
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[125\].u.inv
timestamp 1676382929
transform 1 0 71232 0 -1 14364
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[126\].u.buff
timestamp 1676381911
transform 1 0 69792 0 1 12852
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[126\].u.inv
timestamp 1676382929
transform 1 0 70368 0 -1 12852
box -48 -56 336 834
use sg13g2_buf_1  digitalL.g\[127\].u.buff
timestamp 1676381911
transform 1 0 70656 0 1 12852
box -48 -56 432 834
use sg13g2_inv_1  digitalL.g\[127\].u.inv
timestamp 1676382929
transform 1 0 70752 0 -1 12852
box -48 -56 336 834
use sg13g2_buf_2  fanout21
timestamp 1676381867
transform 1 0 69792 0 -1 27972
box -48 -56 528 834
use sg13g2_buf_1  fanout22
timestamp 1676381911
transform -1 0 71040 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout23
timestamp 1676381911
transform -1 0 70656 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  fanout24
timestamp 1676381911
transform -1 0 74592 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout25
timestamp 1676381911
transform 1 0 74976 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout26
timestamp 1676381911
transform 1 0 77568 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout27
timestamp 1676381911
transform 1 0 77472 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout28
timestamp 1676381911
transform -1 0 74976 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout29
timestamp 1676381911
transform -1 0 81120 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_2  fanout30
timestamp 1676381867
transform 1 0 80256 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_1  fanout31
timestamp 1676381911
transform 1 0 84000 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout32
timestamp 1676381911
transform 1 0 83520 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout33
timestamp 1676381911
transform 1 0 74112 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout34
timestamp 1676381911
transform -1 0 74496 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout35
timestamp 1676381911
transform 1 0 75744 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout36
timestamp 1676381911
transform -1 0 77376 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout37
timestamp 1676381911
transform 1 0 78624 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout38
timestamp 1676381911
transform 1 0 74592 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout39
timestamp 1676381911
transform 1 0 80256 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout40
timestamp 1676381911
transform -1 0 82560 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout41
timestamp 1676381911
transform 1 0 83040 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout42
timestamp 1676381911
transform 1 0 84576 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout43
timestamp 1676381911
transform 1 0 81024 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout44
timestamp 1676381911
transform 1 0 73728 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout45
timestamp 1676381911
transform 1 0 86496 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_2  fanout46
timestamp 1676381867
transform 1 0 86592 0 1 24948
box -48 -56 528 834
use sg13g2_buf_1  fanout47
timestamp 1676381911
transform 1 0 88800 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout48
timestamp 1676381911
transform 1 0 89472 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout49
timestamp 1676381911
transform -1 0 92832 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_2  fanout50
timestamp 1676381867
transform -1 0 92736 0 1 24948
box -48 -56 528 834
use sg13g2_buf_1  fanout51
timestamp 1676381911
transform 1 0 95712 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout52
timestamp 1676381911
transform 1 0 95616 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout53
timestamp 1676381911
transform 1 0 87072 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout54
timestamp 1676381911
transform 1 0 86208 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout55
timestamp 1676381911
transform 1 0 87840 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout56
timestamp 1676381911
transform -1 0 89856 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout57
timestamp 1676381911
transform 1 0 90624 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout58
timestamp 1676381911
transform -1 0 87168 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout59
timestamp 1676381911
transform -1 0 92640 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout60
timestamp 1676381911
transform 1 0 93792 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout61
timestamp 1676381911
transform -1 0 95808 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout62
timestamp 1676381911
transform 1 0 96672 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  fanout63
timestamp 1676381911
transform 1 0 92544 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  fanout64
timestamp 1676381911
transform 1 0 72864 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  fanout65
timestamp 1676381911
transform -1 0 2208 0 1 8316
box -48 -56 432 834
use sg13g2_buf_2  fanout66
timestamp 1676381867
transform 1 0 70176 0 1 12852
box -48 -56 528 834
use sg13g2_buf_2  fanout67
timestamp 1676381867
transform -1 0 71328 0 1 8316
box -48 -56 528 834
use sg13g2_buf_1  fanout68
timestamp 1676381911
transform -1 0 74400 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout69
timestamp 1676381911
transform 1 0 75456 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout70
timestamp 1676381911
transform -1 0 77472 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout71
timestamp 1676381911
transform 1 0 78720 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout72
timestamp 1676381911
transform -1 0 74784 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout73
timestamp 1676381911
transform -1 0 74400 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout74
timestamp 1676381911
transform 1 0 73824 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout75
timestamp 1676381911
transform 1 0 76704 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout76
timestamp 1676381911
transform 1 0 78528 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout77
timestamp 1676381911
transform 1 0 77088 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout78
timestamp 1676381911
transform 1 0 79680 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout79
timestamp 1676381911
transform 1 0 81504 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout80
timestamp 1676381911
transform 1 0 83136 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout81
timestamp 1676381911
transform 1 0 84768 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout82
timestamp 1676381911
transform -1 0 80448 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout83
timestamp 1676381911
transform -1 0 80640 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout84
timestamp 1676381911
transform -1 0 81888 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout85
timestamp 1676381911
transform -1 0 83424 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout86
timestamp 1676381911
transform 1 0 84576 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout87
timestamp 1676381911
transform 1 0 80352 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout88
timestamp 1676381911
transform 1 0 74208 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout89
timestamp 1676381911
transform -1 0 86400 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout90
timestamp 1676381911
transform -1 0 88320 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout91
timestamp 1676381911
transform 1 0 89184 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout92
timestamp 1676381911
transform 1 0 90720 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout93
timestamp 1676381911
transform -1 0 86784 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout94
timestamp 1676381911
transform -1 0 86688 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout95
timestamp 1676381911
transform -1 0 88320 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout96
timestamp 1676381911
transform -1 0 89472 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout97
timestamp 1676381911
transform 1 0 90528 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout98
timestamp 1676381911
transform 1 0 86112 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  fanout99
timestamp 1676381911
transform -1 0 92448 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout100
timestamp 1676381911
transform -1 0 94368 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout101
timestamp 1676381911
transform 1 0 95136 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout102
timestamp 1676381911
transform 1 0 96768 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout103
timestamp 1676381911
transform -1 0 92832 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  fanout104
timestamp 1676381911
transform -1 0 92352 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout105
timestamp 1676381911
transform -1 0 94176 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout106
timestamp 1676381911
transform 1 0 92352 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout107
timestamp 1676381911
transform -1 0 95808 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout108
timestamp 1676381911
transform -1 0 97344 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  fanout109
timestamp 1676381911
transform 1 0 95520 0 1 15876
box -48 -56 432 834
use sg13g2_buf_2  fanout110
timestamp 1676381867
transform -1 0 86976 0 -1 17388
box -48 -56 528 834
use sg13g2_buf_2  fanout111
timestamp 1676381867
transform -1 0 71040 0 -1 14364
box -48 -56 528 834
use sg13g2_buf_1  fanout112
timestamp 1676381911
transform -1 0 2112 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 1920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 2592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 3264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 3936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 4608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 5280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 5952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 6624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 7296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 7968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 8640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 9312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 9984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 10656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 11328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 12000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 12672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 13344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 14016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 14688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 15360 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 16032 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 16704 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 17376 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 18048 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 18720 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 19392 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 20064 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 20736 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 21408 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 22080 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 22752 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 23424 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 24096 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 24768 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 25440 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 26112 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 26784 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 27456 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 28128 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 28800 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 29472 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 30144 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 30816 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 31488 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 32160 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 32832 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 33504 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 34176 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 34848 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 35520 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 36192 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 36864 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 37536 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 38208 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 38880 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 39552 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 40224 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 40896 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 41568 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679581782
transform 1 0 42240 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679581782
transform 1 0 42912 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679581782
transform 1 0 43584 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679581782
transform 1 0 44256 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679581782
transform 1 0 44928 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679581782
transform 1 0 45600 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679581782
transform 1 0 46272 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679581782
transform 1 0 46944 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679581782
transform 1 0 47616 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679581782
transform 1 0 48288 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679581782
transform 1 0 48960 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679581782
transform 1 0 49632 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679581782
transform 1 0 50304 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679581782
transform 1 0 50976 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679581782
transform 1 0 51648 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679581782
transform 1 0 52320 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679581782
transform 1 0 52992 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679581782
transform 1 0 53664 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679581782
transform 1 0 54336 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679581782
transform 1 0 55008 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679581782
transform 1 0 55680 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679581782
transform 1 0 56352 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679581782
transform 1 0 57024 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679581782
transform 1 0 57696 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679581782
transform 1 0 58368 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679581782
transform 1 0 59040 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679581782
transform 1 0 59712 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679581782
transform 1 0 60384 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679581782
transform 1 0 61056 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679581782
transform 1 0 61728 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679581782
transform 1 0 62400 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679581782
transform 1 0 63072 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679581782
transform 1 0 63744 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679581782
transform 1 0 64416 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679581782
transform 1 0 65088 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679581782
transform 1 0 65760 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679581782
transform 1 0 66432 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679581782
transform 1 0 67104 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679581782
transform 1 0 67776 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679581782
transform 1 0 68448 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679581782
transform 1 0 69120 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679581782
transform 1 0 69792 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679581782
transform 1 0 70464 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679581782
transform 1 0 71136 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679581782
transform 1 0 71808 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_749
timestamp 1679581782
transform 1 0 72480 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_756
timestamp 1679581782
transform 1 0 73152 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_763
timestamp 1679581782
transform 1 0 73824 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_770
timestamp 1679581782
transform 1 0 74496 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_777
timestamp 1679581782
transform 1 0 75168 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_784
timestamp 1679581782
transform 1 0 75840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_791
timestamp 1679581782
transform 1 0 76512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_798
timestamp 1679581782
transform 1 0 77184 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_805
timestamp 1679581782
transform 1 0 77856 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_812
timestamp 1679581782
transform 1 0 78528 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_819
timestamp 1679581782
transform 1 0 79200 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_826
timestamp 1679581782
transform 1 0 79872 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_833
timestamp 1679581782
transform 1 0 80544 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_840
timestamp 1679581782
transform 1 0 81216 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_847
timestamp 1679581782
transform 1 0 81888 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_854
timestamp 1679581782
transform 1 0 82560 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_861
timestamp 1679581782
transform 1 0 83232 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_868
timestamp 1679581782
transform 1 0 83904 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_875
timestamp 1679581782
transform 1 0 84576 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_882
timestamp 1679581782
transform 1 0 85248 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_889
timestamp 1679581782
transform 1 0 85920 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_896
timestamp 1679581782
transform 1 0 86592 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_903
timestamp 1679581782
transform 1 0 87264 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_910
timestamp 1679581782
transform 1 0 87936 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_917
timestamp 1679581782
transform 1 0 88608 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_924
timestamp 1679581782
transform 1 0 89280 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_931
timestamp 1679581782
transform 1 0 89952 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_938
timestamp 1679581782
transform 1 0 90624 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_945
timestamp 1679581782
transform 1 0 91296 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_952
timestamp 1679581782
transform 1 0 91968 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_959
timestamp 1679581782
transform 1 0 92640 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_966
timestamp 1679581782
transform 1 0 93312 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_973
timestamp 1679581782
transform 1 0 93984 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_980
timestamp 1679581782
transform 1 0 94656 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_987
timestamp 1679581782
transform 1 0 95328 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_994
timestamp 1679581782
transform 1 0 96000 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1001
timestamp 1679581782
transform 1 0 96672 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1008
timestamp 1679581782
transform 1 0 97344 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1015
timestamp 1679581782
transform 1 0 98016 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_1022
timestamp 1679581782
transform 1 0 98688 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 1920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 2592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 3936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 4608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 5952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 6624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 7968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 8640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 9312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 9984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 10656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 11328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 12000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 12672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 13344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 14016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 14688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15360 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16032 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 16704 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17376 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18048 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 18720 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19392 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20064 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 20736 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679581782
transform 1 0 21408 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679581782
transform 1 0 22080 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 22752 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679581782
transform 1 0 23424 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679581782
transform 1 0 24096 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679581782
transform 1 0 24768 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679581782
transform 1 0 25440 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679581782
transform 1 0 26112 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679581782
transform 1 0 26784 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679581782
transform 1 0 27456 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679581782
transform 1 0 28128 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679581782
transform 1 0 28800 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679581782
transform 1 0 29472 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679581782
transform 1 0 30144 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679581782
transform 1 0 30816 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679581782
transform 1 0 31488 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679581782
transform 1 0 32160 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679581782
transform 1 0 32832 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679581782
transform 1 0 33504 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679581782
transform 1 0 34176 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679581782
transform 1 0 34848 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679581782
transform 1 0 35520 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679581782
transform 1 0 36192 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679581782
transform 1 0 36864 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679581782
transform 1 0 37536 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679581782
transform 1 0 38208 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679581782
transform 1 0 38880 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 39552 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 40224 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 40896 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 41568 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42240 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 42912 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 43584 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 44256 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 44928 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 45600 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 46272 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 46944 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 47616 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679581782
transform 1 0 48288 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679581782
transform 1 0 48960 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679581782
transform 1 0 49632 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679581782
transform 1 0 50304 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 50976 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 51648 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 52320 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679581782
transform 1 0 52992 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679581782
transform 1 0 53664 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679581782
transform 1 0 54336 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679581782
transform 1 0 55008 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679581782
transform 1 0 55680 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679581782
transform 1 0 56352 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679581782
transform 1 0 57024 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_595
timestamp 1679581782
transform 1 0 57696 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_602
timestamp 1679581782
transform 1 0 58368 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679581782
transform 1 0 59040 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_616
timestamp 1679581782
transform 1 0 59712 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_623
timestamp 1679581782
transform 1 0 60384 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_630
timestamp 1679581782
transform 1 0 61056 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_637
timestamp 1679581782
transform 1 0 61728 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_644
timestamp 1679581782
transform 1 0 62400 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_651
timestamp 1679581782
transform 1 0 63072 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_658
timestamp 1679581782
transform 1 0 63744 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_665
timestamp 1679581782
transform 1 0 64416 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_672
timestamp 1679581782
transform 1 0 65088 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_679
timestamp 1679581782
transform 1 0 65760 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_686
timestamp 1679581782
transform 1 0 66432 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_693
timestamp 1679581782
transform 1 0 67104 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_700
timestamp 1679581782
transform 1 0 67776 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_707
timestamp 1679581782
transform 1 0 68448 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_714
timestamp 1679581782
transform 1 0 69120 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_721
timestamp 1679581782
transform 1 0 69792 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_728
timestamp 1679581782
transform 1 0 70464 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_735
timestamp 1679581782
transform 1 0 71136 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_742
timestamp 1679581782
transform 1 0 71808 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_749
timestamp 1679581782
transform 1 0 72480 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_756
timestamp 1679581782
transform 1 0 73152 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_763
timestamp 1679581782
transform 1 0 73824 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_770
timestamp 1679581782
transform 1 0 74496 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_777
timestamp 1679581782
transform 1 0 75168 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_784
timestamp 1679581782
transform 1 0 75840 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_791
timestamp 1679581782
transform 1 0 76512 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_798
timestamp 1679581782
transform 1 0 77184 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_805
timestamp 1679581782
transform 1 0 77856 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_812
timestamp 1679581782
transform 1 0 78528 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_819
timestamp 1679581782
transform 1 0 79200 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_826
timestamp 1679581782
transform 1 0 79872 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_833
timestamp 1679581782
transform 1 0 80544 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_840
timestamp 1679581782
transform 1 0 81216 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_847
timestamp 1679581782
transform 1 0 81888 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_854
timestamp 1679581782
transform 1 0 82560 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_861
timestamp 1679581782
transform 1 0 83232 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_868
timestamp 1679581782
transform 1 0 83904 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_875
timestamp 1679581782
transform 1 0 84576 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_882
timestamp 1679581782
transform 1 0 85248 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_889
timestamp 1679581782
transform 1 0 85920 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_896
timestamp 1679581782
transform 1 0 86592 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_903
timestamp 1679581782
transform 1 0 87264 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_910
timestamp 1679581782
transform 1 0 87936 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_917
timestamp 1679581782
transform 1 0 88608 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_924
timestamp 1679581782
transform 1 0 89280 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_931
timestamp 1679581782
transform 1 0 89952 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_938
timestamp 1679581782
transform 1 0 90624 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_945
timestamp 1679581782
transform 1 0 91296 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_952
timestamp 1679581782
transform 1 0 91968 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_959
timestamp 1679581782
transform 1 0 92640 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_966
timestamp 1679581782
transform 1 0 93312 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_973
timestamp 1679581782
transform 1 0 93984 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_980
timestamp 1679581782
transform 1 0 94656 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_987
timestamp 1679581782
transform 1 0 95328 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_994
timestamp 1679581782
transform 1 0 96000 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1001
timestamp 1679581782
transform 1 0 96672 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1008
timestamp 1679581782
transform 1 0 97344 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1015
timestamp 1679581782
transform 1 0 98016 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_1022
timestamp 1679581782
transform 1 0 98688 0 -1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_4
timestamp 1679581782
transform 1 0 960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_11
timestamp 1679581782
transform 1 0 1632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_18
timestamp 1679581782
transform 1 0 2304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_25
timestamp 1679581782
transform 1 0 2976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_32
timestamp 1679581782
transform 1 0 3648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_39
timestamp 1679581782
transform 1 0 4320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_46
timestamp 1679581782
transform 1 0 4992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_53
timestamp 1679581782
transform 1 0 5664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_60
timestamp 1679581782
transform 1 0 6336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_67
timestamp 1679581782
transform 1 0 7008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_74
timestamp 1679581782
transform 1 0 7680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_81
timestamp 1679581782
transform 1 0 8352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_88
timestamp 1679581782
transform 1 0 9024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_95
timestamp 1679581782
transform 1 0 9696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_102
timestamp 1679581782
transform 1 0 10368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_109
timestamp 1679581782
transform 1 0 11040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_116
timestamp 1679581782
transform 1 0 11712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_123
timestamp 1679581782
transform 1 0 12384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_130
timestamp 1679581782
transform 1 0 13056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_137
timestamp 1679581782
transform 1 0 13728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_144
timestamp 1679581782
transform 1 0 14400 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_151
timestamp 1679581782
transform 1 0 15072 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_158
timestamp 1679581782
transform 1 0 15744 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_165
timestamp 1679581782
transform 1 0 16416 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_172
timestamp 1679581782
transform 1 0 17088 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_179
timestamp 1679581782
transform 1 0 17760 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_186
timestamp 1679581782
transform 1 0 18432 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_193
timestamp 1679581782
transform 1 0 19104 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_200
timestamp 1679581782
transform 1 0 19776 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_207
timestamp 1679581782
transform 1 0 20448 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_214
timestamp 1679581782
transform 1 0 21120 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_221
timestamp 1679581782
transform 1 0 21792 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_228
timestamp 1679581782
transform 1 0 22464 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_235
timestamp 1679581782
transform 1 0 23136 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_242
timestamp 1679581782
transform 1 0 23808 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_249
timestamp 1679581782
transform 1 0 24480 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_256
timestamp 1679581782
transform 1 0 25152 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_263
timestamp 1679581782
transform 1 0 25824 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_270
timestamp 1679581782
transform 1 0 26496 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_277
timestamp 1679581782
transform 1 0 27168 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_284
timestamp 1679581782
transform 1 0 27840 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_291
timestamp 1679581782
transform 1 0 28512 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_298
timestamp 1679581782
transform 1 0 29184 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_305
timestamp 1679581782
transform 1 0 29856 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_312
timestamp 1679581782
transform 1 0 30528 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_319
timestamp 1679581782
transform 1 0 31200 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_326
timestamp 1679581782
transform 1 0 31872 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_333
timestamp 1679581782
transform 1 0 32544 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_340
timestamp 1679581782
transform 1 0 33216 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_347
timestamp 1679581782
transform 1 0 33888 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_354
timestamp 1679581782
transform 1 0 34560 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_361
timestamp 1679581782
transform 1 0 35232 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_368
timestamp 1679581782
transform 1 0 35904 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_375
timestamp 1679581782
transform 1 0 36576 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_382
timestamp 1679581782
transform 1 0 37248 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_389
timestamp 1679581782
transform 1 0 37920 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_396
timestamp 1679581782
transform 1 0 38592 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_403
timestamp 1679581782
transform 1 0 39264 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_410
timestamp 1679581782
transform 1 0 39936 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_417
timestamp 1679581782
transform 1 0 40608 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_424
timestamp 1679581782
transform 1 0 41280 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_431
timestamp 1679581782
transform 1 0 41952 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_438
timestamp 1679581782
transform 1 0 42624 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_445
timestamp 1679581782
transform 1 0 43296 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_452
timestamp 1679581782
transform 1 0 43968 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_459
timestamp 1679581782
transform 1 0 44640 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_466
timestamp 1679581782
transform 1 0 45312 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_473
timestamp 1679581782
transform 1 0 45984 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_480
timestamp 1679581782
transform 1 0 46656 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_487
timestamp 1679581782
transform 1 0 47328 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_494
timestamp 1679581782
transform 1 0 48000 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_501
timestamp 1679581782
transform 1 0 48672 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_508
timestamp 1679581782
transform 1 0 49344 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_515
timestamp 1679581782
transform 1 0 50016 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_522
timestamp 1679581782
transform 1 0 50688 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_529
timestamp 1679581782
transform 1 0 51360 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_536
timestamp 1679581782
transform 1 0 52032 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_543
timestamp 1679581782
transform 1 0 52704 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_550
timestamp 1679581782
transform 1 0 53376 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_557
timestamp 1679581782
transform 1 0 54048 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_564
timestamp 1679581782
transform 1 0 54720 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_571
timestamp 1679581782
transform 1 0 55392 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_578
timestamp 1679581782
transform 1 0 56064 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_585
timestamp 1679581782
transform 1 0 56736 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_592
timestamp 1679581782
transform 1 0 57408 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_599
timestamp 1679581782
transform 1 0 58080 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_606
timestamp 1679581782
transform 1 0 58752 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_613
timestamp 1679581782
transform 1 0 59424 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_620
timestamp 1679581782
transform 1 0 60096 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_627
timestamp 1679581782
transform 1 0 60768 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_634
timestamp 1679581782
transform 1 0 61440 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_641
timestamp 1679581782
transform 1 0 62112 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_648
timestamp 1679581782
transform 1 0 62784 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_655
timestamp 1679581782
transform 1 0 63456 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_662
timestamp 1679581782
transform 1 0 64128 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_669
timestamp 1679581782
transform 1 0 64800 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_676
timestamp 1679581782
transform 1 0 65472 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_683
timestamp 1679581782
transform 1 0 66144 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_690
timestamp 1679581782
transform 1 0 66816 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_697
timestamp 1679581782
transform 1 0 67488 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_704
timestamp 1679581782
transform 1 0 68160 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_711
timestamp 1679581782
transform 1 0 68832 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_718
timestamp 1679581782
transform 1 0 69504 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_725
timestamp 1679581782
transform 1 0 70176 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_732
timestamp 1679581782
transform 1 0 70848 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_739
timestamp 1679581782
transform 1 0 71520 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_746
timestamp 1679581782
transform 1 0 72192 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_753
timestamp 1679581782
transform 1 0 72864 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_760
timestamp 1679581782
transform 1 0 73536 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_767
timestamp 1679581782
transform 1 0 74208 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_774
timestamp 1679581782
transform 1 0 74880 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_781
timestamp 1679581782
transform 1 0 75552 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_788
timestamp 1679581782
transform 1 0 76224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_795
timestamp 1679581782
transform 1 0 76896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_802
timestamp 1679581782
transform 1 0 77568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_809
timestamp 1679581782
transform 1 0 78240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_816
timestamp 1679581782
transform 1 0 78912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_823
timestamp 1679581782
transform 1 0 79584 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_830
timestamp 1679581782
transform 1 0 80256 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_837
timestamp 1679581782
transform 1 0 80928 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_844
timestamp 1679581782
transform 1 0 81600 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_851
timestamp 1679581782
transform 1 0 82272 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_858
timestamp 1679581782
transform 1 0 82944 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_865
timestamp 1679581782
transform 1 0 83616 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_872
timestamp 1679581782
transform 1 0 84288 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_879
timestamp 1679581782
transform 1 0 84960 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_886
timestamp 1679581782
transform 1 0 85632 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_893
timestamp 1679581782
transform 1 0 86304 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_900
timestamp 1679581782
transform 1 0 86976 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_907
timestamp 1679581782
transform 1 0 87648 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_914
timestamp 1679581782
transform 1 0 88320 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_921
timestamp 1679581782
transform 1 0 88992 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_928
timestamp 1679581782
transform 1 0 89664 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_935
timestamp 1679581782
transform 1 0 90336 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_942
timestamp 1679581782
transform 1 0 91008 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_949
timestamp 1679581782
transform 1 0 91680 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_956
timestamp 1679581782
transform 1 0 92352 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_963
timestamp 1679581782
transform 1 0 93024 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_970
timestamp 1679581782
transform 1 0 93696 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_977
timestamp 1679581782
transform 1 0 94368 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_984
timestamp 1679581782
transform 1 0 95040 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_991
timestamp 1679581782
transform 1 0 95712 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_998
timestamp 1679581782
transform 1 0 96384 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1005
timestamp 1679581782
transform 1 0 97056 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1012
timestamp 1679581782
transform 1 0 97728 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_1019
timestamp 1679581782
transform 1 0 98400 0 1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_1026
timestamp 1677580104
transform 1 0 99072 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_1028
timestamp 1677579658
transform 1 0 99264 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_4
timestamp 1679581782
transform 1 0 960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_11
timestamp 1679581782
transform 1 0 1632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_18
timestamp 1679581782
transform 1 0 2304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_25
timestamp 1679581782
transform 1 0 2976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_32
timestamp 1679581782
transform 1 0 3648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_39
timestamp 1679581782
transform 1 0 4320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_46
timestamp 1679581782
transform 1 0 4992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_53
timestamp 1679581782
transform 1 0 5664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_60
timestamp 1679581782
transform 1 0 6336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_67
timestamp 1679581782
transform 1 0 7008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_74
timestamp 1679581782
transform 1 0 7680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_81
timestamp 1679581782
transform 1 0 8352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_88
timestamp 1679581782
transform 1 0 9024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_95
timestamp 1679581782
transform 1 0 9696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_102
timestamp 1679581782
transform 1 0 10368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_109
timestamp 1679581782
transform 1 0 11040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_116
timestamp 1679581782
transform 1 0 11712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_123
timestamp 1679581782
transform 1 0 12384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_130
timestamp 1679581782
transform 1 0 13056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_137
timestamp 1679581782
transform 1 0 13728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_144
timestamp 1679581782
transform 1 0 14400 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_151
timestamp 1679581782
transform 1 0 15072 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_158
timestamp 1679581782
transform 1 0 15744 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_165
timestamp 1679581782
transform 1 0 16416 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_172
timestamp 1679581782
transform 1 0 17088 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_179
timestamp 1679581782
transform 1 0 17760 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_186
timestamp 1679581782
transform 1 0 18432 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_193
timestamp 1679581782
transform 1 0 19104 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_200
timestamp 1679581782
transform 1 0 19776 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_207
timestamp 1679581782
transform 1 0 20448 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_214
timestamp 1679581782
transform 1 0 21120 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_221
timestamp 1679581782
transform 1 0 21792 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_228
timestamp 1679581782
transform 1 0 22464 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_235
timestamp 1679581782
transform 1 0 23136 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_242
timestamp 1679581782
transform 1 0 23808 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_249
timestamp 1679581782
transform 1 0 24480 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_256
timestamp 1679581782
transform 1 0 25152 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_263
timestamp 1679581782
transform 1 0 25824 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_270
timestamp 1679581782
transform 1 0 26496 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_277
timestamp 1679581782
transform 1 0 27168 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_284
timestamp 1679581782
transform 1 0 27840 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_291
timestamp 1679581782
transform 1 0 28512 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_298
timestamp 1679581782
transform 1 0 29184 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_305
timestamp 1679581782
transform 1 0 29856 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_312
timestamp 1679581782
transform 1 0 30528 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_319
timestamp 1679581782
transform 1 0 31200 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_326
timestamp 1679581782
transform 1 0 31872 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_333
timestamp 1679581782
transform 1 0 32544 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_340
timestamp 1679581782
transform 1 0 33216 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_347
timestamp 1679581782
transform 1 0 33888 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_354
timestamp 1679581782
transform 1 0 34560 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_361
timestamp 1679581782
transform 1 0 35232 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_368
timestamp 1679581782
transform 1 0 35904 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_375
timestamp 1679581782
transform 1 0 36576 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_382
timestamp 1679581782
transform 1 0 37248 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_389
timestamp 1679581782
transform 1 0 37920 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_396
timestamp 1679581782
transform 1 0 38592 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_403
timestamp 1679581782
transform 1 0 39264 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_410
timestamp 1679581782
transform 1 0 39936 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_417
timestamp 1679581782
transform 1 0 40608 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_424
timestamp 1679581782
transform 1 0 41280 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_431
timestamp 1679581782
transform 1 0 41952 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_438
timestamp 1679581782
transform 1 0 42624 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_445
timestamp 1679581782
transform 1 0 43296 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_452
timestamp 1679581782
transform 1 0 43968 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_459
timestamp 1679581782
transform 1 0 44640 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_466
timestamp 1679581782
transform 1 0 45312 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_473
timestamp 1679581782
transform 1 0 45984 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_480
timestamp 1679581782
transform 1 0 46656 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_487
timestamp 1679581782
transform 1 0 47328 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_494
timestamp 1679581782
transform 1 0 48000 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_501
timestamp 1679581782
transform 1 0 48672 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_508
timestamp 1679581782
transform 1 0 49344 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_515
timestamp 1679581782
transform 1 0 50016 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_522
timestamp 1679581782
transform 1 0 50688 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_529
timestamp 1679581782
transform 1 0 51360 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_536
timestamp 1679581782
transform 1 0 52032 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_543
timestamp 1679581782
transform 1 0 52704 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_550
timestamp 1679581782
transform 1 0 53376 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_557
timestamp 1679581782
transform 1 0 54048 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_564
timestamp 1679581782
transform 1 0 54720 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_571
timestamp 1679581782
transform 1 0 55392 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_578
timestamp 1679581782
transform 1 0 56064 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_585
timestamp 1679581782
transform 1 0 56736 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_592
timestamp 1679581782
transform 1 0 57408 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_599
timestamp 1679581782
transform 1 0 58080 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_606
timestamp 1679581782
transform 1 0 58752 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_613
timestamp 1679581782
transform 1 0 59424 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_620
timestamp 1679581782
transform 1 0 60096 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_627
timestamp 1679581782
transform 1 0 60768 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_634
timestamp 1679581782
transform 1 0 61440 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_641
timestamp 1679581782
transform 1 0 62112 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_648
timestamp 1679581782
transform 1 0 62784 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_655
timestamp 1679581782
transform 1 0 63456 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_662
timestamp 1679581782
transform 1 0 64128 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_669
timestamp 1679581782
transform 1 0 64800 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_676
timestamp 1679581782
transform 1 0 65472 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_683
timestamp 1679581782
transform 1 0 66144 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_690
timestamp 1679581782
transform 1 0 66816 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_697
timestamp 1679581782
transform 1 0 67488 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_704
timestamp 1679581782
transform 1 0 68160 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_711
timestamp 1679581782
transform 1 0 68832 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_718
timestamp 1679581782
transform 1 0 69504 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_725
timestamp 1679581782
transform 1 0 70176 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_732
timestamp 1679581782
transform 1 0 70848 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_739
timestamp 1679581782
transform 1 0 71520 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_746
timestamp 1679581782
transform 1 0 72192 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_753
timestamp 1679581782
transform 1 0 72864 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_760
timestamp 1679581782
transform 1 0 73536 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_767
timestamp 1679581782
transform 1 0 74208 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_774
timestamp 1679581782
transform 1 0 74880 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_781
timestamp 1679581782
transform 1 0 75552 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_788
timestamp 1679581782
transform 1 0 76224 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_795
timestamp 1679581782
transform 1 0 76896 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_802
timestamp 1679581782
transform 1 0 77568 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_809
timestamp 1679581782
transform 1 0 78240 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_816
timestamp 1679581782
transform 1 0 78912 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_823
timestamp 1679581782
transform 1 0 79584 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_830
timestamp 1679581782
transform 1 0 80256 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_837
timestamp 1679581782
transform 1 0 80928 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_844
timestamp 1679581782
transform 1 0 81600 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_851
timestamp 1679581782
transform 1 0 82272 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_858
timestamp 1679581782
transform 1 0 82944 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_865
timestamp 1679581782
transform 1 0 83616 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_872
timestamp 1679581782
transform 1 0 84288 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_879
timestamp 1679581782
transform 1 0 84960 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_886
timestamp 1679581782
transform 1 0 85632 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_893
timestamp 1679581782
transform 1 0 86304 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_900
timestamp 1679581782
transform 1 0 86976 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_907
timestamp 1679581782
transform 1 0 87648 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_914
timestamp 1679581782
transform 1 0 88320 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_921
timestamp 1679581782
transform 1 0 88992 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_928
timestamp 1679581782
transform 1 0 89664 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_935
timestamp 1679581782
transform 1 0 90336 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_942
timestamp 1679581782
transform 1 0 91008 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_949
timestamp 1679581782
transform 1 0 91680 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_956
timestamp 1679581782
transform 1 0 92352 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_963
timestamp 1679581782
transform 1 0 93024 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_970
timestamp 1679581782
transform 1 0 93696 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_977
timestamp 1679581782
transform 1 0 94368 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_984
timestamp 1679581782
transform 1 0 95040 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_991
timestamp 1679581782
transform 1 0 95712 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_998
timestamp 1679581782
transform 1 0 96384 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1005
timestamp 1679581782
transform 1 0 97056 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1012
timestamp 1679581782
transform 1 0 97728 0 -1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_1019
timestamp 1679581782
transform 1 0 98400 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_1026
timestamp 1677580104
transform 1 0 99072 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_1028
timestamp 1677579658
transform 1 0 99264 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_8
timestamp 1679581782
transform 1 0 1344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_15
timestamp 1679581782
transform 1 0 2016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_22
timestamp 1679581782
transform 1 0 2688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_29
timestamp 1679581782
transform 1 0 3360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_36
timestamp 1679581782
transform 1 0 4032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_43
timestamp 1679581782
transform 1 0 4704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_50
timestamp 1679581782
transform 1 0 5376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_57
timestamp 1679581782
transform 1 0 6048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_64
timestamp 1679581782
transform 1 0 6720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_71
timestamp 1679581782
transform 1 0 7392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_78
timestamp 1679581782
transform 1 0 8064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_85
timestamp 1679581782
transform 1 0 8736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_92
timestamp 1679581782
transform 1 0 9408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_99
timestamp 1679581782
transform 1 0 10080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_106
timestamp 1679581782
transform 1 0 10752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_113
timestamp 1679581782
transform 1 0 11424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_120
timestamp 1679581782
transform 1 0 12096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_127
timestamp 1679581782
transform 1 0 12768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_134
timestamp 1679581782
transform 1 0 13440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_141
timestamp 1679581782
transform 1 0 14112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_148
timestamp 1679581782
transform 1 0 14784 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_155
timestamp 1679581782
transform 1 0 15456 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_162
timestamp 1679581782
transform 1 0 16128 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_169
timestamp 1679581782
transform 1 0 16800 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_176
timestamp 1679581782
transform 1 0 17472 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_183
timestamp 1679581782
transform 1 0 18144 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_190
timestamp 1679581782
transform 1 0 18816 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_197
timestamp 1679581782
transform 1 0 19488 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_204
timestamp 1679581782
transform 1 0 20160 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_211
timestamp 1679581782
transform 1 0 20832 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_218
timestamp 1679581782
transform 1 0 21504 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_225
timestamp 1679581782
transform 1 0 22176 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_232
timestamp 1679581782
transform 1 0 22848 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_239
timestamp 1679581782
transform 1 0 23520 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_246
timestamp 1679581782
transform 1 0 24192 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_253
timestamp 1679581782
transform 1 0 24864 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_260
timestamp 1679581782
transform 1 0 25536 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_267
timestamp 1679581782
transform 1 0 26208 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_274
timestamp 1679581782
transform 1 0 26880 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_281
timestamp 1679581782
transform 1 0 27552 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_288
timestamp 1679581782
transform 1 0 28224 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_295
timestamp 1679581782
transform 1 0 28896 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_302
timestamp 1679581782
transform 1 0 29568 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_309
timestamp 1679581782
transform 1 0 30240 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_316
timestamp 1679581782
transform 1 0 30912 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_323
timestamp 1679581782
transform 1 0 31584 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_330
timestamp 1679581782
transform 1 0 32256 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_337
timestamp 1679581782
transform 1 0 32928 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_344
timestamp 1679581782
transform 1 0 33600 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_351
timestamp 1679581782
transform 1 0 34272 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_358
timestamp 1679581782
transform 1 0 34944 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_365
timestamp 1679581782
transform 1 0 35616 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_372
timestamp 1679581782
transform 1 0 36288 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_379
timestamp 1679581782
transform 1 0 36960 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_386
timestamp 1679581782
transform 1 0 37632 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_393
timestamp 1679581782
transform 1 0 38304 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_400
timestamp 1679581782
transform 1 0 38976 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_407
timestamp 1679581782
transform 1 0 39648 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_414
timestamp 1679581782
transform 1 0 40320 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_421
timestamp 1679581782
transform 1 0 40992 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_428
timestamp 1679581782
transform 1 0 41664 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_435
timestamp 1679581782
transform 1 0 42336 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_442
timestamp 1679581782
transform 1 0 43008 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_449
timestamp 1679581782
transform 1 0 43680 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_456
timestamp 1679581782
transform 1 0 44352 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_463
timestamp 1679581782
transform 1 0 45024 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_470
timestamp 1679581782
transform 1 0 45696 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_477
timestamp 1679581782
transform 1 0 46368 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_484
timestamp 1679581782
transform 1 0 47040 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_491
timestamp 1679581782
transform 1 0 47712 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_498
timestamp 1679581782
transform 1 0 48384 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_505
timestamp 1679581782
transform 1 0 49056 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_512
timestamp 1679581782
transform 1 0 49728 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_519
timestamp 1679581782
transform 1 0 50400 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_526
timestamp 1679581782
transform 1 0 51072 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_533
timestamp 1679581782
transform 1 0 51744 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_540
timestamp 1679581782
transform 1 0 52416 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_547
timestamp 1679581782
transform 1 0 53088 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_554
timestamp 1679581782
transform 1 0 53760 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_561
timestamp 1679581782
transform 1 0 54432 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_568
timestamp 1679581782
transform 1 0 55104 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_575
timestamp 1679581782
transform 1 0 55776 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_582
timestamp 1679581782
transform 1 0 56448 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_589
timestamp 1679581782
transform 1 0 57120 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_596
timestamp 1679581782
transform 1 0 57792 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_603
timestamp 1679581782
transform 1 0 58464 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_610
timestamp 1679581782
transform 1 0 59136 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_617
timestamp 1679581782
transform 1 0 59808 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_624
timestamp 1679581782
transform 1 0 60480 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_631
timestamp 1679581782
transform 1 0 61152 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_638
timestamp 1679581782
transform 1 0 61824 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_645
timestamp 1679581782
transform 1 0 62496 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_652
timestamp 1679581782
transform 1 0 63168 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_659
timestamp 1679581782
transform 1 0 63840 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_666
timestamp 1679581782
transform 1 0 64512 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_673
timestamp 1679581782
transform 1 0 65184 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_680
timestamp 1679581782
transform 1 0 65856 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_687
timestamp 1679581782
transform 1 0 66528 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_694
timestamp 1679581782
transform 1 0 67200 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_701
timestamp 1679581782
transform 1 0 67872 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_708
timestamp 1679581782
transform 1 0 68544 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_715
timestamp 1679581782
transform 1 0 69216 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_722
timestamp 1679581782
transform 1 0 69888 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_729
timestamp 1679581782
transform 1 0 70560 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_736
timestamp 1679581782
transform 1 0 71232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_743
timestamp 1679581782
transform 1 0 71904 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_750
timestamp 1679581782
transform 1 0 72576 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_757
timestamp 1679581782
transform 1 0 73248 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_764
timestamp 1679581782
transform 1 0 73920 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_771
timestamp 1679581782
transform 1 0 74592 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_778
timestamp 1679581782
transform 1 0 75264 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_785
timestamp 1679581782
transform 1 0 75936 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_792
timestamp 1679581782
transform 1 0 76608 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_799
timestamp 1679581782
transform 1 0 77280 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_806
timestamp 1679581782
transform 1 0 77952 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_813
timestamp 1679581782
transform 1 0 78624 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_820
timestamp 1679581782
transform 1 0 79296 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_827
timestamp 1679581782
transform 1 0 79968 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_834
timestamp 1679581782
transform 1 0 80640 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_841
timestamp 1679581782
transform 1 0 81312 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_848
timestamp 1679581782
transform 1 0 81984 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_855
timestamp 1679581782
transform 1 0 82656 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_862
timestamp 1679581782
transform 1 0 83328 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_869
timestamp 1679581782
transform 1 0 84000 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_876
timestamp 1679581782
transform 1 0 84672 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_883
timestamp 1679581782
transform 1 0 85344 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_890
timestamp 1679581782
transform 1 0 86016 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_897
timestamp 1679581782
transform 1 0 86688 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_904
timestamp 1679581782
transform 1 0 87360 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_911
timestamp 1679581782
transform 1 0 88032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_918
timestamp 1679581782
transform 1 0 88704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_925
timestamp 1679581782
transform 1 0 89376 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_932
timestamp 1679581782
transform 1 0 90048 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_939
timestamp 1679581782
transform 1 0 90720 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_946
timestamp 1679581782
transform 1 0 91392 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_953
timestamp 1679581782
transform 1 0 92064 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_960
timestamp 1679581782
transform 1 0 92736 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_967
timestamp 1679581782
transform 1 0 93408 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_974
timestamp 1679581782
transform 1 0 94080 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_981
timestamp 1679581782
transform 1 0 94752 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_988
timestamp 1679581782
transform 1 0 95424 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_995
timestamp 1679581782
transform 1 0 96096 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1002
timestamp 1679581782
transform 1 0 96768 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1009
timestamp 1679581782
transform 1 0 97440 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_1016
timestamp 1679581782
transform 1 0 98112 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_1023
timestamp 1679577901
transform 1 0 98784 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_1027
timestamp 1677580104
transform 1 0 99168 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_0
timestamp 1677580104
transform 1 0 576 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_5_18
timestamp 1679581782
transform 1 0 2304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_25
timestamp 1679581782
transform 1 0 2976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_32
timestamp 1679581782
transform 1 0 3648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_39
timestamp 1679581782
transform 1 0 4320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_46
timestamp 1679581782
transform 1 0 4992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_53
timestamp 1679581782
transform 1 0 5664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_60
timestamp 1679581782
transform 1 0 6336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_67
timestamp 1679581782
transform 1 0 7008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_74
timestamp 1679581782
transform 1 0 7680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_81
timestamp 1679581782
transform 1 0 8352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_88
timestamp 1679581782
transform 1 0 9024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_95
timestamp 1679581782
transform 1 0 9696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_102
timestamp 1679581782
transform 1 0 10368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_109
timestamp 1679581782
transform 1 0 11040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_116
timestamp 1679581782
transform 1 0 11712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_123
timestamp 1679581782
transform 1 0 12384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_130
timestamp 1679581782
transform 1 0 13056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_137
timestamp 1679581782
transform 1 0 13728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_144
timestamp 1679581782
transform 1 0 14400 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_151
timestamp 1679581782
transform 1 0 15072 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_158
timestamp 1679581782
transform 1 0 15744 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_165
timestamp 1679581782
transform 1 0 16416 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_172
timestamp 1679581782
transform 1 0 17088 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_179
timestamp 1679581782
transform 1 0 17760 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_186
timestamp 1679581782
transform 1 0 18432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_193
timestamp 1679581782
transform 1 0 19104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_200
timestamp 1679581782
transform 1 0 19776 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_207
timestamp 1679581782
transform 1 0 20448 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_214
timestamp 1679581782
transform 1 0 21120 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_221
timestamp 1679581782
transform 1 0 21792 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_228
timestamp 1679581782
transform 1 0 22464 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_235
timestamp 1679581782
transform 1 0 23136 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_242
timestamp 1679581782
transform 1 0 23808 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_249
timestamp 1679581782
transform 1 0 24480 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_256
timestamp 1679581782
transform 1 0 25152 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_263
timestamp 1679581782
transform 1 0 25824 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_270
timestamp 1679581782
transform 1 0 26496 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_277
timestamp 1679581782
transform 1 0 27168 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_284
timestamp 1679581782
transform 1 0 27840 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_291
timestamp 1679581782
transform 1 0 28512 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_298
timestamp 1679581782
transform 1 0 29184 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_305
timestamp 1679581782
transform 1 0 29856 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_312
timestamp 1679581782
transform 1 0 30528 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_319
timestamp 1679581782
transform 1 0 31200 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_326
timestamp 1679581782
transform 1 0 31872 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_333
timestamp 1679581782
transform 1 0 32544 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_340
timestamp 1679581782
transform 1 0 33216 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_347
timestamp 1679581782
transform 1 0 33888 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_354
timestamp 1679581782
transform 1 0 34560 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_361
timestamp 1679581782
transform 1 0 35232 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_368
timestamp 1679581782
transform 1 0 35904 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_375
timestamp 1679581782
transform 1 0 36576 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_382
timestamp 1679581782
transform 1 0 37248 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_389
timestamp 1679581782
transform 1 0 37920 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_396
timestamp 1679581782
transform 1 0 38592 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_403
timestamp 1679581782
transform 1 0 39264 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_410
timestamp 1679581782
transform 1 0 39936 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_417
timestamp 1679581782
transform 1 0 40608 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_424
timestamp 1679581782
transform 1 0 41280 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_431
timestamp 1679581782
transform 1 0 41952 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_438
timestamp 1679581782
transform 1 0 42624 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_445
timestamp 1679581782
transform 1 0 43296 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_452
timestamp 1679581782
transform 1 0 43968 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_459
timestamp 1679581782
transform 1 0 44640 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_466
timestamp 1679581782
transform 1 0 45312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_473
timestamp 1679581782
transform 1 0 45984 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_480
timestamp 1679581782
transform 1 0 46656 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_487
timestamp 1679581782
transform 1 0 47328 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_494
timestamp 1679581782
transform 1 0 48000 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_501
timestamp 1679581782
transform 1 0 48672 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_508
timestamp 1679581782
transform 1 0 49344 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_515
timestamp 1679581782
transform 1 0 50016 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_522
timestamp 1679581782
transform 1 0 50688 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_529
timestamp 1679581782
transform 1 0 51360 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_536
timestamp 1679581782
transform 1 0 52032 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_543
timestamp 1679581782
transform 1 0 52704 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_550
timestamp 1679581782
transform 1 0 53376 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_557
timestamp 1679581782
transform 1 0 54048 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_564
timestamp 1679581782
transform 1 0 54720 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_571
timestamp 1679581782
transform 1 0 55392 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_578
timestamp 1679581782
transform 1 0 56064 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_585
timestamp 1679581782
transform 1 0 56736 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_592
timestamp 1679581782
transform 1 0 57408 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_599
timestamp 1679581782
transform 1 0 58080 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_606
timestamp 1679581782
transform 1 0 58752 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_613
timestamp 1679581782
transform 1 0 59424 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_620
timestamp 1679581782
transform 1 0 60096 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_627
timestamp 1679581782
transform 1 0 60768 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_634
timestamp 1679581782
transform 1 0 61440 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_641
timestamp 1679581782
transform 1 0 62112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_648
timestamp 1679581782
transform 1 0 62784 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_655
timestamp 1679581782
transform 1 0 63456 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_662
timestamp 1679581782
transform 1 0 64128 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_669
timestamp 1679581782
transform 1 0 64800 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_676
timestamp 1679581782
transform 1 0 65472 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_683
timestamp 1679581782
transform 1 0 66144 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_690
timestamp 1679581782
transform 1 0 66816 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_697
timestamp 1679581782
transform 1 0 67488 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_704
timestamp 1679581782
transform 1 0 68160 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_711
timestamp 1679581782
transform 1 0 68832 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_718
timestamp 1679581782
transform 1 0 69504 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_725
timestamp 1679581782
transform 1 0 70176 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_732
timestamp 1679581782
transform 1 0 70848 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_739
timestamp 1679581782
transform 1 0 71520 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_746
timestamp 1679581782
transform 1 0 72192 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_753
timestamp 1679581782
transform 1 0 72864 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_760
timestamp 1679581782
transform 1 0 73536 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_767
timestamp 1679581782
transform 1 0 74208 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_774
timestamp 1679581782
transform 1 0 74880 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_781
timestamp 1679581782
transform 1 0 75552 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_788
timestamp 1679581782
transform 1 0 76224 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_795
timestamp 1679581782
transform 1 0 76896 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_802
timestamp 1679581782
transform 1 0 77568 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_809
timestamp 1679581782
transform 1 0 78240 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_816
timestamp 1679581782
transform 1 0 78912 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_823
timestamp 1679581782
transform 1 0 79584 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_830
timestamp 1679581782
transform 1 0 80256 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_837
timestamp 1679581782
transform 1 0 80928 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_844
timestamp 1679581782
transform 1 0 81600 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_851
timestamp 1679581782
transform 1 0 82272 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_858
timestamp 1679581782
transform 1 0 82944 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_865
timestamp 1679581782
transform 1 0 83616 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_872
timestamp 1679581782
transform 1 0 84288 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_879
timestamp 1679581782
transform 1 0 84960 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_886
timestamp 1679581782
transform 1 0 85632 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_893
timestamp 1679581782
transform 1 0 86304 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_900
timestamp 1679581782
transform 1 0 86976 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_907
timestamp 1679581782
transform 1 0 87648 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_914
timestamp 1679581782
transform 1 0 88320 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_921
timestamp 1679581782
transform 1 0 88992 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_928
timestamp 1679581782
transform 1 0 89664 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_935
timestamp 1679581782
transform 1 0 90336 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_942
timestamp 1679581782
transform 1 0 91008 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_949
timestamp 1679581782
transform 1 0 91680 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_956
timestamp 1679581782
transform 1 0 92352 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_963
timestamp 1679581782
transform 1 0 93024 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_970
timestamp 1679581782
transform 1 0 93696 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_977
timestamp 1679581782
transform 1 0 94368 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_984
timestamp 1679581782
transform 1 0 95040 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_991
timestamp 1679581782
transform 1 0 95712 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_998
timestamp 1679581782
transform 1 0 96384 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1005
timestamp 1679581782
transform 1 0 97056 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1012
timestamp 1679581782
transform 1 0 97728 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_1019
timestamp 1679581782
transform 1 0 98400 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_1026
timestamp 1677580104
transform 1 0 99072 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_1028
timestamp 1677579658
transform 1 0 99264 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_4
timestamp 1679581782
transform 1 0 960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_11
timestamp 1679581782
transform 1 0 1632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_18
timestamp 1679581782
transform 1 0 2304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_25
timestamp 1679581782
transform 1 0 2976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_32
timestamp 1679581782
transform 1 0 3648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_39
timestamp 1679581782
transform 1 0 4320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_46
timestamp 1679581782
transform 1 0 4992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_53
timestamp 1679581782
transform 1 0 5664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_60
timestamp 1679581782
transform 1 0 6336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_67
timestamp 1679581782
transform 1 0 7008 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_74
timestamp 1679581782
transform 1 0 7680 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_81
timestamp 1679581782
transform 1 0 8352 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_88
timestamp 1679581782
transform 1 0 9024 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_95
timestamp 1679581782
transform 1 0 9696 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_102
timestamp 1679581782
transform 1 0 10368 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_109
timestamp 1679581782
transform 1 0 11040 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_116
timestamp 1679581782
transform 1 0 11712 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_123
timestamp 1679581782
transform 1 0 12384 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_130
timestamp 1679581782
transform 1 0 13056 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_137
timestamp 1679581782
transform 1 0 13728 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_144
timestamp 1679581782
transform 1 0 14400 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_151
timestamp 1679581782
transform 1 0 15072 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_158
timestamp 1679581782
transform 1 0 15744 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_165
timestamp 1679581782
transform 1 0 16416 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_172
timestamp 1679581782
transform 1 0 17088 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_179
timestamp 1679581782
transform 1 0 17760 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_186
timestamp 1679581782
transform 1 0 18432 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_193
timestamp 1679581782
transform 1 0 19104 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_200
timestamp 1679581782
transform 1 0 19776 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_207
timestamp 1679581782
transform 1 0 20448 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_214
timestamp 1679581782
transform 1 0 21120 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_221
timestamp 1679581782
transform 1 0 21792 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_228
timestamp 1679581782
transform 1 0 22464 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_235
timestamp 1679581782
transform 1 0 23136 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_242
timestamp 1679581782
transform 1 0 23808 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_249
timestamp 1679581782
transform 1 0 24480 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_256
timestamp 1679581782
transform 1 0 25152 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_263
timestamp 1679581782
transform 1 0 25824 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_270
timestamp 1679581782
transform 1 0 26496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_277
timestamp 1679581782
transform 1 0 27168 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_284
timestamp 1679581782
transform 1 0 27840 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_291
timestamp 1679581782
transform 1 0 28512 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_298
timestamp 1679581782
transform 1 0 29184 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_305
timestamp 1679581782
transform 1 0 29856 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_312
timestamp 1679581782
transform 1 0 30528 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_319
timestamp 1679581782
transform 1 0 31200 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_326
timestamp 1679581782
transform 1 0 31872 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_333
timestamp 1679581782
transform 1 0 32544 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_340
timestamp 1679581782
transform 1 0 33216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_347
timestamp 1679581782
transform 1 0 33888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_354
timestamp 1679581782
transform 1 0 34560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_361
timestamp 1679581782
transform 1 0 35232 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_368
timestamp 1679581782
transform 1 0 35904 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_375
timestamp 1679581782
transform 1 0 36576 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_382
timestamp 1679581782
transform 1 0 37248 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_389
timestamp 1679581782
transform 1 0 37920 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_396
timestamp 1679581782
transform 1 0 38592 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_403
timestamp 1679581782
transform 1 0 39264 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_410
timestamp 1679581782
transform 1 0 39936 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_417
timestamp 1679581782
transform 1 0 40608 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_424
timestamp 1679581782
transform 1 0 41280 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_431
timestamp 1679581782
transform 1 0 41952 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_438
timestamp 1679581782
transform 1 0 42624 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_445
timestamp 1679581782
transform 1 0 43296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_452
timestamp 1679581782
transform 1 0 43968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_459
timestamp 1679581782
transform 1 0 44640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_466
timestamp 1679581782
transform 1 0 45312 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_473
timestamp 1679581782
transform 1 0 45984 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_480
timestamp 1679581782
transform 1 0 46656 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_487
timestamp 1679581782
transform 1 0 47328 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_494
timestamp 1679581782
transform 1 0 48000 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_501
timestamp 1679581782
transform 1 0 48672 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_508
timestamp 1679581782
transform 1 0 49344 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_515
timestamp 1679581782
transform 1 0 50016 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_522
timestamp 1679581782
transform 1 0 50688 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_529
timestamp 1679581782
transform 1 0 51360 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_536
timestamp 1679581782
transform 1 0 52032 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_543
timestamp 1679581782
transform 1 0 52704 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_550
timestamp 1679581782
transform 1 0 53376 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_557
timestamp 1679581782
transform 1 0 54048 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_564
timestamp 1679581782
transform 1 0 54720 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_571
timestamp 1679581782
transform 1 0 55392 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_578
timestamp 1679581782
transform 1 0 56064 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_585
timestamp 1679581782
transform 1 0 56736 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_592
timestamp 1679581782
transform 1 0 57408 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_599
timestamp 1679581782
transform 1 0 58080 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_606
timestamp 1679581782
transform 1 0 58752 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_613
timestamp 1679581782
transform 1 0 59424 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_620
timestamp 1679581782
transform 1 0 60096 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_627
timestamp 1679581782
transform 1 0 60768 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_634
timestamp 1679581782
transform 1 0 61440 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_641
timestamp 1679581782
transform 1 0 62112 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_648
timestamp 1679581782
transform 1 0 62784 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_655
timestamp 1679581782
transform 1 0 63456 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_662
timestamp 1679581782
transform 1 0 64128 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_669
timestamp 1679581782
transform 1 0 64800 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_676
timestamp 1679581782
transform 1 0 65472 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_683
timestamp 1679581782
transform 1 0 66144 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_690
timestamp 1679581782
transform 1 0 66816 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_697
timestamp 1679581782
transform 1 0 67488 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_704
timestamp 1679581782
transform 1 0 68160 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_711
timestamp 1679581782
transform 1 0 68832 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_718
timestamp 1679581782
transform 1 0 69504 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_725
timestamp 1679581782
transform 1 0 70176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_732
timestamp 1679581782
transform 1 0 70848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_739
timestamp 1679581782
transform 1 0 71520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_746
timestamp 1679581782
transform 1 0 72192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_753
timestamp 1679581782
transform 1 0 72864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_760
timestamp 1679581782
transform 1 0 73536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_767
timestamp 1679581782
transform 1 0 74208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_774
timestamp 1679581782
transform 1 0 74880 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_781
timestamp 1679581782
transform 1 0 75552 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_788
timestamp 1679581782
transform 1 0 76224 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_795
timestamp 1679581782
transform 1 0 76896 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_802
timestamp 1679581782
transform 1 0 77568 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_809
timestamp 1679581782
transform 1 0 78240 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_816
timestamp 1679581782
transform 1 0 78912 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_823
timestamp 1679581782
transform 1 0 79584 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_830
timestamp 1679577901
transform 1 0 80256 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_834
timestamp 1677580104
transform 1 0 80640 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_840
timestamp 1679581782
transform 1 0 81216 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_847
timestamp 1679581782
transform 1 0 81888 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_854
timestamp 1679581782
transform 1 0 82560 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_865
timestamp 1679581782
transform 1 0 83616 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_872
timestamp 1679581782
transform 1 0 84288 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_879
timestamp 1679581782
transform 1 0 84960 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_886
timestamp 1679581782
transform 1 0 85632 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_893
timestamp 1679581782
transform 1 0 86304 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_900
timestamp 1679581782
transform 1 0 86976 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_907
timestamp 1679581782
transform 1 0 87648 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_914
timestamp 1679581782
transform 1 0 88320 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_921
timestamp 1679581782
transform 1 0 88992 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_928
timestamp 1679581782
transform 1 0 89664 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_935
timestamp 1679581782
transform 1 0 90336 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_945
timestamp 1679581782
transform 1 0 91296 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_952
timestamp 1679581782
transform 1 0 91968 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_959
timestamp 1679581782
transform 1 0 92640 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_966
timestamp 1679577901
transform 1 0 93312 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_970
timestamp 1677580104
transform 1 0 93696 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_975
timestamp 1679581782
transform 1 0 94176 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_982
timestamp 1679581782
transform 1 0 94848 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_989
timestamp 1679581782
transform 1 0 95520 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_996
timestamp 1679581782
transform 1 0 96192 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1003
timestamp 1679581782
transform 1 0 96864 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1010
timestamp 1679581782
transform 1 0 97536 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_1017
timestamp 1679581782
transform 1 0 98208 0 1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_1024
timestamp 1679577901
transform 1 0 98880 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_1028
timestamp 1677579658
transform 1 0 99264 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 576 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_15
timestamp 1679581782
transform 1 0 2016 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_22
timestamp 1679581782
transform 1 0 2688 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_29
timestamp 1679581782
transform 1 0 3360 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_36
timestamp 1679581782
transform 1 0 4032 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_43
timestamp 1679581782
transform 1 0 4704 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_50
timestamp 1679581782
transform 1 0 5376 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_57
timestamp 1679581782
transform 1 0 6048 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_64
timestamp 1679581782
transform 1 0 6720 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_71
timestamp 1679581782
transform 1 0 7392 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_78
timestamp 1679581782
transform 1 0 8064 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_85
timestamp 1679581782
transform 1 0 8736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_92
timestamp 1679581782
transform 1 0 9408 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_99
timestamp 1679581782
transform 1 0 10080 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_106
timestamp 1679581782
transform 1 0 10752 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_113
timestamp 1679581782
transform 1 0 11424 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_120
timestamp 1679581782
transform 1 0 12096 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_127
timestamp 1679581782
transform 1 0 12768 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_134
timestamp 1679581782
transform 1 0 13440 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_141
timestamp 1679581782
transform 1 0 14112 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_148
timestamp 1679581782
transform 1 0 14784 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_155
timestamp 1679581782
transform 1 0 15456 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_162
timestamp 1679581782
transform 1 0 16128 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_169
timestamp 1679581782
transform 1 0 16800 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_176
timestamp 1679581782
transform 1 0 17472 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_183
timestamp 1679581782
transform 1 0 18144 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_190
timestamp 1679581782
transform 1 0 18816 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_197
timestamp 1679581782
transform 1 0 19488 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_204
timestamp 1679581782
transform 1 0 20160 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_211
timestamp 1679581782
transform 1 0 20832 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_218
timestamp 1679581782
transform 1 0 21504 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_225
timestamp 1679581782
transform 1 0 22176 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_232
timestamp 1679581782
transform 1 0 22848 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_239
timestamp 1679581782
transform 1 0 23520 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_246
timestamp 1679581782
transform 1 0 24192 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_253
timestamp 1679581782
transform 1 0 24864 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_260
timestamp 1679581782
transform 1 0 25536 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_267
timestamp 1679581782
transform 1 0 26208 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_274
timestamp 1679581782
transform 1 0 26880 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_281
timestamp 1679581782
transform 1 0 27552 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_288
timestamp 1679581782
transform 1 0 28224 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_295
timestamp 1679581782
transform 1 0 28896 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_302
timestamp 1679581782
transform 1 0 29568 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_309
timestamp 1679581782
transform 1 0 30240 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_316
timestamp 1679581782
transform 1 0 30912 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_323
timestamp 1679581782
transform 1 0 31584 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_330
timestamp 1679581782
transform 1 0 32256 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_337
timestamp 1679581782
transform 1 0 32928 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_344
timestamp 1679581782
transform 1 0 33600 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_351
timestamp 1679581782
transform 1 0 34272 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_358
timestamp 1679581782
transform 1 0 34944 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_365
timestamp 1679581782
transform 1 0 35616 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_372
timestamp 1679581782
transform 1 0 36288 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_379
timestamp 1679581782
transform 1 0 36960 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_386
timestamp 1679581782
transform 1 0 37632 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_393
timestamp 1679581782
transform 1 0 38304 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_400
timestamp 1679581782
transform 1 0 38976 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_407
timestamp 1679581782
transform 1 0 39648 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_414
timestamp 1679581782
transform 1 0 40320 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_421
timestamp 1679581782
transform 1 0 40992 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_428
timestamp 1679581782
transform 1 0 41664 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_435
timestamp 1679581782
transform 1 0 42336 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_442
timestamp 1679581782
transform 1 0 43008 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_449
timestamp 1679581782
transform 1 0 43680 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_456
timestamp 1679581782
transform 1 0 44352 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_463
timestamp 1679581782
transform 1 0 45024 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_470
timestamp 1679581782
transform 1 0 45696 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_477
timestamp 1679581782
transform 1 0 46368 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_484
timestamp 1679581782
transform 1 0 47040 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_491
timestamp 1679581782
transform 1 0 47712 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_498
timestamp 1679581782
transform 1 0 48384 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_505
timestamp 1679581782
transform 1 0 49056 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_512
timestamp 1679581782
transform 1 0 49728 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_519
timestamp 1679581782
transform 1 0 50400 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_526
timestamp 1679581782
transform 1 0 51072 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_533
timestamp 1679581782
transform 1 0 51744 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_540
timestamp 1679581782
transform 1 0 52416 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_547
timestamp 1679581782
transform 1 0 53088 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_554
timestamp 1679581782
transform 1 0 53760 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_561
timestamp 1679581782
transform 1 0 54432 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_568
timestamp 1679581782
transform 1 0 55104 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_575
timestamp 1679581782
transform 1 0 55776 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_582
timestamp 1679581782
transform 1 0 56448 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_589
timestamp 1679581782
transform 1 0 57120 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_596
timestamp 1679581782
transform 1 0 57792 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_603
timestamp 1679581782
transform 1 0 58464 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_610
timestamp 1679581782
transform 1 0 59136 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_617
timestamp 1679581782
transform 1 0 59808 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_624
timestamp 1679581782
transform 1 0 60480 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_631
timestamp 1679581782
transform 1 0 61152 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_638
timestamp 1679581782
transform 1 0 61824 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_645
timestamp 1679581782
transform 1 0 62496 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_652
timestamp 1679581782
transform 1 0 63168 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_659
timestamp 1679581782
transform 1 0 63840 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_666
timestamp 1679581782
transform 1 0 64512 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_673
timestamp 1679581782
transform 1 0 65184 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_680
timestamp 1679581782
transform 1 0 65856 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_687
timestamp 1679581782
transform 1 0 66528 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_694
timestamp 1679581782
transform 1 0 67200 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_701
timestamp 1679581782
transform 1 0 67872 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_708
timestamp 1679581782
transform 1 0 68544 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_715
timestamp 1679581782
transform 1 0 69216 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_722
timestamp 1679581782
transform 1 0 69888 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_729
timestamp 1679581782
transform 1 0 70560 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_736
timestamp 1679581782
transform 1 0 71232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_743
timestamp 1679581782
transform 1 0 71904 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_750
timestamp 1679577901
transform 1 0 72576 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_754
timestamp 1677580104
transform 1 0 72960 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_763
timestamp 1677579658
transform 1 0 73824 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_772
timestamp 1677579658
transform 1 0 74688 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_789
timestamp 1677579658
transform 1 0 76320 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_806
timestamp 1677579658
transform 1 0 77952 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_823
timestamp 1677579658
transform 1 0 79584 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_839
timestamp 1677579658
transform 1 0 81120 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_852
timestamp 1677579658
transform 1 0 82368 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_864
timestamp 1677579658
transform 1 0 83520 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_881
timestamp 1677579658
transform 1 0 85152 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_902
timestamp 1677579658
transform 1 0 87168 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_927
timestamp 1677579658
transform 1 0 89568 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_948
timestamp 1677579658
transform 1 0 91584 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_965
timestamp 1677579658
transform 1 0 93216 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_986
timestamp 1677579658
transform 1 0 95232 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_1003
timestamp 1677579658
transform 1 0 96864 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_1008
timestamp 1677579658
transform 1 0 97344 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_1017
timestamp 1677579658
transform 1 0 98208 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_1021
timestamp 1679581782
transform 1 0 98592 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_1028
timestamp 1677579658
transform 1 0 99264 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_4
timestamp 1679577901
transform 1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_8
timestamp 1677579658
transform 1 0 1344 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_13
timestamp 1679581782
transform 1 0 1824 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_20
timestamp 1679581782
transform 1 0 2496 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_27
timestamp 1679581782
transform 1 0 3168 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_34
timestamp 1679581782
transform 1 0 3840 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_41
timestamp 1679581782
transform 1 0 4512 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_48
timestamp 1679581782
transform 1 0 5184 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_55
timestamp 1679581782
transform 1 0 5856 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_62
timestamp 1679581782
transform 1 0 6528 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_69
timestamp 1679581782
transform 1 0 7200 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_76
timestamp 1679581782
transform 1 0 7872 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_83
timestamp 1679581782
transform 1 0 8544 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_90
timestamp 1679581782
transform 1 0 9216 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_97
timestamp 1679581782
transform 1 0 9888 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_104
timestamp 1679581782
transform 1 0 10560 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_111
timestamp 1679581782
transform 1 0 11232 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_118
timestamp 1679581782
transform 1 0 11904 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_125
timestamp 1679581782
transform 1 0 12576 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_132
timestamp 1679581782
transform 1 0 13248 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_139
timestamp 1679581782
transform 1 0 13920 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_146
timestamp 1679581782
transform 1 0 14592 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_153
timestamp 1679581782
transform 1 0 15264 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_160
timestamp 1679581782
transform 1 0 15936 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_167
timestamp 1679581782
transform 1 0 16608 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_174
timestamp 1679581782
transform 1 0 17280 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_181
timestamp 1679581782
transform 1 0 17952 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_188
timestamp 1679581782
transform 1 0 18624 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_195
timestamp 1679581782
transform 1 0 19296 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_202
timestamp 1679581782
transform 1 0 19968 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_209
timestamp 1679581782
transform 1 0 20640 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_216
timestamp 1679581782
transform 1 0 21312 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_223
timestamp 1679581782
transform 1 0 21984 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_230
timestamp 1679581782
transform 1 0 22656 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_237
timestamp 1679581782
transform 1 0 23328 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_244
timestamp 1679581782
transform 1 0 24000 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_251
timestamp 1679581782
transform 1 0 24672 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_258
timestamp 1679581782
transform 1 0 25344 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_265
timestamp 1679581782
transform 1 0 26016 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_272
timestamp 1679581782
transform 1 0 26688 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_279
timestamp 1679581782
transform 1 0 27360 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_286
timestamp 1679581782
transform 1 0 28032 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_293
timestamp 1679581782
transform 1 0 28704 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_300
timestamp 1679581782
transform 1 0 29376 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_307
timestamp 1679581782
transform 1 0 30048 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_314
timestamp 1679581782
transform 1 0 30720 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_321
timestamp 1679581782
transform 1 0 31392 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_328
timestamp 1679581782
transform 1 0 32064 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_335
timestamp 1679581782
transform 1 0 32736 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_342
timestamp 1679581782
transform 1 0 33408 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_349
timestamp 1679581782
transform 1 0 34080 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_356
timestamp 1679581782
transform 1 0 34752 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_363
timestamp 1679581782
transform 1 0 35424 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_370
timestamp 1679581782
transform 1 0 36096 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_377
timestamp 1679581782
transform 1 0 36768 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_384
timestamp 1679581782
transform 1 0 37440 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_391
timestamp 1679581782
transform 1 0 38112 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_398
timestamp 1679581782
transform 1 0 38784 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_405
timestamp 1679581782
transform 1 0 39456 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_412
timestamp 1679581782
transform 1 0 40128 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_419
timestamp 1679581782
transform 1 0 40800 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_426
timestamp 1679581782
transform 1 0 41472 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_433
timestamp 1679581782
transform 1 0 42144 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_440
timestamp 1679581782
transform 1 0 42816 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_447
timestamp 1679581782
transform 1 0 43488 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_454
timestamp 1679581782
transform 1 0 44160 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_461
timestamp 1679581782
transform 1 0 44832 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_468
timestamp 1679581782
transform 1 0 45504 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_475
timestamp 1679581782
transform 1 0 46176 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_482
timestamp 1679581782
transform 1 0 46848 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_489
timestamp 1679581782
transform 1 0 47520 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_496
timestamp 1679581782
transform 1 0 48192 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_503
timestamp 1679581782
transform 1 0 48864 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_510
timestamp 1679581782
transform 1 0 49536 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_517
timestamp 1679581782
transform 1 0 50208 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_524
timestamp 1679581782
transform 1 0 50880 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_531
timestamp 1679581782
transform 1 0 51552 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_538
timestamp 1679581782
transform 1 0 52224 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_545
timestamp 1679581782
transform 1 0 52896 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_552
timestamp 1679581782
transform 1 0 53568 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_559
timestamp 1679581782
transform 1 0 54240 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_566
timestamp 1679581782
transform 1 0 54912 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_573
timestamp 1679581782
transform 1 0 55584 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_580
timestamp 1679581782
transform 1 0 56256 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_587
timestamp 1679581782
transform 1 0 56928 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_594
timestamp 1679581782
transform 1 0 57600 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_601
timestamp 1679581782
transform 1 0 58272 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_608
timestamp 1679581782
transform 1 0 58944 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_615
timestamp 1679581782
transform 1 0 59616 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_622
timestamp 1679581782
transform 1 0 60288 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_629
timestamp 1679581782
transform 1 0 60960 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_636
timestamp 1679581782
transform 1 0 61632 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_643
timestamp 1679581782
transform 1 0 62304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_650
timestamp 1679581782
transform 1 0 62976 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_657
timestamp 1679581782
transform 1 0 63648 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_664
timestamp 1679581782
transform 1 0 64320 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_671
timestamp 1679581782
transform 1 0 64992 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_678
timestamp 1679581782
transform 1 0 65664 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_685
timestamp 1679581782
transform 1 0 66336 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_692
timestamp 1679581782
transform 1 0 67008 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_699
timestamp 1679581782
transform 1 0 67680 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_706
timestamp 1679581782
transform 1 0 68352 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_713
timestamp 1679581782
transform 1 0 69024 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_720
timestamp 1679581782
transform 1 0 69696 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_727
timestamp 1679581782
transform 1 0 70368 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_734
timestamp 1677580104
transform 1 0 71040 0 1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_739
timestamp 1679577901
transform 1 0 71520 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_743
timestamp 1677579658
transform 1 0 71904 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_751
timestamp 1677580104
transform 1 0 72672 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_763
timestamp 1677580104
transform 1 0 73824 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_779
timestamp 1677579658
transform 1 0 75360 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_796
timestamp 1677579658
transform 1 0 76992 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_813
timestamp 1677579658
transform 1 0 78624 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_841
timestamp 1677580104
transform 1 0 81312 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_859
timestamp 1677579658
transform 1 0 83040 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_876
timestamp 1677579658
transform 1 0 84672 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_952
timestamp 1677579658
transform 1 0 91968 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_983
timestamp 1677580104
transform 1 0 94944 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_1001
timestamp 1677579658
transform 1 0 96672 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_1018
timestamp 1677579658
transform 1 0 98304 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_4
timestamp 1679581782
transform 1 0 960 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_11
timestamp 1679581782
transform 1 0 1632 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_18
timestamp 1679581782
transform 1 0 2304 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_25
timestamp 1679581782
transform 1 0 2976 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_32
timestamp 1679581782
transform 1 0 3648 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_39
timestamp 1679581782
transform 1 0 4320 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_46
timestamp 1679581782
transform 1 0 4992 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_53
timestamp 1679581782
transform 1 0 5664 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_60
timestamp 1679581782
transform 1 0 6336 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_67
timestamp 1679581782
transform 1 0 7008 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_74
timestamp 1679581782
transform 1 0 7680 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_81
timestamp 1679581782
transform 1 0 8352 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_88
timestamp 1679581782
transform 1 0 9024 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_95
timestamp 1679581782
transform 1 0 9696 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_102
timestamp 1679581782
transform 1 0 10368 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_109
timestamp 1679581782
transform 1 0 11040 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_116
timestamp 1679581782
transform 1 0 11712 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_123
timestamp 1679581782
transform 1 0 12384 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_130
timestamp 1679581782
transform 1 0 13056 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_137
timestamp 1679581782
transform 1 0 13728 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_144
timestamp 1679581782
transform 1 0 14400 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_151
timestamp 1679581782
transform 1 0 15072 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_158
timestamp 1679581782
transform 1 0 15744 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_165
timestamp 1679581782
transform 1 0 16416 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_172
timestamp 1679581782
transform 1 0 17088 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_179
timestamp 1679581782
transform 1 0 17760 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_186
timestamp 1679581782
transform 1 0 18432 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_193
timestamp 1679581782
transform 1 0 19104 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_200
timestamp 1679581782
transform 1 0 19776 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_207
timestamp 1679581782
transform 1 0 20448 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_214
timestamp 1679581782
transform 1 0 21120 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_221
timestamp 1679581782
transform 1 0 21792 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_228
timestamp 1679581782
transform 1 0 22464 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_235
timestamp 1679581782
transform 1 0 23136 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_242
timestamp 1679581782
transform 1 0 23808 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_249
timestamp 1679581782
transform 1 0 24480 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_256
timestamp 1679581782
transform 1 0 25152 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_263
timestamp 1679581782
transform 1 0 25824 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_270
timestamp 1679581782
transform 1 0 26496 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_277
timestamp 1679581782
transform 1 0 27168 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_284
timestamp 1679581782
transform 1 0 27840 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_291
timestamp 1679581782
transform 1 0 28512 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_298
timestamp 1679581782
transform 1 0 29184 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_305
timestamp 1679581782
transform 1 0 29856 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_312
timestamp 1679581782
transform 1 0 30528 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_319
timestamp 1679581782
transform 1 0 31200 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_326
timestamp 1679581782
transform 1 0 31872 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_333
timestamp 1679581782
transform 1 0 32544 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_340
timestamp 1679581782
transform 1 0 33216 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_347
timestamp 1679581782
transform 1 0 33888 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_354
timestamp 1679581782
transform 1 0 34560 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_361
timestamp 1679581782
transform 1 0 35232 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_368
timestamp 1679581782
transform 1 0 35904 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_375
timestamp 1679581782
transform 1 0 36576 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_382
timestamp 1679581782
transform 1 0 37248 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_389
timestamp 1679581782
transform 1 0 37920 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_396
timestamp 1679581782
transform 1 0 38592 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_403
timestamp 1679581782
transform 1 0 39264 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_410
timestamp 1679581782
transform 1 0 39936 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_417
timestamp 1679581782
transform 1 0 40608 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_424
timestamp 1679581782
transform 1 0 41280 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_431
timestamp 1679581782
transform 1 0 41952 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_438
timestamp 1679581782
transform 1 0 42624 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_445
timestamp 1679581782
transform 1 0 43296 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_452
timestamp 1679581782
transform 1 0 43968 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_459
timestamp 1679581782
transform 1 0 44640 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_466
timestamp 1679581782
transform 1 0 45312 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_473
timestamp 1679581782
transform 1 0 45984 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_480
timestamp 1679581782
transform 1 0 46656 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_487
timestamp 1679581782
transform 1 0 47328 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_494
timestamp 1679581782
transform 1 0 48000 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_501
timestamp 1679581782
transform 1 0 48672 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_508
timestamp 1679581782
transform 1 0 49344 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_515
timestamp 1679581782
transform 1 0 50016 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_522
timestamp 1679581782
transform 1 0 50688 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_529
timestamp 1679581782
transform 1 0 51360 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_536
timestamp 1679581782
transform 1 0 52032 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_543
timestamp 1679581782
transform 1 0 52704 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_550
timestamp 1679581782
transform 1 0 53376 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_557
timestamp 1679581782
transform 1 0 54048 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_564
timestamp 1679581782
transform 1 0 54720 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_571
timestamp 1679581782
transform 1 0 55392 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_578
timestamp 1679581782
transform 1 0 56064 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_585
timestamp 1679581782
transform 1 0 56736 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_592
timestamp 1679581782
transform 1 0 57408 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_599
timestamp 1679581782
transform 1 0 58080 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_606
timestamp 1679581782
transform 1 0 58752 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_613
timestamp 1679581782
transform 1 0 59424 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_620
timestamp 1679581782
transform 1 0 60096 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_627
timestamp 1679581782
transform 1 0 60768 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_634
timestamp 1679581782
transform 1 0 61440 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_641
timestamp 1679581782
transform 1 0 62112 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_648
timestamp 1679581782
transform 1 0 62784 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_655
timestamp 1679581782
transform 1 0 63456 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_662
timestamp 1679581782
transform 1 0 64128 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_669
timestamp 1679581782
transform 1 0 64800 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_676
timestamp 1679581782
transform 1 0 65472 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_683
timestamp 1679581782
transform 1 0 66144 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_690
timestamp 1679581782
transform 1 0 66816 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_697
timestamp 1679581782
transform 1 0 67488 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_704
timestamp 1679581782
transform 1 0 68160 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_711
timestamp 1679581782
transform 1 0 68832 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_718
timestamp 1679581782
transform 1 0 69504 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_725
timestamp 1679577901
transform 1 0 70176 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_729
timestamp 1677580104
transform 1 0 70560 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_4
timestamp 1677579658
transform 1 0 960 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_17
timestamp 1679581782
transform 1 0 2208 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_24
timestamp 1679581782
transform 1 0 2880 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_31
timestamp 1679581782
transform 1 0 3552 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_38
timestamp 1679581782
transform 1 0 4224 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_45
timestamp 1679581782
transform 1 0 4896 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_52
timestamp 1679581782
transform 1 0 5568 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_59
timestamp 1679581782
transform 1 0 6240 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_66
timestamp 1679581782
transform 1 0 6912 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_73
timestamp 1679581782
transform 1 0 7584 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_80
timestamp 1679581782
transform 1 0 8256 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_87
timestamp 1679581782
transform 1 0 8928 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_94
timestamp 1679581782
transform 1 0 9600 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_101
timestamp 1679581782
transform 1 0 10272 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_108
timestamp 1679581782
transform 1 0 10944 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_115
timestamp 1679581782
transform 1 0 11616 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_122
timestamp 1679581782
transform 1 0 12288 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_129
timestamp 1679581782
transform 1 0 12960 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_136
timestamp 1679581782
transform 1 0 13632 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_143
timestamp 1679581782
transform 1 0 14304 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_150
timestamp 1679581782
transform 1 0 14976 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_157
timestamp 1679581782
transform 1 0 15648 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_164
timestamp 1679581782
transform 1 0 16320 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_171
timestamp 1679581782
transform 1 0 16992 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_178
timestamp 1679581782
transform 1 0 17664 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_185
timestamp 1679581782
transform 1 0 18336 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_192
timestamp 1679581782
transform 1 0 19008 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_199
timestamp 1679581782
transform 1 0 19680 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_206
timestamp 1679581782
transform 1 0 20352 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_213
timestamp 1679581782
transform 1 0 21024 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_220
timestamp 1679581782
transform 1 0 21696 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_227
timestamp 1679581782
transform 1 0 22368 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_234
timestamp 1679581782
transform 1 0 23040 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_241
timestamp 1679581782
transform 1 0 23712 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_248
timestamp 1679581782
transform 1 0 24384 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_255
timestamp 1679581782
transform 1 0 25056 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_262
timestamp 1679581782
transform 1 0 25728 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_269
timestamp 1679581782
transform 1 0 26400 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_276
timestamp 1679581782
transform 1 0 27072 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_283
timestamp 1679581782
transform 1 0 27744 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_290
timestamp 1679581782
transform 1 0 28416 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_297
timestamp 1679581782
transform 1 0 29088 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_304
timestamp 1679581782
transform 1 0 29760 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_311
timestamp 1679581782
transform 1 0 30432 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_318
timestamp 1679581782
transform 1 0 31104 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_325
timestamp 1679581782
transform 1 0 31776 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_332
timestamp 1679581782
transform 1 0 32448 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_339
timestamp 1679581782
transform 1 0 33120 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_346
timestamp 1679581782
transform 1 0 33792 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_353
timestamp 1679581782
transform 1 0 34464 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_360
timestamp 1679581782
transform 1 0 35136 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_367
timestamp 1679581782
transform 1 0 35808 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_374
timestamp 1679581782
transform 1 0 36480 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_381
timestamp 1679581782
transform 1 0 37152 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_388
timestamp 1679581782
transform 1 0 37824 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_395
timestamp 1679581782
transform 1 0 38496 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_402
timestamp 1679581782
transform 1 0 39168 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_409
timestamp 1679581782
transform 1 0 39840 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_416
timestamp 1679581782
transform 1 0 40512 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_423
timestamp 1679581782
transform 1 0 41184 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_430
timestamp 1679581782
transform 1 0 41856 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_437
timestamp 1679581782
transform 1 0 42528 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_444
timestamp 1679581782
transform 1 0 43200 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_451
timestamp 1679581782
transform 1 0 43872 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_458
timestamp 1679581782
transform 1 0 44544 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_465
timestamp 1679581782
transform 1 0 45216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_472
timestamp 1679581782
transform 1 0 45888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_479
timestamp 1679581782
transform 1 0 46560 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_486
timestamp 1679581782
transform 1 0 47232 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_493
timestamp 1679581782
transform 1 0 47904 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_500
timestamp 1679581782
transform 1 0 48576 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_507
timestamp 1679581782
transform 1 0 49248 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_514
timestamp 1679581782
transform 1 0 49920 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_521
timestamp 1679581782
transform 1 0 50592 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_528
timestamp 1679581782
transform 1 0 51264 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_535
timestamp 1679581782
transform 1 0 51936 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_542
timestamp 1679581782
transform 1 0 52608 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_549
timestamp 1679581782
transform 1 0 53280 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_556
timestamp 1679581782
transform 1 0 53952 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_563
timestamp 1679581782
transform 1 0 54624 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_570
timestamp 1679581782
transform 1 0 55296 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_577
timestamp 1679581782
transform 1 0 55968 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_584
timestamp 1679581782
transform 1 0 56640 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_591
timestamp 1679581782
transform 1 0 57312 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_598
timestamp 1679581782
transform 1 0 57984 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_605
timestamp 1679581782
transform 1 0 58656 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_612
timestamp 1679581782
transform 1 0 59328 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_619
timestamp 1679581782
transform 1 0 60000 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_626
timestamp 1679581782
transform 1 0 60672 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_633
timestamp 1679581782
transform 1 0 61344 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_640
timestamp 1679581782
transform 1 0 62016 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_647
timestamp 1679581782
transform 1 0 62688 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_654
timestamp 1679581782
transform 1 0 63360 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_661
timestamp 1679581782
transform 1 0 64032 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_668
timestamp 1679581782
transform 1 0 64704 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_675
timestamp 1679581782
transform 1 0 65376 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_682
timestamp 1679581782
transform 1 0 66048 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_689
timestamp 1679581782
transform 1 0 66720 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_696
timestamp 1679581782
transform 1 0 67392 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_703
timestamp 1679581782
transform 1 0 68064 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_710
timestamp 1679581782
transform 1 0 68736 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_717
timestamp 1679581782
transform 1 0 69408 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_724
timestamp 1679581782
transform 1 0 70080 0 1 8316
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_731
timestamp 1677579658
transform 1 0 70752 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_737
timestamp 1677580104
transform 1 0 71328 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_4
timestamp 1679581782
transform 1 0 960 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_11
timestamp 1679581782
transform 1 0 1632 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_18
timestamp 1679581782
transform 1 0 2304 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_25
timestamp 1679581782
transform 1 0 2976 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_32
timestamp 1679581782
transform 1 0 3648 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_39
timestamp 1679581782
transform 1 0 4320 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_46
timestamp 1679581782
transform 1 0 4992 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_53
timestamp 1679581782
transform 1 0 5664 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_60
timestamp 1679581782
transform 1 0 6336 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_67
timestamp 1679581782
transform 1 0 7008 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_74
timestamp 1679581782
transform 1 0 7680 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_81
timestamp 1679581782
transform 1 0 8352 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_88
timestamp 1679581782
transform 1 0 9024 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_95
timestamp 1679581782
transform 1 0 9696 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_102
timestamp 1679581782
transform 1 0 10368 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_109
timestamp 1679581782
transform 1 0 11040 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_116
timestamp 1679581782
transform 1 0 11712 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_123
timestamp 1679581782
transform 1 0 12384 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_130
timestamp 1679581782
transform 1 0 13056 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_137
timestamp 1679581782
transform 1 0 13728 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_144
timestamp 1679581782
transform 1 0 14400 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_151
timestamp 1679581782
transform 1 0 15072 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_158
timestamp 1679581782
transform 1 0 15744 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_165
timestamp 1679581782
transform 1 0 16416 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_172
timestamp 1679581782
transform 1 0 17088 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_179
timestamp 1679581782
transform 1 0 17760 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_186
timestamp 1679581782
transform 1 0 18432 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_193
timestamp 1679581782
transform 1 0 19104 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_200
timestamp 1679581782
transform 1 0 19776 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_207
timestamp 1679581782
transform 1 0 20448 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_214
timestamp 1679581782
transform 1 0 21120 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_221
timestamp 1679581782
transform 1 0 21792 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_228
timestamp 1679581782
transform 1 0 22464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_235
timestamp 1679581782
transform 1 0 23136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_242
timestamp 1679581782
transform 1 0 23808 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_249
timestamp 1679581782
transform 1 0 24480 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_256
timestamp 1679581782
transform 1 0 25152 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_263
timestamp 1679581782
transform 1 0 25824 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_270
timestamp 1679581782
transform 1 0 26496 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_277
timestamp 1679581782
transform 1 0 27168 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_284
timestamp 1679581782
transform 1 0 27840 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_291
timestamp 1679581782
transform 1 0 28512 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_298
timestamp 1679581782
transform 1 0 29184 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_305
timestamp 1679581782
transform 1 0 29856 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_312
timestamp 1679581782
transform 1 0 30528 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_319
timestamp 1679581782
transform 1 0 31200 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_326
timestamp 1679581782
transform 1 0 31872 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_333
timestamp 1679581782
transform 1 0 32544 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_340
timestamp 1679581782
transform 1 0 33216 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_347
timestamp 1679581782
transform 1 0 33888 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_354
timestamp 1679581782
transform 1 0 34560 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_361
timestamp 1679581782
transform 1 0 35232 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_368
timestamp 1679581782
transform 1 0 35904 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_375
timestamp 1679581782
transform 1 0 36576 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_382
timestamp 1679581782
transform 1 0 37248 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_389
timestamp 1679581782
transform 1 0 37920 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_396
timestamp 1679581782
transform 1 0 38592 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_403
timestamp 1679581782
transform 1 0 39264 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_410
timestamp 1679581782
transform 1 0 39936 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_417
timestamp 1679581782
transform 1 0 40608 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_424
timestamp 1679581782
transform 1 0 41280 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_431
timestamp 1679581782
transform 1 0 41952 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_438
timestamp 1679581782
transform 1 0 42624 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_445
timestamp 1679581782
transform 1 0 43296 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_452
timestamp 1679581782
transform 1 0 43968 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_459
timestamp 1679581782
transform 1 0 44640 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_466
timestamp 1679581782
transform 1 0 45312 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_473
timestamp 1679581782
transform 1 0 45984 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_480
timestamp 1679581782
transform 1 0 46656 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_487
timestamp 1679581782
transform 1 0 47328 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_494
timestamp 1679581782
transform 1 0 48000 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_501
timestamp 1679581782
transform 1 0 48672 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_508
timestamp 1679581782
transform 1 0 49344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_515
timestamp 1679581782
transform 1 0 50016 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_522
timestamp 1679581782
transform 1 0 50688 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_529
timestamp 1679581782
transform 1 0 51360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_536
timestamp 1679581782
transform 1 0 52032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_543
timestamp 1679581782
transform 1 0 52704 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_550
timestamp 1679581782
transform 1 0 53376 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_557
timestamp 1679581782
transform 1 0 54048 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_564
timestamp 1679581782
transform 1 0 54720 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_571
timestamp 1679581782
transform 1 0 55392 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_578
timestamp 1679581782
transform 1 0 56064 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_585
timestamp 1679581782
transform 1 0 56736 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_592
timestamp 1679581782
transform 1 0 57408 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_599
timestamp 1679581782
transform 1 0 58080 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_606
timestamp 1679581782
transform 1 0 58752 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_613
timestamp 1679581782
transform 1 0 59424 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_620
timestamp 1679581782
transform 1 0 60096 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_627
timestamp 1679581782
transform 1 0 60768 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_634
timestamp 1679581782
transform 1 0 61440 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_641
timestamp 1679581782
transform 1 0 62112 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_648
timestamp 1679581782
transform 1 0 62784 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_655
timestamp 1679581782
transform 1 0 63456 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_662
timestamp 1679581782
transform 1 0 64128 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_669
timestamp 1679581782
transform 1 0 64800 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_676
timestamp 1679581782
transform 1 0 65472 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_683
timestamp 1679581782
transform 1 0 66144 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_690
timestamp 1679581782
transform 1 0 66816 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_697
timestamp 1679581782
transform 1 0 67488 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_704
timestamp 1679581782
transform 1 0 68160 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_711
timestamp 1679581782
transform 1 0 68832 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_718
timestamp 1679581782
transform 1 0 69504 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_725
timestamp 1679581782
transform 1 0 70176 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_732
timestamp 1679581782
transform 1 0 70848 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_12
timestamp 1679581782
transform 1 0 1728 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_19
timestamp 1679581782
transform 1 0 2400 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_26
timestamp 1679581782
transform 1 0 3072 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_33
timestamp 1679581782
transform 1 0 3744 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_40
timestamp 1679581782
transform 1 0 4416 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_47
timestamp 1679581782
transform 1 0 5088 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_54
timestamp 1679581782
transform 1 0 5760 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_61
timestamp 1679581782
transform 1 0 6432 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_68
timestamp 1679581782
transform 1 0 7104 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_75
timestamp 1679581782
transform 1 0 7776 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_82
timestamp 1679581782
transform 1 0 8448 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_89
timestamp 1679581782
transform 1 0 9120 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_96
timestamp 1679581782
transform 1 0 9792 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_103
timestamp 1679581782
transform 1 0 10464 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_110
timestamp 1679581782
transform 1 0 11136 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_117
timestamp 1679581782
transform 1 0 11808 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_124
timestamp 1679581782
transform 1 0 12480 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_131
timestamp 1679581782
transform 1 0 13152 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_138
timestamp 1679581782
transform 1 0 13824 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_145
timestamp 1679581782
transform 1 0 14496 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_152
timestamp 1679581782
transform 1 0 15168 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_159
timestamp 1679581782
transform 1 0 15840 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_166
timestamp 1679581782
transform 1 0 16512 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_173
timestamp 1679581782
transform 1 0 17184 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_180
timestamp 1679581782
transform 1 0 17856 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_187
timestamp 1679581782
transform 1 0 18528 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_194
timestamp 1679581782
transform 1 0 19200 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_201
timestamp 1679581782
transform 1 0 19872 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_208
timestamp 1679581782
transform 1 0 20544 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_215
timestamp 1679581782
transform 1 0 21216 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_222
timestamp 1679581782
transform 1 0 21888 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_229
timestamp 1679581782
transform 1 0 22560 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_236
timestamp 1679581782
transform 1 0 23232 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_243
timestamp 1679581782
transform 1 0 23904 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_250
timestamp 1679581782
transform 1 0 24576 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_257
timestamp 1679581782
transform 1 0 25248 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_264
timestamp 1679581782
transform 1 0 25920 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_271
timestamp 1679581782
transform 1 0 26592 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_278
timestamp 1679581782
transform 1 0 27264 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_285
timestamp 1679581782
transform 1 0 27936 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_292
timestamp 1679581782
transform 1 0 28608 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_299
timestamp 1679581782
transform 1 0 29280 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_306
timestamp 1679581782
transform 1 0 29952 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_313
timestamp 1679581782
transform 1 0 30624 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_320
timestamp 1679581782
transform 1 0 31296 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_327
timestamp 1679581782
transform 1 0 31968 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_334
timestamp 1679581782
transform 1 0 32640 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_341
timestamp 1679581782
transform 1 0 33312 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_348
timestamp 1679581782
transform 1 0 33984 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_355
timestamp 1679581782
transform 1 0 34656 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_362
timestamp 1679581782
transform 1 0 35328 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_369
timestamp 1679581782
transform 1 0 36000 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_376
timestamp 1679581782
transform 1 0 36672 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_383
timestamp 1679581782
transform 1 0 37344 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_390
timestamp 1679581782
transform 1 0 38016 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_397
timestamp 1679581782
transform 1 0 38688 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_404
timestamp 1679581782
transform 1 0 39360 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_411
timestamp 1679581782
transform 1 0 40032 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_418
timestamp 1679581782
transform 1 0 40704 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_425
timestamp 1679581782
transform 1 0 41376 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_432
timestamp 1679581782
transform 1 0 42048 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_439
timestamp 1679581782
transform 1 0 42720 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_446
timestamp 1679581782
transform 1 0 43392 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_453
timestamp 1679581782
transform 1 0 44064 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_460
timestamp 1679581782
transform 1 0 44736 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_467
timestamp 1679581782
transform 1 0 45408 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_474
timestamp 1679581782
transform 1 0 46080 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_481
timestamp 1679581782
transform 1 0 46752 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_488
timestamp 1679581782
transform 1 0 47424 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_495
timestamp 1679581782
transform 1 0 48096 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_502
timestamp 1679581782
transform 1 0 48768 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_509
timestamp 1679581782
transform 1 0 49440 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_516
timestamp 1679581782
transform 1 0 50112 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_523
timestamp 1679581782
transform 1 0 50784 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_530
timestamp 1679581782
transform 1 0 51456 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_537
timestamp 1679581782
transform 1 0 52128 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_544
timestamp 1679581782
transform 1 0 52800 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_551
timestamp 1679581782
transform 1 0 53472 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_558
timestamp 1679581782
transform 1 0 54144 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_565
timestamp 1679581782
transform 1 0 54816 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_572
timestamp 1679581782
transform 1 0 55488 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_579
timestamp 1679581782
transform 1 0 56160 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_586
timestamp 1679581782
transform 1 0 56832 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_593
timestamp 1679581782
transform 1 0 57504 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_600
timestamp 1679581782
transform 1 0 58176 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_607
timestamp 1679581782
transform 1 0 58848 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_614
timestamp 1679581782
transform 1 0 59520 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_621
timestamp 1679581782
transform 1 0 60192 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_628
timestamp 1679581782
transform 1 0 60864 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_635
timestamp 1679581782
transform 1 0 61536 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_642
timestamp 1679581782
transform 1 0 62208 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_649
timestamp 1679581782
transform 1 0 62880 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_656
timestamp 1679581782
transform 1 0 63552 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_663
timestamp 1679581782
transform 1 0 64224 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_670
timestamp 1679581782
transform 1 0 64896 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_677
timestamp 1679581782
transform 1 0 65568 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_684
timestamp 1679581782
transform 1 0 66240 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_691
timestamp 1679581782
transform 1 0 66912 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_698
timestamp 1679581782
transform 1 0 67584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_705
timestamp 1679581782
transform 1 0 68256 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_712
timestamp 1679581782
transform 1 0 68928 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_719
timestamp 1679581782
transform 1 0 69600 0 1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_726
timestamp 1679581782
transform 1 0 70272 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_733
timestamp 1679577901
transform 1 0 70944 0 1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_12_737
timestamp 1677580104
transform 1 0 71328 0 1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_13_4
timestamp 1677580104
transform 1 0 960 0 -1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_13_10
timestamp 1679581782
transform 1 0 1536 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_17
timestamp 1679581782
transform 1 0 2208 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_24
timestamp 1679581782
transform 1 0 2880 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_31
timestamp 1679581782
transform 1 0 3552 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_38
timestamp 1679581782
transform 1 0 4224 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_45
timestamp 1679581782
transform 1 0 4896 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_52
timestamp 1679581782
transform 1 0 5568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_59
timestamp 1679581782
transform 1 0 6240 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_66
timestamp 1679581782
transform 1 0 6912 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_73
timestamp 1679581782
transform 1 0 7584 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_80
timestamp 1679581782
transform 1 0 8256 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_87
timestamp 1679581782
transform 1 0 8928 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_94
timestamp 1679581782
transform 1 0 9600 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_101
timestamp 1679581782
transform 1 0 10272 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_108
timestamp 1679581782
transform 1 0 10944 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_115
timestamp 1679581782
transform 1 0 11616 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_122
timestamp 1679581782
transform 1 0 12288 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_129
timestamp 1679581782
transform 1 0 12960 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_136
timestamp 1679581782
transform 1 0 13632 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_143
timestamp 1679581782
transform 1 0 14304 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_150
timestamp 1679581782
transform 1 0 14976 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_157
timestamp 1679581782
transform 1 0 15648 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_164
timestamp 1679581782
transform 1 0 16320 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_171
timestamp 1679581782
transform 1 0 16992 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_178
timestamp 1679581782
transform 1 0 17664 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_185
timestamp 1679581782
transform 1 0 18336 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_192
timestamp 1679581782
transform 1 0 19008 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_199
timestamp 1679581782
transform 1 0 19680 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_206
timestamp 1679581782
transform 1 0 20352 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_213
timestamp 1679581782
transform 1 0 21024 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_220
timestamp 1679581782
transform 1 0 21696 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_227
timestamp 1679581782
transform 1 0 22368 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_234
timestamp 1679581782
transform 1 0 23040 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_241
timestamp 1679581782
transform 1 0 23712 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_248
timestamp 1679581782
transform 1 0 24384 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_255
timestamp 1679581782
transform 1 0 25056 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_262
timestamp 1679581782
transform 1 0 25728 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_269
timestamp 1679581782
transform 1 0 26400 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_276
timestamp 1679581782
transform 1 0 27072 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_283
timestamp 1679581782
transform 1 0 27744 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_290
timestamp 1679581782
transform 1 0 28416 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_297
timestamp 1679581782
transform 1 0 29088 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_304
timestamp 1679581782
transform 1 0 29760 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_311
timestamp 1679581782
transform 1 0 30432 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_318
timestamp 1679581782
transform 1 0 31104 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_325
timestamp 1679581782
transform 1 0 31776 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_332
timestamp 1679581782
transform 1 0 32448 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_339
timestamp 1679581782
transform 1 0 33120 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_346
timestamp 1679581782
transform 1 0 33792 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_353
timestamp 1679581782
transform 1 0 34464 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_360
timestamp 1679581782
transform 1 0 35136 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_367
timestamp 1679581782
transform 1 0 35808 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_374
timestamp 1679581782
transform 1 0 36480 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_381
timestamp 1679581782
transform 1 0 37152 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_388
timestamp 1679581782
transform 1 0 37824 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_395
timestamp 1679581782
transform 1 0 38496 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_402
timestamp 1679581782
transform 1 0 39168 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_409
timestamp 1679581782
transform 1 0 39840 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_416
timestamp 1679581782
transform 1 0 40512 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_423
timestamp 1679581782
transform 1 0 41184 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_430
timestamp 1679581782
transform 1 0 41856 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_437
timestamp 1679581782
transform 1 0 42528 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_444
timestamp 1679581782
transform 1 0 43200 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_451
timestamp 1679581782
transform 1 0 43872 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_458
timestamp 1679581782
transform 1 0 44544 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_465
timestamp 1679581782
transform 1 0 45216 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_472
timestamp 1679581782
transform 1 0 45888 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_479
timestamp 1679581782
transform 1 0 46560 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_486
timestamp 1679581782
transform 1 0 47232 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_493
timestamp 1679581782
transform 1 0 47904 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_500
timestamp 1679581782
transform 1 0 48576 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_507
timestamp 1679581782
transform 1 0 49248 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_514
timestamp 1679581782
transform 1 0 49920 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_521
timestamp 1679581782
transform 1 0 50592 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_528
timestamp 1679581782
transform 1 0 51264 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_535
timestamp 1679581782
transform 1 0 51936 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_542
timestamp 1679581782
transform 1 0 52608 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_549
timestamp 1679581782
transform 1 0 53280 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_556
timestamp 1679581782
transform 1 0 53952 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_563
timestamp 1679581782
transform 1 0 54624 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_570
timestamp 1679581782
transform 1 0 55296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_577
timestamp 1679581782
transform 1 0 55968 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_584
timestamp 1679581782
transform 1 0 56640 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_591
timestamp 1679581782
transform 1 0 57312 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_598
timestamp 1679581782
transform 1 0 57984 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_605
timestamp 1679581782
transform 1 0 58656 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_612
timestamp 1679581782
transform 1 0 59328 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_619
timestamp 1679581782
transform 1 0 60000 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_626
timestamp 1679581782
transform 1 0 60672 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_633
timestamp 1679581782
transform 1 0 61344 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_640
timestamp 1679581782
transform 1 0 62016 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_647
timestamp 1679581782
transform 1 0 62688 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_654
timestamp 1679581782
transform 1 0 63360 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_661
timestamp 1679581782
transform 1 0 64032 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_668
timestamp 1679581782
transform 1 0 64704 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_675
timestamp 1679581782
transform 1 0 65376 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_682
timestamp 1679581782
transform 1 0 66048 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_689
timestamp 1679581782
transform 1 0 66720 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_696
timestamp 1679581782
transform 1 0 67392 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_703
timestamp 1679581782
transform 1 0 68064 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_710
timestamp 1679581782
transform 1 0 68736 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_717
timestamp 1679581782
transform 1 0 69408 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_724
timestamp 1679581782
transform 1 0 70080 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_731
timestamp 1679581782
transform 1 0 70752 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_738
timestamp 1677579658
transform 1 0 71424 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_4
timestamp 1679581782
transform 1 0 960 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_11
timestamp 1679581782
transform 1 0 1632 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_18
timestamp 1679581782
transform 1 0 2304 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_25
timestamp 1679581782
transform 1 0 2976 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_32
timestamp 1679581782
transform 1 0 3648 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_39
timestamp 1679581782
transform 1 0 4320 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_46
timestamp 1679581782
transform 1 0 4992 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_53
timestamp 1679581782
transform 1 0 5664 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_60
timestamp 1679581782
transform 1 0 6336 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_67
timestamp 1679581782
transform 1 0 7008 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_74
timestamp 1679581782
transform 1 0 7680 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_81
timestamp 1679581782
transform 1 0 8352 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_88
timestamp 1679581782
transform 1 0 9024 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_95
timestamp 1679581782
transform 1 0 9696 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_102
timestamp 1679581782
transform 1 0 10368 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_109
timestamp 1679581782
transform 1 0 11040 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_116
timestamp 1679581782
transform 1 0 11712 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_123
timestamp 1679581782
transform 1 0 12384 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_130
timestamp 1679581782
transform 1 0 13056 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_137
timestamp 1679581782
transform 1 0 13728 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_144
timestamp 1679581782
transform 1 0 14400 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_151
timestamp 1679581782
transform 1 0 15072 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_158
timestamp 1679581782
transform 1 0 15744 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_165
timestamp 1679581782
transform 1 0 16416 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_172
timestamp 1679581782
transform 1 0 17088 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_179
timestamp 1679581782
transform 1 0 17760 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_186
timestamp 1679581782
transform 1 0 18432 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_193
timestamp 1679581782
transform 1 0 19104 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_200
timestamp 1679581782
transform 1 0 19776 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_207
timestamp 1679581782
transform 1 0 20448 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_214
timestamp 1679581782
transform 1 0 21120 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_221
timestamp 1679581782
transform 1 0 21792 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_228
timestamp 1679581782
transform 1 0 22464 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_235
timestamp 1679581782
transform 1 0 23136 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_242
timestamp 1679581782
transform 1 0 23808 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_249
timestamp 1679581782
transform 1 0 24480 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_256
timestamp 1679581782
transform 1 0 25152 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_263
timestamp 1679581782
transform 1 0 25824 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_270
timestamp 1679581782
transform 1 0 26496 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_277
timestamp 1679581782
transform 1 0 27168 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_284
timestamp 1679581782
transform 1 0 27840 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_291
timestamp 1679581782
transform 1 0 28512 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_298
timestamp 1679581782
transform 1 0 29184 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_305
timestamp 1679581782
transform 1 0 29856 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_312
timestamp 1679581782
transform 1 0 30528 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_319
timestamp 1679581782
transform 1 0 31200 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_326
timestamp 1679581782
transform 1 0 31872 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_333
timestamp 1679581782
transform 1 0 32544 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_340
timestamp 1679581782
transform 1 0 33216 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_347
timestamp 1679581782
transform 1 0 33888 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_354
timestamp 1679581782
transform 1 0 34560 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_361
timestamp 1679581782
transform 1 0 35232 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_368
timestamp 1679581782
transform 1 0 35904 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_375
timestamp 1679581782
transform 1 0 36576 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_382
timestamp 1679581782
transform 1 0 37248 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_389
timestamp 1679581782
transform 1 0 37920 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_396
timestamp 1679581782
transform 1 0 38592 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_403
timestamp 1679581782
transform 1 0 39264 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_410
timestamp 1679581782
transform 1 0 39936 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_417
timestamp 1679581782
transform 1 0 40608 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_424
timestamp 1679581782
transform 1 0 41280 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_431
timestamp 1679581782
transform 1 0 41952 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_438
timestamp 1679581782
transform 1 0 42624 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_445
timestamp 1679581782
transform 1 0 43296 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_452
timestamp 1679581782
transform 1 0 43968 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_459
timestamp 1679581782
transform 1 0 44640 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_466
timestamp 1679581782
transform 1 0 45312 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_473
timestamp 1679581782
transform 1 0 45984 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_480
timestamp 1679581782
transform 1 0 46656 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_487
timestamp 1679581782
transform 1 0 47328 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_494
timestamp 1679581782
transform 1 0 48000 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_501
timestamp 1679581782
transform 1 0 48672 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_508
timestamp 1679581782
transform 1 0 49344 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_515
timestamp 1679581782
transform 1 0 50016 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_522
timestamp 1679581782
transform 1 0 50688 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_529
timestamp 1679581782
transform 1 0 51360 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_536
timestamp 1679581782
transform 1 0 52032 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_543
timestamp 1679581782
transform 1 0 52704 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_550
timestamp 1679581782
transform 1 0 53376 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_557
timestamp 1679581782
transform 1 0 54048 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_564
timestamp 1679581782
transform 1 0 54720 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_571
timestamp 1679581782
transform 1 0 55392 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_578
timestamp 1679581782
transform 1 0 56064 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_585
timestamp 1679581782
transform 1 0 56736 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_592
timestamp 1679581782
transform 1 0 57408 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_599
timestamp 1679581782
transform 1 0 58080 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_606
timestamp 1679581782
transform 1 0 58752 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_613
timestamp 1679581782
transform 1 0 59424 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_620
timestamp 1679581782
transform 1 0 60096 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_627
timestamp 1679581782
transform 1 0 60768 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_634
timestamp 1679581782
transform 1 0 61440 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_641
timestamp 1679581782
transform 1 0 62112 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_648
timestamp 1679581782
transform 1 0 62784 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_655
timestamp 1679581782
transform 1 0 63456 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_662
timestamp 1679581782
transform 1 0 64128 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_669
timestamp 1679581782
transform 1 0 64800 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_676
timestamp 1679581782
transform 1 0 65472 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_683
timestamp 1679581782
transform 1 0 66144 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_690
timestamp 1679581782
transform 1 0 66816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_697
timestamp 1679581782
transform 1 0 67488 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_704
timestamp 1679581782
transform 1 0 68160 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_711
timestamp 1679581782
transform 1 0 68832 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_718
timestamp 1679581782
transform 1 0 69504 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_725
timestamp 1679581782
transform 1 0 70176 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_732
timestamp 1679581782
transform 1 0 70848 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_4
timestamp 1677580104
transform 1 0 960 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_15_10
timestamp 1679581782
transform 1 0 1536 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_17
timestamp 1679581782
transform 1 0 2208 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_24
timestamp 1679581782
transform 1 0 2880 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_31
timestamp 1679581782
transform 1 0 3552 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_38
timestamp 1679581782
transform 1 0 4224 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_45
timestamp 1679581782
transform 1 0 4896 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_52
timestamp 1679581782
transform 1 0 5568 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_59
timestamp 1679581782
transform 1 0 6240 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_66
timestamp 1679581782
transform 1 0 6912 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_73
timestamp 1679581782
transform 1 0 7584 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_80
timestamp 1679581782
transform 1 0 8256 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_87
timestamp 1679581782
transform 1 0 8928 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_94
timestamp 1679581782
transform 1 0 9600 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_101
timestamp 1679581782
transform 1 0 10272 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_108
timestamp 1679581782
transform 1 0 10944 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_115
timestamp 1679581782
transform 1 0 11616 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_122
timestamp 1679581782
transform 1 0 12288 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_129
timestamp 1679581782
transform 1 0 12960 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_136
timestamp 1679581782
transform 1 0 13632 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_143
timestamp 1679581782
transform 1 0 14304 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_150
timestamp 1679581782
transform 1 0 14976 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_157
timestamp 1679581782
transform 1 0 15648 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_164
timestamp 1679581782
transform 1 0 16320 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_171
timestamp 1679581782
transform 1 0 16992 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_178
timestamp 1679581782
transform 1 0 17664 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_185
timestamp 1679581782
transform 1 0 18336 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_192
timestamp 1679581782
transform 1 0 19008 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_199
timestamp 1679581782
transform 1 0 19680 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_206
timestamp 1679581782
transform 1 0 20352 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_213
timestamp 1679581782
transform 1 0 21024 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_220
timestamp 1679581782
transform 1 0 21696 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_227
timestamp 1679581782
transform 1 0 22368 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_234
timestamp 1679581782
transform 1 0 23040 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_241
timestamp 1679581782
transform 1 0 23712 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_248
timestamp 1679581782
transform 1 0 24384 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_255
timestamp 1679581782
transform 1 0 25056 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_262
timestamp 1679581782
transform 1 0 25728 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_269
timestamp 1679581782
transform 1 0 26400 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_276
timestamp 1679581782
transform 1 0 27072 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_283
timestamp 1679581782
transform 1 0 27744 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_290
timestamp 1679581782
transform 1 0 28416 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_297
timestamp 1679581782
transform 1 0 29088 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_304
timestamp 1679581782
transform 1 0 29760 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_311
timestamp 1679581782
transform 1 0 30432 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_318
timestamp 1679581782
transform 1 0 31104 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_325
timestamp 1679581782
transform 1 0 31776 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_332
timestamp 1679581782
transform 1 0 32448 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_339
timestamp 1679581782
transform 1 0 33120 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_346
timestamp 1679581782
transform 1 0 33792 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_353
timestamp 1679581782
transform 1 0 34464 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_360
timestamp 1679581782
transform 1 0 35136 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_367
timestamp 1679581782
transform 1 0 35808 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_374
timestamp 1679581782
transform 1 0 36480 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_381
timestamp 1679581782
transform 1 0 37152 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_388
timestamp 1679581782
transform 1 0 37824 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_395
timestamp 1679581782
transform 1 0 38496 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_402
timestamp 1679581782
transform 1 0 39168 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_409
timestamp 1679581782
transform 1 0 39840 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_416
timestamp 1679581782
transform 1 0 40512 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_423
timestamp 1679581782
transform 1 0 41184 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_430
timestamp 1679581782
transform 1 0 41856 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_437
timestamp 1679581782
transform 1 0 42528 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_444
timestamp 1679581782
transform 1 0 43200 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_451
timestamp 1679581782
transform 1 0 43872 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_458
timestamp 1679581782
transform 1 0 44544 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_465
timestamp 1679581782
transform 1 0 45216 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_472
timestamp 1679581782
transform 1 0 45888 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_479
timestamp 1679581782
transform 1 0 46560 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_486
timestamp 1679581782
transform 1 0 47232 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_493
timestamp 1679581782
transform 1 0 47904 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_500
timestamp 1679581782
transform 1 0 48576 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_507
timestamp 1679581782
transform 1 0 49248 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_514
timestamp 1679581782
transform 1 0 49920 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_521
timestamp 1679581782
transform 1 0 50592 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_528
timestamp 1679581782
transform 1 0 51264 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_535
timestamp 1679581782
transform 1 0 51936 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_542
timestamp 1679581782
transform 1 0 52608 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_549
timestamp 1679581782
transform 1 0 53280 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_556
timestamp 1679581782
transform 1 0 53952 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_563
timestamp 1679581782
transform 1 0 54624 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_570
timestamp 1679581782
transform 1 0 55296 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_577
timestamp 1679581782
transform 1 0 55968 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_584
timestamp 1679581782
transform 1 0 56640 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_591
timestamp 1679581782
transform 1 0 57312 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_598
timestamp 1679581782
transform 1 0 57984 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_605
timestamp 1679581782
transform 1 0 58656 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_612
timestamp 1679581782
transform 1 0 59328 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_619
timestamp 1679581782
transform 1 0 60000 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_626
timestamp 1679581782
transform 1 0 60672 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_633
timestamp 1679581782
transform 1 0 61344 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_640
timestamp 1679581782
transform 1 0 62016 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_647
timestamp 1679581782
transform 1 0 62688 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_654
timestamp 1679581782
transform 1 0 63360 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_661
timestamp 1679581782
transform 1 0 64032 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_668
timestamp 1679581782
transform 1 0 64704 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_675
timestamp 1679581782
transform 1 0 65376 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_682
timestamp 1679581782
transform 1 0 66048 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_689
timestamp 1679581782
transform 1 0 66720 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_696
timestamp 1679581782
transform 1 0 67392 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_703
timestamp 1679581782
transform 1 0 68064 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_710
timestamp 1679581782
transform 1 0 68736 0 -1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_717
timestamp 1679581782
transform 1 0 69408 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_724
timestamp 1677580104
transform 1 0 70080 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_726
timestamp 1677579658
transform 1 0 70272 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_730
timestamp 1677579658
transform 1 0 70656 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_737
timestamp 1677580104
transform 1 0 71328 0 -1 12852
box -48 -56 240 834
use sg13g2_decap_4  FILLER_16_4
timestamp 1679577901
transform 1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_16_8
timestamp 1677580104
transform 1 0 1344 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_14
timestamp 1679581782
transform 1 0 1920 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_21
timestamp 1679581782
transform 1 0 2592 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_28
timestamp 1679581782
transform 1 0 3264 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_35
timestamp 1679581782
transform 1 0 3936 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_42
timestamp 1679581782
transform 1 0 4608 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_49
timestamp 1679581782
transform 1 0 5280 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_56
timestamp 1679581782
transform 1 0 5952 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_63
timestamp 1679581782
transform 1 0 6624 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_70
timestamp 1679581782
transform 1 0 7296 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_77
timestamp 1679581782
transform 1 0 7968 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_84
timestamp 1679581782
transform 1 0 8640 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_91
timestamp 1679581782
transform 1 0 9312 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_98
timestamp 1679581782
transform 1 0 9984 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_105
timestamp 1679581782
transform 1 0 10656 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_112
timestamp 1679581782
transform 1 0 11328 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_119
timestamp 1679581782
transform 1 0 12000 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_126
timestamp 1679581782
transform 1 0 12672 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_133
timestamp 1679581782
transform 1 0 13344 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_140
timestamp 1679581782
transform 1 0 14016 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_147
timestamp 1679581782
transform 1 0 14688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_154
timestamp 1679581782
transform 1 0 15360 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_161
timestamp 1679581782
transform 1 0 16032 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_168
timestamp 1679581782
transform 1 0 16704 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_175
timestamp 1679581782
transform 1 0 17376 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_182
timestamp 1679581782
transform 1 0 18048 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_189
timestamp 1679581782
transform 1 0 18720 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_196
timestamp 1679581782
transform 1 0 19392 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_203
timestamp 1679581782
transform 1 0 20064 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_210
timestamp 1679581782
transform 1 0 20736 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_217
timestamp 1679581782
transform 1 0 21408 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_224
timestamp 1679581782
transform 1 0 22080 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_231
timestamp 1679581782
transform 1 0 22752 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_238
timestamp 1679581782
transform 1 0 23424 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_245
timestamp 1679581782
transform 1 0 24096 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_252
timestamp 1679581782
transform 1 0 24768 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_259
timestamp 1679581782
transform 1 0 25440 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_266
timestamp 1679581782
transform 1 0 26112 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_273
timestamp 1679581782
transform 1 0 26784 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_280
timestamp 1679581782
transform 1 0 27456 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_287
timestamp 1679581782
transform 1 0 28128 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_294
timestamp 1679581782
transform 1 0 28800 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_301
timestamp 1679581782
transform 1 0 29472 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_308
timestamp 1679581782
transform 1 0 30144 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_315
timestamp 1679581782
transform 1 0 30816 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_322
timestamp 1679581782
transform 1 0 31488 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_329
timestamp 1679581782
transform 1 0 32160 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_336
timestamp 1679581782
transform 1 0 32832 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_343
timestamp 1679581782
transform 1 0 33504 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_350
timestamp 1679581782
transform 1 0 34176 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_357
timestamp 1679581782
transform 1 0 34848 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_364
timestamp 1679581782
transform 1 0 35520 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_371
timestamp 1679581782
transform 1 0 36192 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_378
timestamp 1679581782
transform 1 0 36864 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_385
timestamp 1679581782
transform 1 0 37536 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_392
timestamp 1679581782
transform 1 0 38208 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_399
timestamp 1679581782
transform 1 0 38880 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_406
timestamp 1679581782
transform 1 0 39552 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_413
timestamp 1679581782
transform 1 0 40224 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_420
timestamp 1679581782
transform 1 0 40896 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_427
timestamp 1679581782
transform 1 0 41568 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_434
timestamp 1679581782
transform 1 0 42240 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_441
timestamp 1679581782
transform 1 0 42912 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_448
timestamp 1679581782
transform 1 0 43584 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_455
timestamp 1679581782
transform 1 0 44256 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_462
timestamp 1679581782
transform 1 0 44928 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_469
timestamp 1679581782
transform 1 0 45600 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_476
timestamp 1679581782
transform 1 0 46272 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_483
timestamp 1679581782
transform 1 0 46944 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_490
timestamp 1679581782
transform 1 0 47616 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_497
timestamp 1679581782
transform 1 0 48288 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_504
timestamp 1679581782
transform 1 0 48960 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_511
timestamp 1679581782
transform 1 0 49632 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_518
timestamp 1679581782
transform 1 0 50304 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_525
timestamp 1679581782
transform 1 0 50976 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_532
timestamp 1679581782
transform 1 0 51648 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_539
timestamp 1679581782
transform 1 0 52320 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_546
timestamp 1679581782
transform 1 0 52992 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_553
timestamp 1679581782
transform 1 0 53664 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_560
timestamp 1679581782
transform 1 0 54336 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_567
timestamp 1679581782
transform 1 0 55008 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_574
timestamp 1679581782
transform 1 0 55680 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_581
timestamp 1679581782
transform 1 0 56352 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_588
timestamp 1679581782
transform 1 0 57024 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_595
timestamp 1679581782
transform 1 0 57696 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_602
timestamp 1679581782
transform 1 0 58368 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_609
timestamp 1679581782
transform 1 0 59040 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_616
timestamp 1679581782
transform 1 0 59712 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_623
timestamp 1679581782
transform 1 0 60384 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_630
timestamp 1679581782
transform 1 0 61056 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_637
timestamp 1679581782
transform 1 0 61728 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_644
timestamp 1679581782
transform 1 0 62400 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_651
timestamp 1679581782
transform 1 0 63072 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_658
timestamp 1679581782
transform 1 0 63744 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_665
timestamp 1679581782
transform 1 0 64416 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_672
timestamp 1679581782
transform 1 0 65088 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_679
timestamp 1679581782
transform 1 0 65760 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_686
timestamp 1679581782
transform 1 0 66432 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_693
timestamp 1679581782
transform 1 0 67104 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_700
timestamp 1679581782
transform 1 0 67776 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_707
timestamp 1679581782
transform 1 0 68448 0 1 12852
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_714
timestamp 1679581782
transform 1 0 69120 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_738
timestamp 1677579658
transform 1 0 71424 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_17_0
timestamp 1679577901
transform 1 0 576 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_8
timestamp 1679581782
transform 1 0 1344 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_15
timestamp 1679581782
transform 1 0 2016 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_22
timestamp 1679581782
transform 1 0 2688 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_29
timestamp 1679581782
transform 1 0 3360 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_36
timestamp 1679581782
transform 1 0 4032 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_43
timestamp 1679581782
transform 1 0 4704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_50
timestamp 1679581782
transform 1 0 5376 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_57
timestamp 1679581782
transform 1 0 6048 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_64
timestamp 1679581782
transform 1 0 6720 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_71
timestamp 1679581782
transform 1 0 7392 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_78
timestamp 1679581782
transform 1 0 8064 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_85
timestamp 1679581782
transform 1 0 8736 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_92
timestamp 1679581782
transform 1 0 9408 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_99
timestamp 1679581782
transform 1 0 10080 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_106
timestamp 1679581782
transform 1 0 10752 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_113
timestamp 1679581782
transform 1 0 11424 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_120
timestamp 1679581782
transform 1 0 12096 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_127
timestamp 1679581782
transform 1 0 12768 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_134
timestamp 1679581782
transform 1 0 13440 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_141
timestamp 1679581782
transform 1 0 14112 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_148
timestamp 1679581782
transform 1 0 14784 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_155
timestamp 1679581782
transform 1 0 15456 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_162
timestamp 1679581782
transform 1 0 16128 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_169
timestamp 1679581782
transform 1 0 16800 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_176
timestamp 1679581782
transform 1 0 17472 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_183
timestamp 1679581782
transform 1 0 18144 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_190
timestamp 1679581782
transform 1 0 18816 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_197
timestamp 1679581782
transform 1 0 19488 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_204
timestamp 1679581782
transform 1 0 20160 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_211
timestamp 1679581782
transform 1 0 20832 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_218
timestamp 1679581782
transform 1 0 21504 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_225
timestamp 1679581782
transform 1 0 22176 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_232
timestamp 1679581782
transform 1 0 22848 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_239
timestamp 1679581782
transform 1 0 23520 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_246
timestamp 1679581782
transform 1 0 24192 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_253
timestamp 1679581782
transform 1 0 24864 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_260
timestamp 1679581782
transform 1 0 25536 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_267
timestamp 1679581782
transform 1 0 26208 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_274
timestamp 1679581782
transform 1 0 26880 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_281
timestamp 1679581782
transform 1 0 27552 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_288
timestamp 1679581782
transform 1 0 28224 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_295
timestamp 1679581782
transform 1 0 28896 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_302
timestamp 1679581782
transform 1 0 29568 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_309
timestamp 1679581782
transform 1 0 30240 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_316
timestamp 1679581782
transform 1 0 30912 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_323
timestamp 1679581782
transform 1 0 31584 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_330
timestamp 1679581782
transform 1 0 32256 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_337
timestamp 1679581782
transform 1 0 32928 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_344
timestamp 1679581782
transform 1 0 33600 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_351
timestamp 1679581782
transform 1 0 34272 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_358
timestamp 1679581782
transform 1 0 34944 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_365
timestamp 1679581782
transform 1 0 35616 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_372
timestamp 1679581782
transform 1 0 36288 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_379
timestamp 1679581782
transform 1 0 36960 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_386
timestamp 1679581782
transform 1 0 37632 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_393
timestamp 1679581782
transform 1 0 38304 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_400
timestamp 1679581782
transform 1 0 38976 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_407
timestamp 1679581782
transform 1 0 39648 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_414
timestamp 1679581782
transform 1 0 40320 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_421
timestamp 1679581782
transform 1 0 40992 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_428
timestamp 1679581782
transform 1 0 41664 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_435
timestamp 1679581782
transform 1 0 42336 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_442
timestamp 1679581782
transform 1 0 43008 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_449
timestamp 1679581782
transform 1 0 43680 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_456
timestamp 1679581782
transform 1 0 44352 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_463
timestamp 1679581782
transform 1 0 45024 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_470
timestamp 1679581782
transform 1 0 45696 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_477
timestamp 1679581782
transform 1 0 46368 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_484
timestamp 1679581782
transform 1 0 47040 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_491
timestamp 1679581782
transform 1 0 47712 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_498
timestamp 1679581782
transform 1 0 48384 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_505
timestamp 1679581782
transform 1 0 49056 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_512
timestamp 1679581782
transform 1 0 49728 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_519
timestamp 1679581782
transform 1 0 50400 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_526
timestamp 1679581782
transform 1 0 51072 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_533
timestamp 1679581782
transform 1 0 51744 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_540
timestamp 1679581782
transform 1 0 52416 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_547
timestamp 1679581782
transform 1 0 53088 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_554
timestamp 1679581782
transform 1 0 53760 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_561
timestamp 1679581782
transform 1 0 54432 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_568
timestamp 1679581782
transform 1 0 55104 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_575
timestamp 1679581782
transform 1 0 55776 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_582
timestamp 1679581782
transform 1 0 56448 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_589
timestamp 1679581782
transform 1 0 57120 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_596
timestamp 1679581782
transform 1 0 57792 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_603
timestamp 1679581782
transform 1 0 58464 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_610
timestamp 1679581782
transform 1 0 59136 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_617
timestamp 1679581782
transform 1 0 59808 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_624
timestamp 1679581782
transform 1 0 60480 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_631
timestamp 1679581782
transform 1 0 61152 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_638
timestamp 1679581782
transform 1 0 61824 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_645
timestamp 1679581782
transform 1 0 62496 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_652
timestamp 1679581782
transform 1 0 63168 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_659
timestamp 1679581782
transform 1 0 63840 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_666
timestamp 1679581782
transform 1 0 64512 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_673
timestamp 1679581782
transform 1 0 65184 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_680
timestamp 1679581782
transform 1 0 65856 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_687
timestamp 1679581782
transform 1 0 66528 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_694
timestamp 1679581782
transform 1 0 67200 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_701
timestamp 1679581782
transform 1 0 67872 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_708
timestamp 1679581782
transform 1 0 68544 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_715
timestamp 1679581782
transform 1 0 69216 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_722
timestamp 1679581782
transform 1 0 69888 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_734
timestamp 1677580104
transform 1 0 71040 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_18_4
timestamp 1679577901
transform 1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_decap_8  FILLER_18_16
timestamp 1679581782
transform 1 0 2112 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_23
timestamp 1679581782
transform 1 0 2784 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_30
timestamp 1679581782
transform 1 0 3456 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_37
timestamp 1679581782
transform 1 0 4128 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_44
timestamp 1679581782
transform 1 0 4800 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_51
timestamp 1679581782
transform 1 0 5472 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_58
timestamp 1679581782
transform 1 0 6144 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_65
timestamp 1679581782
transform 1 0 6816 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_72
timestamp 1679581782
transform 1 0 7488 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_79
timestamp 1679581782
transform 1 0 8160 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_86
timestamp 1679581782
transform 1 0 8832 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_93
timestamp 1679581782
transform 1 0 9504 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_100
timestamp 1679581782
transform 1 0 10176 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_107
timestamp 1679581782
transform 1 0 10848 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_114
timestamp 1679581782
transform 1 0 11520 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_121
timestamp 1679581782
transform 1 0 12192 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_128
timestamp 1679581782
transform 1 0 12864 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_135
timestamp 1679581782
transform 1 0 13536 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_142
timestamp 1679581782
transform 1 0 14208 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_149
timestamp 1679581782
transform 1 0 14880 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_156
timestamp 1679581782
transform 1 0 15552 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_163
timestamp 1679581782
transform 1 0 16224 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_170
timestamp 1679581782
transform 1 0 16896 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_177
timestamp 1679581782
transform 1 0 17568 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_184
timestamp 1679581782
transform 1 0 18240 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_191
timestamp 1679581782
transform 1 0 18912 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_198
timestamp 1679581782
transform 1 0 19584 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_205
timestamp 1679581782
transform 1 0 20256 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_212
timestamp 1679581782
transform 1 0 20928 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_219
timestamp 1679581782
transform 1 0 21600 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_226
timestamp 1679581782
transform 1 0 22272 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_233
timestamp 1679581782
transform 1 0 22944 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_240
timestamp 1679581782
transform 1 0 23616 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_247
timestamp 1679581782
transform 1 0 24288 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_254
timestamp 1679581782
transform 1 0 24960 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_261
timestamp 1679581782
transform 1 0 25632 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_268
timestamp 1679581782
transform 1 0 26304 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_275
timestamp 1679581782
transform 1 0 26976 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_282
timestamp 1679581782
transform 1 0 27648 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_289
timestamp 1679581782
transform 1 0 28320 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_296
timestamp 1679581782
transform 1 0 28992 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_303
timestamp 1679581782
transform 1 0 29664 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_310
timestamp 1679581782
transform 1 0 30336 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_317
timestamp 1679581782
transform 1 0 31008 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_324
timestamp 1679581782
transform 1 0 31680 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_331
timestamp 1679581782
transform 1 0 32352 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_338
timestamp 1679581782
transform 1 0 33024 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_345
timestamp 1679581782
transform 1 0 33696 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_352
timestamp 1679581782
transform 1 0 34368 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_359
timestamp 1679581782
transform 1 0 35040 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_366
timestamp 1679581782
transform 1 0 35712 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_373
timestamp 1679581782
transform 1 0 36384 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_380
timestamp 1679581782
transform 1 0 37056 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_387
timestamp 1679581782
transform 1 0 37728 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_394
timestamp 1679581782
transform 1 0 38400 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_401
timestamp 1679581782
transform 1 0 39072 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_408
timestamp 1679581782
transform 1 0 39744 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_415
timestamp 1679581782
transform 1 0 40416 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_422
timestamp 1679581782
transform 1 0 41088 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_429
timestamp 1679581782
transform 1 0 41760 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_436
timestamp 1679581782
transform 1 0 42432 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_443
timestamp 1679581782
transform 1 0 43104 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_450
timestamp 1679581782
transform 1 0 43776 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_457
timestamp 1679581782
transform 1 0 44448 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_464
timestamp 1679581782
transform 1 0 45120 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_471
timestamp 1679581782
transform 1 0 45792 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_478
timestamp 1679581782
transform 1 0 46464 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_485
timestamp 1679581782
transform 1 0 47136 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_492
timestamp 1679581782
transform 1 0 47808 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_499
timestamp 1679581782
transform 1 0 48480 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_506
timestamp 1679581782
transform 1 0 49152 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_513
timestamp 1679581782
transform 1 0 49824 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_520
timestamp 1679581782
transform 1 0 50496 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_527
timestamp 1679581782
transform 1 0 51168 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_534
timestamp 1679581782
transform 1 0 51840 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_541
timestamp 1679581782
transform 1 0 52512 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_548
timestamp 1679581782
transform 1 0 53184 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_555
timestamp 1679581782
transform 1 0 53856 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_562
timestamp 1679581782
transform 1 0 54528 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_569
timestamp 1679581782
transform 1 0 55200 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_576
timestamp 1679581782
transform 1 0 55872 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_583
timestamp 1679581782
transform 1 0 56544 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_590
timestamp 1679581782
transform 1 0 57216 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_597
timestamp 1679581782
transform 1 0 57888 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_604
timestamp 1679581782
transform 1 0 58560 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_611
timestamp 1679581782
transform 1 0 59232 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_618
timestamp 1679581782
transform 1 0 59904 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_625
timestamp 1679581782
transform 1 0 60576 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_632
timestamp 1679581782
transform 1 0 61248 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_639
timestamp 1679581782
transform 1 0 61920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_646
timestamp 1679581782
transform 1 0 62592 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_653
timestamp 1679581782
transform 1 0 63264 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_660
timestamp 1679581782
transform 1 0 63936 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_667
timestamp 1679581782
transform 1 0 64608 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_674
timestamp 1679581782
transform 1 0 65280 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_681
timestamp 1679581782
transform 1 0 65952 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_688
timestamp 1679581782
transform 1 0 66624 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_695
timestamp 1679581782
transform 1 0 67296 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_702
timestamp 1679581782
transform 1 0 67968 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_709
timestamp 1679581782
transform 1 0 68640 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_716
timestamp 1679581782
transform 1 0 69312 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_723
timestamp 1679581782
transform 1 0 69984 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_730
timestamp 1679581782
transform 1 0 70656 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_737
timestamp 1679581782
transform 1 0 71328 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_744
timestamp 1679581782
transform 1 0 72000 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_758
timestamp 1677579658
transform 1 0 73344 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_776
timestamp 1677580104
transform 1 0 75072 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_781
timestamp 1677580104
transform 1 0 75552 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_789
timestamp 1677580104
transform 1 0 76320 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_794
timestamp 1677579658
transform 1 0 76800 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_798
timestamp 1677579658
transform 1 0 77184 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_802
timestamp 1677580104
transform 1 0 77568 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_810
timestamp 1677580104
transform 1 0 78336 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_819
timestamp 1677579658
transform 1 0 79200 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_826
timestamp 1677580104
transform 1 0 79872 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_840
timestamp 1677579658
transform 1 0 81216 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_844
timestamp 1677580104
transform 1 0 81600 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_846
timestamp 1677579658
transform 1 0 81792 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_857
timestamp 1677579658
transform 1 0 82848 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_861
timestamp 1677579658
transform 1 0 83232 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_865
timestamp 1677579658
transform 1 0 83616 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_869
timestamp 1679577901
transform 1 0 84000 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_873
timestamp 1677579658
transform 1 0 84384 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_877
timestamp 1677580104
transform 1 0 84768 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_882
timestamp 1677579658
transform 1 0 85248 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_886
timestamp 1677579658
transform 1 0 85632 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_890
timestamp 1677580104
transform 1 0 86016 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_895
timestamp 1677579658
transform 1 0 86496 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_899
timestamp 1677579658
transform 1 0 86880 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_903
timestamp 1679577901
transform 1 0 87264 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_907
timestamp 1677579658
transform 1 0 87648 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_911
timestamp 1677579658
transform 1 0 88032 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_915
timestamp 1677579658
transform 1 0 88416 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_919
timestamp 1677579658
transform 1 0 88800 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_923
timestamp 1677580104
transform 1 0 89184 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_925
timestamp 1677579658
transform 1 0 89376 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_929
timestamp 1677579658
transform 1 0 89760 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_936
timestamp 1677579658
transform 1 0 90432 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_940
timestamp 1677580104
transform 1 0 90816 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_952
timestamp 1677579658
transform 1 0 91968 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_969
timestamp 1677580104
transform 1 0 93600 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_974
timestamp 1677579658
transform 1 0 94080 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_978
timestamp 1677579658
transform 1 0 94464 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_982
timestamp 1677579658
transform 1 0 94848 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_986
timestamp 1677579658
transform 1 0 95232 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_990
timestamp 1677580104
transform 1 0 95616 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_995
timestamp 1677579658
transform 1 0 96096 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_999
timestamp 1677579658
transform 1 0 96480 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_1007
timestamp 1677579658
transform 1 0 97248 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_1014
timestamp 1677580104
transform 1 0 97920 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_1016
timestamp 1677579658
transform 1 0 98112 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_1024
timestamp 1679577901
transform 1 0 98880 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_1028
timestamp 1677579658
transform 1 0 99264 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_4
timestamp 1679581782
transform 1 0 960 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_11
timestamp 1679581782
transform 1 0 1632 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_18
timestamp 1679581782
transform 1 0 2304 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_25
timestamp 1679581782
transform 1 0 2976 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_32
timestamp 1679581782
transform 1 0 3648 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_39
timestamp 1679581782
transform 1 0 4320 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_46
timestamp 1679581782
transform 1 0 4992 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_53
timestamp 1679581782
transform 1 0 5664 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_60
timestamp 1679581782
transform 1 0 6336 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_67
timestamp 1679581782
transform 1 0 7008 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_74
timestamp 1679581782
transform 1 0 7680 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_81
timestamp 1679581782
transform 1 0 8352 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_88
timestamp 1679581782
transform 1 0 9024 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_95
timestamp 1679581782
transform 1 0 9696 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_102
timestamp 1679581782
transform 1 0 10368 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_109
timestamp 1679581782
transform 1 0 11040 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_116
timestamp 1679581782
transform 1 0 11712 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_123
timestamp 1679581782
transform 1 0 12384 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_130
timestamp 1679581782
transform 1 0 13056 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_137
timestamp 1679581782
transform 1 0 13728 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_144
timestamp 1679581782
transform 1 0 14400 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_151
timestamp 1679581782
transform 1 0 15072 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_158
timestamp 1679581782
transform 1 0 15744 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_165
timestamp 1679581782
transform 1 0 16416 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_172
timestamp 1679581782
transform 1 0 17088 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_179
timestamp 1679581782
transform 1 0 17760 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_186
timestamp 1679581782
transform 1 0 18432 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_193
timestamp 1679581782
transform 1 0 19104 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_200
timestamp 1679581782
transform 1 0 19776 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_207
timestamp 1679581782
transform 1 0 20448 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_214
timestamp 1679581782
transform 1 0 21120 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_221
timestamp 1679581782
transform 1 0 21792 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_228
timestamp 1679581782
transform 1 0 22464 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_235
timestamp 1679581782
transform 1 0 23136 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_242
timestamp 1679581782
transform 1 0 23808 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_249
timestamp 1679581782
transform 1 0 24480 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_256
timestamp 1679581782
transform 1 0 25152 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_263
timestamp 1679581782
transform 1 0 25824 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_270
timestamp 1679581782
transform 1 0 26496 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_277
timestamp 1679581782
transform 1 0 27168 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_284
timestamp 1679581782
transform 1 0 27840 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_291
timestamp 1679581782
transform 1 0 28512 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_298
timestamp 1679581782
transform 1 0 29184 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_305
timestamp 1679581782
transform 1 0 29856 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_312
timestamp 1679581782
transform 1 0 30528 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_319
timestamp 1679581782
transform 1 0 31200 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_326
timestamp 1679581782
transform 1 0 31872 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_333
timestamp 1679581782
transform 1 0 32544 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_340
timestamp 1679581782
transform 1 0 33216 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_347
timestamp 1679581782
transform 1 0 33888 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_354
timestamp 1679581782
transform 1 0 34560 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_361
timestamp 1679581782
transform 1 0 35232 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_368
timestamp 1679581782
transform 1 0 35904 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_375
timestamp 1679581782
transform 1 0 36576 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_382
timestamp 1679581782
transform 1 0 37248 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_389
timestamp 1679581782
transform 1 0 37920 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_396
timestamp 1679581782
transform 1 0 38592 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_403
timestamp 1679581782
transform 1 0 39264 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_410
timestamp 1679581782
transform 1 0 39936 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_417
timestamp 1679581782
transform 1 0 40608 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_424
timestamp 1679581782
transform 1 0 41280 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_431
timestamp 1679581782
transform 1 0 41952 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_438
timestamp 1679581782
transform 1 0 42624 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_445
timestamp 1679581782
transform 1 0 43296 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_452
timestamp 1679581782
transform 1 0 43968 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_459
timestamp 1679581782
transform 1 0 44640 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_466
timestamp 1679581782
transform 1 0 45312 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_473
timestamp 1679581782
transform 1 0 45984 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_480
timestamp 1679581782
transform 1 0 46656 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_487
timestamp 1679581782
transform 1 0 47328 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_494
timestamp 1679581782
transform 1 0 48000 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_501
timestamp 1679581782
transform 1 0 48672 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_508
timestamp 1679581782
transform 1 0 49344 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_515
timestamp 1679581782
transform 1 0 50016 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_522
timestamp 1679581782
transform 1 0 50688 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_529
timestamp 1679581782
transform 1 0 51360 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_536
timestamp 1679581782
transform 1 0 52032 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_543
timestamp 1679581782
transform 1 0 52704 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_550
timestamp 1679581782
transform 1 0 53376 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_557
timestamp 1679581782
transform 1 0 54048 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_564
timestamp 1679581782
transform 1 0 54720 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_571
timestamp 1679581782
transform 1 0 55392 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_578
timestamp 1679581782
transform 1 0 56064 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_585
timestamp 1679581782
transform 1 0 56736 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_592
timestamp 1679581782
transform 1 0 57408 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_599
timestamp 1679581782
transform 1 0 58080 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_606
timestamp 1679581782
transform 1 0 58752 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_613
timestamp 1679581782
transform 1 0 59424 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_620
timestamp 1679581782
transform 1 0 60096 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_627
timestamp 1679581782
transform 1 0 60768 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_634
timestamp 1679581782
transform 1 0 61440 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_641
timestamp 1679581782
transform 1 0 62112 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_648
timestamp 1679581782
transform 1 0 62784 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_655
timestamp 1679581782
transform 1 0 63456 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_662
timestamp 1679581782
transform 1 0 64128 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_669
timestamp 1679581782
transform 1 0 64800 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_676
timestamp 1679581782
transform 1 0 65472 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_683
timestamp 1679581782
transform 1 0 66144 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_690
timestamp 1679581782
transform 1 0 66816 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_697
timestamp 1679581782
transform 1 0 67488 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_704
timestamp 1679581782
transform 1 0 68160 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_711
timestamp 1679581782
transform 1 0 68832 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_718
timestamp 1679581782
transform 1 0 69504 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_725
timestamp 1679581782
transform 1 0 70176 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_732
timestamp 1679581782
transform 1 0 70848 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_739
timestamp 1679581782
transform 1 0 71520 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_746
timestamp 1679581782
transform 1 0 72192 0 -1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_753
timestamp 1679581782
transform 1 0 72864 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_760
timestamp 1677579658
transform 1 0 73536 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_769
timestamp 1679577901
transform 1 0 74400 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_777
timestamp 1677579658
transform 1 0 75168 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_782
timestamp 1677579658
transform 1 0 75648 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_811
timestamp 1677579658
transform 1 0 78432 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_828
timestamp 1677579658
transform 1 0 80064 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_833
timestamp 1677579658
transform 1 0 80544 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_842
timestamp 1677580104
transform 1 0 81408 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_844
timestamp 1677579658
transform 1 0 81600 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_848
timestamp 1679581782
transform 1 0 81984 0 -1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_19_855
timestamp 1677580104
transform 1 0 82656 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_857
timestamp 1677579658
transform 1 0 82848 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_866
timestamp 1677579658
transform 1 0 83712 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_878
timestamp 1677579658
transform 1 0 84864 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_899
timestamp 1677579658
transform 1 0 86880 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_907
timestamp 1677580104
transform 1 0 87648 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_933
timestamp 1677580104
transform 1 0 90144 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_935
timestamp 1677579658
transform 1 0 90336 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_944
timestamp 1677580104
transform 1 0 91200 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_950
timestamp 1677579658
transform 1 0 91776 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_963
timestamp 1677580104
transform 1 0 93024 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_965
timestamp 1677579658
transform 1 0 93216 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_974
timestamp 1677579658
transform 1 0 94080 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_987
timestamp 1677579658
transform 1 0 95328 0 -1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_1023
timestamp 1679577901
transform 1 0 98784 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_1027
timestamp 1677580104
transform 1 0 99168 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_4
timestamp 1679581782
transform 1 0 960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_11
timestamp 1679581782
transform 1 0 1632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_18
timestamp 1679581782
transform 1 0 2304 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_25
timestamp 1679581782
transform 1 0 2976 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_32
timestamp 1679581782
transform 1 0 3648 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_39
timestamp 1679581782
transform 1 0 4320 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_46
timestamp 1679581782
transform 1 0 4992 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_53
timestamp 1679581782
transform 1 0 5664 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_60
timestamp 1679581782
transform 1 0 6336 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_67
timestamp 1679581782
transform 1 0 7008 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_74
timestamp 1679581782
transform 1 0 7680 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_81
timestamp 1679581782
transform 1 0 8352 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_88
timestamp 1679581782
transform 1 0 9024 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_95
timestamp 1679581782
transform 1 0 9696 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_102
timestamp 1679581782
transform 1 0 10368 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_109
timestamp 1679581782
transform 1 0 11040 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_116
timestamp 1679581782
transform 1 0 11712 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_123
timestamp 1679581782
transform 1 0 12384 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_130
timestamp 1679581782
transform 1 0 13056 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_137
timestamp 1679581782
transform 1 0 13728 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_144
timestamp 1679581782
transform 1 0 14400 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_151
timestamp 1679581782
transform 1 0 15072 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_158
timestamp 1679581782
transform 1 0 15744 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_165
timestamp 1679581782
transform 1 0 16416 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_172
timestamp 1679581782
transform 1 0 17088 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_179
timestamp 1679581782
transform 1 0 17760 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_186
timestamp 1679581782
transform 1 0 18432 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_193
timestamp 1679581782
transform 1 0 19104 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_200
timestamp 1679581782
transform 1 0 19776 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_207
timestamp 1679581782
transform 1 0 20448 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_214
timestamp 1679581782
transform 1 0 21120 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_221
timestamp 1679581782
transform 1 0 21792 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_228
timestamp 1679581782
transform 1 0 22464 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_235
timestamp 1679581782
transform 1 0 23136 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_242
timestamp 1679581782
transform 1 0 23808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_249
timestamp 1679581782
transform 1 0 24480 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_256
timestamp 1679581782
transform 1 0 25152 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_263
timestamp 1679581782
transform 1 0 25824 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_270
timestamp 1679581782
transform 1 0 26496 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_277
timestamp 1679581782
transform 1 0 27168 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_284
timestamp 1679581782
transform 1 0 27840 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_291
timestamp 1679581782
transform 1 0 28512 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_298
timestamp 1679581782
transform 1 0 29184 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_305
timestamp 1679581782
transform 1 0 29856 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_312
timestamp 1679581782
transform 1 0 30528 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_319
timestamp 1679581782
transform 1 0 31200 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_326
timestamp 1679581782
transform 1 0 31872 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_333
timestamp 1679581782
transform 1 0 32544 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_340
timestamp 1679581782
transform 1 0 33216 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_347
timestamp 1679581782
transform 1 0 33888 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_354
timestamp 1679581782
transform 1 0 34560 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_361
timestamp 1679581782
transform 1 0 35232 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_368
timestamp 1679581782
transform 1 0 35904 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_375
timestamp 1679581782
transform 1 0 36576 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_382
timestamp 1679581782
transform 1 0 37248 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_389
timestamp 1679581782
transform 1 0 37920 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_396
timestamp 1679581782
transform 1 0 38592 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_403
timestamp 1679581782
transform 1 0 39264 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_410
timestamp 1679581782
transform 1 0 39936 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_417
timestamp 1679581782
transform 1 0 40608 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_424
timestamp 1679581782
transform 1 0 41280 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_431
timestamp 1679581782
transform 1 0 41952 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_438
timestamp 1679581782
transform 1 0 42624 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_445
timestamp 1679581782
transform 1 0 43296 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_452
timestamp 1679581782
transform 1 0 43968 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_459
timestamp 1679581782
transform 1 0 44640 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_466
timestamp 1679581782
transform 1 0 45312 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_473
timestamp 1679581782
transform 1 0 45984 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_480
timestamp 1679581782
transform 1 0 46656 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_487
timestamp 1679581782
transform 1 0 47328 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_494
timestamp 1679581782
transform 1 0 48000 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_501
timestamp 1679581782
transform 1 0 48672 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_508
timestamp 1679581782
transform 1 0 49344 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_515
timestamp 1679581782
transform 1 0 50016 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_522
timestamp 1679581782
transform 1 0 50688 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_529
timestamp 1679581782
transform 1 0 51360 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_536
timestamp 1679581782
transform 1 0 52032 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_543
timestamp 1679581782
transform 1 0 52704 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_550
timestamp 1679581782
transform 1 0 53376 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_557
timestamp 1679581782
transform 1 0 54048 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_564
timestamp 1679581782
transform 1 0 54720 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_571
timestamp 1679581782
transform 1 0 55392 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_578
timestamp 1679581782
transform 1 0 56064 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_585
timestamp 1679581782
transform 1 0 56736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_592
timestamp 1679581782
transform 1 0 57408 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_599
timestamp 1679581782
transform 1 0 58080 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_606
timestamp 1679581782
transform 1 0 58752 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_613
timestamp 1679581782
transform 1 0 59424 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_620
timestamp 1679581782
transform 1 0 60096 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_627
timestamp 1679581782
transform 1 0 60768 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_634
timestamp 1679581782
transform 1 0 61440 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_641
timestamp 1679581782
transform 1 0 62112 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_648
timestamp 1679581782
transform 1 0 62784 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_655
timestamp 1679581782
transform 1 0 63456 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_662
timestamp 1679581782
transform 1 0 64128 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_669
timestamp 1679581782
transform 1 0 64800 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_676
timestamp 1679581782
transform 1 0 65472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_683
timestamp 1679581782
transform 1 0 66144 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_690
timestamp 1679581782
transform 1 0 66816 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_697
timestamp 1679581782
transform 1 0 67488 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_704
timestamp 1679581782
transform 1 0 68160 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_711
timestamp 1679581782
transform 1 0 68832 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_718
timestamp 1679581782
transform 1 0 69504 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_725
timestamp 1679581782
transform 1 0 70176 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_732
timestamp 1679581782
transform 1 0 70848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_739
timestamp 1679581782
transform 1 0 71520 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_746
timestamp 1679581782
transform 1 0 72192 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_753
timestamp 1679581782
transform 1 0 72864 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_760
timestamp 1677580104
transform 1 0 73536 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_762
timestamp 1677579658
transform 1 0 73728 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_771
timestamp 1679581782
transform 1 0 74592 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_778
timestamp 1679581782
transform 1 0 75264 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_785
timestamp 1679581782
transform 1 0 75936 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_792
timestamp 1677579658
transform 1 0 76608 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_801
timestamp 1679581782
transform 1 0 77472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_808
timestamp 1679581782
transform 1 0 78144 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_815
timestamp 1679581782
transform 1 0 78816 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_822
timestamp 1679581782
transform 1 0 79488 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_829
timestamp 1677579658
transform 1 0 80160 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_834
timestamp 1679577901
transform 1 0 80640 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_838
timestamp 1677579658
transform 1 0 81024 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_851
timestamp 1677580104
transform 1 0 82272 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_857
timestamp 1677580104
transform 1 0 82848 0 1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_20_863
timestamp 1677580104
transform 1 0 83424 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_865
timestamp 1677579658
transform 1 0 83616 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_870
timestamp 1679577901
transform 1 0 84096 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_874
timestamp 1677579658
transform 1 0 84480 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_879
timestamp 1679581782
transform 1 0 84960 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_886
timestamp 1679581782
transform 1 0 85632 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_897
timestamp 1679581782
transform 1 0 86688 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_908
timestamp 1677580104
transform 1 0 87744 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_914
timestamp 1679581782
transform 1 0 88320 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_921
timestamp 1677579658
transform 1 0 88992 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_926
timestamp 1679581782
transform 1 0 89472 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_933
timestamp 1679577901
transform 1 0 90144 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_944
timestamp 1679581782
transform 1 0 91200 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_951
timestamp 1677579658
transform 1 0 91872 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_960
timestamp 1679581782
transform 1 0 92736 0 1 15876
box -48 -56 720 834
use sg13g2_decap_4  FILLER_20_967
timestamp 1679577901
transform 1 0 93408 0 1 15876
box -48 -56 432 834
use sg13g2_decap_8  FILLER_20_975
timestamp 1679581782
transform 1 0 94176 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_982
timestamp 1679581782
transform 1 0 94848 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_993
timestamp 1679581782
transform 1 0 95904 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1000
timestamp 1679581782
transform 1 0 96576 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1007
timestamp 1679581782
transform 1 0 97248 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1014
timestamp 1679581782
transform 1 0 97920 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_1021
timestamp 1679581782
transform 1 0 98592 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_1028
timestamp 1677579658
transform 1 0 99264 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_4
timestamp 1679581782
transform 1 0 960 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_11
timestamp 1679581782
transform 1 0 1632 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_18
timestamp 1679581782
transform 1 0 2304 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_25
timestamp 1679581782
transform 1 0 2976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_32
timestamp 1679581782
transform 1 0 3648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_39
timestamp 1679581782
transform 1 0 4320 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_46
timestamp 1679581782
transform 1 0 4992 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_53
timestamp 1679581782
transform 1 0 5664 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_60
timestamp 1679581782
transform 1 0 6336 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_67
timestamp 1679581782
transform 1 0 7008 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_74
timestamp 1679581782
transform 1 0 7680 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_81
timestamp 1679581782
transform 1 0 8352 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_88
timestamp 1679581782
transform 1 0 9024 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_95
timestamp 1679581782
transform 1 0 9696 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_102
timestamp 1679581782
transform 1 0 10368 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_109
timestamp 1679581782
transform 1 0 11040 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_116
timestamp 1679581782
transform 1 0 11712 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_123
timestamp 1679581782
transform 1 0 12384 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_130
timestamp 1679581782
transform 1 0 13056 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_137
timestamp 1679581782
transform 1 0 13728 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_144
timestamp 1679581782
transform 1 0 14400 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_151
timestamp 1679581782
transform 1 0 15072 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_158
timestamp 1679581782
transform 1 0 15744 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_165
timestamp 1679581782
transform 1 0 16416 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_172
timestamp 1679581782
transform 1 0 17088 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_179
timestamp 1679581782
transform 1 0 17760 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_186
timestamp 1679581782
transform 1 0 18432 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_193
timestamp 1679581782
transform 1 0 19104 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_200
timestamp 1679581782
transform 1 0 19776 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_207
timestamp 1679581782
transform 1 0 20448 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_214
timestamp 1679581782
transform 1 0 21120 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_221
timestamp 1679581782
transform 1 0 21792 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_228
timestamp 1679581782
transform 1 0 22464 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_235
timestamp 1679581782
transform 1 0 23136 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_242
timestamp 1679581782
transform 1 0 23808 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_249
timestamp 1679581782
transform 1 0 24480 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_256
timestamp 1679581782
transform 1 0 25152 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_263
timestamp 1679581782
transform 1 0 25824 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_270
timestamp 1679581782
transform 1 0 26496 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_277
timestamp 1679581782
transform 1 0 27168 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_284
timestamp 1679581782
transform 1 0 27840 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_291
timestamp 1679581782
transform 1 0 28512 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_298
timestamp 1679581782
transform 1 0 29184 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_305
timestamp 1679581782
transform 1 0 29856 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_312
timestamp 1679581782
transform 1 0 30528 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_319
timestamp 1679581782
transform 1 0 31200 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_326
timestamp 1679581782
transform 1 0 31872 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_333
timestamp 1679581782
transform 1 0 32544 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_340
timestamp 1679581782
transform 1 0 33216 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_347
timestamp 1679581782
transform 1 0 33888 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_354
timestamp 1679581782
transform 1 0 34560 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_361
timestamp 1679581782
transform 1 0 35232 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_368
timestamp 1679581782
transform 1 0 35904 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_375
timestamp 1679581782
transform 1 0 36576 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_382
timestamp 1679581782
transform 1 0 37248 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_389
timestamp 1679581782
transform 1 0 37920 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_396
timestamp 1679581782
transform 1 0 38592 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_403
timestamp 1679581782
transform 1 0 39264 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_410
timestamp 1679581782
transform 1 0 39936 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_417
timestamp 1679581782
transform 1 0 40608 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_424
timestamp 1679581782
transform 1 0 41280 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_431
timestamp 1679581782
transform 1 0 41952 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_438
timestamp 1679581782
transform 1 0 42624 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_445
timestamp 1679581782
transform 1 0 43296 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_452
timestamp 1679581782
transform 1 0 43968 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_459
timestamp 1679581782
transform 1 0 44640 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_466
timestamp 1679581782
transform 1 0 45312 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_473
timestamp 1679581782
transform 1 0 45984 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_480
timestamp 1679581782
transform 1 0 46656 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_487
timestamp 1679581782
transform 1 0 47328 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_494
timestamp 1679581782
transform 1 0 48000 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_501
timestamp 1679581782
transform 1 0 48672 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_508
timestamp 1679581782
transform 1 0 49344 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_515
timestamp 1679581782
transform 1 0 50016 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_522
timestamp 1679581782
transform 1 0 50688 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_529
timestamp 1679581782
transform 1 0 51360 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_536
timestamp 1679581782
transform 1 0 52032 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_543
timestamp 1679581782
transform 1 0 52704 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_550
timestamp 1679581782
transform 1 0 53376 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_557
timestamp 1679581782
transform 1 0 54048 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_564
timestamp 1679581782
transform 1 0 54720 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_571
timestamp 1679581782
transform 1 0 55392 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_578
timestamp 1679581782
transform 1 0 56064 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_585
timestamp 1679581782
transform 1 0 56736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_592
timestamp 1679581782
transform 1 0 57408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_599
timestamp 1679581782
transform 1 0 58080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_606
timestamp 1679581782
transform 1 0 58752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_613
timestamp 1679581782
transform 1 0 59424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_620
timestamp 1679581782
transform 1 0 60096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_627
timestamp 1679581782
transform 1 0 60768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_634
timestamp 1679581782
transform 1 0 61440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_641
timestamp 1679581782
transform 1 0 62112 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_648
timestamp 1679581782
transform 1 0 62784 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_655
timestamp 1679581782
transform 1 0 63456 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_662
timestamp 1679581782
transform 1 0 64128 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_669
timestamp 1679581782
transform 1 0 64800 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_676
timestamp 1679581782
transform 1 0 65472 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_683
timestamp 1679581782
transform 1 0 66144 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_690
timestamp 1679581782
transform 1 0 66816 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_697
timestamp 1679581782
transform 1 0 67488 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_704
timestamp 1679581782
transform 1 0 68160 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_711
timestamp 1679581782
transform 1 0 68832 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_718
timestamp 1679581782
transform 1 0 69504 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_725
timestamp 1679581782
transform 1 0 70176 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_732
timestamp 1679581782
transform 1 0 70848 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_739
timestamp 1679581782
transform 1 0 71520 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_746
timestamp 1679581782
transform 1 0 72192 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_753
timestamp 1679581782
transform 1 0 72864 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_760
timestamp 1679581782
transform 1 0 73536 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_767
timestamp 1679581782
transform 1 0 74208 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_774
timestamp 1679581782
transform 1 0 74880 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_781
timestamp 1679581782
transform 1 0 75552 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_788
timestamp 1679581782
transform 1 0 76224 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_795
timestamp 1679581782
transform 1 0 76896 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_802
timestamp 1679581782
transform 1 0 77568 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_809
timestamp 1679581782
transform 1 0 78240 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_816
timestamp 1679581782
transform 1 0 78912 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_823
timestamp 1679581782
transform 1 0 79584 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_830
timestamp 1677579658
transform 1 0 80256 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_835
timestamp 1679581782
transform 1 0 80736 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_842
timestamp 1679581782
transform 1 0 81408 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_849
timestamp 1679581782
transform 1 0 82080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_856
timestamp 1679581782
transform 1 0 82752 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_863
timestamp 1679581782
transform 1 0 83424 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_870
timestamp 1679581782
transform 1 0 84096 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_877
timestamp 1679581782
transform 1 0 84768 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_884
timestamp 1679581782
transform 1 0 85440 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_900
timestamp 1679581782
transform 1 0 86976 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_907
timestamp 1679581782
transform 1 0 87648 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_914
timestamp 1679581782
transform 1 0 88320 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_921
timestamp 1679581782
transform 1 0 88992 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_928
timestamp 1679581782
transform 1 0 89664 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_935
timestamp 1679581782
transform 1 0 90336 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_942
timestamp 1679581782
transform 1 0 91008 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_949
timestamp 1679581782
transform 1 0 91680 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_956
timestamp 1679581782
transform 1 0 92352 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_963
timestamp 1679581782
transform 1 0 93024 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_970
timestamp 1679581782
transform 1 0 93696 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_977
timestamp 1679581782
transform 1 0 94368 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_984
timestamp 1679581782
transform 1 0 95040 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_991
timestamp 1679581782
transform 1 0 95712 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_998
timestamp 1679581782
transform 1 0 96384 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1005
timestamp 1679581782
transform 1 0 97056 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1012
timestamp 1679581782
transform 1 0 97728 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_1019
timestamp 1679581782
transform 1 0 98400 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_1026
timestamp 1677580104
transform 1 0 99072 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_1028
timestamp 1677579658
transform 1 0 99264 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_4
timestamp 1679581782
transform 1 0 960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_11
timestamp 1679581782
transform 1 0 1632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_18
timestamp 1679581782
transform 1 0 2304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_25
timestamp 1679581782
transform 1 0 2976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_32
timestamp 1679581782
transform 1 0 3648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_39
timestamp 1679581782
transform 1 0 4320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_46
timestamp 1679581782
transform 1 0 4992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_53
timestamp 1679581782
transform 1 0 5664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_60
timestamp 1679581782
transform 1 0 6336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_67
timestamp 1679581782
transform 1 0 7008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_74
timestamp 1679581782
transform 1 0 7680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_81
timestamp 1679581782
transform 1 0 8352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_88
timestamp 1679581782
transform 1 0 9024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_95
timestamp 1679581782
transform 1 0 9696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_102
timestamp 1679581782
transform 1 0 10368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_109
timestamp 1679581782
transform 1 0 11040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_116
timestamp 1679581782
transform 1 0 11712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_123
timestamp 1679581782
transform 1 0 12384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_130
timestamp 1679581782
transform 1 0 13056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_137
timestamp 1679581782
transform 1 0 13728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_144
timestamp 1679581782
transform 1 0 14400 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_151
timestamp 1679581782
transform 1 0 15072 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_158
timestamp 1679581782
transform 1 0 15744 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_165
timestamp 1679581782
transform 1 0 16416 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_172
timestamp 1679581782
transform 1 0 17088 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_179
timestamp 1679581782
transform 1 0 17760 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_186
timestamp 1679581782
transform 1 0 18432 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_193
timestamp 1679581782
transform 1 0 19104 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_200
timestamp 1679581782
transform 1 0 19776 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_207
timestamp 1679581782
transform 1 0 20448 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_214
timestamp 1679581782
transform 1 0 21120 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_221
timestamp 1679581782
transform 1 0 21792 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_228
timestamp 1679581782
transform 1 0 22464 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_235
timestamp 1679581782
transform 1 0 23136 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_242
timestamp 1679581782
transform 1 0 23808 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_249
timestamp 1679581782
transform 1 0 24480 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_256
timestamp 1679581782
transform 1 0 25152 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_263
timestamp 1679581782
transform 1 0 25824 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_270
timestamp 1679581782
transform 1 0 26496 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_277
timestamp 1679581782
transform 1 0 27168 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_284
timestamp 1679581782
transform 1 0 27840 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_291
timestamp 1679581782
transform 1 0 28512 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_298
timestamp 1679581782
transform 1 0 29184 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_305
timestamp 1679581782
transform 1 0 29856 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_312
timestamp 1679581782
transform 1 0 30528 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_319
timestamp 1679581782
transform 1 0 31200 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_326
timestamp 1679581782
transform 1 0 31872 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_333
timestamp 1679581782
transform 1 0 32544 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_340
timestamp 1679581782
transform 1 0 33216 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_347
timestamp 1679581782
transform 1 0 33888 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_354
timestamp 1679581782
transform 1 0 34560 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_361
timestamp 1679581782
transform 1 0 35232 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_368
timestamp 1679581782
transform 1 0 35904 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_375
timestamp 1679581782
transform 1 0 36576 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_382
timestamp 1679581782
transform 1 0 37248 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_389
timestamp 1679581782
transform 1 0 37920 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_396
timestamp 1679581782
transform 1 0 38592 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_403
timestamp 1679581782
transform 1 0 39264 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_410
timestamp 1679581782
transform 1 0 39936 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_417
timestamp 1679581782
transform 1 0 40608 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_424
timestamp 1679581782
transform 1 0 41280 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_431
timestamp 1679581782
transform 1 0 41952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_438
timestamp 1679581782
transform 1 0 42624 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_445
timestamp 1679581782
transform 1 0 43296 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_452
timestamp 1679581782
transform 1 0 43968 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_459
timestamp 1679581782
transform 1 0 44640 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_466
timestamp 1679581782
transform 1 0 45312 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_473
timestamp 1679581782
transform 1 0 45984 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_480
timestamp 1679581782
transform 1 0 46656 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_487
timestamp 1679581782
transform 1 0 47328 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_494
timestamp 1679581782
transform 1 0 48000 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_501
timestamp 1679581782
transform 1 0 48672 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_508
timestamp 1679581782
transform 1 0 49344 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_515
timestamp 1679581782
transform 1 0 50016 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_522
timestamp 1679581782
transform 1 0 50688 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_529
timestamp 1679581782
transform 1 0 51360 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_536
timestamp 1679581782
transform 1 0 52032 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_543
timestamp 1679581782
transform 1 0 52704 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_550
timestamp 1679581782
transform 1 0 53376 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_557
timestamp 1679581782
transform 1 0 54048 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_564
timestamp 1679581782
transform 1 0 54720 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_571
timestamp 1679581782
transform 1 0 55392 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_578
timestamp 1679581782
transform 1 0 56064 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_585
timestamp 1679581782
transform 1 0 56736 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_592
timestamp 1679581782
transform 1 0 57408 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_599
timestamp 1679581782
transform 1 0 58080 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_606
timestamp 1679581782
transform 1 0 58752 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_613
timestamp 1679581782
transform 1 0 59424 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_620
timestamp 1679581782
transform 1 0 60096 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_627
timestamp 1679581782
transform 1 0 60768 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_634
timestamp 1679581782
transform 1 0 61440 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_641
timestamp 1679581782
transform 1 0 62112 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_648
timestamp 1679581782
transform 1 0 62784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_655
timestamp 1679581782
transform 1 0 63456 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_662
timestamp 1679581782
transform 1 0 64128 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_669
timestamp 1679581782
transform 1 0 64800 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_676
timestamp 1679581782
transform 1 0 65472 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_683
timestamp 1679581782
transform 1 0 66144 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_690
timestamp 1679581782
transform 1 0 66816 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_697
timestamp 1679581782
transform 1 0 67488 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_704
timestamp 1679581782
transform 1 0 68160 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_711
timestamp 1679581782
transform 1 0 68832 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_718
timestamp 1679581782
transform 1 0 69504 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_725
timestamp 1679581782
transform 1 0 70176 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_732
timestamp 1679581782
transform 1 0 70848 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_739
timestamp 1679581782
transform 1 0 71520 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_746
timestamp 1679581782
transform 1 0 72192 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_753
timestamp 1679581782
transform 1 0 72864 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_760
timestamp 1679581782
transform 1 0 73536 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_767
timestamp 1679581782
transform 1 0 74208 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_774
timestamp 1679581782
transform 1 0 74880 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_781
timestamp 1679581782
transform 1 0 75552 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_788
timestamp 1679581782
transform 1 0 76224 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_795
timestamp 1679581782
transform 1 0 76896 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_802
timestamp 1679581782
transform 1 0 77568 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_809
timestamp 1679581782
transform 1 0 78240 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_816
timestamp 1679581782
transform 1 0 78912 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_823
timestamp 1679581782
transform 1 0 79584 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_830
timestamp 1679581782
transform 1 0 80256 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_837
timestamp 1679581782
transform 1 0 80928 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_844
timestamp 1679581782
transform 1 0 81600 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_851
timestamp 1679581782
transform 1 0 82272 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_858
timestamp 1679581782
transform 1 0 82944 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_865
timestamp 1679581782
transform 1 0 83616 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_872
timestamp 1679581782
transform 1 0 84288 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_879
timestamp 1679581782
transform 1 0 84960 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_886
timestamp 1679581782
transform 1 0 85632 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_893
timestamp 1679581782
transform 1 0 86304 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_900
timestamp 1679581782
transform 1 0 86976 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_907
timestamp 1679581782
transform 1 0 87648 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_914
timestamp 1679581782
transform 1 0 88320 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_921
timestamp 1679581782
transform 1 0 88992 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_928
timestamp 1679581782
transform 1 0 89664 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_935
timestamp 1679581782
transform 1 0 90336 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_942
timestamp 1679581782
transform 1 0 91008 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_949
timestamp 1679581782
transform 1 0 91680 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_956
timestamp 1679581782
transform 1 0 92352 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_963
timestamp 1679581782
transform 1 0 93024 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_970
timestamp 1679581782
transform 1 0 93696 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_977
timestamp 1679581782
transform 1 0 94368 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_984
timestamp 1679581782
transform 1 0 95040 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_991
timestamp 1679581782
transform 1 0 95712 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_998
timestamp 1679581782
transform 1 0 96384 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1005
timestamp 1679581782
transform 1 0 97056 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1012
timestamp 1679581782
transform 1 0 97728 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_1019
timestamp 1679581782
transform 1 0 98400 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_1026
timestamp 1677580104
transform 1 0 99072 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_1028
timestamp 1677579658
transform 1 0 99264 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_4
timestamp 1679581782
transform 1 0 960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_11
timestamp 1679581782
transform 1 0 1632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_18
timestamp 1679581782
transform 1 0 2304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_25
timestamp 1679581782
transform 1 0 2976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_32
timestamp 1679581782
transform 1 0 3648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_39
timestamp 1679581782
transform 1 0 4320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_46
timestamp 1679581782
transform 1 0 4992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_53
timestamp 1679581782
transform 1 0 5664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_60
timestamp 1679581782
transform 1 0 6336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_67
timestamp 1679581782
transform 1 0 7008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_74
timestamp 1679581782
transform 1 0 7680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_81
timestamp 1679581782
transform 1 0 8352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_88
timestamp 1679581782
transform 1 0 9024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_95
timestamp 1679581782
transform 1 0 9696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_102
timestamp 1679581782
transform 1 0 10368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_109
timestamp 1679581782
transform 1 0 11040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_116
timestamp 1679581782
transform 1 0 11712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_123
timestamp 1679581782
transform 1 0 12384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_130
timestamp 1679581782
transform 1 0 13056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_137
timestamp 1679581782
transform 1 0 13728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_144
timestamp 1679581782
transform 1 0 14400 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_151
timestamp 1679581782
transform 1 0 15072 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_158
timestamp 1679581782
transform 1 0 15744 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_165
timestamp 1679581782
transform 1 0 16416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_172
timestamp 1679581782
transform 1 0 17088 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_179
timestamp 1679581782
transform 1 0 17760 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_186
timestamp 1679581782
transform 1 0 18432 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_193
timestamp 1679581782
transform 1 0 19104 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_200
timestamp 1679581782
transform 1 0 19776 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_207
timestamp 1679581782
transform 1 0 20448 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_214
timestamp 1679581782
transform 1 0 21120 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_221
timestamp 1679581782
transform 1 0 21792 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_228
timestamp 1679581782
transform 1 0 22464 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_235
timestamp 1679581782
transform 1 0 23136 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_242
timestamp 1679581782
transform 1 0 23808 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_249
timestamp 1679581782
transform 1 0 24480 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_256
timestamp 1679581782
transform 1 0 25152 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_263
timestamp 1679581782
transform 1 0 25824 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_270
timestamp 1679581782
transform 1 0 26496 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_277
timestamp 1679581782
transform 1 0 27168 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_284
timestamp 1679581782
transform 1 0 27840 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_291
timestamp 1679581782
transform 1 0 28512 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_298
timestamp 1679581782
transform 1 0 29184 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_305
timestamp 1679581782
transform 1 0 29856 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_312
timestamp 1679581782
transform 1 0 30528 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_319
timestamp 1679581782
transform 1 0 31200 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_326
timestamp 1679581782
transform 1 0 31872 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_333
timestamp 1679581782
transform 1 0 32544 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_340
timestamp 1679581782
transform 1 0 33216 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_347
timestamp 1679581782
transform 1 0 33888 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_354
timestamp 1679581782
transform 1 0 34560 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_361
timestamp 1679581782
transform 1 0 35232 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_368
timestamp 1679581782
transform 1 0 35904 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_375
timestamp 1679581782
transform 1 0 36576 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_382
timestamp 1679581782
transform 1 0 37248 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_389
timestamp 1679581782
transform 1 0 37920 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_396
timestamp 1679581782
transform 1 0 38592 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_403
timestamp 1679581782
transform 1 0 39264 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_410
timestamp 1679581782
transform 1 0 39936 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_417
timestamp 1679581782
transform 1 0 40608 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_424
timestamp 1679581782
transform 1 0 41280 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_431
timestamp 1679581782
transform 1 0 41952 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_438
timestamp 1679581782
transform 1 0 42624 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_445
timestamp 1679581782
transform 1 0 43296 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_452
timestamp 1679581782
transform 1 0 43968 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_459
timestamp 1679581782
transform 1 0 44640 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_466
timestamp 1679581782
transform 1 0 45312 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_473
timestamp 1679581782
transform 1 0 45984 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_480
timestamp 1679581782
transform 1 0 46656 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_487
timestamp 1679581782
transform 1 0 47328 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_494
timestamp 1679581782
transform 1 0 48000 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_501
timestamp 1679581782
transform 1 0 48672 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_508
timestamp 1679581782
transform 1 0 49344 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_515
timestamp 1679581782
transform 1 0 50016 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_522
timestamp 1679581782
transform 1 0 50688 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_529
timestamp 1679581782
transform 1 0 51360 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_536
timestamp 1679581782
transform 1 0 52032 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_543
timestamp 1679581782
transform 1 0 52704 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_550
timestamp 1679581782
transform 1 0 53376 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_557
timestamp 1679581782
transform 1 0 54048 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_564
timestamp 1679581782
transform 1 0 54720 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_571
timestamp 1679581782
transform 1 0 55392 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_578
timestamp 1679581782
transform 1 0 56064 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_585
timestamp 1679581782
transform 1 0 56736 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_592
timestamp 1679581782
transform 1 0 57408 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_599
timestamp 1679581782
transform 1 0 58080 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_606
timestamp 1679581782
transform 1 0 58752 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_613
timestamp 1679581782
transform 1 0 59424 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_620
timestamp 1679581782
transform 1 0 60096 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_627
timestamp 1679581782
transform 1 0 60768 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_634
timestamp 1679581782
transform 1 0 61440 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_641
timestamp 1679581782
transform 1 0 62112 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_648
timestamp 1679581782
transform 1 0 62784 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_655
timestamp 1679581782
transform 1 0 63456 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_662
timestamp 1679581782
transform 1 0 64128 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_669
timestamp 1679581782
transform 1 0 64800 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_676
timestamp 1679581782
transform 1 0 65472 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_683
timestamp 1679581782
transform 1 0 66144 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_690
timestamp 1679581782
transform 1 0 66816 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_697
timestamp 1679581782
transform 1 0 67488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_704
timestamp 1679581782
transform 1 0 68160 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_711
timestamp 1679581782
transform 1 0 68832 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_718
timestamp 1679581782
transform 1 0 69504 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_725
timestamp 1679581782
transform 1 0 70176 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_732
timestamp 1679581782
transform 1 0 70848 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_739
timestamp 1679581782
transform 1 0 71520 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_746
timestamp 1679581782
transform 1 0 72192 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_753
timestamp 1679581782
transform 1 0 72864 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_760
timestamp 1679581782
transform 1 0 73536 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_767
timestamp 1679581782
transform 1 0 74208 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_774
timestamp 1679581782
transform 1 0 74880 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_781
timestamp 1679581782
transform 1 0 75552 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_788
timestamp 1679581782
transform 1 0 76224 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_795
timestamp 1679581782
transform 1 0 76896 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_802
timestamp 1679581782
transform 1 0 77568 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_809
timestamp 1679581782
transform 1 0 78240 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_816
timestamp 1679581782
transform 1 0 78912 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_823
timestamp 1679581782
transform 1 0 79584 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_830
timestamp 1679581782
transform 1 0 80256 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_837
timestamp 1679581782
transform 1 0 80928 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_844
timestamp 1679581782
transform 1 0 81600 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_851
timestamp 1679581782
transform 1 0 82272 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_858
timestamp 1679581782
transform 1 0 82944 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_865
timestamp 1679581782
transform 1 0 83616 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_872
timestamp 1679581782
transform 1 0 84288 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_879
timestamp 1679581782
transform 1 0 84960 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_886
timestamp 1679581782
transform 1 0 85632 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_893
timestamp 1679581782
transform 1 0 86304 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_900
timestamp 1679581782
transform 1 0 86976 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_907
timestamp 1679581782
transform 1 0 87648 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_914
timestamp 1679581782
transform 1 0 88320 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_921
timestamp 1679581782
transform 1 0 88992 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_928
timestamp 1679581782
transform 1 0 89664 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_935
timestamp 1679581782
transform 1 0 90336 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_942
timestamp 1679581782
transform 1 0 91008 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_949
timestamp 1679581782
transform 1 0 91680 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_956
timestamp 1679581782
transform 1 0 92352 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_963
timestamp 1679581782
transform 1 0 93024 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_970
timestamp 1679581782
transform 1 0 93696 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_977
timestamp 1679581782
transform 1 0 94368 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_984
timestamp 1679581782
transform 1 0 95040 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_991
timestamp 1679581782
transform 1 0 95712 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_998
timestamp 1679581782
transform 1 0 96384 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1005
timestamp 1679581782
transform 1 0 97056 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1012
timestamp 1679581782
transform 1 0 97728 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_1019
timestamp 1679581782
transform 1 0 98400 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_1026
timestamp 1677580104
transform 1 0 99072 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_1028
timestamp 1677579658
transform 1 0 99264 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_4
timestamp 1679581782
transform 1 0 960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_11
timestamp 1679581782
transform 1 0 1632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_18
timestamp 1679581782
transform 1 0 2304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_25
timestamp 1679581782
transform 1 0 2976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_32
timestamp 1679581782
transform 1 0 3648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_39
timestamp 1679581782
transform 1 0 4320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_46
timestamp 1679581782
transform 1 0 4992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_53
timestamp 1679581782
transform 1 0 5664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_60
timestamp 1679581782
transform 1 0 6336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_67
timestamp 1679581782
transform 1 0 7008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_74
timestamp 1679581782
transform 1 0 7680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_81
timestamp 1679581782
transform 1 0 8352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_88
timestamp 1679581782
transform 1 0 9024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_95
timestamp 1679581782
transform 1 0 9696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_102
timestamp 1679581782
transform 1 0 10368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_109
timestamp 1679581782
transform 1 0 11040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_116
timestamp 1679581782
transform 1 0 11712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_123
timestamp 1679581782
transform 1 0 12384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_130
timestamp 1679581782
transform 1 0 13056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_137
timestamp 1679581782
transform 1 0 13728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_144
timestamp 1679581782
transform 1 0 14400 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_151
timestamp 1679581782
transform 1 0 15072 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_158
timestamp 1679581782
transform 1 0 15744 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_165
timestamp 1679581782
transform 1 0 16416 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_172
timestamp 1679581782
transform 1 0 17088 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_179
timestamp 1679581782
transform 1 0 17760 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_186
timestamp 1679581782
transform 1 0 18432 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_193
timestamp 1679581782
transform 1 0 19104 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_200
timestamp 1679581782
transform 1 0 19776 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_207
timestamp 1679581782
transform 1 0 20448 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_214
timestamp 1679581782
transform 1 0 21120 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_221
timestamp 1679581782
transform 1 0 21792 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_228
timestamp 1679581782
transform 1 0 22464 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_235
timestamp 1679581782
transform 1 0 23136 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_242
timestamp 1679581782
transform 1 0 23808 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_249
timestamp 1679581782
transform 1 0 24480 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_256
timestamp 1679581782
transform 1 0 25152 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_263
timestamp 1679581782
transform 1 0 25824 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_270
timestamp 1679581782
transform 1 0 26496 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_277
timestamp 1679581782
transform 1 0 27168 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_284
timestamp 1679581782
transform 1 0 27840 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_291
timestamp 1679581782
transform 1 0 28512 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_298
timestamp 1679581782
transform 1 0 29184 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_305
timestamp 1679581782
transform 1 0 29856 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_312
timestamp 1679581782
transform 1 0 30528 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_319
timestamp 1679581782
transform 1 0 31200 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_326
timestamp 1679581782
transform 1 0 31872 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_333
timestamp 1679581782
transform 1 0 32544 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_340
timestamp 1679581782
transform 1 0 33216 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_347
timestamp 1679581782
transform 1 0 33888 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_354
timestamp 1679581782
transform 1 0 34560 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_361
timestamp 1679581782
transform 1 0 35232 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_368
timestamp 1679581782
transform 1 0 35904 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_375
timestamp 1679581782
transform 1 0 36576 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_382
timestamp 1679581782
transform 1 0 37248 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_389
timestamp 1679581782
transform 1 0 37920 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_396
timestamp 1679581782
transform 1 0 38592 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_403
timestamp 1679581782
transform 1 0 39264 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_410
timestamp 1679581782
transform 1 0 39936 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_417
timestamp 1679581782
transform 1 0 40608 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_424
timestamp 1679581782
transform 1 0 41280 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_431
timestamp 1679581782
transform 1 0 41952 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_438
timestamp 1679581782
transform 1 0 42624 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_445
timestamp 1679581782
transform 1 0 43296 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_452
timestamp 1679581782
transform 1 0 43968 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_459
timestamp 1679581782
transform 1 0 44640 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_466
timestamp 1679581782
transform 1 0 45312 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_473
timestamp 1679581782
transform 1 0 45984 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_480
timestamp 1679581782
transform 1 0 46656 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_487
timestamp 1679581782
transform 1 0 47328 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_494
timestamp 1679581782
transform 1 0 48000 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_501
timestamp 1679581782
transform 1 0 48672 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_508
timestamp 1679581782
transform 1 0 49344 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_515
timestamp 1679581782
transform 1 0 50016 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_522
timestamp 1679581782
transform 1 0 50688 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_529
timestamp 1679581782
transform 1 0 51360 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_536
timestamp 1679581782
transform 1 0 52032 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_543
timestamp 1679581782
transform 1 0 52704 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_550
timestamp 1679581782
transform 1 0 53376 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_557
timestamp 1679581782
transform 1 0 54048 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_564
timestamp 1679581782
transform 1 0 54720 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_571
timestamp 1679581782
transform 1 0 55392 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_578
timestamp 1679581782
transform 1 0 56064 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_585
timestamp 1679581782
transform 1 0 56736 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_592
timestamp 1679581782
transform 1 0 57408 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_599
timestamp 1679581782
transform 1 0 58080 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_606
timestamp 1679581782
transform 1 0 58752 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_613
timestamp 1679581782
transform 1 0 59424 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_620
timestamp 1679581782
transform 1 0 60096 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_627
timestamp 1679581782
transform 1 0 60768 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_634
timestamp 1679581782
transform 1 0 61440 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_641
timestamp 1679581782
transform 1 0 62112 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_648
timestamp 1679581782
transform 1 0 62784 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_655
timestamp 1679581782
transform 1 0 63456 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_662
timestamp 1679581782
transform 1 0 64128 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_669
timestamp 1679581782
transform 1 0 64800 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_676
timestamp 1679581782
transform 1 0 65472 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_683
timestamp 1679581782
transform 1 0 66144 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_690
timestamp 1679581782
transform 1 0 66816 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_697
timestamp 1679581782
transform 1 0 67488 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_704
timestamp 1679581782
transform 1 0 68160 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_711
timestamp 1679581782
transform 1 0 68832 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_718
timestamp 1679581782
transform 1 0 69504 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_725
timestamp 1679581782
transform 1 0 70176 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_732
timestamp 1679581782
transform 1 0 70848 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_739
timestamp 1679581782
transform 1 0 71520 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_746
timestamp 1679581782
transform 1 0 72192 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_753
timestamp 1679581782
transform 1 0 72864 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_760
timestamp 1679581782
transform 1 0 73536 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_767
timestamp 1679581782
transform 1 0 74208 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_774
timestamp 1679581782
transform 1 0 74880 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_781
timestamp 1679581782
transform 1 0 75552 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_788
timestamp 1679581782
transform 1 0 76224 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_795
timestamp 1679581782
transform 1 0 76896 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_802
timestamp 1679581782
transform 1 0 77568 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_809
timestamp 1679581782
transform 1 0 78240 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_816
timestamp 1679581782
transform 1 0 78912 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_823
timestamp 1679581782
transform 1 0 79584 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_830
timestamp 1679581782
transform 1 0 80256 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_837
timestamp 1679581782
transform 1 0 80928 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_844
timestamp 1679581782
transform 1 0 81600 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_851
timestamp 1679581782
transform 1 0 82272 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_858
timestamp 1679581782
transform 1 0 82944 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_865
timestamp 1679581782
transform 1 0 83616 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_872
timestamp 1679581782
transform 1 0 84288 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_879
timestamp 1679581782
transform 1 0 84960 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_886
timestamp 1679581782
transform 1 0 85632 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_893
timestamp 1679581782
transform 1 0 86304 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_900
timestamp 1679581782
transform 1 0 86976 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_907
timestamp 1679581782
transform 1 0 87648 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_914
timestamp 1679581782
transform 1 0 88320 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_921
timestamp 1679581782
transform 1 0 88992 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_928
timestamp 1679581782
transform 1 0 89664 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_935
timestamp 1679581782
transform 1 0 90336 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_942
timestamp 1679581782
transform 1 0 91008 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_949
timestamp 1679581782
transform 1 0 91680 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_956
timestamp 1679581782
transform 1 0 92352 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_963
timestamp 1679581782
transform 1 0 93024 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_970
timestamp 1679581782
transform 1 0 93696 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_977
timestamp 1679581782
transform 1 0 94368 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_984
timestamp 1679581782
transform 1 0 95040 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_991
timestamp 1679581782
transform 1 0 95712 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_998
timestamp 1679581782
transform 1 0 96384 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1005
timestamp 1679581782
transform 1 0 97056 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1012
timestamp 1679581782
transform 1 0 97728 0 1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_1019
timestamp 1679581782
transform 1 0 98400 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_1026
timestamp 1677580104
transform 1 0 99072 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_1028
timestamp 1677579658
transform 1 0 99264 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_4
timestamp 1679581782
transform 1 0 960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_11
timestamp 1679581782
transform 1 0 1632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_18
timestamp 1679581782
transform 1 0 2304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_25
timestamp 1679581782
transform 1 0 2976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_32
timestamp 1679581782
transform 1 0 3648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_39
timestamp 1679581782
transform 1 0 4320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_46
timestamp 1679581782
transform 1 0 4992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_53
timestamp 1679581782
transform 1 0 5664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_60
timestamp 1679581782
transform 1 0 6336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_67
timestamp 1679581782
transform 1 0 7008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_74
timestamp 1679581782
transform 1 0 7680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_81
timestamp 1679581782
transform 1 0 8352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_88
timestamp 1679581782
transform 1 0 9024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_95
timestamp 1679581782
transform 1 0 9696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_102
timestamp 1679581782
transform 1 0 10368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_109
timestamp 1679581782
transform 1 0 11040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_116
timestamp 1679581782
transform 1 0 11712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_123
timestamp 1679581782
transform 1 0 12384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_130
timestamp 1679581782
transform 1 0 13056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_137
timestamp 1679581782
transform 1 0 13728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_144
timestamp 1679581782
transform 1 0 14400 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_151
timestamp 1679581782
transform 1 0 15072 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_158
timestamp 1679581782
transform 1 0 15744 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_165
timestamp 1679581782
transform 1 0 16416 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_172
timestamp 1679581782
transform 1 0 17088 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_179
timestamp 1679581782
transform 1 0 17760 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_186
timestamp 1679581782
transform 1 0 18432 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_193
timestamp 1679581782
transform 1 0 19104 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_200
timestamp 1679581782
transform 1 0 19776 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_207
timestamp 1679581782
transform 1 0 20448 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_214
timestamp 1679581782
transform 1 0 21120 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_221
timestamp 1679581782
transform 1 0 21792 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_228
timestamp 1679581782
transform 1 0 22464 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_235
timestamp 1679581782
transform 1 0 23136 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_242
timestamp 1679581782
transform 1 0 23808 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_249
timestamp 1679581782
transform 1 0 24480 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_256
timestamp 1679581782
transform 1 0 25152 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_263
timestamp 1679581782
transform 1 0 25824 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_270
timestamp 1679581782
transform 1 0 26496 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_277
timestamp 1679581782
transform 1 0 27168 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_284
timestamp 1679581782
transform 1 0 27840 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_291
timestamp 1679581782
transform 1 0 28512 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_298
timestamp 1679581782
transform 1 0 29184 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_305
timestamp 1679581782
transform 1 0 29856 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_312
timestamp 1679581782
transform 1 0 30528 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_319
timestamp 1679581782
transform 1 0 31200 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_326
timestamp 1679581782
transform 1 0 31872 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_333
timestamp 1679581782
transform 1 0 32544 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_340
timestamp 1679581782
transform 1 0 33216 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_347
timestamp 1679581782
transform 1 0 33888 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_354
timestamp 1679581782
transform 1 0 34560 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_361
timestamp 1679581782
transform 1 0 35232 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_368
timestamp 1679581782
transform 1 0 35904 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_375
timestamp 1679581782
transform 1 0 36576 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_382
timestamp 1679581782
transform 1 0 37248 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_389
timestamp 1679581782
transform 1 0 37920 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_396
timestamp 1679581782
transform 1 0 38592 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_403
timestamp 1679581782
transform 1 0 39264 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_410
timestamp 1679581782
transform 1 0 39936 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_417
timestamp 1679581782
transform 1 0 40608 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_424
timestamp 1679581782
transform 1 0 41280 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_431
timestamp 1679581782
transform 1 0 41952 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_438
timestamp 1679581782
transform 1 0 42624 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_445
timestamp 1679581782
transform 1 0 43296 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_452
timestamp 1679581782
transform 1 0 43968 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_459
timestamp 1679581782
transform 1 0 44640 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_466
timestamp 1679581782
transform 1 0 45312 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_473
timestamp 1679581782
transform 1 0 45984 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_480
timestamp 1679581782
transform 1 0 46656 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_487
timestamp 1679581782
transform 1 0 47328 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_494
timestamp 1679581782
transform 1 0 48000 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_501
timestamp 1679581782
transform 1 0 48672 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_508
timestamp 1679581782
transform 1 0 49344 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_515
timestamp 1679581782
transform 1 0 50016 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_522
timestamp 1679581782
transform 1 0 50688 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_529
timestamp 1679581782
transform 1 0 51360 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_536
timestamp 1679581782
transform 1 0 52032 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_543
timestamp 1679581782
transform 1 0 52704 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_550
timestamp 1679581782
transform 1 0 53376 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_557
timestamp 1679581782
transform 1 0 54048 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_564
timestamp 1679581782
transform 1 0 54720 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_571
timestamp 1679581782
transform 1 0 55392 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_578
timestamp 1679581782
transform 1 0 56064 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_585
timestamp 1679581782
transform 1 0 56736 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_592
timestamp 1679581782
transform 1 0 57408 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_599
timestamp 1679581782
transform 1 0 58080 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_606
timestamp 1679581782
transform 1 0 58752 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_613
timestamp 1679581782
transform 1 0 59424 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_620
timestamp 1679581782
transform 1 0 60096 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_627
timestamp 1679581782
transform 1 0 60768 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_634
timestamp 1679581782
transform 1 0 61440 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_641
timestamp 1679581782
transform 1 0 62112 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_648
timestamp 1679581782
transform 1 0 62784 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_655
timestamp 1679581782
transform 1 0 63456 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_662
timestamp 1679581782
transform 1 0 64128 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_669
timestamp 1679581782
transform 1 0 64800 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_676
timestamp 1679581782
transform 1 0 65472 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_683
timestamp 1679581782
transform 1 0 66144 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_690
timestamp 1679581782
transform 1 0 66816 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_697
timestamp 1679581782
transform 1 0 67488 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_704
timestamp 1679581782
transform 1 0 68160 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_711
timestamp 1679581782
transform 1 0 68832 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_718
timestamp 1679581782
transform 1 0 69504 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_725
timestamp 1679581782
transform 1 0 70176 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_732
timestamp 1679581782
transform 1 0 70848 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_739
timestamp 1679581782
transform 1 0 71520 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_746
timestamp 1679581782
transform 1 0 72192 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_753
timestamp 1679581782
transform 1 0 72864 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_760
timestamp 1679581782
transform 1 0 73536 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_767
timestamp 1679581782
transform 1 0 74208 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_774
timestamp 1679581782
transform 1 0 74880 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_781
timestamp 1679581782
transform 1 0 75552 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_788
timestamp 1679581782
transform 1 0 76224 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_795
timestamp 1679581782
transform 1 0 76896 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_802
timestamp 1679581782
transform 1 0 77568 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_809
timestamp 1679581782
transform 1 0 78240 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_816
timestamp 1679581782
transform 1 0 78912 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_823
timestamp 1679581782
transform 1 0 79584 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_830
timestamp 1679581782
transform 1 0 80256 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_837
timestamp 1679581782
transform 1 0 80928 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_844
timestamp 1679581782
transform 1 0 81600 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_851
timestamp 1679581782
transform 1 0 82272 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_858
timestamp 1679581782
transform 1 0 82944 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_865
timestamp 1679581782
transform 1 0 83616 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_872
timestamp 1679581782
transform 1 0 84288 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_879
timestamp 1679581782
transform 1 0 84960 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_886
timestamp 1679581782
transform 1 0 85632 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_893
timestamp 1679581782
transform 1 0 86304 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_900
timestamp 1679581782
transform 1 0 86976 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_907
timestamp 1679581782
transform 1 0 87648 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_914
timestamp 1679581782
transform 1 0 88320 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_921
timestamp 1679581782
transform 1 0 88992 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_928
timestamp 1679581782
transform 1 0 89664 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_935
timestamp 1679581782
transform 1 0 90336 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_942
timestamp 1679581782
transform 1 0 91008 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_949
timestamp 1679581782
transform 1 0 91680 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_956
timestamp 1679581782
transform 1 0 92352 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_963
timestamp 1679581782
transform 1 0 93024 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_970
timestamp 1679581782
transform 1 0 93696 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_977
timestamp 1679581782
transform 1 0 94368 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_984
timestamp 1679581782
transform 1 0 95040 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_991
timestamp 1679581782
transform 1 0 95712 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_998
timestamp 1679581782
transform 1 0 96384 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1005
timestamp 1679581782
transform 1 0 97056 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1012
timestamp 1679581782
transform 1 0 97728 0 -1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_1019
timestamp 1679581782
transform 1 0 98400 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_1026
timestamp 1677580104
transform 1 0 99072 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_1028
timestamp 1677579658
transform 1 0 99264 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_4
timestamp 1679581782
transform 1 0 960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_11
timestamp 1679581782
transform 1 0 1632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_18
timestamp 1679581782
transform 1 0 2304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_25
timestamp 1679581782
transform 1 0 2976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_32
timestamp 1679581782
transform 1 0 3648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_39
timestamp 1679581782
transform 1 0 4320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_46
timestamp 1679581782
transform 1 0 4992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_53
timestamp 1679581782
transform 1 0 5664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_60
timestamp 1679581782
transform 1 0 6336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_67
timestamp 1679581782
transform 1 0 7008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_74
timestamp 1679581782
transform 1 0 7680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_81
timestamp 1679581782
transform 1 0 8352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_88
timestamp 1679581782
transform 1 0 9024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_95
timestamp 1679581782
transform 1 0 9696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_102
timestamp 1679581782
transform 1 0 10368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_109
timestamp 1679581782
transform 1 0 11040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_116
timestamp 1679581782
transform 1 0 11712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_123
timestamp 1679581782
transform 1 0 12384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_130
timestamp 1679581782
transform 1 0 13056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_137
timestamp 1679581782
transform 1 0 13728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_144
timestamp 1679581782
transform 1 0 14400 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_151
timestamp 1679581782
transform 1 0 15072 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_158
timestamp 1679581782
transform 1 0 15744 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_165
timestamp 1679581782
transform 1 0 16416 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_172
timestamp 1679581782
transform 1 0 17088 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_179
timestamp 1679581782
transform 1 0 17760 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_186
timestamp 1679581782
transform 1 0 18432 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_193
timestamp 1679581782
transform 1 0 19104 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_200
timestamp 1679581782
transform 1 0 19776 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_207
timestamp 1679581782
transform 1 0 20448 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_214
timestamp 1679581782
transform 1 0 21120 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_221
timestamp 1679581782
transform 1 0 21792 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_228
timestamp 1679581782
transform 1 0 22464 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_235
timestamp 1679581782
transform 1 0 23136 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_242
timestamp 1679581782
transform 1 0 23808 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_249
timestamp 1679581782
transform 1 0 24480 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_256
timestamp 1679581782
transform 1 0 25152 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_263
timestamp 1679581782
transform 1 0 25824 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_270
timestamp 1679581782
transform 1 0 26496 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_277
timestamp 1679581782
transform 1 0 27168 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_284
timestamp 1679581782
transform 1 0 27840 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_291
timestamp 1679581782
transform 1 0 28512 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_298
timestamp 1679581782
transform 1 0 29184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_305
timestamp 1679581782
transform 1 0 29856 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_312
timestamp 1679581782
transform 1 0 30528 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_319
timestamp 1679581782
transform 1 0 31200 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_326
timestamp 1679581782
transform 1 0 31872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_333
timestamp 1679581782
transform 1 0 32544 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_340
timestamp 1679581782
transform 1 0 33216 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_347
timestamp 1679581782
transform 1 0 33888 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_354
timestamp 1679581782
transform 1 0 34560 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_361
timestamp 1679581782
transform 1 0 35232 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_368
timestamp 1679581782
transform 1 0 35904 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_375
timestamp 1679581782
transform 1 0 36576 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_382
timestamp 1679581782
transform 1 0 37248 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_389
timestamp 1679581782
transform 1 0 37920 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_396
timestamp 1679581782
transform 1 0 38592 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_403
timestamp 1679581782
transform 1 0 39264 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_410
timestamp 1679581782
transform 1 0 39936 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_417
timestamp 1679581782
transform 1 0 40608 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_424
timestamp 1679581782
transform 1 0 41280 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_431
timestamp 1679581782
transform 1 0 41952 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_438
timestamp 1679581782
transform 1 0 42624 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_445
timestamp 1679581782
transform 1 0 43296 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_452
timestamp 1679581782
transform 1 0 43968 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_459
timestamp 1679581782
transform 1 0 44640 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_466
timestamp 1679581782
transform 1 0 45312 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_473
timestamp 1679581782
transform 1 0 45984 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_480
timestamp 1679581782
transform 1 0 46656 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_487
timestamp 1679581782
transform 1 0 47328 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_494
timestamp 1679581782
transform 1 0 48000 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_501
timestamp 1679581782
transform 1 0 48672 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_508
timestamp 1679581782
transform 1 0 49344 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_515
timestamp 1679581782
transform 1 0 50016 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_522
timestamp 1679581782
transform 1 0 50688 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_529
timestamp 1679581782
transform 1 0 51360 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_536
timestamp 1679581782
transform 1 0 52032 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_543
timestamp 1679581782
transform 1 0 52704 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_550
timestamp 1679581782
transform 1 0 53376 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_557
timestamp 1679581782
transform 1 0 54048 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_564
timestamp 1679581782
transform 1 0 54720 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_571
timestamp 1679581782
transform 1 0 55392 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_578
timestamp 1679581782
transform 1 0 56064 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_585
timestamp 1679581782
transform 1 0 56736 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_592
timestamp 1679581782
transform 1 0 57408 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_599
timestamp 1679581782
transform 1 0 58080 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_606
timestamp 1679581782
transform 1 0 58752 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_613
timestamp 1679581782
transform 1 0 59424 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_620
timestamp 1679581782
transform 1 0 60096 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_627
timestamp 1679581782
transform 1 0 60768 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_634
timestamp 1679581782
transform 1 0 61440 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_641
timestamp 1679581782
transform 1 0 62112 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_648
timestamp 1679581782
transform 1 0 62784 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_655
timestamp 1679581782
transform 1 0 63456 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_662
timestamp 1679581782
transform 1 0 64128 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_669
timestamp 1679581782
transform 1 0 64800 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_676
timestamp 1679581782
transform 1 0 65472 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_683
timestamp 1679581782
transform 1 0 66144 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_690
timestamp 1679581782
transform 1 0 66816 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_697
timestamp 1679581782
transform 1 0 67488 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_704
timestamp 1679581782
transform 1 0 68160 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_711
timestamp 1679581782
transform 1 0 68832 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_718
timestamp 1679581782
transform 1 0 69504 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_725
timestamp 1679581782
transform 1 0 70176 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_732
timestamp 1679581782
transform 1 0 70848 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_739
timestamp 1679581782
transform 1 0 71520 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_746
timestamp 1679581782
transform 1 0 72192 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_753
timestamp 1679581782
transform 1 0 72864 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_760
timestamp 1679581782
transform 1 0 73536 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_767
timestamp 1679581782
transform 1 0 74208 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_774
timestamp 1679581782
transform 1 0 74880 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_781
timestamp 1679581782
transform 1 0 75552 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_788
timestamp 1679581782
transform 1 0 76224 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_795
timestamp 1679581782
transform 1 0 76896 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_802
timestamp 1679581782
transform 1 0 77568 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_809
timestamp 1679581782
transform 1 0 78240 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_816
timestamp 1679581782
transform 1 0 78912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_823
timestamp 1679581782
transform 1 0 79584 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_830
timestamp 1679581782
transform 1 0 80256 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_837
timestamp 1679581782
transform 1 0 80928 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_844
timestamp 1679581782
transform 1 0 81600 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_851
timestamp 1679581782
transform 1 0 82272 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_858
timestamp 1679581782
transform 1 0 82944 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_865
timestamp 1679581782
transform 1 0 83616 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_872
timestamp 1679581782
transform 1 0 84288 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_879
timestamp 1679581782
transform 1 0 84960 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_886
timestamp 1679581782
transform 1 0 85632 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_893
timestamp 1679581782
transform 1 0 86304 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_900
timestamp 1679581782
transform 1 0 86976 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_907
timestamp 1679581782
transform 1 0 87648 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_914
timestamp 1679581782
transform 1 0 88320 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_921
timestamp 1679581782
transform 1 0 88992 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_928
timestamp 1679581782
transform 1 0 89664 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_935
timestamp 1679581782
transform 1 0 90336 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_942
timestamp 1679581782
transform 1 0 91008 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_949
timestamp 1679581782
transform 1 0 91680 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_956
timestamp 1679581782
transform 1 0 92352 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_963
timestamp 1679581782
transform 1 0 93024 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_970
timestamp 1679581782
transform 1 0 93696 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_977
timestamp 1679581782
transform 1 0 94368 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_984
timestamp 1679581782
transform 1 0 95040 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_991
timestamp 1679581782
transform 1 0 95712 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_998
timestamp 1679581782
transform 1 0 96384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1005
timestamp 1679581782
transform 1 0 97056 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1012
timestamp 1679581782
transform 1 0 97728 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_1019
timestamp 1679581782
transform 1 0 98400 0 1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_1026
timestamp 1677580104
transform 1 0 99072 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_1028
timestamp 1677579658
transform 1 0 99264 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 1248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 1920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679581782
transform 1 0 2592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_28
timestamp 1679581782
transform 1 0 3264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_35
timestamp 1679581782
transform 1 0 3936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_42
timestamp 1679581782
transform 1 0 4608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_49
timestamp 1679581782
transform 1 0 5280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_56
timestamp 1679581782
transform 1 0 5952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_63
timestamp 1679581782
transform 1 0 6624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_70
timestamp 1679581782
transform 1 0 7296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_77
timestamp 1679581782
transform 1 0 7968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_84
timestamp 1679581782
transform 1 0 8640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_91
timestamp 1679581782
transform 1 0 9312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_98
timestamp 1679581782
transform 1 0 9984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_105
timestamp 1679581782
transform 1 0 10656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_112
timestamp 1679581782
transform 1 0 11328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_119
timestamp 1679581782
transform 1 0 12000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_126
timestamp 1679581782
transform 1 0 12672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_133
timestamp 1679581782
transform 1 0 13344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_140
timestamp 1679581782
transform 1 0 14016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_147
timestamp 1679581782
transform 1 0 14688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_154
timestamp 1679581782
transform 1 0 15360 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_161
timestamp 1679581782
transform 1 0 16032 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_168
timestamp 1679581782
transform 1 0 16704 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_175
timestamp 1679581782
transform 1 0 17376 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_182
timestamp 1679581782
transform 1 0 18048 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_189
timestamp 1679581782
transform 1 0 18720 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_196
timestamp 1679581782
transform 1 0 19392 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_203
timestamp 1679581782
transform 1 0 20064 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_210
timestamp 1679581782
transform 1 0 20736 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_217
timestamp 1679581782
transform 1 0 21408 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_224
timestamp 1679581782
transform 1 0 22080 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_231
timestamp 1679581782
transform 1 0 22752 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_238
timestamp 1679581782
transform 1 0 23424 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_245
timestamp 1679581782
transform 1 0 24096 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_252
timestamp 1679581782
transform 1 0 24768 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_259
timestamp 1679581782
transform 1 0 25440 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_266
timestamp 1679581782
transform 1 0 26112 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_273
timestamp 1679581782
transform 1 0 26784 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_280
timestamp 1679581782
transform 1 0 27456 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_287
timestamp 1679581782
transform 1 0 28128 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_294
timestamp 1679581782
transform 1 0 28800 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_301
timestamp 1679581782
transform 1 0 29472 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_308
timestamp 1679581782
transform 1 0 30144 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_315
timestamp 1679581782
transform 1 0 30816 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_322
timestamp 1679581782
transform 1 0 31488 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_329
timestamp 1679581782
transform 1 0 32160 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_336
timestamp 1679581782
transform 1 0 32832 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_343
timestamp 1679581782
transform 1 0 33504 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_350
timestamp 1679581782
transform 1 0 34176 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_357
timestamp 1679581782
transform 1 0 34848 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_364
timestamp 1679581782
transform 1 0 35520 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_371
timestamp 1679581782
transform 1 0 36192 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_378
timestamp 1679581782
transform 1 0 36864 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_385
timestamp 1679581782
transform 1 0 37536 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_392
timestamp 1679581782
transform 1 0 38208 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_399
timestamp 1679581782
transform 1 0 38880 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_406
timestamp 1679581782
transform 1 0 39552 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_413
timestamp 1679581782
transform 1 0 40224 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_420
timestamp 1679581782
transform 1 0 40896 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_427
timestamp 1679581782
transform 1 0 41568 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_434
timestamp 1679581782
transform 1 0 42240 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_441
timestamp 1679581782
transform 1 0 42912 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_448
timestamp 1679581782
transform 1 0 43584 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_455
timestamp 1679581782
transform 1 0 44256 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_462
timestamp 1679581782
transform 1 0 44928 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_469
timestamp 1679581782
transform 1 0 45600 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_476
timestamp 1679581782
transform 1 0 46272 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_483
timestamp 1679581782
transform 1 0 46944 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_490
timestamp 1679581782
transform 1 0 47616 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_497
timestamp 1679581782
transform 1 0 48288 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_504
timestamp 1679581782
transform 1 0 48960 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_511
timestamp 1679581782
transform 1 0 49632 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_518
timestamp 1679581782
transform 1 0 50304 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_525
timestamp 1679581782
transform 1 0 50976 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_532
timestamp 1679581782
transform 1 0 51648 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_539
timestamp 1679581782
transform 1 0 52320 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_546
timestamp 1679581782
transform 1 0 52992 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_553
timestamp 1679581782
transform 1 0 53664 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_560
timestamp 1679581782
transform 1 0 54336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_567
timestamp 1679581782
transform 1 0 55008 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_574
timestamp 1679581782
transform 1 0 55680 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_581
timestamp 1679581782
transform 1 0 56352 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_588
timestamp 1679581782
transform 1 0 57024 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_595
timestamp 1679581782
transform 1 0 57696 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_602
timestamp 1679581782
transform 1 0 58368 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_609
timestamp 1679581782
transform 1 0 59040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_616
timestamp 1679581782
transform 1 0 59712 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_623
timestamp 1679581782
transform 1 0 60384 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_630
timestamp 1679581782
transform 1 0 61056 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_637
timestamp 1679581782
transform 1 0 61728 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_644
timestamp 1679581782
transform 1 0 62400 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_651
timestamp 1679581782
transform 1 0 63072 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_658
timestamp 1679581782
transform 1 0 63744 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_665
timestamp 1679581782
transform 1 0 64416 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_672
timestamp 1679581782
transform 1 0 65088 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_679
timestamp 1679581782
transform 1 0 65760 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_686
timestamp 1679581782
transform 1 0 66432 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_693
timestamp 1679581782
transform 1 0 67104 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_700
timestamp 1679581782
transform 1 0 67776 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_707
timestamp 1679581782
transform 1 0 68448 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_714
timestamp 1679581782
transform 1 0 69120 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_721
timestamp 1679581782
transform 1 0 69792 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_728
timestamp 1679581782
transform 1 0 70464 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_735
timestamp 1679581782
transform 1 0 71136 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_742
timestamp 1679581782
transform 1 0 71808 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_749
timestamp 1679581782
transform 1 0 72480 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_756
timestamp 1679581782
transform 1 0 73152 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_763
timestamp 1679581782
transform 1 0 73824 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_770
timestamp 1679581782
transform 1 0 74496 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_777
timestamp 1679581782
transform 1 0 75168 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_784
timestamp 1679581782
transform 1 0 75840 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_791
timestamp 1679581782
transform 1 0 76512 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_798
timestamp 1679581782
transform 1 0 77184 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_805
timestamp 1679581782
transform 1 0 77856 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_812
timestamp 1679581782
transform 1 0 78528 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_819
timestamp 1679581782
transform 1 0 79200 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_826
timestamp 1679581782
transform 1 0 79872 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_833
timestamp 1679581782
transform 1 0 80544 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_840
timestamp 1679581782
transform 1 0 81216 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_847
timestamp 1679581782
transform 1 0 81888 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_854
timestamp 1679581782
transform 1 0 82560 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_861
timestamp 1679581782
transform 1 0 83232 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_868
timestamp 1679581782
transform 1 0 83904 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_875
timestamp 1679581782
transform 1 0 84576 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_882
timestamp 1679581782
transform 1 0 85248 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_889
timestamp 1679581782
transform 1 0 85920 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_896
timestamp 1679581782
transform 1 0 86592 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_903
timestamp 1679581782
transform 1 0 87264 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_910
timestamp 1679581782
transform 1 0 87936 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_917
timestamp 1679581782
transform 1 0 88608 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_924
timestamp 1679581782
transform 1 0 89280 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_931
timestamp 1679581782
transform 1 0 89952 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_938
timestamp 1679581782
transform 1 0 90624 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_945
timestamp 1679581782
transform 1 0 91296 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_952
timestamp 1679581782
transform 1 0 91968 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_959
timestamp 1679581782
transform 1 0 92640 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_966
timestamp 1679581782
transform 1 0 93312 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_973
timestamp 1679581782
transform 1 0 93984 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_980
timestamp 1679581782
transform 1 0 94656 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_987
timestamp 1679581782
transform 1 0 95328 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_994
timestamp 1679581782
transform 1 0 96000 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1001
timestamp 1679581782
transform 1 0 96672 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1008
timestamp 1679581782
transform 1 0 97344 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1015
timestamp 1679581782
transform 1 0 98016 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_1022
timestamp 1679581782
transform 1 0 98688 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_4
timestamp 1679581782
transform 1 0 960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_11
timestamp 1679581782
transform 1 0 1632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_18
timestamp 1679581782
transform 1 0 2304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_25
timestamp 1679581782
transform 1 0 2976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_32
timestamp 1679581782
transform 1 0 3648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_39
timestamp 1679581782
transform 1 0 4320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_46
timestamp 1679581782
transform 1 0 4992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_53
timestamp 1679581782
transform 1 0 5664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_60
timestamp 1679581782
transform 1 0 6336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_67
timestamp 1679581782
transform 1 0 7008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_74
timestamp 1679581782
transform 1 0 7680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_81
timestamp 1679581782
transform 1 0 8352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_88
timestamp 1679581782
transform 1 0 9024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_95
timestamp 1679581782
transform 1 0 9696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_102
timestamp 1679581782
transform 1 0 10368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_109
timestamp 1679581782
transform 1 0 11040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_116
timestamp 1679581782
transform 1 0 11712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_123
timestamp 1679581782
transform 1 0 12384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_130
timestamp 1679581782
transform 1 0 13056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_137
timestamp 1679581782
transform 1 0 13728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_144
timestamp 1679581782
transform 1 0 14400 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_151
timestamp 1679581782
transform 1 0 15072 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_158
timestamp 1679581782
transform 1 0 15744 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_165
timestamp 1679581782
transform 1 0 16416 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_172
timestamp 1679581782
transform 1 0 17088 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_179
timestamp 1679581782
transform 1 0 17760 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_186
timestamp 1679581782
transform 1 0 18432 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_193
timestamp 1679581782
transform 1 0 19104 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_200
timestamp 1679581782
transform 1 0 19776 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_207
timestamp 1679581782
transform 1 0 20448 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_214
timestamp 1679581782
transform 1 0 21120 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_221
timestamp 1679581782
transform 1 0 21792 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_228
timestamp 1679581782
transform 1 0 22464 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_235
timestamp 1679581782
transform 1 0 23136 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_242
timestamp 1679581782
transform 1 0 23808 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_249
timestamp 1679581782
transform 1 0 24480 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_256
timestamp 1679581782
transform 1 0 25152 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_263
timestamp 1679581782
transform 1 0 25824 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_270
timestamp 1679581782
transform 1 0 26496 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_277
timestamp 1679581782
transform 1 0 27168 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_284
timestamp 1679581782
transform 1 0 27840 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_291
timestamp 1679581782
transform 1 0 28512 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_298
timestamp 1679581782
transform 1 0 29184 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_305
timestamp 1679581782
transform 1 0 29856 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_312
timestamp 1679581782
transform 1 0 30528 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_319
timestamp 1679581782
transform 1 0 31200 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_326
timestamp 1679581782
transform 1 0 31872 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_333
timestamp 1679581782
transform 1 0 32544 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_340
timestamp 1679581782
transform 1 0 33216 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_347
timestamp 1679581782
transform 1 0 33888 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_354
timestamp 1679581782
transform 1 0 34560 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_361
timestamp 1679581782
transform 1 0 35232 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_368
timestamp 1679581782
transform 1 0 35904 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_375
timestamp 1679581782
transform 1 0 36576 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_382
timestamp 1679581782
transform 1 0 37248 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_389
timestamp 1679581782
transform 1 0 37920 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_396
timestamp 1679581782
transform 1 0 38592 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_403
timestamp 1679581782
transform 1 0 39264 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_410
timestamp 1679581782
transform 1 0 39936 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_417
timestamp 1679581782
transform 1 0 40608 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_424
timestamp 1679581782
transform 1 0 41280 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_431
timestamp 1679581782
transform 1 0 41952 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_438
timestamp 1679581782
transform 1 0 42624 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_445
timestamp 1679581782
transform 1 0 43296 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_452
timestamp 1679581782
transform 1 0 43968 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_459
timestamp 1679581782
transform 1 0 44640 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_466
timestamp 1679581782
transform 1 0 45312 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_473
timestamp 1679581782
transform 1 0 45984 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_480
timestamp 1679581782
transform 1 0 46656 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_487
timestamp 1679581782
transform 1 0 47328 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_494
timestamp 1679581782
transform 1 0 48000 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_501
timestamp 1679581782
transform 1 0 48672 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_508
timestamp 1679581782
transform 1 0 49344 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_515
timestamp 1679581782
transform 1 0 50016 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_522
timestamp 1679581782
transform 1 0 50688 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_529
timestamp 1679581782
transform 1 0 51360 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_536
timestamp 1679581782
transform 1 0 52032 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_543
timestamp 1679581782
transform 1 0 52704 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_550
timestamp 1679581782
transform 1 0 53376 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_557
timestamp 1679581782
transform 1 0 54048 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_564
timestamp 1679581782
transform 1 0 54720 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_571
timestamp 1679581782
transform 1 0 55392 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_578
timestamp 1679581782
transform 1 0 56064 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_585
timestamp 1679581782
transform 1 0 56736 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_592
timestamp 1679581782
transform 1 0 57408 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_599
timestamp 1679581782
transform 1 0 58080 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_606
timestamp 1679581782
transform 1 0 58752 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_613
timestamp 1679581782
transform 1 0 59424 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_620
timestamp 1679581782
transform 1 0 60096 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_627
timestamp 1679581782
transform 1 0 60768 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_634
timestamp 1679581782
transform 1 0 61440 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_641
timestamp 1679581782
transform 1 0 62112 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_648
timestamp 1679581782
transform 1 0 62784 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_655
timestamp 1679581782
transform 1 0 63456 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_662
timestamp 1679581782
transform 1 0 64128 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_669
timestamp 1679581782
transform 1 0 64800 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_676
timestamp 1679581782
transform 1 0 65472 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_683
timestamp 1679581782
transform 1 0 66144 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_690
timestamp 1679581782
transform 1 0 66816 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_697
timestamp 1679581782
transform 1 0 67488 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_704
timestamp 1679581782
transform 1 0 68160 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_711
timestamp 1679581782
transform 1 0 68832 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_718
timestamp 1679581782
transform 1 0 69504 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_725
timestamp 1679581782
transform 1 0 70176 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_732
timestamp 1679581782
transform 1 0 70848 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_739
timestamp 1679581782
transform 1 0 71520 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_746
timestamp 1679581782
transform 1 0 72192 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_753
timestamp 1679581782
transform 1 0 72864 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_760
timestamp 1679581782
transform 1 0 73536 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_767
timestamp 1679581782
transform 1 0 74208 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_774
timestamp 1679581782
transform 1 0 74880 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_781
timestamp 1679581782
transform 1 0 75552 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_788
timestamp 1679581782
transform 1 0 76224 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_795
timestamp 1679581782
transform 1 0 76896 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_802
timestamp 1679581782
transform 1 0 77568 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_809
timestamp 1679581782
transform 1 0 78240 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_816
timestamp 1679581782
transform 1 0 78912 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_823
timestamp 1679581782
transform 1 0 79584 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_830
timestamp 1679581782
transform 1 0 80256 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_837
timestamp 1679581782
transform 1 0 80928 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_844
timestamp 1679581782
transform 1 0 81600 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_851
timestamp 1679581782
transform 1 0 82272 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_858
timestamp 1679581782
transform 1 0 82944 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_865
timestamp 1679581782
transform 1 0 83616 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_872
timestamp 1679581782
transform 1 0 84288 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_879
timestamp 1679581782
transform 1 0 84960 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_886
timestamp 1679581782
transform 1 0 85632 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_893
timestamp 1679581782
transform 1 0 86304 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_900
timestamp 1679581782
transform 1 0 86976 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_907
timestamp 1679581782
transform 1 0 87648 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_914
timestamp 1679581782
transform 1 0 88320 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_921
timestamp 1679581782
transform 1 0 88992 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_928
timestamp 1679581782
transform 1 0 89664 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_935
timestamp 1679581782
transform 1 0 90336 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_942
timestamp 1679581782
transform 1 0 91008 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_949
timestamp 1679581782
transform 1 0 91680 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_956
timestamp 1679581782
transform 1 0 92352 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_963
timestamp 1679581782
transform 1 0 93024 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_970
timestamp 1679581782
transform 1 0 93696 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_977
timestamp 1679581782
transform 1 0 94368 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_984
timestamp 1679581782
transform 1 0 95040 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_991
timestamp 1679581782
transform 1 0 95712 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_998
timestamp 1679581782
transform 1 0 96384 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1005
timestamp 1679581782
transform 1 0 97056 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1012
timestamp 1679581782
transform 1 0 97728 0 1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_1019
timestamp 1679581782
transform 1 0 98400 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_1026
timestamp 1677580104
transform 1 0 99072 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_1028
timestamp 1677579658
transform 1 0 99264 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_5
timestamp 1679581782
transform 1 0 1056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_12
timestamp 1679581782
transform 1 0 1728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_19
timestamp 1679581782
transform 1 0 2400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_26
timestamp 1679581782
transform 1 0 3072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_33
timestamp 1679581782
transform 1 0 3744 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_40
timestamp 1679581782
transform 1 0 4416 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_47
timestamp 1679581782
transform 1 0 5088 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_54
timestamp 1679581782
transform 1 0 5760 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_61
timestamp 1679581782
transform 1 0 6432 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_68
timestamp 1679581782
transform 1 0 7104 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_75
timestamp 1679581782
transform 1 0 7776 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_82
timestamp 1679581782
transform 1 0 8448 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_89
timestamp 1679581782
transform 1 0 9120 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_96
timestamp 1679581782
transform 1 0 9792 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_103
timestamp 1679581782
transform 1 0 10464 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_110
timestamp 1679581782
transform 1 0 11136 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_117
timestamp 1679581782
transform 1 0 11808 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_124
timestamp 1679581782
transform 1 0 12480 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_131
timestamp 1679581782
transform 1 0 13152 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_138
timestamp 1679581782
transform 1 0 13824 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_145
timestamp 1679581782
transform 1 0 14496 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_152
timestamp 1679581782
transform 1 0 15168 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_159
timestamp 1679581782
transform 1 0 15840 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_166
timestamp 1679581782
transform 1 0 16512 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_173
timestamp 1679581782
transform 1 0 17184 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_180
timestamp 1679581782
transform 1 0 17856 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_187
timestamp 1679581782
transform 1 0 18528 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_194
timestamp 1679581782
transform 1 0 19200 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_201
timestamp 1679581782
transform 1 0 19872 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_208
timestamp 1679581782
transform 1 0 20544 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_215
timestamp 1679581782
transform 1 0 21216 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_222
timestamp 1679581782
transform 1 0 21888 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_229
timestamp 1679581782
transform 1 0 22560 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_236
timestamp 1679581782
transform 1 0 23232 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_243
timestamp 1679581782
transform 1 0 23904 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_250
timestamp 1679581782
transform 1 0 24576 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_257
timestamp 1679581782
transform 1 0 25248 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_264
timestamp 1679581782
transform 1 0 25920 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_271
timestamp 1679581782
transform 1 0 26592 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_278
timestamp 1679581782
transform 1 0 27264 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_285
timestamp 1679581782
transform 1 0 27936 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_292
timestamp 1679581782
transform 1 0 28608 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_299
timestamp 1679581782
transform 1 0 29280 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_306
timestamp 1679581782
transform 1 0 29952 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_313
timestamp 1679581782
transform 1 0 30624 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_320
timestamp 1679581782
transform 1 0 31296 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_327
timestamp 1679581782
transform 1 0 31968 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_334
timestamp 1679581782
transform 1 0 32640 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_341
timestamp 1679581782
transform 1 0 33312 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_348
timestamp 1679581782
transform 1 0 33984 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_355
timestamp 1679581782
transform 1 0 34656 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_362
timestamp 1679581782
transform 1 0 35328 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_369
timestamp 1679581782
transform 1 0 36000 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_376
timestamp 1679581782
transform 1 0 36672 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_383
timestamp 1679581782
transform 1 0 37344 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_390
timestamp 1679581782
transform 1 0 38016 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_397
timestamp 1679581782
transform 1 0 38688 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_404
timestamp 1679581782
transform 1 0 39360 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_411
timestamp 1679581782
transform 1 0 40032 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_418
timestamp 1679581782
transform 1 0 40704 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_425
timestamp 1679581782
transform 1 0 41376 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_432
timestamp 1679581782
transform 1 0 42048 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_439
timestamp 1679581782
transform 1 0 42720 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_446
timestamp 1679581782
transform 1 0 43392 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_453
timestamp 1679581782
transform 1 0 44064 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_460
timestamp 1679581782
transform 1 0 44736 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_467
timestamp 1679581782
transform 1 0 45408 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_474
timestamp 1679581782
transform 1 0 46080 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_481
timestamp 1679581782
transform 1 0 46752 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_488
timestamp 1679581782
transform 1 0 47424 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_495
timestamp 1679581782
transform 1 0 48096 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_502
timestamp 1679581782
transform 1 0 48768 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_509
timestamp 1679581782
transform 1 0 49440 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_516
timestamp 1679581782
transform 1 0 50112 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_523
timestamp 1679581782
transform 1 0 50784 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_530
timestamp 1679581782
transform 1 0 51456 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_537
timestamp 1679581782
transform 1 0 52128 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_544
timestamp 1679581782
transform 1 0 52800 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_551
timestamp 1679581782
transform 1 0 53472 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_558
timestamp 1679581782
transform 1 0 54144 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_565
timestamp 1679581782
transform 1 0 54816 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_572
timestamp 1679581782
transform 1 0 55488 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_579
timestamp 1679581782
transform 1 0 56160 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_586
timestamp 1679581782
transform 1 0 56832 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_593
timestamp 1679581782
transform 1 0 57504 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_600
timestamp 1679581782
transform 1 0 58176 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_607
timestamp 1679581782
transform 1 0 58848 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_614
timestamp 1679581782
transform 1 0 59520 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_621
timestamp 1679581782
transform 1 0 60192 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_628
timestamp 1679581782
transform 1 0 60864 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_635
timestamp 1679581782
transform 1 0 61536 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_642
timestamp 1679581782
transform 1 0 62208 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_649
timestamp 1679581782
transform 1 0 62880 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_656
timestamp 1679581782
transform 1 0 63552 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_663
timestamp 1679581782
transform 1 0 64224 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_670
timestamp 1679581782
transform 1 0 64896 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_677
timestamp 1679581782
transform 1 0 65568 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_684
timestamp 1679581782
transform 1 0 66240 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_691
timestamp 1679581782
transform 1 0 66912 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_698
timestamp 1679581782
transform 1 0 67584 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_705
timestamp 1679581782
transform 1 0 68256 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_712
timestamp 1679581782
transform 1 0 68928 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_719
timestamp 1679581782
transform 1 0 69600 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_726
timestamp 1679581782
transform 1 0 70272 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_733
timestamp 1679581782
transform 1 0 70944 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_740
timestamp 1679581782
transform 1 0 71616 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_747
timestamp 1679581782
transform 1 0 72288 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_754
timestamp 1679581782
transform 1 0 72960 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_761
timestamp 1679581782
transform 1 0 73632 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_768
timestamp 1679581782
transform 1 0 74304 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_775
timestamp 1679581782
transform 1 0 74976 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_782
timestamp 1679581782
transform 1 0 75648 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_789
timestamp 1679581782
transform 1 0 76320 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_796
timestamp 1679581782
transform 1 0 76992 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_803
timestamp 1679581782
transform 1 0 77664 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_810
timestamp 1679581782
transform 1 0 78336 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_817
timestamp 1679581782
transform 1 0 79008 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_824
timestamp 1679581782
transform 1 0 79680 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_831
timestamp 1679581782
transform 1 0 80352 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_838
timestamp 1679581782
transform 1 0 81024 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_845
timestamp 1679581782
transform 1 0 81696 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_852
timestamp 1679581782
transform 1 0 82368 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_859
timestamp 1679581782
transform 1 0 83040 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_866
timestamp 1679581782
transform 1 0 83712 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_873
timestamp 1679581782
transform 1 0 84384 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_880
timestamp 1679581782
transform 1 0 85056 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_887
timestamp 1679581782
transform 1 0 85728 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_894
timestamp 1679581782
transform 1 0 86400 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_901
timestamp 1679581782
transform 1 0 87072 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_908
timestamp 1679581782
transform 1 0 87744 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_915
timestamp 1679581782
transform 1 0 88416 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_922
timestamp 1679581782
transform 1 0 89088 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_929
timestamp 1679581782
transform 1 0 89760 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_936
timestamp 1679581782
transform 1 0 90432 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_943
timestamp 1679581782
transform 1 0 91104 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_950
timestamp 1679581782
transform 1 0 91776 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_957
timestamp 1679581782
transform 1 0 92448 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_964
timestamp 1679581782
transform 1 0 93120 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_971
timestamp 1679581782
transform 1 0 93792 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_978
timestamp 1679581782
transform 1 0 94464 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_985
timestamp 1679581782
transform 1 0 95136 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_992
timestamp 1679581782
transform 1 0 95808 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_999
timestamp 1679581782
transform 1 0 96480 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1006
timestamp 1679581782
transform 1 0 97152 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1013
timestamp 1679581782
transform 1 0 97824 0 -1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_1020
timestamp 1679581782
transform 1 0 98496 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_1027
timestamp 1677580104
transform 1 0 99168 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_5
timestamp 1679581782
transform 1 0 1056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_12
timestamp 1679581782
transform 1 0 1728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_19
timestamp 1679581782
transform 1 0 2400 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_26
timestamp 1679581782
transform 1 0 3072 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_33
timestamp 1679581782
transform 1 0 3744 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_40
timestamp 1679581782
transform 1 0 4416 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_47
timestamp 1679581782
transform 1 0 5088 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_54
timestamp 1679581782
transform 1 0 5760 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_61
timestamp 1679581782
transform 1 0 6432 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_68
timestamp 1679581782
transform 1 0 7104 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_75
timestamp 1679581782
transform 1 0 7776 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_82
timestamp 1679581782
transform 1 0 8448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_89
timestamp 1679581782
transform 1 0 9120 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_96
timestamp 1679581782
transform 1 0 9792 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_103
timestamp 1679581782
transform 1 0 10464 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_110
timestamp 1679581782
transform 1 0 11136 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_117
timestamp 1679581782
transform 1 0 11808 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_124
timestamp 1679581782
transform 1 0 12480 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_131
timestamp 1679581782
transform 1 0 13152 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_138
timestamp 1679581782
transform 1 0 13824 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_145
timestamp 1679581782
transform 1 0 14496 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_152
timestamp 1679581782
transform 1 0 15168 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_159
timestamp 1679581782
transform 1 0 15840 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_166
timestamp 1679581782
transform 1 0 16512 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_173
timestamp 1679581782
transform 1 0 17184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_180
timestamp 1679581782
transform 1 0 17856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_187
timestamp 1679581782
transform 1 0 18528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_194
timestamp 1679581782
transform 1 0 19200 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_201
timestamp 1679581782
transform 1 0 19872 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_208
timestamp 1679581782
transform 1 0 20544 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_215
timestamp 1679581782
transform 1 0 21216 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_222
timestamp 1679581782
transform 1 0 21888 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_229
timestamp 1679581782
transform 1 0 22560 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_236
timestamp 1679581782
transform 1 0 23232 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_243
timestamp 1679581782
transform 1 0 23904 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_250
timestamp 1679581782
transform 1 0 24576 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_257
timestamp 1679581782
transform 1 0 25248 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_264
timestamp 1679581782
transform 1 0 25920 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_271
timestamp 1679581782
transform 1 0 26592 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_278
timestamp 1679581782
transform 1 0 27264 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_285
timestamp 1679581782
transform 1 0 27936 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_292
timestamp 1679581782
transform 1 0 28608 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_299
timestamp 1679581782
transform 1 0 29280 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_306
timestamp 1679581782
transform 1 0 29952 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_313
timestamp 1679581782
transform 1 0 30624 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_320
timestamp 1679581782
transform 1 0 31296 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_327
timestamp 1679581782
transform 1 0 31968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_334
timestamp 1679581782
transform 1 0 32640 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_341
timestamp 1679581782
transform 1 0 33312 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_348
timestamp 1679581782
transform 1 0 33984 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_355
timestamp 1679581782
transform 1 0 34656 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_362
timestamp 1679581782
transform 1 0 35328 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_369
timestamp 1679581782
transform 1 0 36000 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_376
timestamp 1679581782
transform 1 0 36672 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_383
timestamp 1679581782
transform 1 0 37344 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_390
timestamp 1679581782
transform 1 0 38016 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_397
timestamp 1679581782
transform 1 0 38688 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_404
timestamp 1679581782
transform 1 0 39360 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_411
timestamp 1679581782
transform 1 0 40032 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_418
timestamp 1679581782
transform 1 0 40704 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_425
timestamp 1679581782
transform 1 0 41376 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_432
timestamp 1679581782
transform 1 0 42048 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_439
timestamp 1679581782
transform 1 0 42720 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_446
timestamp 1679581782
transform 1 0 43392 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_453
timestamp 1679581782
transform 1 0 44064 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_460
timestamp 1679581782
transform 1 0 44736 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_467
timestamp 1679581782
transform 1 0 45408 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_474
timestamp 1679581782
transform 1 0 46080 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_481
timestamp 1679581782
transform 1 0 46752 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_488
timestamp 1679581782
transform 1 0 47424 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_495
timestamp 1679581782
transform 1 0 48096 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_502
timestamp 1679581782
transform 1 0 48768 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_509
timestamp 1679581782
transform 1 0 49440 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_516
timestamp 1679581782
transform 1 0 50112 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_523
timestamp 1679581782
transform 1 0 50784 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_530
timestamp 1679581782
transform 1 0 51456 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_537
timestamp 1679581782
transform 1 0 52128 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_544
timestamp 1679581782
transform 1 0 52800 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_551
timestamp 1679581782
transform 1 0 53472 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_558
timestamp 1679581782
transform 1 0 54144 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_565
timestamp 1679581782
transform 1 0 54816 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_572
timestamp 1679581782
transform 1 0 55488 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_579
timestamp 1679581782
transform 1 0 56160 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_586
timestamp 1679581782
transform 1 0 56832 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_593
timestamp 1679581782
transform 1 0 57504 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_600
timestamp 1679581782
transform 1 0 58176 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_607
timestamp 1679581782
transform 1 0 58848 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_614
timestamp 1679581782
transform 1 0 59520 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_621
timestamp 1679581782
transform 1 0 60192 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_628
timestamp 1679581782
transform 1 0 60864 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_635
timestamp 1679581782
transform 1 0 61536 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_642
timestamp 1679581782
transform 1 0 62208 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_649
timestamp 1679581782
transform 1 0 62880 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_656
timestamp 1679581782
transform 1 0 63552 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_663
timestamp 1679581782
transform 1 0 64224 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_670
timestamp 1679581782
transform 1 0 64896 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_677
timestamp 1679581782
transform 1 0 65568 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_684
timestamp 1679581782
transform 1 0 66240 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_691
timestamp 1679581782
transform 1 0 66912 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_698
timestamp 1679581782
transform 1 0 67584 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_705
timestamp 1679581782
transform 1 0 68256 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_712
timestamp 1679581782
transform 1 0 68928 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_719
timestamp 1679581782
transform 1 0 69600 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_726
timestamp 1679581782
transform 1 0 70272 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_733
timestamp 1679581782
transform 1 0 70944 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_740
timestamp 1679581782
transform 1 0 71616 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_747
timestamp 1679581782
transform 1 0 72288 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_754
timestamp 1679581782
transform 1 0 72960 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_761
timestamp 1679581782
transform 1 0 73632 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_768
timestamp 1679581782
transform 1 0 74304 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_775
timestamp 1679581782
transform 1 0 74976 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_782
timestamp 1679581782
transform 1 0 75648 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_789
timestamp 1679581782
transform 1 0 76320 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_796
timestamp 1679581782
transform 1 0 76992 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_803
timestamp 1679581782
transform 1 0 77664 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_810
timestamp 1679581782
transform 1 0 78336 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_817
timestamp 1679581782
transform 1 0 79008 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_824
timestamp 1679577901
transform 1 0 79680 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_832
timestamp 1679581782
transform 1 0 80448 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_839
timestamp 1679577901
transform 1 0 81120 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_843
timestamp 1677579658
transform 1 0 81504 0 1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_848
timestamp 1679577901
transform 1 0 81984 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_856
timestamp 1679581782
transform 1 0 82752 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_863
timestamp 1679581782
transform 1 0 83424 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_870
timestamp 1679581782
transform 1 0 84096 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_877
timestamp 1677579658
transform 1 0 84768 0 1 23436
box -48 -56 144 834
use sg13g2_decap_4  FILLER_30_882
timestamp 1679577901
transform 1 0 85248 0 1 23436
box -48 -56 432 834
use sg13g2_decap_4  FILLER_30_890
timestamp 1679577901
transform 1 0 86016 0 1 23436
box -48 -56 432 834
use sg13g2_decap_8  FILLER_30_898
timestamp 1679581782
transform 1 0 86784 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_905
timestamp 1677580104
transform 1 0 87456 0 1 23436
box -48 -56 240 834
use sg13g2_decap_8  FILLER_30_911
timestamp 1679581782
transform 1 0 88032 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_918
timestamp 1677579658
transform 1 0 88704 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_923
timestamp 1679581782
transform 1 0 89184 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_930
timestamp 1679581782
transform 1 0 89856 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_937
timestamp 1679581782
transform 1 0 90528 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_948
timestamp 1679581782
transform 1 0 91584 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_958
timestamp 1679581782
transform 1 0 92544 0 1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_965
timestamp 1677579658
transform 1 0 93216 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_970
timestamp 1679581782
transform 1 0 93696 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_977
timestamp 1679581782
transform 1 0 94368 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_984
timestamp 1679581782
transform 1 0 95040 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_991
timestamp 1679581782
transform 1 0 95712 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_998
timestamp 1679581782
transform 1 0 96384 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1005
timestamp 1679581782
transform 1 0 97056 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1012
timestamp 1679581782
transform 1 0 97728 0 1 23436
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_1019
timestamp 1679581782
transform 1 0 98400 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_1026
timestamp 1677580104
transform 1 0 99072 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_1028
timestamp 1677579658
transform 1 0 99264 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_5
timestamp 1679581782
transform 1 0 1056 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_12
timestamp 1679581782
transform 1 0 1728 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_19
timestamp 1679581782
transform 1 0 2400 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_26
timestamp 1679581782
transform 1 0 3072 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_33
timestamp 1679581782
transform 1 0 3744 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_40
timestamp 1679581782
transform 1 0 4416 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_47
timestamp 1679581782
transform 1 0 5088 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_54
timestamp 1679581782
transform 1 0 5760 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_61
timestamp 1679581782
transform 1 0 6432 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_68
timestamp 1679581782
transform 1 0 7104 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_75
timestamp 1679581782
transform 1 0 7776 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_82
timestamp 1679581782
transform 1 0 8448 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_89
timestamp 1679581782
transform 1 0 9120 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_96
timestamp 1679581782
transform 1 0 9792 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_103
timestamp 1679581782
transform 1 0 10464 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_110
timestamp 1679581782
transform 1 0 11136 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_117
timestamp 1679581782
transform 1 0 11808 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_124
timestamp 1679581782
transform 1 0 12480 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_131
timestamp 1679581782
transform 1 0 13152 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_138
timestamp 1679581782
transform 1 0 13824 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_145
timestamp 1679581782
transform 1 0 14496 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_152
timestamp 1679581782
transform 1 0 15168 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_159
timestamp 1679581782
transform 1 0 15840 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_166
timestamp 1679581782
transform 1 0 16512 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_173
timestamp 1679581782
transform 1 0 17184 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_180
timestamp 1679581782
transform 1 0 17856 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_187
timestamp 1679581782
transform 1 0 18528 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_194
timestamp 1679581782
transform 1 0 19200 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_201
timestamp 1679581782
transform 1 0 19872 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_208
timestamp 1679581782
transform 1 0 20544 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_215
timestamp 1679581782
transform 1 0 21216 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_222
timestamp 1679581782
transform 1 0 21888 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_229
timestamp 1679581782
transform 1 0 22560 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_236
timestamp 1679581782
transform 1 0 23232 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_243
timestamp 1679581782
transform 1 0 23904 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_250
timestamp 1679581782
transform 1 0 24576 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_257
timestamp 1679581782
transform 1 0 25248 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_264
timestamp 1679581782
transform 1 0 25920 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_271
timestamp 1679581782
transform 1 0 26592 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_278
timestamp 1679581782
transform 1 0 27264 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_285
timestamp 1679581782
transform 1 0 27936 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_292
timestamp 1679581782
transform 1 0 28608 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_299
timestamp 1679581782
transform 1 0 29280 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_306
timestamp 1679581782
transform 1 0 29952 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_313
timestamp 1679581782
transform 1 0 30624 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_320
timestamp 1679581782
transform 1 0 31296 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_327
timestamp 1679581782
transform 1 0 31968 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_334
timestamp 1679581782
transform 1 0 32640 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_341
timestamp 1679581782
transform 1 0 33312 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_348
timestamp 1679581782
transform 1 0 33984 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_355
timestamp 1679581782
transform 1 0 34656 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_362
timestamp 1679581782
transform 1 0 35328 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_369
timestamp 1679581782
transform 1 0 36000 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_376
timestamp 1679581782
transform 1 0 36672 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_383
timestamp 1679581782
transform 1 0 37344 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_390
timestamp 1679581782
transform 1 0 38016 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_397
timestamp 1679581782
transform 1 0 38688 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_404
timestamp 1679581782
transform 1 0 39360 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_411
timestamp 1679581782
transform 1 0 40032 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_418
timestamp 1679581782
transform 1 0 40704 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_425
timestamp 1679581782
transform 1 0 41376 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_432
timestamp 1679581782
transform 1 0 42048 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_439
timestamp 1679581782
transform 1 0 42720 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_446
timestamp 1679581782
transform 1 0 43392 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_453
timestamp 1679581782
transform 1 0 44064 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_460
timestamp 1679581782
transform 1 0 44736 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_467
timestamp 1679581782
transform 1 0 45408 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_474
timestamp 1679581782
transform 1 0 46080 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_481
timestamp 1679581782
transform 1 0 46752 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_488
timestamp 1679581782
transform 1 0 47424 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_495
timestamp 1679581782
transform 1 0 48096 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_502
timestamp 1679581782
transform 1 0 48768 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_509
timestamp 1679581782
transform 1 0 49440 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_516
timestamp 1679581782
transform 1 0 50112 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_523
timestamp 1679581782
transform 1 0 50784 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_530
timestamp 1679581782
transform 1 0 51456 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_537
timestamp 1679581782
transform 1 0 52128 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_544
timestamp 1679581782
transform 1 0 52800 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_551
timestamp 1679581782
transform 1 0 53472 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_558
timestamp 1679581782
transform 1 0 54144 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_565
timestamp 1679581782
transform 1 0 54816 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_572
timestamp 1679581782
transform 1 0 55488 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_579
timestamp 1679581782
transform 1 0 56160 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_586
timestamp 1679581782
transform 1 0 56832 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_593
timestamp 1679581782
transform 1 0 57504 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_600
timestamp 1679581782
transform 1 0 58176 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_607
timestamp 1679581782
transform 1 0 58848 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_614
timestamp 1679581782
transform 1 0 59520 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_621
timestamp 1679581782
transform 1 0 60192 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_628
timestamp 1679581782
transform 1 0 60864 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_635
timestamp 1679581782
transform 1 0 61536 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_642
timestamp 1679581782
transform 1 0 62208 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_649
timestamp 1679581782
transform 1 0 62880 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_656
timestamp 1679581782
transform 1 0 63552 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_663
timestamp 1679581782
transform 1 0 64224 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_670
timestamp 1679581782
transform 1 0 64896 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_677
timestamp 1679581782
transform 1 0 65568 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_684
timestamp 1679581782
transform 1 0 66240 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_691
timestamp 1679581782
transform 1 0 66912 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_698
timestamp 1679581782
transform 1 0 67584 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_705
timestamp 1679581782
transform 1 0 68256 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_712
timestamp 1679581782
transform 1 0 68928 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_719
timestamp 1679581782
transform 1 0 69600 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_726
timestamp 1679581782
transform 1 0 70272 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_733
timestamp 1679581782
transform 1 0 70944 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_740
timestamp 1679581782
transform 1 0 71616 0 -1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_747
timestamp 1679581782
transform 1 0 72288 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_754
timestamp 1677580104
transform 1 0 72960 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_770
timestamp 1677579658
transform 1 0 74496 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_775
timestamp 1677580104
transform 1 0 74976 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_784
timestamp 1677579658
transform 1 0 75840 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_793
timestamp 1677579658
transform 1 0 76704 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_855
timestamp 1677580104
transform 1 0 82656 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_881
timestamp 1677579658
transform 1 0 85152 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_31_886
timestamp 1679577901
transform 1 0 85632 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_894
timestamp 1677579658
transform 1 0 86400 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_910
timestamp 1677579658
transform 1 0 87936 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_927
timestamp 1677579658
transform 1 0 89568 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_940
timestamp 1677579658
transform 1 0 90816 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_945
timestamp 1677580104
transform 1 0 91296 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_947
timestamp 1677579658
transform 1 0 91488 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_952
timestamp 1677579658
transform 1 0 91968 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_969
timestamp 1677579658
transform 1 0 93600 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_986
timestamp 1677579658
transform 1 0 95232 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_1019
timestamp 1679581782
transform 1 0 98400 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_31_1026
timestamp 1677580104
transform 1 0 99072 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_1028
timestamp 1677579658
transform 1 0 99264 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_5
timestamp 1679581782
transform 1 0 1056 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_12
timestamp 1679581782
transform 1 0 1728 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_19
timestamp 1679581782
transform 1 0 2400 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_26
timestamp 1679581782
transform 1 0 3072 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_33
timestamp 1679581782
transform 1 0 3744 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_40
timestamp 1679581782
transform 1 0 4416 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_47
timestamp 1679581782
transform 1 0 5088 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_54
timestamp 1679581782
transform 1 0 5760 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_61
timestamp 1679581782
transform 1 0 6432 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_68
timestamp 1679581782
transform 1 0 7104 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_75
timestamp 1679581782
transform 1 0 7776 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_82
timestamp 1679581782
transform 1 0 8448 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_89
timestamp 1679581782
transform 1 0 9120 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_96
timestamp 1679581782
transform 1 0 9792 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_103
timestamp 1679581782
transform 1 0 10464 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_110
timestamp 1679581782
transform 1 0 11136 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_117
timestamp 1679581782
transform 1 0 11808 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_124
timestamp 1679581782
transform 1 0 12480 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_131
timestamp 1679581782
transform 1 0 13152 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_138
timestamp 1679581782
transform 1 0 13824 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_145
timestamp 1679581782
transform 1 0 14496 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_152
timestamp 1679581782
transform 1 0 15168 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_159
timestamp 1679581782
transform 1 0 15840 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_166
timestamp 1679581782
transform 1 0 16512 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_173
timestamp 1679581782
transform 1 0 17184 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_180
timestamp 1679581782
transform 1 0 17856 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_187
timestamp 1679581782
transform 1 0 18528 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_194
timestamp 1679581782
transform 1 0 19200 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_201
timestamp 1679581782
transform 1 0 19872 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_208
timestamp 1679581782
transform 1 0 20544 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_215
timestamp 1679581782
transform 1 0 21216 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_222
timestamp 1679581782
transform 1 0 21888 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_229
timestamp 1679581782
transform 1 0 22560 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_236
timestamp 1679581782
transform 1 0 23232 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_243
timestamp 1679581782
transform 1 0 23904 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_250
timestamp 1679581782
transform 1 0 24576 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_257
timestamp 1679581782
transform 1 0 25248 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_264
timestamp 1679581782
transform 1 0 25920 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_271
timestamp 1679581782
transform 1 0 26592 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_278
timestamp 1679581782
transform 1 0 27264 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_285
timestamp 1679581782
transform 1 0 27936 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_292
timestamp 1679581782
transform 1 0 28608 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_299
timestamp 1679581782
transform 1 0 29280 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_306
timestamp 1679581782
transform 1 0 29952 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_313
timestamp 1679581782
transform 1 0 30624 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_320
timestamp 1679581782
transform 1 0 31296 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_327
timestamp 1679581782
transform 1 0 31968 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_334
timestamp 1679581782
transform 1 0 32640 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_341
timestamp 1679581782
transform 1 0 33312 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_348
timestamp 1679581782
transform 1 0 33984 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_355
timestamp 1679581782
transform 1 0 34656 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_362
timestamp 1679581782
transform 1 0 35328 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_369
timestamp 1679581782
transform 1 0 36000 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_376
timestamp 1679581782
transform 1 0 36672 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_383
timestamp 1679581782
transform 1 0 37344 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_390
timestamp 1679581782
transform 1 0 38016 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_397
timestamp 1679581782
transform 1 0 38688 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_404
timestamp 1679581782
transform 1 0 39360 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_411
timestamp 1679581782
transform 1 0 40032 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_418
timestamp 1679581782
transform 1 0 40704 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_425
timestamp 1679581782
transform 1 0 41376 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_432
timestamp 1679581782
transform 1 0 42048 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_439
timestamp 1679581782
transform 1 0 42720 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_446
timestamp 1679581782
transform 1 0 43392 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_453
timestamp 1679581782
transform 1 0 44064 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_460
timestamp 1679581782
transform 1 0 44736 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_467
timestamp 1679581782
transform 1 0 45408 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_474
timestamp 1679581782
transform 1 0 46080 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_481
timestamp 1679581782
transform 1 0 46752 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_488
timestamp 1679581782
transform 1 0 47424 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_495
timestamp 1679581782
transform 1 0 48096 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_502
timestamp 1679581782
transform 1 0 48768 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_509
timestamp 1679581782
transform 1 0 49440 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_516
timestamp 1679581782
transform 1 0 50112 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_523
timestamp 1679581782
transform 1 0 50784 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_530
timestamp 1679581782
transform 1 0 51456 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_537
timestamp 1679581782
transform 1 0 52128 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_544
timestamp 1679581782
transform 1 0 52800 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_551
timestamp 1679581782
transform 1 0 53472 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_558
timestamp 1679581782
transform 1 0 54144 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_565
timestamp 1679581782
transform 1 0 54816 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_572
timestamp 1679581782
transform 1 0 55488 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_579
timestamp 1679581782
transform 1 0 56160 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_586
timestamp 1679581782
transform 1 0 56832 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_593
timestamp 1679581782
transform 1 0 57504 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_600
timestamp 1679581782
transform 1 0 58176 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_607
timestamp 1679581782
transform 1 0 58848 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_614
timestamp 1679581782
transform 1 0 59520 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_621
timestamp 1679581782
transform 1 0 60192 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_628
timestamp 1679581782
transform 1 0 60864 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_635
timestamp 1679581782
transform 1 0 61536 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_642
timestamp 1679581782
transform 1 0 62208 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_649
timestamp 1679581782
transform 1 0 62880 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_656
timestamp 1679581782
transform 1 0 63552 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_663
timestamp 1679581782
transform 1 0 64224 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_670
timestamp 1679581782
transform 1 0 64896 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_677
timestamp 1679581782
transform 1 0 65568 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_684
timestamp 1679581782
transform 1 0 66240 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_691
timestamp 1679581782
transform 1 0 66912 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_698
timestamp 1679581782
transform 1 0 67584 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_705
timestamp 1679581782
transform 1 0 68256 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_712
timestamp 1679581782
transform 1 0 68928 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_719
timestamp 1679581782
transform 1 0 69600 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_726
timestamp 1679581782
transform 1 0 70272 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_733
timestamp 1679581782
transform 1 0 70944 0 1 24948
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_740
timestamp 1679581782
transform 1 0 71616 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_747
timestamp 1677580104
transform 1 0 72288 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_749
timestamp 1677579658
transform 1 0 72480 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_761
timestamp 1677580104
transform 1 0 73632 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_779
timestamp 1677579658
transform 1 0 75360 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_799
timestamp 1677580104
transform 1 0 77280 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_820
timestamp 1677579658
transform 1 0 79296 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_833
timestamp 1677579658
transform 1 0 80544 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_837
timestamp 1677579658
transform 1 0 80928 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_841
timestamp 1677579658
transform 1 0 81312 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_845
timestamp 1677580104
transform 1 0 81696 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_853
timestamp 1677579658
transform 1 0 82464 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_857
timestamp 1677580104
transform 1 0 82848 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_862
timestamp 1677580104
transform 1 0 83328 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_883
timestamp 1677579658
transform 1 0 85344 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_887
timestamp 1677579658
transform 1 0 85728 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_891
timestamp 1677580104
transform 1 0 86112 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_920
timestamp 1677579658
transform 1 0 88896 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_924
timestamp 1677580104
transform 1 0 89280 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_942
timestamp 1677579658
transform 1 0 91008 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_949
timestamp 1677580104
transform 1 0 91680 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_954
timestamp 1677579658
transform 1 0 92160 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_966
timestamp 1677580104
transform 1 0 93312 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_971
timestamp 1677579658
transform 1 0 93792 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_978
timestamp 1677580104
transform 1 0 94464 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_980
timestamp 1677579658
transform 1 0 94656 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_984
timestamp 1677579658
transform 1 0 95040 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_988
timestamp 1677580104
transform 1 0 95424 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_1000
timestamp 1677579658
transform 1 0 96576 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_1004
timestamp 1677579658
transform 1 0 96960 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_32_1017
timestamp 1677579658
transform 1 0 98208 0 1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_1025
timestamp 1679577901
transform 1 0 98976 0 1 24948
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679581782
transform 1 0 576 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1679581782
transform 1 0 1248 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1679581782
transform 1 0 1920 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_21
timestamp 1679581782
transform 1 0 2592 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_28
timestamp 1679581782
transform 1 0 3264 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_35
timestamp 1679581782
transform 1 0 3936 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_42
timestamp 1679581782
transform 1 0 4608 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_49
timestamp 1679581782
transform 1 0 5280 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_56
timestamp 1679581782
transform 1 0 5952 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_63
timestamp 1679581782
transform 1 0 6624 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_70
timestamp 1679581782
transform 1 0 7296 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_77
timestamp 1679581782
transform 1 0 7968 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_84
timestamp 1679581782
transform 1 0 8640 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_91
timestamp 1679581782
transform 1 0 9312 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_98
timestamp 1679581782
transform 1 0 9984 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_105
timestamp 1679581782
transform 1 0 10656 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_112
timestamp 1679581782
transform 1 0 11328 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_119
timestamp 1679581782
transform 1 0 12000 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_126
timestamp 1679581782
transform 1 0 12672 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_133
timestamp 1679581782
transform 1 0 13344 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_140
timestamp 1679581782
transform 1 0 14016 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_147
timestamp 1679581782
transform 1 0 14688 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_154
timestamp 1679581782
transform 1 0 15360 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_161
timestamp 1679581782
transform 1 0 16032 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_168
timestamp 1679581782
transform 1 0 16704 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_175
timestamp 1679581782
transform 1 0 17376 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_182
timestamp 1679581782
transform 1 0 18048 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_189
timestamp 1679581782
transform 1 0 18720 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_196
timestamp 1679581782
transform 1 0 19392 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_203
timestamp 1679581782
transform 1 0 20064 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_210
timestamp 1679581782
transform 1 0 20736 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_217
timestamp 1679581782
transform 1 0 21408 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_224
timestamp 1679581782
transform 1 0 22080 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_231
timestamp 1679581782
transform 1 0 22752 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_238
timestamp 1679581782
transform 1 0 23424 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_245
timestamp 1679581782
transform 1 0 24096 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_252
timestamp 1679581782
transform 1 0 24768 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_259
timestamp 1679581782
transform 1 0 25440 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_266
timestamp 1679581782
transform 1 0 26112 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_273
timestamp 1679581782
transform 1 0 26784 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_280
timestamp 1679581782
transform 1 0 27456 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_287
timestamp 1679581782
transform 1 0 28128 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_294
timestamp 1679581782
transform 1 0 28800 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_301
timestamp 1679581782
transform 1 0 29472 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_308
timestamp 1679581782
transform 1 0 30144 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_315
timestamp 1679581782
transform 1 0 30816 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_322
timestamp 1679581782
transform 1 0 31488 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_329
timestamp 1679581782
transform 1 0 32160 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_336
timestamp 1679581782
transform 1 0 32832 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_343
timestamp 1679581782
transform 1 0 33504 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_350
timestamp 1679581782
transform 1 0 34176 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_357
timestamp 1679581782
transform 1 0 34848 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_364
timestamp 1679581782
transform 1 0 35520 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_371
timestamp 1679581782
transform 1 0 36192 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_378
timestamp 1679581782
transform 1 0 36864 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_385
timestamp 1679581782
transform 1 0 37536 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_392
timestamp 1679581782
transform 1 0 38208 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_399
timestamp 1679581782
transform 1 0 38880 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_406
timestamp 1679581782
transform 1 0 39552 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_413
timestamp 1679581782
transform 1 0 40224 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_420
timestamp 1679581782
transform 1 0 40896 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_427
timestamp 1679581782
transform 1 0 41568 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_434
timestamp 1679581782
transform 1 0 42240 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_441
timestamp 1679581782
transform 1 0 42912 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_448
timestamp 1679581782
transform 1 0 43584 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_455
timestamp 1679581782
transform 1 0 44256 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_462
timestamp 1679581782
transform 1 0 44928 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_469
timestamp 1679581782
transform 1 0 45600 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_476
timestamp 1679581782
transform 1 0 46272 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_483
timestamp 1679581782
transform 1 0 46944 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_490
timestamp 1679581782
transform 1 0 47616 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_497
timestamp 1679581782
transform 1 0 48288 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_504
timestamp 1679581782
transform 1 0 48960 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_511
timestamp 1679581782
transform 1 0 49632 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_518
timestamp 1679581782
transform 1 0 50304 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_525
timestamp 1679581782
transform 1 0 50976 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_532
timestamp 1679581782
transform 1 0 51648 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_539
timestamp 1679581782
transform 1 0 52320 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_546
timestamp 1679581782
transform 1 0 52992 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_553
timestamp 1679581782
transform 1 0 53664 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_560
timestamp 1679581782
transform 1 0 54336 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_567
timestamp 1679581782
transform 1 0 55008 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_574
timestamp 1679581782
transform 1 0 55680 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_581
timestamp 1679581782
transform 1 0 56352 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_588
timestamp 1679581782
transform 1 0 57024 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_595
timestamp 1679581782
transform 1 0 57696 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_602
timestamp 1679581782
transform 1 0 58368 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_609
timestamp 1679581782
transform 1 0 59040 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_616
timestamp 1679581782
transform 1 0 59712 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_623
timestamp 1679581782
transform 1 0 60384 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_630
timestamp 1679581782
transform 1 0 61056 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_637
timestamp 1679581782
transform 1 0 61728 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_644
timestamp 1679581782
transform 1 0 62400 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_651
timestamp 1679581782
transform 1 0 63072 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_658
timestamp 1679581782
transform 1 0 63744 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_665
timestamp 1679581782
transform 1 0 64416 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_672
timestamp 1679581782
transform 1 0 65088 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_679
timestamp 1679581782
transform 1 0 65760 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_686
timestamp 1679581782
transform 1 0 66432 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_693
timestamp 1679581782
transform 1 0 67104 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_700
timestamp 1679581782
transform 1 0 67776 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_707
timestamp 1679581782
transform 1 0 68448 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_714
timestamp 1679581782
transform 1 0 69120 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_721
timestamp 1679581782
transform 1 0 69792 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_33_728
timestamp 1679577901
transform 1 0 70464 0 -1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_33_735
timestamp 1677579658
transform 1 0 71136 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 576 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679581782
transform 1 0 1248 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679581782
transform 1 0 1920 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679581782
transform 1 0 2592 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679581782
transform 1 0 3264 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_35
timestamp 1679581782
transform 1 0 3936 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_42
timestamp 1679581782
transform 1 0 4608 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679581782
transform 1 0 5280 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_56
timestamp 1679581782
transform 1 0 5952 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_63
timestamp 1679581782
transform 1 0 6624 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_70
timestamp 1679581782
transform 1 0 7296 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_77
timestamp 1679581782
transform 1 0 7968 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_84
timestamp 1679581782
transform 1 0 8640 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_91
timestamp 1679581782
transform 1 0 9312 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_98
timestamp 1679581782
transform 1 0 9984 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_105
timestamp 1679581782
transform 1 0 10656 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_112
timestamp 1679581782
transform 1 0 11328 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_119
timestamp 1679581782
transform 1 0 12000 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_126
timestamp 1679581782
transform 1 0 12672 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_133
timestamp 1679581782
transform 1 0 13344 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_140
timestamp 1679581782
transform 1 0 14016 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_147
timestamp 1679581782
transform 1 0 14688 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_154
timestamp 1679581782
transform 1 0 15360 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_161
timestamp 1679581782
transform 1 0 16032 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_168
timestamp 1679581782
transform 1 0 16704 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_175
timestamp 1679581782
transform 1 0 17376 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_182
timestamp 1679581782
transform 1 0 18048 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_189
timestamp 1679581782
transform 1 0 18720 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_196
timestamp 1679581782
transform 1 0 19392 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_203
timestamp 1679581782
transform 1 0 20064 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_210
timestamp 1679581782
transform 1 0 20736 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_217
timestamp 1679581782
transform 1 0 21408 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_224
timestamp 1679581782
transform 1 0 22080 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_231
timestamp 1679581782
transform 1 0 22752 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_238
timestamp 1679581782
transform 1 0 23424 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_245
timestamp 1679581782
transform 1 0 24096 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_252
timestamp 1679581782
transform 1 0 24768 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_259
timestamp 1679581782
transform 1 0 25440 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_266
timestamp 1679581782
transform 1 0 26112 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_273
timestamp 1679581782
transform 1 0 26784 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_280
timestamp 1679581782
transform 1 0 27456 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_287
timestamp 1679581782
transform 1 0 28128 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_294
timestamp 1679581782
transform 1 0 28800 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_301
timestamp 1679581782
transform 1 0 29472 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_308
timestamp 1679581782
transform 1 0 30144 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_315
timestamp 1679581782
transform 1 0 30816 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_322
timestamp 1679581782
transform 1 0 31488 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_329
timestamp 1679581782
transform 1 0 32160 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_336
timestamp 1679581782
transform 1 0 32832 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_343
timestamp 1679581782
transform 1 0 33504 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_350
timestamp 1679581782
transform 1 0 34176 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_357
timestamp 1679581782
transform 1 0 34848 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_364
timestamp 1679581782
transform 1 0 35520 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_371
timestamp 1679581782
transform 1 0 36192 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_378
timestamp 1679581782
transform 1 0 36864 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_385
timestamp 1679581782
transform 1 0 37536 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_392
timestamp 1679581782
transform 1 0 38208 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_399
timestamp 1679581782
transform 1 0 38880 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_406
timestamp 1679581782
transform 1 0 39552 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_413
timestamp 1679581782
transform 1 0 40224 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_420
timestamp 1679581782
transform 1 0 40896 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_427
timestamp 1679581782
transform 1 0 41568 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_434
timestamp 1679581782
transform 1 0 42240 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_441
timestamp 1679581782
transform 1 0 42912 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_448
timestamp 1679581782
transform 1 0 43584 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_455
timestamp 1679581782
transform 1 0 44256 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_462
timestamp 1679581782
transform 1 0 44928 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_469
timestamp 1679581782
transform 1 0 45600 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_476
timestamp 1679581782
transform 1 0 46272 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_483
timestamp 1679581782
transform 1 0 46944 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_490
timestamp 1679581782
transform 1 0 47616 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_497
timestamp 1679581782
transform 1 0 48288 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_504
timestamp 1679581782
transform 1 0 48960 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_511
timestamp 1679581782
transform 1 0 49632 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_518
timestamp 1679581782
transform 1 0 50304 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_525
timestamp 1679581782
transform 1 0 50976 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_532
timestamp 1679581782
transform 1 0 51648 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_539
timestamp 1679581782
transform 1 0 52320 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_546
timestamp 1679581782
transform 1 0 52992 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_553
timestamp 1679581782
transform 1 0 53664 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_560
timestamp 1679581782
transform 1 0 54336 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_567
timestamp 1679581782
transform 1 0 55008 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_574
timestamp 1679581782
transform 1 0 55680 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_581
timestamp 1679581782
transform 1 0 56352 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_588
timestamp 1679581782
transform 1 0 57024 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_595
timestamp 1679581782
transform 1 0 57696 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_602
timestamp 1679581782
transform 1 0 58368 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_609
timestamp 1679581782
transform 1 0 59040 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_616
timestamp 1679581782
transform 1 0 59712 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_623
timestamp 1679581782
transform 1 0 60384 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_630
timestamp 1679581782
transform 1 0 61056 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_637
timestamp 1679581782
transform 1 0 61728 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_644
timestamp 1679581782
transform 1 0 62400 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_651
timestamp 1679581782
transform 1 0 63072 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_658
timestamp 1679581782
transform 1 0 63744 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_665
timestamp 1679581782
transform 1 0 64416 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_672
timestamp 1679581782
transform 1 0 65088 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_679
timestamp 1679581782
transform 1 0 65760 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_686
timestamp 1679581782
transform 1 0 66432 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_693
timestamp 1679581782
transform 1 0 67104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_700
timestamp 1679581782
transform 1 0 67776 0 1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_707
timestamp 1679581782
transform 1 0 68448 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_714
timestamp 1679577901
transform 1 0 69120 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_718
timestamp 1677580104
transform 1 0 69504 0 1 26460
box -48 -56 240 834
use sg13g2_fill_2  FILLER_34_724
timestamp 1677580104
transform 1 0 70080 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_738
timestamp 1677579658
transform 1 0 71424 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 576 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679581782
transform 1 0 1248 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679581782
transform 1 0 1920 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679581782
transform 1 0 2592 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_28
timestamp 1679581782
transform 1 0 3264 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_35
timestamp 1679581782
transform 1 0 3936 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_42
timestamp 1679581782
transform 1 0 4608 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_49
timestamp 1679581782
transform 1 0 5280 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_56
timestamp 1679581782
transform 1 0 5952 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_63
timestamp 1679581782
transform 1 0 6624 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_70
timestamp 1679581782
transform 1 0 7296 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_77
timestamp 1679581782
transform 1 0 7968 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_84
timestamp 1679581782
transform 1 0 8640 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_91
timestamp 1679581782
transform 1 0 9312 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_98
timestamp 1679581782
transform 1 0 9984 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_105
timestamp 1679581782
transform 1 0 10656 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_112
timestamp 1679581782
transform 1 0 11328 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_119
timestamp 1679581782
transform 1 0 12000 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_126
timestamp 1679581782
transform 1 0 12672 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_133
timestamp 1679581782
transform 1 0 13344 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_140
timestamp 1679581782
transform 1 0 14016 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_147
timestamp 1679581782
transform 1 0 14688 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_154
timestamp 1679581782
transform 1 0 15360 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_161
timestamp 1679581782
transform 1 0 16032 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_168
timestamp 1679581782
transform 1 0 16704 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_175
timestamp 1679581782
transform 1 0 17376 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_182
timestamp 1679581782
transform 1 0 18048 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_189
timestamp 1679581782
transform 1 0 18720 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_196
timestamp 1679581782
transform 1 0 19392 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_203
timestamp 1679581782
transform 1 0 20064 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_210
timestamp 1679581782
transform 1 0 20736 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_217
timestamp 1679581782
transform 1 0 21408 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_224
timestamp 1679581782
transform 1 0 22080 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_231
timestamp 1679581782
transform 1 0 22752 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_238
timestamp 1679581782
transform 1 0 23424 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_245
timestamp 1679581782
transform 1 0 24096 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_252
timestamp 1679581782
transform 1 0 24768 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_259
timestamp 1679581782
transform 1 0 25440 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_266
timestamp 1679581782
transform 1 0 26112 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_273
timestamp 1679581782
transform 1 0 26784 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_280
timestamp 1679581782
transform 1 0 27456 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_287
timestamp 1679581782
transform 1 0 28128 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_294
timestamp 1679581782
transform 1 0 28800 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_301
timestamp 1679581782
transform 1 0 29472 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_308
timestamp 1679581782
transform 1 0 30144 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_315
timestamp 1679581782
transform 1 0 30816 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_322
timestamp 1679581782
transform 1 0 31488 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_329
timestamp 1679581782
transform 1 0 32160 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_336
timestamp 1679581782
transform 1 0 32832 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_343
timestamp 1679581782
transform 1 0 33504 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_350
timestamp 1679581782
transform 1 0 34176 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_357
timestamp 1679581782
transform 1 0 34848 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_364
timestamp 1679581782
transform 1 0 35520 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_371
timestamp 1679581782
transform 1 0 36192 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_378
timestamp 1679581782
transform 1 0 36864 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_385
timestamp 1679581782
transform 1 0 37536 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_392
timestamp 1679581782
transform 1 0 38208 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_399
timestamp 1679581782
transform 1 0 38880 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_406
timestamp 1679581782
transform 1 0 39552 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_413
timestamp 1679581782
transform 1 0 40224 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_420
timestamp 1679581782
transform 1 0 40896 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_427
timestamp 1679581782
transform 1 0 41568 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_434
timestamp 1679581782
transform 1 0 42240 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_441
timestamp 1679581782
transform 1 0 42912 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_448
timestamp 1679581782
transform 1 0 43584 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_455
timestamp 1679581782
transform 1 0 44256 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_462
timestamp 1679581782
transform 1 0 44928 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_469
timestamp 1679581782
transform 1 0 45600 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_476
timestamp 1679581782
transform 1 0 46272 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_483
timestamp 1679581782
transform 1 0 46944 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_490
timestamp 1679581782
transform 1 0 47616 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_497
timestamp 1679581782
transform 1 0 48288 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_504
timestamp 1679581782
transform 1 0 48960 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_511
timestamp 1679581782
transform 1 0 49632 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_518
timestamp 1679581782
transform 1 0 50304 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_525
timestamp 1679581782
transform 1 0 50976 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_532
timestamp 1679581782
transform 1 0 51648 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_539
timestamp 1679581782
transform 1 0 52320 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_546
timestamp 1679581782
transform 1 0 52992 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_553
timestamp 1679581782
transform 1 0 53664 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_560
timestamp 1679581782
transform 1 0 54336 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_567
timestamp 1679581782
transform 1 0 55008 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_574
timestamp 1679581782
transform 1 0 55680 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_581
timestamp 1679581782
transform 1 0 56352 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_588
timestamp 1679581782
transform 1 0 57024 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_595
timestamp 1679581782
transform 1 0 57696 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_602
timestamp 1679581782
transform 1 0 58368 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_609
timestamp 1679581782
transform 1 0 59040 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_616
timestamp 1679581782
transform 1 0 59712 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_623
timestamp 1679581782
transform 1 0 60384 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_630
timestamp 1679581782
transform 1 0 61056 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_637
timestamp 1679581782
transform 1 0 61728 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_644
timestamp 1679581782
transform 1 0 62400 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_651
timestamp 1679581782
transform 1 0 63072 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_658
timestamp 1679581782
transform 1 0 63744 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_665
timestamp 1679581782
transform 1 0 64416 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_672
timestamp 1679581782
transform 1 0 65088 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_679
timestamp 1679581782
transform 1 0 65760 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_686
timestamp 1679581782
transform 1 0 66432 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_693
timestamp 1679581782
transform 1 0 67104 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_700
timestamp 1679581782
transform 1 0 67776 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_707
timestamp 1679581782
transform 1 0 68448 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_714
timestamp 1679581782
transform 1 0 69120 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_730
timestamp 1677580104
transform 1 0 70656 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 576 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679581782
transform 1 0 1248 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679581782
transform 1 0 1920 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679581782
transform 1 0 2592 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679581782
transform 1 0 3264 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679581782
transform 1 0 3936 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679581782
transform 1 0 4608 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679581782
transform 1 0 5280 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_56
timestamp 1679581782
transform 1 0 5952 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_63
timestamp 1679581782
transform 1 0 6624 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_70
timestamp 1679581782
transform 1 0 7296 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_77
timestamp 1679581782
transform 1 0 7968 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_84
timestamp 1679581782
transform 1 0 8640 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_91
timestamp 1679581782
transform 1 0 9312 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_98
timestamp 1679581782
transform 1 0 9984 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_105
timestamp 1679581782
transform 1 0 10656 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_112
timestamp 1679581782
transform 1 0 11328 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_119
timestamp 1679581782
transform 1 0 12000 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679581782
transform 1 0 12672 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_133
timestamp 1679581782
transform 1 0 13344 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_140
timestamp 1679581782
transform 1 0 14016 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_147
timestamp 1679581782
transform 1 0 14688 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_154
timestamp 1679581782
transform 1 0 15360 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_161
timestamp 1679581782
transform 1 0 16032 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_168
timestamp 1679581782
transform 1 0 16704 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_175
timestamp 1679581782
transform 1 0 17376 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_182
timestamp 1679581782
transform 1 0 18048 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_189
timestamp 1679581782
transform 1 0 18720 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_196
timestamp 1679581782
transform 1 0 19392 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_203
timestamp 1679581782
transform 1 0 20064 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_210
timestamp 1679581782
transform 1 0 20736 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_217
timestamp 1679581782
transform 1 0 21408 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_224
timestamp 1679581782
transform 1 0 22080 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_231
timestamp 1679581782
transform 1 0 22752 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_238
timestamp 1679581782
transform 1 0 23424 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_245
timestamp 1679581782
transform 1 0 24096 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_252
timestamp 1679581782
transform 1 0 24768 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_259
timestamp 1679581782
transform 1 0 25440 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_266
timestamp 1679581782
transform 1 0 26112 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_273
timestamp 1679581782
transform 1 0 26784 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_280
timestamp 1679581782
transform 1 0 27456 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_287
timestamp 1679581782
transform 1 0 28128 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_294
timestamp 1679581782
transform 1 0 28800 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_301
timestamp 1679581782
transform 1 0 29472 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_308
timestamp 1679581782
transform 1 0 30144 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_315
timestamp 1679581782
transform 1 0 30816 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_322
timestamp 1679581782
transform 1 0 31488 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_329
timestamp 1679581782
transform 1 0 32160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_336
timestamp 1679581782
transform 1 0 32832 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_343
timestamp 1679581782
transform 1 0 33504 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_350
timestamp 1679581782
transform 1 0 34176 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_357
timestamp 1679581782
transform 1 0 34848 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_364
timestamp 1679581782
transform 1 0 35520 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_371
timestamp 1679581782
transform 1 0 36192 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_378
timestamp 1679581782
transform 1 0 36864 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_385
timestamp 1679581782
transform 1 0 37536 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_392
timestamp 1679581782
transform 1 0 38208 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_399
timestamp 1679581782
transform 1 0 38880 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_406
timestamp 1679581782
transform 1 0 39552 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_413
timestamp 1679581782
transform 1 0 40224 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_420
timestamp 1679581782
transform 1 0 40896 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_427
timestamp 1679581782
transform 1 0 41568 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_434
timestamp 1679581782
transform 1 0 42240 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_441
timestamp 1679581782
transform 1 0 42912 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_448
timestamp 1679581782
transform 1 0 43584 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_455
timestamp 1679581782
transform 1 0 44256 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_462
timestamp 1679581782
transform 1 0 44928 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_469
timestamp 1679581782
transform 1 0 45600 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_476
timestamp 1679581782
transform 1 0 46272 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_483
timestamp 1679581782
transform 1 0 46944 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_490
timestamp 1679581782
transform 1 0 47616 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_497
timestamp 1679581782
transform 1 0 48288 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_504
timestamp 1679581782
transform 1 0 48960 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_511
timestamp 1679581782
transform 1 0 49632 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_518
timestamp 1679581782
transform 1 0 50304 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_525
timestamp 1679581782
transform 1 0 50976 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_532
timestamp 1679581782
transform 1 0 51648 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_539
timestamp 1679581782
transform 1 0 52320 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_546
timestamp 1679581782
transform 1 0 52992 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_553
timestamp 1679581782
transform 1 0 53664 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_560
timestamp 1679581782
transform 1 0 54336 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_567
timestamp 1679581782
transform 1 0 55008 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_574
timestamp 1679581782
transform 1 0 55680 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_581
timestamp 1679581782
transform 1 0 56352 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_588
timestamp 1679581782
transform 1 0 57024 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_595
timestamp 1679581782
transform 1 0 57696 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_602
timestamp 1679581782
transform 1 0 58368 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_609
timestamp 1679581782
transform 1 0 59040 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_616
timestamp 1679581782
transform 1 0 59712 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_623
timestamp 1679581782
transform 1 0 60384 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_630
timestamp 1679581782
transform 1 0 61056 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_637
timestamp 1679581782
transform 1 0 61728 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_644
timestamp 1679581782
transform 1 0 62400 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_651
timestamp 1679581782
transform 1 0 63072 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_658
timestamp 1679581782
transform 1 0 63744 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_665
timestamp 1679581782
transform 1 0 64416 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_672
timestamp 1679581782
transform 1 0 65088 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_679
timestamp 1679581782
transform 1 0 65760 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_686
timestamp 1679581782
transform 1 0 66432 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_693
timestamp 1679581782
transform 1 0 67104 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_700
timestamp 1679581782
transform 1 0 67776 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_707
timestamp 1679581782
transform 1 0 68448 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_714
timestamp 1679581782
transform 1 0 69120 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_721
timestamp 1679581782
transform 1 0 69792 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_728
timestamp 1679581782
transform 1 0 70464 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_735
timestamp 1679577901
transform 1 0 71136 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 576 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679581782
transform 1 0 1248 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679581782
transform 1 0 1920 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679581782
transform 1 0 2592 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679581782
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679581782
transform 1 0 3936 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679581782
transform 1 0 4608 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679581782
transform 1 0 5280 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679581782
transform 1 0 5952 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679581782
transform 1 0 6624 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_70
timestamp 1679581782
transform 1 0 7296 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_77
timestamp 1679581782
transform 1 0 7968 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_84
timestamp 1679581782
transform 1 0 8640 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_91
timestamp 1679581782
transform 1 0 9312 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679581782
transform 1 0 9984 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679581782
transform 1 0 10656 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679581782
transform 1 0 11328 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679581782
transform 1 0 12000 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679581782
transform 1 0 12672 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679581782
transform 1 0 13344 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679581782
transform 1 0 14016 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_147
timestamp 1679581782
transform 1 0 14688 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_154
timestamp 1679581782
transform 1 0 15360 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_161
timestamp 1679581782
transform 1 0 16032 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_168
timestamp 1679581782
transform 1 0 16704 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_175
timestamp 1679581782
transform 1 0 17376 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_182
timestamp 1679581782
transform 1 0 18048 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_189
timestamp 1679581782
transform 1 0 18720 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_196
timestamp 1679581782
transform 1 0 19392 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_203
timestamp 1679581782
transform 1 0 20064 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_210
timestamp 1679581782
transform 1 0 20736 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_217
timestamp 1679581782
transform 1 0 21408 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_224
timestamp 1679581782
transform 1 0 22080 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_231
timestamp 1679581782
transform 1 0 22752 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_238
timestamp 1679581782
transform 1 0 23424 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_245
timestamp 1679581782
transform 1 0 24096 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_252
timestamp 1679581782
transform 1 0 24768 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_259
timestamp 1679581782
transform 1 0 25440 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_266
timestamp 1679581782
transform 1 0 26112 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_273
timestamp 1679581782
transform 1 0 26784 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_280
timestamp 1679581782
transform 1 0 27456 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_287
timestamp 1679581782
transform 1 0 28128 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_294
timestamp 1679581782
transform 1 0 28800 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_301
timestamp 1679581782
transform 1 0 29472 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_308
timestamp 1679581782
transform 1 0 30144 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_315
timestamp 1679581782
transform 1 0 30816 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_322
timestamp 1679581782
transform 1 0 31488 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_329
timestamp 1679581782
transform 1 0 32160 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_336
timestamp 1679581782
transform 1 0 32832 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_343
timestamp 1679581782
transform 1 0 33504 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_350
timestamp 1679581782
transform 1 0 34176 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_357
timestamp 1679581782
transform 1 0 34848 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_364
timestamp 1679581782
transform 1 0 35520 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_371
timestamp 1679581782
transform 1 0 36192 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_378
timestamp 1679581782
transform 1 0 36864 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_385
timestamp 1679581782
transform 1 0 37536 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_392
timestamp 1679581782
transform 1 0 38208 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_399
timestamp 1679581782
transform 1 0 38880 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_406
timestamp 1679581782
transform 1 0 39552 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_413
timestamp 1679581782
transform 1 0 40224 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_420
timestamp 1679581782
transform 1 0 40896 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_427
timestamp 1679581782
transform 1 0 41568 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_434
timestamp 1679581782
transform 1 0 42240 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_441
timestamp 1679581782
transform 1 0 42912 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_448
timestamp 1679581782
transform 1 0 43584 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_455
timestamp 1679581782
transform 1 0 44256 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_462
timestamp 1679581782
transform 1 0 44928 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_469
timestamp 1679581782
transform 1 0 45600 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_476
timestamp 1679581782
transform 1 0 46272 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_483
timestamp 1679581782
transform 1 0 46944 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_490
timestamp 1679581782
transform 1 0 47616 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_497
timestamp 1679581782
transform 1 0 48288 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_504
timestamp 1679581782
transform 1 0 48960 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_511
timestamp 1679581782
transform 1 0 49632 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_518
timestamp 1679581782
transform 1 0 50304 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_525
timestamp 1679581782
transform 1 0 50976 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_532
timestamp 1679581782
transform 1 0 51648 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_539
timestamp 1679581782
transform 1 0 52320 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_546
timestamp 1679581782
transform 1 0 52992 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_553
timestamp 1679581782
transform 1 0 53664 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_560
timestamp 1679581782
transform 1 0 54336 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_567
timestamp 1679581782
transform 1 0 55008 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_574
timestamp 1679581782
transform 1 0 55680 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_581
timestamp 1679581782
transform 1 0 56352 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_588
timestamp 1679581782
transform 1 0 57024 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_595
timestamp 1679581782
transform 1 0 57696 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_602
timestamp 1679581782
transform 1 0 58368 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_609
timestamp 1679581782
transform 1 0 59040 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_616
timestamp 1679581782
transform 1 0 59712 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_623
timestamp 1679581782
transform 1 0 60384 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_630
timestamp 1679581782
transform 1 0 61056 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_637
timestamp 1679581782
transform 1 0 61728 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_644
timestamp 1679581782
transform 1 0 62400 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_651
timestamp 1679581782
transform 1 0 63072 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_658
timestamp 1679581782
transform 1 0 63744 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_665
timestamp 1679581782
transform 1 0 64416 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_672
timestamp 1679581782
transform 1 0 65088 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_679
timestamp 1679581782
transform 1 0 65760 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_686
timestamp 1679581782
transform 1 0 66432 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_693
timestamp 1679581782
transform 1 0 67104 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_700
timestamp 1679581782
transform 1 0 67776 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_707
timestamp 1679581782
transform 1 0 68448 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_714
timestamp 1679581782
transform 1 0 69120 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_721
timestamp 1679581782
transform 1 0 69792 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_728
timestamp 1679581782
transform 1 0 70464 0 -1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_735
timestamp 1679577901
transform 1 0 71136 0 -1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 576 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679581782
transform 1 0 1248 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679581782
transform 1 0 1920 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679581782
transform 1 0 2592 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679581782
transform 1 0 3264 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679581782
transform 1 0 3936 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679581782
transform 1 0 4608 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679581782
transform 1 0 5280 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_56
timestamp 1679581782
transform 1 0 5952 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_63
timestamp 1679581782
transform 1 0 6624 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_70
timestamp 1679581782
transform 1 0 7296 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_77
timestamp 1679581782
transform 1 0 7968 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_84
timestamp 1679581782
transform 1 0 8640 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_91
timestamp 1679581782
transform 1 0 9312 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_98
timestamp 1679581782
transform 1 0 9984 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_105
timestamp 1679581782
transform 1 0 10656 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_112
timestamp 1679581782
transform 1 0 11328 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_119
timestamp 1679581782
transform 1 0 12000 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_126
timestamp 1679581782
transform 1 0 12672 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_133
timestamp 1679581782
transform 1 0 13344 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_140
timestamp 1679581782
transform 1 0 14016 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_147
timestamp 1679581782
transform 1 0 14688 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_154
timestamp 1679581782
transform 1 0 15360 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_161
timestamp 1679581782
transform 1 0 16032 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_168
timestamp 1679581782
transform 1 0 16704 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_175
timestamp 1679581782
transform 1 0 17376 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_182
timestamp 1679581782
transform 1 0 18048 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_189
timestamp 1679581782
transform 1 0 18720 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_196
timestamp 1679581782
transform 1 0 19392 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_203
timestamp 1679581782
transform 1 0 20064 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_210
timestamp 1679581782
transform 1 0 20736 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_217
timestamp 1679581782
transform 1 0 21408 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_224
timestamp 1679581782
transform 1 0 22080 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_231
timestamp 1679581782
transform 1 0 22752 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_238
timestamp 1679581782
transform 1 0 23424 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_245
timestamp 1679581782
transform 1 0 24096 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_252
timestamp 1679581782
transform 1 0 24768 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_259
timestamp 1679581782
transform 1 0 25440 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_266
timestamp 1679581782
transform 1 0 26112 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_273
timestamp 1679581782
transform 1 0 26784 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_280
timestamp 1679581782
transform 1 0 27456 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_287
timestamp 1679581782
transform 1 0 28128 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_294
timestamp 1679581782
transform 1 0 28800 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_301
timestamp 1679581782
transform 1 0 29472 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_308
timestamp 1679581782
transform 1 0 30144 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_315
timestamp 1679581782
transform 1 0 30816 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_322
timestamp 1679581782
transform 1 0 31488 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_329
timestamp 1679581782
transform 1 0 32160 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_336
timestamp 1679581782
transform 1 0 32832 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_343
timestamp 1679581782
transform 1 0 33504 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_350
timestamp 1679581782
transform 1 0 34176 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_357
timestamp 1679581782
transform 1 0 34848 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_364
timestamp 1679581782
transform 1 0 35520 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_371
timestamp 1679581782
transform 1 0 36192 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_378
timestamp 1679581782
transform 1 0 36864 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_385
timestamp 1679581782
transform 1 0 37536 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_392
timestamp 1679581782
transform 1 0 38208 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_399
timestamp 1679581782
transform 1 0 38880 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_406
timestamp 1679581782
transform 1 0 39552 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_413
timestamp 1679581782
transform 1 0 40224 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_420
timestamp 1679581782
transform 1 0 40896 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_427
timestamp 1679581782
transform 1 0 41568 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_434
timestamp 1679581782
transform 1 0 42240 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_441
timestamp 1679581782
transform 1 0 42912 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_448
timestamp 1679581782
transform 1 0 43584 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_455
timestamp 1679581782
transform 1 0 44256 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_462
timestamp 1679581782
transform 1 0 44928 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_469
timestamp 1679581782
transform 1 0 45600 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_476
timestamp 1679581782
transform 1 0 46272 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_483
timestamp 1679581782
transform 1 0 46944 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_490
timestamp 1679581782
transform 1 0 47616 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_497
timestamp 1679581782
transform 1 0 48288 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_504
timestamp 1679581782
transform 1 0 48960 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_511
timestamp 1679581782
transform 1 0 49632 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_518
timestamp 1679581782
transform 1 0 50304 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_525
timestamp 1679581782
transform 1 0 50976 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_532
timestamp 1679581782
transform 1 0 51648 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_539
timestamp 1679581782
transform 1 0 52320 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_546
timestamp 1679581782
transform 1 0 52992 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_553
timestamp 1679581782
transform 1 0 53664 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_560
timestamp 1679581782
transform 1 0 54336 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_567
timestamp 1679581782
transform 1 0 55008 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_574
timestamp 1679581782
transform 1 0 55680 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_581
timestamp 1679581782
transform 1 0 56352 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_588
timestamp 1679581782
transform 1 0 57024 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_595
timestamp 1679581782
transform 1 0 57696 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_602
timestamp 1679581782
transform 1 0 58368 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_609
timestamp 1679581782
transform 1 0 59040 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_616
timestamp 1679581782
transform 1 0 59712 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_623
timestamp 1679581782
transform 1 0 60384 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_630
timestamp 1679581782
transform 1 0 61056 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_637
timestamp 1679581782
transform 1 0 61728 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_644
timestamp 1679581782
transform 1 0 62400 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_651
timestamp 1679581782
transform 1 0 63072 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_658
timestamp 1679581782
transform 1 0 63744 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_665
timestamp 1679581782
transform 1 0 64416 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_672
timestamp 1679581782
transform 1 0 65088 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_679
timestamp 1679581782
transform 1 0 65760 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_686
timestamp 1679581782
transform 1 0 66432 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_693
timestamp 1679581782
transform 1 0 67104 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_700
timestamp 1679581782
transform 1 0 67776 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_707
timestamp 1679581782
transform 1 0 68448 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_714
timestamp 1679581782
transform 1 0 69120 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_721
timestamp 1679581782
transform 1 0 69792 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_728
timestamp 1679581782
transform 1 0 70464 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_735
timestamp 1679577901
transform 1 0 71136 0 1 29484
box -48 -56 432 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 576 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679581782
transform 1 0 1248 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679581782
transform 1 0 1920 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679581782
transform 1 0 2592 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_28
timestamp 1679581782
transform 1 0 3264 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_35
timestamp 1679581782
transform 1 0 3936 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_42
timestamp 1679581782
transform 1 0 4608 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_49
timestamp 1679581782
transform 1 0 5280 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_56
timestamp 1679581782
transform 1 0 5952 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_63
timestamp 1679581782
transform 1 0 6624 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_70
timestamp 1679581782
transform 1 0 7296 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_77
timestamp 1679581782
transform 1 0 7968 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_84
timestamp 1679581782
transform 1 0 8640 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_91
timestamp 1679581782
transform 1 0 9312 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_98
timestamp 1679581782
transform 1 0 9984 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_105
timestamp 1679581782
transform 1 0 10656 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_112
timestamp 1679581782
transform 1 0 11328 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_119
timestamp 1679581782
transform 1 0 12000 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_126
timestamp 1679581782
transform 1 0 12672 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_133
timestamp 1679581782
transform 1 0 13344 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_140
timestamp 1679581782
transform 1 0 14016 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_147
timestamp 1679581782
transform 1 0 14688 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_154
timestamp 1679581782
transform 1 0 15360 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_161
timestamp 1679581782
transform 1 0 16032 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_168
timestamp 1679581782
transform 1 0 16704 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_175
timestamp 1679581782
transform 1 0 17376 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_182
timestamp 1679581782
transform 1 0 18048 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_189
timestamp 1679581782
transform 1 0 18720 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_196
timestamp 1679581782
transform 1 0 19392 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_203
timestamp 1679581782
transform 1 0 20064 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_210
timestamp 1679581782
transform 1 0 20736 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_217
timestamp 1679581782
transform 1 0 21408 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_224
timestamp 1679581782
transform 1 0 22080 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_231
timestamp 1679581782
transform 1 0 22752 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_238
timestamp 1679581782
transform 1 0 23424 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_245
timestamp 1679581782
transform 1 0 24096 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_252
timestamp 1679581782
transform 1 0 24768 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_259
timestamp 1679581782
transform 1 0 25440 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_266
timestamp 1679581782
transform 1 0 26112 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_273
timestamp 1679581782
transform 1 0 26784 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_280
timestamp 1679581782
transform 1 0 27456 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_287
timestamp 1679581782
transform 1 0 28128 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_294
timestamp 1679581782
transform 1 0 28800 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_301
timestamp 1679581782
transform 1 0 29472 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_308
timestamp 1679581782
transform 1 0 30144 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_315
timestamp 1679581782
transform 1 0 30816 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_322
timestamp 1679581782
transform 1 0 31488 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_329
timestamp 1679581782
transform 1 0 32160 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_336
timestamp 1679581782
transform 1 0 32832 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_343
timestamp 1679581782
transform 1 0 33504 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_350
timestamp 1679581782
transform 1 0 34176 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_357
timestamp 1679581782
transform 1 0 34848 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_364
timestamp 1679581782
transform 1 0 35520 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_371
timestamp 1679581782
transform 1 0 36192 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_378
timestamp 1679581782
transform 1 0 36864 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_385
timestamp 1679581782
transform 1 0 37536 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_392
timestamp 1679581782
transform 1 0 38208 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_399
timestamp 1679581782
transform 1 0 38880 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_406
timestamp 1679581782
transform 1 0 39552 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_413
timestamp 1679581782
transform 1 0 40224 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_420
timestamp 1679581782
transform 1 0 40896 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_427
timestamp 1679581782
transform 1 0 41568 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_434
timestamp 1679581782
transform 1 0 42240 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_441
timestamp 1679581782
transform 1 0 42912 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_448
timestamp 1679581782
transform 1 0 43584 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_455
timestamp 1679581782
transform 1 0 44256 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_462
timestamp 1679581782
transform 1 0 44928 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_469
timestamp 1679581782
transform 1 0 45600 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_476
timestamp 1679581782
transform 1 0 46272 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_483
timestamp 1679581782
transform 1 0 46944 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_490
timestamp 1679581782
transform 1 0 47616 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_497
timestamp 1679581782
transform 1 0 48288 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_504
timestamp 1679581782
transform 1 0 48960 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_511
timestamp 1679581782
transform 1 0 49632 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_518
timestamp 1679581782
transform 1 0 50304 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_525
timestamp 1679581782
transform 1 0 50976 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_532
timestamp 1679581782
transform 1 0 51648 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_539
timestamp 1679581782
transform 1 0 52320 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_546
timestamp 1679581782
transform 1 0 52992 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_553
timestamp 1679581782
transform 1 0 53664 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_560
timestamp 1679581782
transform 1 0 54336 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_567
timestamp 1679581782
transform 1 0 55008 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_574
timestamp 1679581782
transform 1 0 55680 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_581
timestamp 1679581782
transform 1 0 56352 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_588
timestamp 1679581782
transform 1 0 57024 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_595
timestamp 1679581782
transform 1 0 57696 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_602
timestamp 1679581782
transform 1 0 58368 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_609
timestamp 1679581782
transform 1 0 59040 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_616
timestamp 1679581782
transform 1 0 59712 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_623
timestamp 1679581782
transform 1 0 60384 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_630
timestamp 1679581782
transform 1 0 61056 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_637
timestamp 1679581782
transform 1 0 61728 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_644
timestamp 1679581782
transform 1 0 62400 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_651
timestamp 1679581782
transform 1 0 63072 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_658
timestamp 1679581782
transform 1 0 63744 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_665
timestamp 1679581782
transform 1 0 64416 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_672
timestamp 1679581782
transform 1 0 65088 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_679
timestamp 1679581782
transform 1 0 65760 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_686
timestamp 1679581782
transform 1 0 66432 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_693
timestamp 1679581782
transform 1 0 67104 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_700
timestamp 1679581782
transform 1 0 67776 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_707
timestamp 1679581782
transform 1 0 68448 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_714
timestamp 1679581782
transform 1 0 69120 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_721
timestamp 1679581782
transform 1 0 69792 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_728
timestamp 1679581782
transform 1 0 70464 0 -1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_39_735
timestamp 1679577901
transform 1 0 71136 0 -1 30996
box -48 -56 432 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 576 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679581782
transform 1 0 1248 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679581782
transform 1 0 1920 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679581782
transform 1 0 2592 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_28
timestamp 1679581782
transform 1 0 3264 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_35
timestamp 1679581782
transform 1 0 3936 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_42
timestamp 1679581782
transform 1 0 4608 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_49
timestamp 1679581782
transform 1 0 5280 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_56
timestamp 1679581782
transform 1 0 5952 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_63
timestamp 1679581782
transform 1 0 6624 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_70
timestamp 1679581782
transform 1 0 7296 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_77
timestamp 1679581782
transform 1 0 7968 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_84
timestamp 1679581782
transform 1 0 8640 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_91
timestamp 1679581782
transform 1 0 9312 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_98
timestamp 1679581782
transform 1 0 9984 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_105
timestamp 1679581782
transform 1 0 10656 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_112
timestamp 1679581782
transform 1 0 11328 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_119
timestamp 1679581782
transform 1 0 12000 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_126
timestamp 1679581782
transform 1 0 12672 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_133
timestamp 1679581782
transform 1 0 13344 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_140
timestamp 1679581782
transform 1 0 14016 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_147
timestamp 1679581782
transform 1 0 14688 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_154
timestamp 1679581782
transform 1 0 15360 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_161
timestamp 1679581782
transform 1 0 16032 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_168
timestamp 1679581782
transform 1 0 16704 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_175
timestamp 1679581782
transform 1 0 17376 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_182
timestamp 1679581782
transform 1 0 18048 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_189
timestamp 1679581782
transform 1 0 18720 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_196
timestamp 1679581782
transform 1 0 19392 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_203
timestamp 1679581782
transform 1 0 20064 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_210
timestamp 1679581782
transform 1 0 20736 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_217
timestamp 1679581782
transform 1 0 21408 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_224
timestamp 1679581782
transform 1 0 22080 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_231
timestamp 1679581782
transform 1 0 22752 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_238
timestamp 1679581782
transform 1 0 23424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_245
timestamp 1679581782
transform 1 0 24096 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_252
timestamp 1679581782
transform 1 0 24768 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_259
timestamp 1679581782
transform 1 0 25440 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_266
timestamp 1679581782
transform 1 0 26112 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_273
timestamp 1679581782
transform 1 0 26784 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_280
timestamp 1679581782
transform 1 0 27456 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_287
timestamp 1679581782
transform 1 0 28128 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_294
timestamp 1679581782
transform 1 0 28800 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_301
timestamp 1679581782
transform 1 0 29472 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_308
timestamp 1679581782
transform 1 0 30144 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_315
timestamp 1679581782
transform 1 0 30816 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_322
timestamp 1679581782
transform 1 0 31488 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_329
timestamp 1679581782
transform 1 0 32160 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_336
timestamp 1679581782
transform 1 0 32832 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_343
timestamp 1679581782
transform 1 0 33504 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_350
timestamp 1679581782
transform 1 0 34176 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_357
timestamp 1679581782
transform 1 0 34848 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_364
timestamp 1679581782
transform 1 0 35520 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_371
timestamp 1679581782
transform 1 0 36192 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_378
timestamp 1679581782
transform 1 0 36864 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_385
timestamp 1679581782
transform 1 0 37536 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_392
timestamp 1679581782
transform 1 0 38208 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_399
timestamp 1679581782
transform 1 0 38880 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_406
timestamp 1679581782
transform 1 0 39552 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_413
timestamp 1679581782
transform 1 0 40224 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_420
timestamp 1679581782
transform 1 0 40896 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_427
timestamp 1679581782
transform 1 0 41568 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_434
timestamp 1679581782
transform 1 0 42240 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_441
timestamp 1679581782
transform 1 0 42912 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_448
timestamp 1679581782
transform 1 0 43584 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_455
timestamp 1679581782
transform 1 0 44256 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_462
timestamp 1679581782
transform 1 0 44928 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_469
timestamp 1679581782
transform 1 0 45600 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_476
timestamp 1679581782
transform 1 0 46272 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_483
timestamp 1679581782
transform 1 0 46944 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_490
timestamp 1679581782
transform 1 0 47616 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_497
timestamp 1679581782
transform 1 0 48288 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_504
timestamp 1679581782
transform 1 0 48960 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_511
timestamp 1679581782
transform 1 0 49632 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_518
timestamp 1679581782
transform 1 0 50304 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_525
timestamp 1679581782
transform 1 0 50976 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_532
timestamp 1679581782
transform 1 0 51648 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_539
timestamp 1679581782
transform 1 0 52320 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_546
timestamp 1679581782
transform 1 0 52992 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_553
timestamp 1679581782
transform 1 0 53664 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_560
timestamp 1679581782
transform 1 0 54336 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_567
timestamp 1679581782
transform 1 0 55008 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_574
timestamp 1679581782
transform 1 0 55680 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_581
timestamp 1679581782
transform 1 0 56352 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_588
timestamp 1679581782
transform 1 0 57024 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_595
timestamp 1679581782
transform 1 0 57696 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_602
timestamp 1679581782
transform 1 0 58368 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_609
timestamp 1679581782
transform 1 0 59040 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_616
timestamp 1679581782
transform 1 0 59712 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_623
timestamp 1679581782
transform 1 0 60384 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_630
timestamp 1679581782
transform 1 0 61056 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_637
timestamp 1679581782
transform 1 0 61728 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_644
timestamp 1679581782
transform 1 0 62400 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_651
timestamp 1679581782
transform 1 0 63072 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_658
timestamp 1679581782
transform 1 0 63744 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_665
timestamp 1679581782
transform 1 0 64416 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_672
timestamp 1679581782
transform 1 0 65088 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_679
timestamp 1679581782
transform 1 0 65760 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_686
timestamp 1679581782
transform 1 0 66432 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_693
timestamp 1679581782
transform 1 0 67104 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_700
timestamp 1679581782
transform 1 0 67776 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_707
timestamp 1679581782
transform 1 0 68448 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_714
timestamp 1679581782
transform 1 0 69120 0 1 30996
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_721
timestamp 1679581782
transform 1 0 69792 0 1 30996
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_728
timestamp 1677579658
transform 1 0 70464 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_736
timestamp 1677580104
transform 1 0 71232 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_738
timestamp 1677579658
transform 1 0 71424 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 576 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679581782
transform 1 0 1248 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679581782
transform 1 0 1920 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679581782
transform 1 0 2592 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679581782
transform 1 0 3264 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679581782
transform 1 0 3936 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679581782
transform 1 0 4608 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679581782
transform 1 0 5280 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679581782
transform 1 0 5952 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_63
timestamp 1679581782
transform 1 0 6624 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_70
timestamp 1679581782
transform 1 0 7296 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_77
timestamp 1679581782
transform 1 0 7968 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_84
timestamp 1679581782
transform 1 0 8640 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_91
timestamp 1679581782
transform 1 0 9312 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_98
timestamp 1679581782
transform 1 0 9984 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_105
timestamp 1679581782
transform 1 0 10656 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_112
timestamp 1679581782
transform 1 0 11328 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_119
timestamp 1679581782
transform 1 0 12000 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_126
timestamp 1679581782
transform 1 0 12672 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_133
timestamp 1679581782
transform 1 0 13344 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_140
timestamp 1679581782
transform 1 0 14016 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_147
timestamp 1679581782
transform 1 0 14688 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_154
timestamp 1679581782
transform 1 0 15360 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679581782
transform 1 0 16032 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_168
timestamp 1679581782
transform 1 0 16704 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_175
timestamp 1679581782
transform 1 0 17376 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_182
timestamp 1679581782
transform 1 0 18048 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_189
timestamp 1679581782
transform 1 0 18720 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_196
timestamp 1679581782
transform 1 0 19392 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_203
timestamp 1679581782
transform 1 0 20064 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_210
timestamp 1679581782
transform 1 0 20736 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_217
timestamp 1679581782
transform 1 0 21408 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_224
timestamp 1679581782
transform 1 0 22080 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_231
timestamp 1679581782
transform 1 0 22752 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_238
timestamp 1679581782
transform 1 0 23424 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_245
timestamp 1679581782
transform 1 0 24096 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_252
timestamp 1679581782
transform 1 0 24768 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_259
timestamp 1679581782
transform 1 0 25440 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_266
timestamp 1679581782
transform 1 0 26112 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_273
timestamp 1679581782
transform 1 0 26784 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_280
timestamp 1679581782
transform 1 0 27456 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_287
timestamp 1679581782
transform 1 0 28128 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_294
timestamp 1679581782
transform 1 0 28800 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_301
timestamp 1679581782
transform 1 0 29472 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_308
timestamp 1679581782
transform 1 0 30144 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_315
timestamp 1679581782
transform 1 0 30816 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_322
timestamp 1679581782
transform 1 0 31488 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_329
timestamp 1679581782
transform 1 0 32160 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_336
timestamp 1679581782
transform 1 0 32832 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_343
timestamp 1679581782
transform 1 0 33504 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_350
timestamp 1679581782
transform 1 0 34176 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_357
timestamp 1679581782
transform 1 0 34848 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_364
timestamp 1679581782
transform 1 0 35520 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_371
timestamp 1679581782
transform 1 0 36192 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_378
timestamp 1679581782
transform 1 0 36864 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_385
timestamp 1679581782
transform 1 0 37536 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_392
timestamp 1679581782
transform 1 0 38208 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_399
timestamp 1679581782
transform 1 0 38880 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_406
timestamp 1679581782
transform 1 0 39552 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_413
timestamp 1679581782
transform 1 0 40224 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_420
timestamp 1679581782
transform 1 0 40896 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_427
timestamp 1679581782
transform 1 0 41568 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_434
timestamp 1679581782
transform 1 0 42240 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_441
timestamp 1679581782
transform 1 0 42912 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_448
timestamp 1679581782
transform 1 0 43584 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_455
timestamp 1679581782
transform 1 0 44256 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_462
timestamp 1679581782
transform 1 0 44928 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_469
timestamp 1679581782
transform 1 0 45600 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_476
timestamp 1679581782
transform 1 0 46272 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_483
timestamp 1679581782
transform 1 0 46944 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_490
timestamp 1679581782
transform 1 0 47616 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_497
timestamp 1679581782
transform 1 0 48288 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_504
timestamp 1679581782
transform 1 0 48960 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_511
timestamp 1679581782
transform 1 0 49632 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_518
timestamp 1679581782
transform 1 0 50304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_525
timestamp 1679581782
transform 1 0 50976 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_532
timestamp 1679581782
transform 1 0 51648 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_539
timestamp 1679581782
transform 1 0 52320 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_546
timestamp 1679581782
transform 1 0 52992 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_553
timestamp 1679581782
transform 1 0 53664 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_560
timestamp 1679581782
transform 1 0 54336 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_567
timestamp 1679581782
transform 1 0 55008 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_574
timestamp 1679581782
transform 1 0 55680 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_581
timestamp 1679581782
transform 1 0 56352 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_588
timestamp 1679581782
transform 1 0 57024 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_595
timestamp 1679581782
transform 1 0 57696 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_602
timestamp 1679581782
transform 1 0 58368 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_609
timestamp 1679581782
transform 1 0 59040 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_616
timestamp 1679581782
transform 1 0 59712 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_623
timestamp 1679581782
transform 1 0 60384 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_630
timestamp 1679581782
transform 1 0 61056 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_637
timestamp 1679581782
transform 1 0 61728 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_644
timestamp 1679581782
transform 1 0 62400 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_651
timestamp 1679581782
transform 1 0 63072 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_658
timestamp 1679581782
transform 1 0 63744 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_665
timestamp 1679581782
transform 1 0 64416 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_672
timestamp 1679581782
transform 1 0 65088 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_679
timestamp 1679581782
transform 1 0 65760 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_686
timestamp 1679581782
transform 1 0 66432 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_693
timestamp 1679581782
transform 1 0 67104 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_700
timestamp 1679581782
transform 1 0 67776 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_707
timestamp 1679581782
transform 1 0 68448 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_714
timestamp 1679581782
transform 1 0 69120 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_721
timestamp 1679581782
transform 1 0 69792 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_728
timestamp 1677580104
transform 1 0 70464 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_734
timestamp 1677579658
transform 1 0 71040 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 1248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679581782
transform 1 0 1920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679581782
transform 1 0 2592 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679581782
transform 1 0 3264 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679581782
transform 1 0 3936 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679581782
transform 1 0 4608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_49
timestamp 1679581782
transform 1 0 5280 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_56
timestamp 1679581782
transform 1 0 5952 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_63
timestamp 1679581782
transform 1 0 6624 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_70
timestamp 1679581782
transform 1 0 7296 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_77
timestamp 1679581782
transform 1 0 7968 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_84
timestamp 1679581782
transform 1 0 8640 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_91
timestamp 1679581782
transform 1 0 9312 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_98
timestamp 1679581782
transform 1 0 9984 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_105
timestamp 1679581782
transform 1 0 10656 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_112
timestamp 1679581782
transform 1 0 11328 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_119
timestamp 1679581782
transform 1 0 12000 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_126
timestamp 1679581782
transform 1 0 12672 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_133
timestamp 1679581782
transform 1 0 13344 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_140
timestamp 1679581782
transform 1 0 14016 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_147
timestamp 1679581782
transform 1 0 14688 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_154
timestamp 1679581782
transform 1 0 15360 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_161
timestamp 1679581782
transform 1 0 16032 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_168
timestamp 1679581782
transform 1 0 16704 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_175
timestamp 1679581782
transform 1 0 17376 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_182
timestamp 1679581782
transform 1 0 18048 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_189
timestamp 1679581782
transform 1 0 18720 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_196
timestamp 1679581782
transform 1 0 19392 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_203
timestamp 1679581782
transform 1 0 20064 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_210
timestamp 1679581782
transform 1 0 20736 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_217
timestamp 1679581782
transform 1 0 21408 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_224
timestamp 1679581782
transform 1 0 22080 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_231
timestamp 1679581782
transform 1 0 22752 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_238
timestamp 1679581782
transform 1 0 23424 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_245
timestamp 1679581782
transform 1 0 24096 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_252
timestamp 1679581782
transform 1 0 24768 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_259
timestamp 1679581782
transform 1 0 25440 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_266
timestamp 1679581782
transform 1 0 26112 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_273
timestamp 1679581782
transform 1 0 26784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_280
timestamp 1679581782
transform 1 0 27456 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_287
timestamp 1679581782
transform 1 0 28128 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_294
timestamp 1679581782
transform 1 0 28800 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_301
timestamp 1679581782
transform 1 0 29472 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_308
timestamp 1679581782
transform 1 0 30144 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_315
timestamp 1679581782
transform 1 0 30816 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_322
timestamp 1679581782
transform 1 0 31488 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_329
timestamp 1679581782
transform 1 0 32160 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_336
timestamp 1679581782
transform 1 0 32832 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_343
timestamp 1679581782
transform 1 0 33504 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_350
timestamp 1679581782
transform 1 0 34176 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_357
timestamp 1679581782
transform 1 0 34848 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_364
timestamp 1679581782
transform 1 0 35520 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_371
timestamp 1679581782
transform 1 0 36192 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_378
timestamp 1679581782
transform 1 0 36864 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_385
timestamp 1679581782
transform 1 0 37536 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_392
timestamp 1679581782
transform 1 0 38208 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_399
timestamp 1679581782
transform 1 0 38880 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_406
timestamp 1679581782
transform 1 0 39552 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_413
timestamp 1679581782
transform 1 0 40224 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_420
timestamp 1679581782
transform 1 0 40896 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_427
timestamp 1679581782
transform 1 0 41568 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_434
timestamp 1679581782
transform 1 0 42240 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_441
timestamp 1679581782
transform 1 0 42912 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_448
timestamp 1679581782
transform 1 0 43584 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_455
timestamp 1679581782
transform 1 0 44256 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_462
timestamp 1679581782
transform 1 0 44928 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_469
timestamp 1679581782
transform 1 0 45600 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_476
timestamp 1679581782
transform 1 0 46272 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_483
timestamp 1679581782
transform 1 0 46944 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_490
timestamp 1679581782
transform 1 0 47616 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_497
timestamp 1679581782
transform 1 0 48288 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_504
timestamp 1679581782
transform 1 0 48960 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_511
timestamp 1679581782
transform 1 0 49632 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_518
timestamp 1679581782
transform 1 0 50304 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_525
timestamp 1679581782
transform 1 0 50976 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_532
timestamp 1679581782
transform 1 0 51648 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_539
timestamp 1679581782
transform 1 0 52320 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_546
timestamp 1679581782
transform 1 0 52992 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_553
timestamp 1679581782
transform 1 0 53664 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_560
timestamp 1679581782
transform 1 0 54336 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_567
timestamp 1679581782
transform 1 0 55008 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_574
timestamp 1679581782
transform 1 0 55680 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_581
timestamp 1679581782
transform 1 0 56352 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_588
timestamp 1679581782
transform 1 0 57024 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_595
timestamp 1679581782
transform 1 0 57696 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_602
timestamp 1679581782
transform 1 0 58368 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_609
timestamp 1679581782
transform 1 0 59040 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_616
timestamp 1679581782
transform 1 0 59712 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_623
timestamp 1679581782
transform 1 0 60384 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_630
timestamp 1679581782
transform 1 0 61056 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_637
timestamp 1679581782
transform 1 0 61728 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_644
timestamp 1679581782
transform 1 0 62400 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_651
timestamp 1679581782
transform 1 0 63072 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_658
timestamp 1679581782
transform 1 0 63744 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_665
timestamp 1679581782
transform 1 0 64416 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_672
timestamp 1679581782
transform 1 0 65088 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_679
timestamp 1679581782
transform 1 0 65760 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_686
timestamp 1679581782
transform 1 0 66432 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_693
timestamp 1679581782
transform 1 0 67104 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_700
timestamp 1679581782
transform 1 0 67776 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_707
timestamp 1679581782
transform 1 0 68448 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_714
timestamp 1679581782
transform 1 0 69120 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_721
timestamp 1679581782
transform 1 0 69792 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_728
timestamp 1679581782
transform 1 0 70464 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_735
timestamp 1677580104
transform 1 0 71136 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_737
timestamp 1677579658
transform 1 0 71328 0 1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_42_741
timestamp 1679577901
transform 1 0 71712 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_745
timestamp 1677580104
transform 1 0 72096 0 1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_42_757
timestamp 1677580104
transform 1 0 73248 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_759
timestamp 1677579658
transform 1 0 73440 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_770
timestamp 1677579658
transform 1 0 74496 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_781
timestamp 1677580104
transform 1 0 75552 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_812
timestamp 1677579658
transform 1 0 78528 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_832
timestamp 1677579658
transform 1 0 80448 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_891
timestamp 1677579658
transform 1 0 86112 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_908
timestamp 1677579658
transform 1 0 87744 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_919
timestamp 1677579658
transform 1 0 88800 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_936
timestamp 1677580104
transform 1 0 90432 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_954
timestamp 1677579658
transform 1 0 92160 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_999
timestamp 1677580104
transform 1 0 96480 0 1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_42_1017
timestamp 1677580104
transform 1 0 98208 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 576 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 1248 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679581782
transform 1 0 1920 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679581782
transform 1 0 2592 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679581782
transform 1 0 3264 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679581782
transform 1 0 3936 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679581782
transform 1 0 4608 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679581782
transform 1 0 5280 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679581782
transform 1 0 5952 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679581782
transform 1 0 6624 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679581782
transform 1 0 7296 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679581782
transform 1 0 7968 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679581782
transform 1 0 8640 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679581782
transform 1 0 9312 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679581782
transform 1 0 9984 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679581782
transform 1 0 10656 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_112
timestamp 1679581782
transform 1 0 11328 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_119
timestamp 1679581782
transform 1 0 12000 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_126
timestamp 1679581782
transform 1 0 12672 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_133
timestamp 1679581782
transform 1 0 13344 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_140
timestamp 1679581782
transform 1 0 14016 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_147
timestamp 1679581782
transform 1 0 14688 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_154
timestamp 1679581782
transform 1 0 15360 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_161
timestamp 1679581782
transform 1 0 16032 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_168
timestamp 1679581782
transform 1 0 16704 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_175
timestamp 1679581782
transform 1 0 17376 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_182
timestamp 1679581782
transform 1 0 18048 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_189
timestamp 1679581782
transform 1 0 18720 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_196
timestamp 1679581782
transform 1 0 19392 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_203
timestamp 1679581782
transform 1 0 20064 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_210
timestamp 1679581782
transform 1 0 20736 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_217
timestamp 1679581782
transform 1 0 21408 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_224
timestamp 1679581782
transform 1 0 22080 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_231
timestamp 1679581782
transform 1 0 22752 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_238
timestamp 1679581782
transform 1 0 23424 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_245
timestamp 1679581782
transform 1 0 24096 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_252
timestamp 1679581782
transform 1 0 24768 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_259
timestamp 1679581782
transform 1 0 25440 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_266
timestamp 1679581782
transform 1 0 26112 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_273
timestamp 1679581782
transform 1 0 26784 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_280
timestamp 1679581782
transform 1 0 27456 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_287
timestamp 1679581782
transform 1 0 28128 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_294
timestamp 1679581782
transform 1 0 28800 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_301
timestamp 1679581782
transform 1 0 29472 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_308
timestamp 1679581782
transform 1 0 30144 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_315
timestamp 1679581782
transform 1 0 30816 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_322
timestamp 1679581782
transform 1 0 31488 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_329
timestamp 1679581782
transform 1 0 32160 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_336
timestamp 1679581782
transform 1 0 32832 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_343
timestamp 1679581782
transform 1 0 33504 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_350
timestamp 1679581782
transform 1 0 34176 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_357
timestamp 1679581782
transform 1 0 34848 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_364
timestamp 1679581782
transform 1 0 35520 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_371
timestamp 1679581782
transform 1 0 36192 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_378
timestamp 1679581782
transform 1 0 36864 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_385
timestamp 1679581782
transform 1 0 37536 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_392
timestamp 1679581782
transform 1 0 38208 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_399
timestamp 1679581782
transform 1 0 38880 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_406
timestamp 1679581782
transform 1 0 39552 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_413
timestamp 1679581782
transform 1 0 40224 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_420
timestamp 1679581782
transform 1 0 40896 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_427
timestamp 1679581782
transform 1 0 41568 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_434
timestamp 1679581782
transform 1 0 42240 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_441
timestamp 1679581782
transform 1 0 42912 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_448
timestamp 1679581782
transform 1 0 43584 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_455
timestamp 1679581782
transform 1 0 44256 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_462
timestamp 1679581782
transform 1 0 44928 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_469
timestamp 1679581782
transform 1 0 45600 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_476
timestamp 1679581782
transform 1 0 46272 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_483
timestamp 1679581782
transform 1 0 46944 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_490
timestamp 1679581782
transform 1 0 47616 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_497
timestamp 1679581782
transform 1 0 48288 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_504
timestamp 1679581782
transform 1 0 48960 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_511
timestamp 1679581782
transform 1 0 49632 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_518
timestamp 1679581782
transform 1 0 50304 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_525
timestamp 1679581782
transform 1 0 50976 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_532
timestamp 1679581782
transform 1 0 51648 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_539
timestamp 1679581782
transform 1 0 52320 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_546
timestamp 1679581782
transform 1 0 52992 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_553
timestamp 1679581782
transform 1 0 53664 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_560
timestamp 1679581782
transform 1 0 54336 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_567
timestamp 1679581782
transform 1 0 55008 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_574
timestamp 1679581782
transform 1 0 55680 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_581
timestamp 1679581782
transform 1 0 56352 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_588
timestamp 1679581782
transform 1 0 57024 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_595
timestamp 1679581782
transform 1 0 57696 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_602
timestamp 1679581782
transform 1 0 58368 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_609
timestamp 1679581782
transform 1 0 59040 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_616
timestamp 1679581782
transform 1 0 59712 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_623
timestamp 1679581782
transform 1 0 60384 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_630
timestamp 1679581782
transform 1 0 61056 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_637
timestamp 1679581782
transform 1 0 61728 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_644
timestamp 1679581782
transform 1 0 62400 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_651
timestamp 1679581782
transform 1 0 63072 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_658
timestamp 1679581782
transform 1 0 63744 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_665
timestamp 1679581782
transform 1 0 64416 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_672
timestamp 1679581782
transform 1 0 65088 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_679
timestamp 1679581782
transform 1 0 65760 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_686
timestamp 1679581782
transform 1 0 66432 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_693
timestamp 1679581782
transform 1 0 67104 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_700
timestamp 1679581782
transform 1 0 67776 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_707
timestamp 1679581782
transform 1 0 68448 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_714
timestamp 1679581782
transform 1 0 69120 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_721
timestamp 1679581782
transform 1 0 69792 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_728
timestamp 1679581782
transform 1 0 70464 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_735
timestamp 1679581782
transform 1 0 71136 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_742
timestamp 1679581782
transform 1 0 71808 0 -1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_749
timestamp 1679581782
transform 1 0 72480 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_764
timestamp 1677579658
transform 1 0 73920 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_777
timestamp 1677579658
transform 1 0 75168 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_782
timestamp 1677579658
transform 1 0 75648 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_799
timestamp 1677579658
transform 1 0 77280 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_828
timestamp 1677580104
transform 1 0 80064 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_970
timestamp 1677579658
transform 1 0 93696 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_983
timestamp 1677579658
transform 1 0 94944 0 -1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_1020
timestamp 1679581782
transform 1 0 98496 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_1027
timestamp 1677580104
transform 1 0 99168 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679581782
transform 1 0 1248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679581782
transform 1 0 1920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679581782
transform 1 0 2592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679581782
transform 1 0 3264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679581782
transform 1 0 3936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679581782
transform 1 0 4608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679581782
transform 1 0 5280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679581782
transform 1 0 5952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_63
timestamp 1679581782
transform 1 0 6624 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_70
timestamp 1679581782
transform 1 0 7296 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_77
timestamp 1679581782
transform 1 0 7968 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_84
timestamp 1679581782
transform 1 0 8640 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_91
timestamp 1679581782
transform 1 0 9312 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_98
timestamp 1679581782
transform 1 0 9984 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_105
timestamp 1679581782
transform 1 0 10656 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_112
timestamp 1679581782
transform 1 0 11328 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_119
timestamp 1679581782
transform 1 0 12000 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_126
timestamp 1679581782
transform 1 0 12672 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_133
timestamp 1679581782
transform 1 0 13344 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_140
timestamp 1679581782
transform 1 0 14016 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_147
timestamp 1679581782
transform 1 0 14688 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_154
timestamp 1679581782
transform 1 0 15360 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_161
timestamp 1679581782
transform 1 0 16032 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_168
timestamp 1679581782
transform 1 0 16704 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_175
timestamp 1679581782
transform 1 0 17376 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_182
timestamp 1679581782
transform 1 0 18048 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_189
timestamp 1679581782
transform 1 0 18720 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_196
timestamp 1679581782
transform 1 0 19392 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_203
timestamp 1679581782
transform 1 0 20064 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_210
timestamp 1679581782
transform 1 0 20736 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_217
timestamp 1679581782
transform 1 0 21408 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_224
timestamp 1679581782
transform 1 0 22080 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_231
timestamp 1679581782
transform 1 0 22752 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_238
timestamp 1679581782
transform 1 0 23424 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_245
timestamp 1679581782
transform 1 0 24096 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_252
timestamp 1679581782
transform 1 0 24768 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_259
timestamp 1679581782
transform 1 0 25440 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_266
timestamp 1679581782
transform 1 0 26112 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_273
timestamp 1679581782
transform 1 0 26784 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_280
timestamp 1679581782
transform 1 0 27456 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_287
timestamp 1679581782
transform 1 0 28128 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_294
timestamp 1679581782
transform 1 0 28800 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_301
timestamp 1679581782
transform 1 0 29472 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_308
timestamp 1679581782
transform 1 0 30144 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_315
timestamp 1679581782
transform 1 0 30816 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_322
timestamp 1679581782
transform 1 0 31488 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_329
timestamp 1679581782
transform 1 0 32160 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_336
timestamp 1679581782
transform 1 0 32832 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_343
timestamp 1679581782
transform 1 0 33504 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_350
timestamp 1679581782
transform 1 0 34176 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_357
timestamp 1679581782
transform 1 0 34848 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_364
timestamp 1679581782
transform 1 0 35520 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_371
timestamp 1679581782
transform 1 0 36192 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_378
timestamp 1679581782
transform 1 0 36864 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_385
timestamp 1679581782
transform 1 0 37536 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_392
timestamp 1679581782
transform 1 0 38208 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_399
timestamp 1679581782
transform 1 0 38880 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_406
timestamp 1679581782
transform 1 0 39552 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_413
timestamp 1679581782
transform 1 0 40224 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_420
timestamp 1679581782
transform 1 0 40896 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_427
timestamp 1679581782
transform 1 0 41568 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_434
timestamp 1679581782
transform 1 0 42240 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_441
timestamp 1679581782
transform 1 0 42912 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_448
timestamp 1679581782
transform 1 0 43584 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_455
timestamp 1679581782
transform 1 0 44256 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_462
timestamp 1679581782
transform 1 0 44928 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_469
timestamp 1679581782
transform 1 0 45600 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_476
timestamp 1679581782
transform 1 0 46272 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_483
timestamp 1679581782
transform 1 0 46944 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_490
timestamp 1679581782
transform 1 0 47616 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_497
timestamp 1679581782
transform 1 0 48288 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_504
timestamp 1679581782
transform 1 0 48960 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_511
timestamp 1679581782
transform 1 0 49632 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_518
timestamp 1679581782
transform 1 0 50304 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_525
timestamp 1679581782
transform 1 0 50976 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_532
timestamp 1679581782
transform 1 0 51648 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_539
timestamp 1679581782
transform 1 0 52320 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_546
timestamp 1679581782
transform 1 0 52992 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_553
timestamp 1679581782
transform 1 0 53664 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_560
timestamp 1679581782
transform 1 0 54336 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_567
timestamp 1679581782
transform 1 0 55008 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_574
timestamp 1679581782
transform 1 0 55680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_581
timestamp 1679581782
transform 1 0 56352 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_588
timestamp 1679581782
transform 1 0 57024 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_595
timestamp 1679581782
transform 1 0 57696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_602
timestamp 1679581782
transform 1 0 58368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_609
timestamp 1679581782
transform 1 0 59040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_616
timestamp 1679581782
transform 1 0 59712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_623
timestamp 1679581782
transform 1 0 60384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_630
timestamp 1679581782
transform 1 0 61056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_637
timestamp 1679581782
transform 1 0 61728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_644
timestamp 1679581782
transform 1 0 62400 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_651
timestamp 1679581782
transform 1 0 63072 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_658
timestamp 1679581782
transform 1 0 63744 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_665
timestamp 1679581782
transform 1 0 64416 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_672
timestamp 1679581782
transform 1 0 65088 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_679
timestamp 1679581782
transform 1 0 65760 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_686
timestamp 1679581782
transform 1 0 66432 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_693
timestamp 1679581782
transform 1 0 67104 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_700
timestamp 1679581782
transform 1 0 67776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_707
timestamp 1679581782
transform 1 0 68448 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_714
timestamp 1679581782
transform 1 0 69120 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_721
timestamp 1679581782
transform 1 0 69792 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_728
timestamp 1679581782
transform 1 0 70464 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_735
timestamp 1679581782
transform 1 0 71136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_742
timestamp 1679581782
transform 1 0 71808 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_749
timestamp 1679581782
transform 1 0 72480 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_756
timestamp 1679581782
transform 1 0 73152 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_763
timestamp 1679581782
transform 1 0 73824 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_770
timestamp 1679581782
transform 1 0 74496 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_777
timestamp 1679581782
transform 1 0 75168 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_784
timestamp 1679581782
transform 1 0 75840 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_791
timestamp 1679581782
transform 1 0 76512 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_798
timestamp 1679581782
transform 1 0 77184 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_805
timestamp 1679581782
transform 1 0 77856 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_812
timestamp 1679581782
transform 1 0 78528 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_819
timestamp 1679581782
transform 1 0 79200 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_826
timestamp 1679581782
transform 1 0 79872 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_833
timestamp 1679581782
transform 1 0 80544 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_840
timestamp 1679581782
transform 1 0 81216 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_847
timestamp 1679581782
transform 1 0 81888 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_854
timestamp 1679581782
transform 1 0 82560 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_861
timestamp 1679581782
transform 1 0 83232 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_868
timestamp 1679581782
transform 1 0 83904 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_875
timestamp 1679581782
transform 1 0 84576 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_882
timestamp 1679581782
transform 1 0 85248 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_889
timestamp 1679581782
transform 1 0 85920 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_896
timestamp 1679581782
transform 1 0 86592 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_903
timestamp 1679581782
transform 1 0 87264 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_910
timestamp 1679581782
transform 1 0 87936 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_917
timestamp 1679581782
transform 1 0 88608 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_924
timestamp 1679581782
transform 1 0 89280 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_931
timestamp 1679581782
transform 1 0 89952 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_938
timestamp 1679581782
transform 1 0 90624 0 1 34020
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_945
timestamp 1677579658
transform 1 0 91296 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_950
timestamp 1679581782
transform 1 0 91776 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_957
timestamp 1679581782
transform 1 0 92448 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_964
timestamp 1677580104
transform 1 0 93120 0 1 34020
box -48 -56 240 834
use sg13g2_decap_8  FILLER_44_970
timestamp 1679581782
transform 1 0 93696 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_977
timestamp 1679581782
transform 1 0 94368 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_984
timestamp 1679581782
transform 1 0 95040 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_991
timestamp 1679581782
transform 1 0 95712 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_998
timestamp 1679581782
transform 1 0 96384 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1005
timestamp 1679581782
transform 1 0 97056 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1012
timestamp 1679581782
transform 1 0 97728 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_1019
timestamp 1679581782
transform 1 0 98400 0 1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_44_1026
timestamp 1677580104
transform 1 0 99072 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_1028
timestamp 1677579658
transform 1 0 99264 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 1248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 1920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 2592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 3936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679581782
transform 1 0 4608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679581782
transform 1 0 5280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679581782
transform 1 0 5952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679581782
transform 1 0 6624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679581782
transform 1 0 7296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679581782
transform 1 0 7968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679581782
transform 1 0 8640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679581782
transform 1 0 9312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679581782
transform 1 0 9984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679581782
transform 1 0 10656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679581782
transform 1 0 11328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_119
timestamp 1679581782
transform 1 0 12000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_126
timestamp 1679581782
transform 1 0 12672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_133
timestamp 1679581782
transform 1 0 13344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_140
timestamp 1679581782
transform 1 0 14016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_147
timestamp 1679581782
transform 1 0 14688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_154
timestamp 1679581782
transform 1 0 15360 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_161
timestamp 1679581782
transform 1 0 16032 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_168
timestamp 1679581782
transform 1 0 16704 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_175
timestamp 1679581782
transform 1 0 17376 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_182
timestamp 1679581782
transform 1 0 18048 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_189
timestamp 1679581782
transform 1 0 18720 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_196
timestamp 1679581782
transform 1 0 19392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_203
timestamp 1679581782
transform 1 0 20064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_210
timestamp 1679581782
transform 1 0 20736 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_217
timestamp 1679581782
transform 1 0 21408 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_224
timestamp 1679581782
transform 1 0 22080 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_231
timestamp 1679581782
transform 1 0 22752 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_238
timestamp 1679581782
transform 1 0 23424 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_245
timestamp 1679581782
transform 1 0 24096 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_252
timestamp 1679581782
transform 1 0 24768 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_259
timestamp 1679581782
transform 1 0 25440 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_266
timestamp 1679581782
transform 1 0 26112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_273
timestamp 1679581782
transform 1 0 26784 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_280
timestamp 1679581782
transform 1 0 27456 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_287
timestamp 1679581782
transform 1 0 28128 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_294
timestamp 1679581782
transform 1 0 28800 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_301
timestamp 1679581782
transform 1 0 29472 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_308
timestamp 1679581782
transform 1 0 30144 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_315
timestamp 1679581782
transform 1 0 30816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_322
timestamp 1679581782
transform 1 0 31488 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_329
timestamp 1679581782
transform 1 0 32160 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_336
timestamp 1679581782
transform 1 0 32832 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_343
timestamp 1679581782
transform 1 0 33504 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_350
timestamp 1679581782
transform 1 0 34176 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_357
timestamp 1679581782
transform 1 0 34848 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_364
timestamp 1679581782
transform 1 0 35520 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_371
timestamp 1679581782
transform 1 0 36192 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_378
timestamp 1679581782
transform 1 0 36864 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_385
timestamp 1679581782
transform 1 0 37536 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_392
timestamp 1679581782
transform 1 0 38208 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_399
timestamp 1679581782
transform 1 0 38880 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_406
timestamp 1679581782
transform 1 0 39552 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_413
timestamp 1679581782
transform 1 0 40224 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_420
timestamp 1679581782
transform 1 0 40896 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_427
timestamp 1679581782
transform 1 0 41568 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_434
timestamp 1679581782
transform 1 0 42240 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_441
timestamp 1679581782
transform 1 0 42912 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_448
timestamp 1679581782
transform 1 0 43584 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_455
timestamp 1679581782
transform 1 0 44256 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_462
timestamp 1679581782
transform 1 0 44928 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_469
timestamp 1679581782
transform 1 0 45600 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_476
timestamp 1679581782
transform 1 0 46272 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_483
timestamp 1679581782
transform 1 0 46944 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_490
timestamp 1679581782
transform 1 0 47616 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_497
timestamp 1679581782
transform 1 0 48288 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_504
timestamp 1679581782
transform 1 0 48960 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_511
timestamp 1679581782
transform 1 0 49632 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_518
timestamp 1679581782
transform 1 0 50304 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_525
timestamp 1679581782
transform 1 0 50976 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_532
timestamp 1679581782
transform 1 0 51648 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_539
timestamp 1679581782
transform 1 0 52320 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_546
timestamp 1679581782
transform 1 0 52992 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_553
timestamp 1679581782
transform 1 0 53664 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_560
timestamp 1679581782
transform 1 0 54336 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_567
timestamp 1679581782
transform 1 0 55008 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_574
timestamp 1679581782
transform 1 0 55680 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_581
timestamp 1679581782
transform 1 0 56352 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_588
timestamp 1679581782
transform 1 0 57024 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_595
timestamp 1679581782
transform 1 0 57696 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_602
timestamp 1679581782
transform 1 0 58368 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_609
timestamp 1679581782
transform 1 0 59040 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_616
timestamp 1679581782
transform 1 0 59712 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_623
timestamp 1679581782
transform 1 0 60384 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_630
timestamp 1679581782
transform 1 0 61056 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_637
timestamp 1679581782
transform 1 0 61728 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_644
timestamp 1679581782
transform 1 0 62400 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_651
timestamp 1679581782
transform 1 0 63072 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_658
timestamp 1679581782
transform 1 0 63744 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_665
timestamp 1679581782
transform 1 0 64416 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_672
timestamp 1679581782
transform 1 0 65088 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_679
timestamp 1679581782
transform 1 0 65760 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_686
timestamp 1679581782
transform 1 0 66432 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_693
timestamp 1679581782
transform 1 0 67104 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_700
timestamp 1679581782
transform 1 0 67776 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_707
timestamp 1679581782
transform 1 0 68448 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_714
timestamp 1679581782
transform 1 0 69120 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_721
timestamp 1679581782
transform 1 0 69792 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_728
timestamp 1679581782
transform 1 0 70464 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_735
timestamp 1679581782
transform 1 0 71136 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_742
timestamp 1679581782
transform 1 0 71808 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_749
timestamp 1679581782
transform 1 0 72480 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_756
timestamp 1679581782
transform 1 0 73152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_763
timestamp 1679581782
transform 1 0 73824 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_770
timestamp 1679581782
transform 1 0 74496 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_777
timestamp 1679581782
transform 1 0 75168 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_784
timestamp 1679581782
transform 1 0 75840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_791
timestamp 1679581782
transform 1 0 76512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_798
timestamp 1679581782
transform 1 0 77184 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_805
timestamp 1679581782
transform 1 0 77856 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_812
timestamp 1679581782
transform 1 0 78528 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_819
timestamp 1679581782
transform 1 0 79200 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_826
timestamp 1679581782
transform 1 0 79872 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_833
timestamp 1679581782
transform 1 0 80544 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_840
timestamp 1679581782
transform 1 0 81216 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_847
timestamp 1679581782
transform 1 0 81888 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_854
timestamp 1679581782
transform 1 0 82560 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_861
timestamp 1679581782
transform 1 0 83232 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_868
timestamp 1679581782
transform 1 0 83904 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_875
timestamp 1679581782
transform 1 0 84576 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_882
timestamp 1679581782
transform 1 0 85248 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_889
timestamp 1679581782
transform 1 0 85920 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_896
timestamp 1679581782
transform 1 0 86592 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_903
timestamp 1679581782
transform 1 0 87264 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_910
timestamp 1679581782
transform 1 0 87936 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_917
timestamp 1679581782
transform 1 0 88608 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_924
timestamp 1679581782
transform 1 0 89280 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_931
timestamp 1679581782
transform 1 0 89952 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_938
timestamp 1679581782
transform 1 0 90624 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_945
timestamp 1679581782
transform 1 0 91296 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_952
timestamp 1679581782
transform 1 0 91968 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_959
timestamp 1679581782
transform 1 0 92640 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_966
timestamp 1679581782
transform 1 0 93312 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_973
timestamp 1679581782
transform 1 0 93984 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_980
timestamp 1679581782
transform 1 0 94656 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_987
timestamp 1679581782
transform 1 0 95328 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_994
timestamp 1679581782
transform 1 0 96000 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1001
timestamp 1679581782
transform 1 0 96672 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1008
timestamp 1679581782
transform 1 0 97344 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1015
timestamp 1679581782
transform 1 0 98016 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_1022
timestamp 1679581782
transform 1 0 98688 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 1248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 1920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 2592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 3264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 3936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 4608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 5280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 5952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 6624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 7296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 7968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 8640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 9312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 9984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 10656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 11328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679581782
transform 1 0 12000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679581782
transform 1 0 12672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679581782
transform 1 0 13344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679581782
transform 1 0 14016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679581782
transform 1 0 14688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679581782
transform 1 0 15360 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679581782
transform 1 0 16032 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679581782
transform 1 0 16704 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679581782
transform 1 0 17376 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_182
timestamp 1679581782
transform 1 0 18048 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_189
timestamp 1679581782
transform 1 0 18720 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_196
timestamp 1679581782
transform 1 0 19392 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679581782
transform 1 0 20064 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_210
timestamp 1679581782
transform 1 0 20736 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_217
timestamp 1679581782
transform 1 0 21408 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679581782
transform 1 0 22080 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679581782
transform 1 0 22752 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679581782
transform 1 0 23424 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679581782
transform 1 0 24096 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679581782
transform 1 0 24768 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679581782
transform 1 0 25440 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_266
timestamp 1679581782
transform 1 0 26112 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_273
timestamp 1679581782
transform 1 0 26784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_280
timestamp 1679581782
transform 1 0 27456 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679581782
transform 1 0 28128 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679581782
transform 1 0 28800 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679581782
transform 1 0 29472 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679581782
transform 1 0 30144 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_315
timestamp 1679581782
transform 1 0 30816 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_322
timestamp 1679581782
transform 1 0 31488 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_329
timestamp 1679581782
transform 1 0 32160 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_336
timestamp 1679581782
transform 1 0 32832 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_343
timestamp 1679581782
transform 1 0 33504 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_350
timestamp 1679581782
transform 1 0 34176 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_357
timestamp 1679581782
transform 1 0 34848 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_364
timestamp 1679581782
transform 1 0 35520 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_371
timestamp 1679581782
transform 1 0 36192 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_378
timestamp 1679581782
transform 1 0 36864 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_385
timestamp 1679581782
transform 1 0 37536 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_392
timestamp 1679581782
transform 1 0 38208 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_399
timestamp 1679581782
transform 1 0 38880 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_406
timestamp 1679581782
transform 1 0 39552 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_413
timestamp 1679581782
transform 1 0 40224 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_420
timestamp 1679581782
transform 1 0 40896 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679581782
transform 1 0 41568 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679581782
transform 1 0 42240 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679581782
transform 1 0 42912 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679581782
transform 1 0 43584 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679581782
transform 1 0 44256 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679581782
transform 1 0 44928 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679581782
transform 1 0 45600 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679581782
transform 1 0 46272 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679581782
transform 1 0 46944 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679581782
transform 1 0 47616 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_497
timestamp 1679581782
transform 1 0 48288 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_504
timestamp 1679581782
transform 1 0 48960 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_511
timestamp 1679581782
transform 1 0 49632 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_518
timestamp 1679581782
transform 1 0 50304 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_525
timestamp 1679581782
transform 1 0 50976 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_532
timestamp 1679581782
transform 1 0 51648 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_539
timestamp 1679581782
transform 1 0 52320 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_546
timestamp 1679581782
transform 1 0 52992 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_553
timestamp 1679581782
transform 1 0 53664 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_560
timestamp 1679581782
transform 1 0 54336 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_567
timestamp 1679581782
transform 1 0 55008 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_574
timestamp 1679581782
transform 1 0 55680 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_581
timestamp 1679581782
transform 1 0 56352 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_588
timestamp 1679581782
transform 1 0 57024 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_595
timestamp 1679581782
transform 1 0 57696 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_602
timestamp 1679581782
transform 1 0 58368 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_609
timestamp 1679581782
transform 1 0 59040 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_616
timestamp 1679581782
transform 1 0 59712 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_623
timestamp 1679581782
transform 1 0 60384 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_630
timestamp 1679581782
transform 1 0 61056 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_637
timestamp 1679581782
transform 1 0 61728 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_644
timestamp 1679581782
transform 1 0 62400 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_651
timestamp 1679581782
transform 1 0 63072 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_658
timestamp 1679581782
transform 1 0 63744 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_665
timestamp 1679581782
transform 1 0 64416 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_672
timestamp 1679581782
transform 1 0 65088 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_679
timestamp 1679581782
transform 1 0 65760 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_686
timestamp 1679581782
transform 1 0 66432 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_693
timestamp 1679581782
transform 1 0 67104 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_700
timestamp 1679581782
transform 1 0 67776 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_707
timestamp 1679581782
transform 1 0 68448 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_714
timestamp 1679581782
transform 1 0 69120 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_721
timestamp 1679581782
transform 1 0 69792 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_728
timestamp 1679581782
transform 1 0 70464 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_735
timestamp 1679581782
transform 1 0 71136 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_742
timestamp 1679581782
transform 1 0 71808 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_749
timestamp 1679581782
transform 1 0 72480 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_756
timestamp 1679581782
transform 1 0 73152 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_763
timestamp 1679581782
transform 1 0 73824 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_770
timestamp 1679581782
transform 1 0 74496 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_777
timestamp 1679581782
transform 1 0 75168 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_784
timestamp 1679581782
transform 1 0 75840 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_791
timestamp 1679581782
transform 1 0 76512 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_798
timestamp 1679581782
transform 1 0 77184 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_805
timestamp 1679581782
transform 1 0 77856 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_812
timestamp 1679581782
transform 1 0 78528 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_819
timestamp 1679581782
transform 1 0 79200 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_826
timestamp 1679581782
transform 1 0 79872 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_833
timestamp 1679581782
transform 1 0 80544 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_840
timestamp 1679581782
transform 1 0 81216 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_847
timestamp 1679581782
transform 1 0 81888 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_854
timestamp 1679581782
transform 1 0 82560 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_861
timestamp 1679581782
transform 1 0 83232 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_868
timestamp 1679581782
transform 1 0 83904 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_875
timestamp 1679581782
transform 1 0 84576 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_882
timestamp 1679581782
transform 1 0 85248 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_889
timestamp 1679581782
transform 1 0 85920 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_896
timestamp 1679581782
transform 1 0 86592 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_903
timestamp 1679581782
transform 1 0 87264 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_910
timestamp 1679581782
transform 1 0 87936 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_917
timestamp 1679581782
transform 1 0 88608 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_924
timestamp 1679581782
transform 1 0 89280 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_931
timestamp 1679581782
transform 1 0 89952 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_938
timestamp 1679581782
transform 1 0 90624 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_945
timestamp 1679581782
transform 1 0 91296 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_952
timestamp 1679581782
transform 1 0 91968 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_959
timestamp 1679581782
transform 1 0 92640 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_966
timestamp 1679581782
transform 1 0 93312 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_973
timestamp 1679581782
transform 1 0 93984 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_980
timestamp 1679581782
transform 1 0 94656 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_987
timestamp 1679581782
transform 1 0 95328 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_994
timestamp 1679581782
transform 1 0 96000 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1001
timestamp 1679581782
transform 1 0 96672 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1008
timestamp 1679581782
transform 1 0 97344 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1015
timestamp 1679581782
transform 1 0 98016 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_1022
timestamp 1679581782
transform 1 0 98688 0 1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 1248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 1920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 2592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 3264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 3936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 4608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 5280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 5952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 6624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 7296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 7968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 8640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 9312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 9984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 10656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 11328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 12000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 12672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 13344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 14688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 15360 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 16032 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 16704 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 17376 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679581782
transform 1 0 18048 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679581782
transform 1 0 18720 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679581782
transform 1 0 19392 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679581782
transform 1 0 20064 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679581782
transform 1 0 20736 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679581782
transform 1 0 21408 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679581782
transform 1 0 22080 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679581782
transform 1 0 22752 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679581782
transform 1 0 23424 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679581782
transform 1 0 24096 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679581782
transform 1 0 24768 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679581782
transform 1 0 25440 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679581782
transform 1 0 26112 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679581782
transform 1 0 26784 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679581782
transform 1 0 27456 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679581782
transform 1 0 28128 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679581782
transform 1 0 28800 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679581782
transform 1 0 29472 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679581782
transform 1 0 30144 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679581782
transform 1 0 30816 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679581782
transform 1 0 31488 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679581782
transform 1 0 32160 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679581782
transform 1 0 32832 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679581782
transform 1 0 33504 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679581782
transform 1 0 34176 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679581782
transform 1 0 34848 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679581782
transform 1 0 35520 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679581782
transform 1 0 36192 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679581782
transform 1 0 36864 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679581782
transform 1 0 37536 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679581782
transform 1 0 38208 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679581782
transform 1 0 38880 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679581782
transform 1 0 39552 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679581782
transform 1 0 40224 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679581782
transform 1 0 40896 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679581782
transform 1 0 41568 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679581782
transform 1 0 42240 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679581782
transform 1 0 42912 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 43584 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679581782
transform 1 0 44256 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679581782
transform 1 0 44928 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 45600 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 46272 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 46944 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 47616 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 48288 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 48960 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 49632 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 50304 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 50976 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 51648 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679581782
transform 1 0 52320 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679581782
transform 1 0 52992 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679581782
transform 1 0 53664 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679581782
transform 1 0 54336 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679581782
transform 1 0 55008 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679581782
transform 1 0 55680 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679581782
transform 1 0 56352 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679581782
transform 1 0 57024 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679581782
transform 1 0 57696 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679581782
transform 1 0 58368 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679581782
transform 1 0 59040 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679581782
transform 1 0 59712 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679581782
transform 1 0 60384 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679581782
transform 1 0 61056 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679581782
transform 1 0 61728 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679581782
transform 1 0 62400 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679581782
transform 1 0 63072 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679581782
transform 1 0 63744 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679581782
transform 1 0 64416 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679581782
transform 1 0 65088 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679581782
transform 1 0 65760 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679581782
transform 1 0 66432 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679581782
transform 1 0 67104 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679581782
transform 1 0 67776 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679581782
transform 1 0 68448 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679581782
transform 1 0 69120 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679581782
transform 1 0 69792 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679581782
transform 1 0 70464 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679581782
transform 1 0 71136 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679581782
transform 1 0 71808 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679581782
transform 1 0 72480 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_756
timestamp 1679581782
transform 1 0 73152 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_763
timestamp 1679581782
transform 1 0 73824 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_770
timestamp 1679581782
transform 1 0 74496 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_777
timestamp 1679581782
transform 1 0 75168 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_784
timestamp 1679581782
transform 1 0 75840 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_791
timestamp 1679581782
transform 1 0 76512 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_798
timestamp 1679581782
transform 1 0 77184 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_805
timestamp 1679581782
transform 1 0 77856 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_812
timestamp 1679581782
transform 1 0 78528 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_819
timestamp 1679581782
transform 1 0 79200 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_826
timestamp 1679581782
transform 1 0 79872 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_833
timestamp 1679581782
transform 1 0 80544 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_840
timestamp 1679581782
transform 1 0 81216 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_847
timestamp 1679581782
transform 1 0 81888 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_854
timestamp 1679581782
transform 1 0 82560 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_861
timestamp 1679581782
transform 1 0 83232 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_868
timestamp 1679581782
transform 1 0 83904 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_875
timestamp 1679581782
transform 1 0 84576 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_882
timestamp 1679581782
transform 1 0 85248 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_889
timestamp 1679581782
transform 1 0 85920 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_896
timestamp 1679581782
transform 1 0 86592 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_903
timestamp 1679581782
transform 1 0 87264 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_910
timestamp 1679581782
transform 1 0 87936 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_917
timestamp 1679581782
transform 1 0 88608 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_924
timestamp 1679581782
transform 1 0 89280 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_931
timestamp 1679581782
transform 1 0 89952 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_938
timestamp 1679581782
transform 1 0 90624 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_945
timestamp 1679581782
transform 1 0 91296 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_952
timestamp 1679581782
transform 1 0 91968 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_959
timestamp 1679581782
transform 1 0 92640 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_966
timestamp 1679581782
transform 1 0 93312 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_973
timestamp 1679581782
transform 1 0 93984 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_980
timestamp 1679581782
transform 1 0 94656 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_987
timestamp 1679581782
transform 1 0 95328 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_994
timestamp 1679581782
transform 1 0 96000 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1001
timestamp 1679581782
transform 1 0 96672 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1008
timestamp 1679581782
transform 1 0 97344 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1015
timestamp 1679581782
transform 1 0 98016 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_1022
timestamp 1679581782
transform 1 0 98688 0 -1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 1248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 1920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 2592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 3264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 3936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 4608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 5280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 5952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 6624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 7296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 7968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 8640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 9312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 9984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 10656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 11328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 12000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 12672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 13344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 14016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 14688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 15360 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 16032 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 16704 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 17376 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 18048 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 18720 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 19392 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 20064 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 20736 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 21408 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 22080 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 22752 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 23424 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 24096 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 24768 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 25440 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 26112 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 26784 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679581782
transform 1 0 27456 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 28128 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 28800 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 29472 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 30144 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679581782
transform 1 0 30816 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679581782
transform 1 0 31488 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679581782
transform 1 0 32160 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679581782
transform 1 0 32832 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679581782
transform 1 0 33504 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679581782
transform 1 0 34176 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679581782
transform 1 0 34848 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679581782
transform 1 0 35520 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679581782
transform 1 0 36192 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679581782
transform 1 0 36864 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679581782
transform 1 0 37536 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679581782
transform 1 0 38208 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679581782
transform 1 0 38880 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679581782
transform 1 0 39552 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679581782
transform 1 0 40224 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679581782
transform 1 0 40896 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679581782
transform 1 0 41568 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679581782
transform 1 0 42240 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679581782
transform 1 0 42912 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679581782
transform 1 0 43584 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679581782
transform 1 0 44256 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679581782
transform 1 0 44928 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679581782
transform 1 0 45600 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679581782
transform 1 0 46272 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679581782
transform 1 0 46944 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679581782
transform 1 0 47616 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679581782
transform 1 0 48288 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679581782
transform 1 0 48960 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679581782
transform 1 0 49632 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679581782
transform 1 0 50304 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679581782
transform 1 0 50976 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679581782
transform 1 0 51648 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679581782
transform 1 0 52320 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679581782
transform 1 0 52992 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679581782
transform 1 0 53664 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679581782
transform 1 0 54336 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_567
timestamp 1679581782
transform 1 0 55008 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_574
timestamp 1679581782
transform 1 0 55680 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_581
timestamp 1679581782
transform 1 0 56352 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_588
timestamp 1679581782
transform 1 0 57024 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_595
timestamp 1679581782
transform 1 0 57696 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_602
timestamp 1679581782
transform 1 0 58368 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_609
timestamp 1679581782
transform 1 0 59040 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_616
timestamp 1679581782
transform 1 0 59712 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_623
timestamp 1679581782
transform 1 0 60384 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_630
timestamp 1679581782
transform 1 0 61056 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_637
timestamp 1679581782
transform 1 0 61728 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_644
timestamp 1679581782
transform 1 0 62400 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_651
timestamp 1679581782
transform 1 0 63072 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_658
timestamp 1679581782
transform 1 0 63744 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_665
timestamp 1679581782
transform 1 0 64416 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_672
timestamp 1679581782
transform 1 0 65088 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_679
timestamp 1679581782
transform 1 0 65760 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_686
timestamp 1679581782
transform 1 0 66432 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_693
timestamp 1679581782
transform 1 0 67104 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_700
timestamp 1679581782
transform 1 0 67776 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_707
timestamp 1679581782
transform 1 0 68448 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_714
timestamp 1679581782
transform 1 0 69120 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_721
timestamp 1679581782
transform 1 0 69792 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_728
timestamp 1679581782
transform 1 0 70464 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_735
timestamp 1679581782
transform 1 0 71136 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_742
timestamp 1679581782
transform 1 0 71808 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_749
timestamp 1679581782
transform 1 0 72480 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_756
timestamp 1679581782
transform 1 0 73152 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_763
timestamp 1679581782
transform 1 0 73824 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_770
timestamp 1679581782
transform 1 0 74496 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_777
timestamp 1679581782
transform 1 0 75168 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_784
timestamp 1679581782
transform 1 0 75840 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_791
timestamp 1679581782
transform 1 0 76512 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_798
timestamp 1679581782
transform 1 0 77184 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_805
timestamp 1679581782
transform 1 0 77856 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_812
timestamp 1679581782
transform 1 0 78528 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_819
timestamp 1679581782
transform 1 0 79200 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_826
timestamp 1679581782
transform 1 0 79872 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_833
timestamp 1679581782
transform 1 0 80544 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_840
timestamp 1679581782
transform 1 0 81216 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_847
timestamp 1679581782
transform 1 0 81888 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_854
timestamp 1679581782
transform 1 0 82560 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_861
timestamp 1679581782
transform 1 0 83232 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_868
timestamp 1679581782
transform 1 0 83904 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_875
timestamp 1679581782
transform 1 0 84576 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_882
timestamp 1679581782
transform 1 0 85248 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_889
timestamp 1679581782
transform 1 0 85920 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_896
timestamp 1679581782
transform 1 0 86592 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_903
timestamp 1679581782
transform 1 0 87264 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_910
timestamp 1679581782
transform 1 0 87936 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_917
timestamp 1679581782
transform 1 0 88608 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_924
timestamp 1679581782
transform 1 0 89280 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_931
timestamp 1679581782
transform 1 0 89952 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_938
timestamp 1679581782
transform 1 0 90624 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_945
timestamp 1679581782
transform 1 0 91296 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_952
timestamp 1679581782
transform 1 0 91968 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_959
timestamp 1679581782
transform 1 0 92640 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_966
timestamp 1679581782
transform 1 0 93312 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_973
timestamp 1679581782
transform 1 0 93984 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_980
timestamp 1679581782
transform 1 0 94656 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_987
timestamp 1679581782
transform 1 0 95328 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_994
timestamp 1679581782
transform 1 0 96000 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1001
timestamp 1679581782
transform 1 0 96672 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1008
timestamp 1679581782
transform 1 0 97344 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1015
timestamp 1679581782
transform 1 0 98016 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_1022
timestamp 1679581782
transform 1 0 98688 0 1 37044
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_0
timestamp 1679581782
transform 1 0 576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_7
timestamp 1679581782
transform 1 0 1248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_14
timestamp 1679581782
transform 1 0 1920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679581782
transform 1 0 2592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_28
timestamp 1679581782
transform 1 0 3264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_35
timestamp 1679581782
transform 1 0 3936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_42
timestamp 1679581782
transform 1 0 4608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_49
timestamp 1679581782
transform 1 0 5280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_56
timestamp 1679581782
transform 1 0 5952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_63
timestamp 1679581782
transform 1 0 6624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_70
timestamp 1679581782
transform 1 0 7296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_77
timestamp 1679581782
transform 1 0 7968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_84
timestamp 1679581782
transform 1 0 8640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_91
timestamp 1679581782
transform 1 0 9312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_98
timestamp 1679581782
transform 1 0 9984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_105
timestamp 1679581782
transform 1 0 10656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_112
timestamp 1679581782
transform 1 0 11328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_119
timestamp 1679581782
transform 1 0 12000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_126
timestamp 1679581782
transform 1 0 12672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_133
timestamp 1679581782
transform 1 0 13344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_140
timestamp 1679581782
transform 1 0 14016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_147
timestamp 1679581782
transform 1 0 14688 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_154
timestamp 1679581782
transform 1 0 15360 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_161
timestamp 1679581782
transform 1 0 16032 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_168
timestamp 1679581782
transform 1 0 16704 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_175
timestamp 1679581782
transform 1 0 17376 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_182
timestamp 1679581782
transform 1 0 18048 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_189
timestamp 1679581782
transform 1 0 18720 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_196
timestamp 1679581782
transform 1 0 19392 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_203
timestamp 1679581782
transform 1 0 20064 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_210
timestamp 1679581782
transform 1 0 20736 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_217
timestamp 1679581782
transform 1 0 21408 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_224
timestamp 1679581782
transform 1 0 22080 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_231
timestamp 1679581782
transform 1 0 22752 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_238
timestamp 1679581782
transform 1 0 23424 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_245
timestamp 1679581782
transform 1 0 24096 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_252
timestamp 1679581782
transform 1 0 24768 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_259
timestamp 1679581782
transform 1 0 25440 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_266
timestamp 1679581782
transform 1 0 26112 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_273
timestamp 1679581782
transform 1 0 26784 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_280
timestamp 1679581782
transform 1 0 27456 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_287
timestamp 1679581782
transform 1 0 28128 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_294
timestamp 1679581782
transform 1 0 28800 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_301
timestamp 1679581782
transform 1 0 29472 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_308
timestamp 1679581782
transform 1 0 30144 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_315
timestamp 1679581782
transform 1 0 30816 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_322
timestamp 1679581782
transform 1 0 31488 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_329
timestamp 1679581782
transform 1 0 32160 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_336
timestamp 1679581782
transform 1 0 32832 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_343
timestamp 1679581782
transform 1 0 33504 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_350
timestamp 1679581782
transform 1 0 34176 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_357
timestamp 1679581782
transform 1 0 34848 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_364
timestamp 1679581782
transform 1 0 35520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_371
timestamp 1679581782
transform 1 0 36192 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_378
timestamp 1679581782
transform 1 0 36864 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_385
timestamp 1679581782
transform 1 0 37536 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_392
timestamp 1679581782
transform 1 0 38208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_399
timestamp 1679581782
transform 1 0 38880 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_406
timestamp 1679581782
transform 1 0 39552 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_413
timestamp 1679581782
transform 1 0 40224 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_420
timestamp 1679581782
transform 1 0 40896 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_427
timestamp 1679581782
transform 1 0 41568 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_434
timestamp 1679581782
transform 1 0 42240 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_441
timestamp 1679581782
transform 1 0 42912 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_448
timestamp 1679581782
transform 1 0 43584 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_455
timestamp 1679581782
transform 1 0 44256 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_462
timestamp 1679581782
transform 1 0 44928 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_469
timestamp 1679581782
transform 1 0 45600 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_476
timestamp 1679581782
transform 1 0 46272 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_483
timestamp 1679581782
transform 1 0 46944 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_490
timestamp 1679581782
transform 1 0 47616 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_497
timestamp 1679581782
transform 1 0 48288 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_504
timestamp 1679581782
transform 1 0 48960 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_511
timestamp 1679581782
transform 1 0 49632 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_518
timestamp 1679581782
transform 1 0 50304 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_525
timestamp 1679581782
transform 1 0 50976 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_532
timestamp 1679581782
transform 1 0 51648 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_539
timestamp 1679581782
transform 1 0 52320 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_546
timestamp 1679581782
transform 1 0 52992 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_553
timestamp 1679581782
transform 1 0 53664 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_560
timestamp 1679581782
transform 1 0 54336 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_567
timestamp 1679581782
transform 1 0 55008 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_574
timestamp 1679581782
transform 1 0 55680 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_581
timestamp 1679581782
transform 1 0 56352 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_588
timestamp 1679581782
transform 1 0 57024 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_595
timestamp 1679581782
transform 1 0 57696 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_602
timestamp 1679581782
transform 1 0 58368 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_609
timestamp 1679581782
transform 1 0 59040 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_616
timestamp 1679581782
transform 1 0 59712 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_623
timestamp 1679581782
transform 1 0 60384 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_630
timestamp 1679581782
transform 1 0 61056 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_637
timestamp 1679581782
transform 1 0 61728 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_644
timestamp 1679581782
transform 1 0 62400 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_651
timestamp 1679581782
transform 1 0 63072 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_658
timestamp 1679581782
transform 1 0 63744 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_665
timestamp 1679581782
transform 1 0 64416 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_672
timestamp 1679581782
transform 1 0 65088 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_679
timestamp 1679581782
transform 1 0 65760 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_686
timestamp 1679581782
transform 1 0 66432 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_693
timestamp 1679581782
transform 1 0 67104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_700
timestamp 1679581782
transform 1 0 67776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_707
timestamp 1679581782
transform 1 0 68448 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_714
timestamp 1679581782
transform 1 0 69120 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_721
timestamp 1679581782
transform 1 0 69792 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_728
timestamp 1679581782
transform 1 0 70464 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_735
timestamp 1679581782
transform 1 0 71136 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_742
timestamp 1679581782
transform 1 0 71808 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_749
timestamp 1679581782
transform 1 0 72480 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_756
timestamp 1679581782
transform 1 0 73152 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_763
timestamp 1679581782
transform 1 0 73824 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_770
timestamp 1679581782
transform 1 0 74496 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_777
timestamp 1679581782
transform 1 0 75168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_784
timestamp 1679581782
transform 1 0 75840 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_791
timestamp 1679581782
transform 1 0 76512 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_798
timestamp 1679581782
transform 1 0 77184 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_805
timestamp 1679581782
transform 1 0 77856 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_812
timestamp 1679581782
transform 1 0 78528 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_819
timestamp 1679581782
transform 1 0 79200 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_826
timestamp 1679581782
transform 1 0 79872 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_833
timestamp 1679581782
transform 1 0 80544 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_840
timestamp 1679581782
transform 1 0 81216 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_847
timestamp 1679581782
transform 1 0 81888 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_854
timestamp 1679581782
transform 1 0 82560 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_861
timestamp 1679581782
transform 1 0 83232 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_868
timestamp 1679581782
transform 1 0 83904 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_875
timestamp 1679581782
transform 1 0 84576 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_882
timestamp 1679581782
transform 1 0 85248 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_889
timestamp 1679581782
transform 1 0 85920 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_896
timestamp 1679581782
transform 1 0 86592 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_903
timestamp 1679581782
transform 1 0 87264 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_910
timestamp 1679581782
transform 1 0 87936 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_917
timestamp 1679581782
transform 1 0 88608 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_924
timestamp 1679581782
transform 1 0 89280 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_931
timestamp 1679581782
transform 1 0 89952 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_938
timestamp 1679581782
transform 1 0 90624 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_945
timestamp 1679581782
transform 1 0 91296 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_952
timestamp 1679581782
transform 1 0 91968 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_959
timestamp 1679581782
transform 1 0 92640 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_966
timestamp 1679581782
transform 1 0 93312 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_973
timestamp 1679581782
transform 1 0 93984 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_980
timestamp 1679581782
transform 1 0 94656 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_987
timestamp 1679581782
transform 1 0 95328 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_994
timestamp 1679581782
transform 1 0 96000 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1001
timestamp 1679581782
transform 1 0 96672 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1008
timestamp 1679581782
transform 1 0 97344 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1015
timestamp 1679581782
transform 1 0 98016 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_1022
timestamp 1679581782
transform 1 0 98688 0 -1 38556
box -48 -56 720 834
use sg13g2_tiehi  heichips25_pudding_113
timestamp 1680000651
transform -1 0 960 0 1 15876
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_114
timestamp 1680000651
transform -1 0 960 0 -1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_115
timestamp 1680000651
transform -1 0 960 0 1 17388
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_116
timestamp 1680000651
transform -1 0 960 0 -1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_117
timestamp 1680000651
transform -1 0 960 0 1 18900
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_118
timestamp 1680000651
transform -1 0 960 0 -1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_119
timestamp 1680000651
transform -1 0 960 0 1 20412
box -48 -56 432 834
use sg13g2_tiehi  heichips25_pudding_120
timestamp 1680000651
transform -1 0 960 0 1 21924
box -48 -56 432 834
use sg13g2_buf_2  input1
timestamp 1676381867
transform -1 0 1056 0 -1 23436
box -48 -56 528 834
use sg13g2_buf_2  input2
timestamp 1676381867
transform -1 0 1056 0 1 23436
box -48 -56 528 834
use sg13g2_buf_2  input3
timestamp 1676381867
transform -1 0 1056 0 -1 24948
box -48 -56 528 834
use sg13g2_buf_2  input4
timestamp 1676381867
transform -1 0 1056 0 1 24948
box -48 -56 528 834
use sg13g2_buf_1  output5
timestamp 1676381911
transform -1 0 960 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  output6
timestamp 1676381911
transform -1 0 960 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  output7
timestamp 1676381911
transform -1 0 960 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  output8
timestamp 1676381911
transform -1 0 960 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  output9
timestamp 1676381911
transform -1 0 960 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  output10
timestamp 1676381911
transform -1 0 960 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  output11
timestamp 1676381911
transform -1 0 960 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  output12
timestamp 1676381911
transform -1 0 960 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  output13
timestamp 1676381911
transform -1 0 960 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  output14
timestamp 1676381911
transform -1 0 960 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  output15
timestamp 1676381911
transform -1 0 1344 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output16
timestamp 1676381911
transform -1 0 960 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  output17
timestamp 1676381911
transform -1 0 960 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  output18
timestamp 1676381911
transform -1 0 960 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  output19
timestamp 1676381911
transform -1 0 960 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  output20
timestamp 1676381911
transform -1 0 960 0 1 8316
box -48 -56 432 834
<< labels >>
flabel metal6 s 4316 630 4756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 8316 630 8756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 12316 630 12756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 16316 630 16756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 20316 630 20756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 24316 630 24756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 28316 630 28756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 32316 630 32756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 36316 630 36756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 40316 630 40756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 44316 630 44756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 48316 630 48756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 52316 630 52756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 56316 630 56756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 60316 630 60756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 64316 630 64756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 68316 630 68756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 72316 630 72756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 76316 630 76756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 80316 630 80756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 84316 630 84756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 88316 630 88756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 92316 630 92756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 96316 630 96756 38682 0 FreeSans 2624 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 4496 99404 4936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 8496 99404 8936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 12496 99404 12936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 16496 99404 16936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 20496 99404 20936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 24496 99404 24936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 28496 99404 28936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 32496 99404 32936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal7 s 532 36496 99404 36936 0 FreeSans 3200 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal6 s 3076 712 3516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 7076 712 7516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 11076 712 11516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 15076 712 15516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 19076 712 19516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 23076 712 23516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 27076 712 27516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 31076 712 31516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 35076 712 35516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 39076 712 39516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 43076 712 43516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 47076 712 47516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 51076 712 51516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 55076 712 55516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 59076 712 59516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 63076 712 63516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 67076 712 67516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 71076 712 71516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 75076 712 75516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 79076 712 79516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 83076 712 83516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 87076 712 87516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 91076 712 91516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 95076 712 95516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal6 s 99076 712 99516 38600 0 FreeSans 2624 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 3256 99516 3696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 7256 99516 7696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 11256 99516 11696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 15256 99516 15696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 19256 99516 19696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 23256 99516 23696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 27256 99516 27696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 31256 99516 31696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal7 s 532 35256 99516 35696 0 FreeSans 3200 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 35828 80 35908 0 FreeSans 320 0 0 0 ena
port 3 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 rst_n
port 4 nsew signal input
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 ui_in[0]
port 5 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 ui_in[1]
port 6 nsew signal input
flabel metal3 s 0 24068 80 24148 0 FreeSans 320 0 0 0 ui_in[2]
port 7 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 ui_in[3]
port 8 nsew signal input
flabel metal3 s 0 25748 80 25828 0 FreeSans 320 0 0 0 ui_in[4]
port 9 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 ui_in[5]
port 10 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 ui_in[6]
port 11 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 ui_in[7]
port 12 nsew signal input
flabel metal3 s 0 29108 80 29188 0 FreeSans 320 0 0 0 uio_in[0]
port 13 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 uio_in[1]
port 14 nsew signal input
flabel metal3 s 0 30788 80 30868 0 FreeSans 320 0 0 0 uio_in[2]
port 15 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 uio_in[3]
port 16 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 uio_in[4]
port 17 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 uio_in[5]
port 18 nsew signal input
flabel metal3 s 0 34148 80 34228 0 FreeSans 320 0 0 0 uio_in[6]
port 19 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 uio_in[7]
port 20 nsew signal input
flabel metal3 s 0 15668 80 15748 0 FreeSans 320 0 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal3 s 0 19028 80 19108 0 FreeSans 320 0 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 20708 80 20788 0 FreeSans 320 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal3 s 0 8948 80 9028 0 FreeSans 320 0 0 0 uio_out[0]
port 29 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 uio_out[1]
port 30 nsew signal output
flabel metal3 s 0 10628 80 10708 0 FreeSans 320 0 0 0 uio_out[2]
port 31 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 uio_out[5]
port 34 nsew signal output
flabel metal3 s 0 13988 80 14068 0 FreeSans 320 0 0 0 uio_out[6]
port 35 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 uio_out[7]
port 36 nsew signal output
flabel metal3 s 0 2228 80 2308 0 FreeSans 320 0 0 0 uo_out[0]
port 37 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 uo_out[1]
port 38 nsew signal output
flabel metal3 s 0 3908 80 3988 0 FreeSans 320 0 0 0 uo_out[2]
port 39 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 uo_out[3]
port 40 nsew signal output
flabel metal3 s 0 5588 80 5668 0 FreeSans 320 0 0 0 uo_out[4]
port 41 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 uo_out[5]
port 42 nsew signal output
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 uo_out[6]
port 43 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 uo_out[7]
port 44 nsew signal output
rlabel via6 96536 12716 96536 12716 0 VGND
rlabel via6 95296 11476 95296 11476 0 VPWR
rlabel metal3 71952 26292 71952 26292 0 digitalH.g\[0\].u.OUTN
rlabel metal2 71328 26586 71328 26586 0 digitalH.g\[0\].u.OUTP
rlabel metal2 83525 32140 83525 32140 0 digitalH.g\[100\].u.OUTN
rlabel metal2 83760 33432 83760 33432 0 digitalH.g\[100\].u.OUTP
rlabel metal3 83472 32844 83472 32844 0 digitalH.g\[101\].u.OUTN
rlabel metal2 83235 32014 83235 32014 0 digitalH.g\[101\].u.OUTP
rlabel metal3 83136 32928 83136 32928 0 digitalH.g\[102\].u.OUTN
rlabel metal2 82835 32056 82835 32056 0 digitalH.g\[102\].u.OUTP
rlabel metal2 82325 32140 82325 32140 0 digitalH.g\[103\].u.OUTN
rlabel metal2 82560 33432 82560 33432 0 digitalH.g\[103\].u.OUTP
rlabel metal2 81925 32014 81925 32014 0 digitalH.g\[104\].u.OUTN
rlabel metal2 81888 32466 81888 32466 0 digitalH.g\[104\].u.OUTP
rlabel metal3 82032 32844 82032 32844 0 digitalH.g\[105\].u.OUTN
rlabel metal2 81840 33432 81840 33432 0 digitalH.g\[105\].u.OUTP
rlabel metal2 81125 32098 81125 32098 0 digitalH.g\[106\].u.OUTN
rlabel metal2 81312 33096 81312 33096 0 digitalH.g\[106\].u.OUTP
rlabel metal2 80725 32140 80725 32140 0 digitalH.g\[107\].u.OUTN
rlabel metal2 80832 32382 80832 32382 0 digitalH.g\[107\].u.OUTP
rlabel metal3 80640 32844 80640 32844 0 digitalH.g\[108\].u.OUTN
rlabel metal2 80736 33096 80736 33096 0 digitalH.g\[108\].u.OUTP
rlabel metal2 79925 32014 79925 32014 0 digitalH.g\[109\].u.OUTN
rlabel metal2 79920 33432 79920 33432 0 digitalH.g\[109\].u.OUTP
rlabel metal2 76800 25956 76800 25956 0 digitalH.g\[10\].u.OUTN
rlabel metal2 76656 24780 76656 24780 0 digitalH.g\[10\].u.OUTP
rlabel metal2 79525 32014 79525 32014 0 digitalH.g\[110\].u.OUTN
rlabel metal2 79609 32172 79609 32172 0 digitalH.g\[110\].u.OUTP
rlabel metal3 79344 32844 79344 32844 0 digitalH.g\[111\].u.OUTN
rlabel metal2 79248 33432 79248 33432 0 digitalH.g\[111\].u.OUTP
rlabel metal3 78768 32844 78768 32844 0 digitalH.g\[112\].u.OUTN
rlabel metal2 78825 32172 78825 32172 0 digitalH.g\[112\].u.OUTP
rlabel metal2 78325 32098 78325 32098 0 digitalH.g\[113\].u.OUTN
rlabel metal2 78480 33432 78480 33432 0 digitalH.g\[113\].u.OUTP
rlabel metal3 78096 32844 78096 32844 0 digitalH.g\[114\].u.OUTN
rlabel metal2 78000 33432 78000 33432 0 digitalH.g\[114\].u.OUTP
rlabel metal2 77525 32140 77525 32140 0 digitalH.g\[115\].u.OUTN
rlabel metal2 77635 32014 77635 32014 0 digitalH.g\[115\].u.OUTP
rlabel metal2 77125 32014 77125 32014 0 digitalH.g\[116\].u.OUTN
rlabel metal2 77209 32172 77209 32172 0 digitalH.g\[116\].u.OUTP
rlabel metal2 76725 32014 76725 32014 0 digitalH.g\[117\].u.OUTN
rlabel metal2 76752 33432 76752 33432 0 digitalH.g\[117\].u.OUTP
rlabel metal2 76325 32014 76325 32014 0 digitalH.g\[118\].u.OUTN
rlabel metal2 76425 32172 76425 32172 0 digitalH.g\[118\].u.OUTP
rlabel metal2 75925 32098 75925 32098 0 digitalH.g\[119\].u.OUTN
rlabel metal2 76080 33432 76080 33432 0 digitalH.g\[119\].u.OUTP
rlabel metal2 78528 25998 78528 25998 0 digitalH.g\[11\].u.OUTN
rlabel metal2 77040 24780 77040 24780 0 digitalH.g\[11\].u.OUTP
rlabel metal3 75840 32844 75840 32844 0 digitalH.g\[120\].u.OUTN
rlabel metal2 75593 32256 75593 32256 0 digitalH.g\[120\].u.OUTP
rlabel metal2 75125 32014 75125 32014 0 digitalH.g\[121\].u.OUTN
rlabel metal2 75168 33432 75168 33432 0 digitalH.g\[121\].u.OUTP
rlabel metal2 74725 32014 74725 32014 0 digitalH.g\[122\].u.OUTN
rlabel metal2 74736 33432 74736 33432 0 digitalH.g\[122\].u.OUTP
rlabel metal2 74325 32014 74325 32014 0 digitalH.g\[123\].u.OUTN
rlabel metal2 74369 32172 74369 32172 0 digitalH.g\[123\].u.OUTP
rlabel metal2 73925 32014 73925 32014 0 digitalH.g\[124\].u.OUTN
rlabel metal2 73968 33432 73968 33432 0 digitalH.g\[124\].u.OUTP
rlabel metal2 73525 32014 73525 32014 0 digitalH.g\[125\].u.OUTN
rlabel metal2 73537 32172 73537 32172 0 digitalH.g\[125\].u.OUTP
rlabel metal2 73125 32014 73125 32014 0 digitalH.g\[126\].u.OUTN
rlabel metal2 72864 32508 72864 32508 0 digitalH.g\[126\].u.OUTP
rlabel metal2 71136 31794 71136 31794 0 digitalH.g\[127\].u.OUTN
rlabel metal2 70848 31878 70848 31878 0 digitalH.g\[127\].u.OUTP
rlabel metal3 77808 25536 77808 25536 0 digitalH.g\[12\].u.OUTN
rlabel metal2 77472 25578 77472 25578 0 digitalH.g\[12\].u.OUTP
rlabel metal2 78240 25956 78240 25956 0 digitalH.g\[13\].u.OUTN
rlabel metal2 78000 24780 78000 24780 0 digitalH.g\[13\].u.OUTP
rlabel metal3 79200 25536 79200 25536 0 digitalH.g\[14\].u.OUTN
rlabel metal2 78432 25578 78432 25578 0 digitalH.g\[14\].u.OUTP
rlabel metal2 78816 25956 78816 25956 0 digitalH.g\[15\].u.OUTN
rlabel metal2 78768 24780 78768 24780 0 digitalH.g\[15\].u.OUTP
rlabel metal2 79200 25956 79200 25956 0 digitalH.g\[16\].u.OUTN
rlabel metal2 79200 25074 79200 25074 0 digitalH.g\[16\].u.OUTP
rlabel metal2 79584 25956 79584 25956 0 digitalH.g\[17\].u.OUTN
rlabel metal2 79584 25074 79584 25074 0 digitalH.g\[17\].u.OUTP
rlabel metal2 80160 25998 80160 25998 0 digitalH.g\[18\].u.OUTN
rlabel metal2 79968 25578 79968 25578 0 digitalH.g\[18\].u.OUTP
rlabel metal2 80352 25956 80352 25956 0 digitalH.g\[19\].u.OUTN
rlabel metal2 80208 23940 80208 23940 0 digitalH.g\[19\].u.OUTP
rlabel metal3 73008 25536 73008 25536 0 digitalH.g\[1\].u.OUTN
rlabel metal2 70560 26502 70560 26502 0 digitalH.g\[1\].u.OUTP
rlabel metal2 80832 25956 80832 25956 0 digitalH.g\[20\].u.OUTN
rlabel metal2 81120 24780 81120 24780 0 digitalH.g\[20\].u.OUTP
rlabel metal2 81216 25956 81216 25956 0 digitalH.g\[21\].u.OUTN
rlabel metal2 81600 25074 81600 25074 0 digitalH.g\[21\].u.OUTP
rlabel metal2 81600 25956 81600 25956 0 digitalH.g\[22\].u.OUTN
rlabel metal2 81408 25620 81408 25620 0 digitalH.g\[22\].u.OUTP
rlabel metal2 82080 25956 82080 25956 0 digitalH.g\[23\].u.OUTN
rlabel metal2 81888 24738 81888 24738 0 digitalH.g\[23\].u.OUTP
rlabel metal2 82368 25956 82368 25956 0 digitalH.g\[24\].u.OUTN
rlabel metal2 82368 25074 82368 25074 0 digitalH.g\[24\].u.OUTP
rlabel metal2 82752 25956 82752 25956 0 digitalH.g\[25\].u.OUTN
rlabel metal2 82656 24528 82656 24528 0 digitalH.g\[25\].u.OUTP
rlabel metal2 83184 25536 83184 25536 0 digitalH.g\[26\].u.OUTN
rlabel metal2 83088 24780 83088 24780 0 digitalH.g\[26\].u.OUTP
rlabel metal3 83856 25536 83856 25536 0 digitalH.g\[27\].u.OUTN
rlabel metal2 83520 25578 83520 25578 0 digitalH.g\[27\].u.OUTP
rlabel metal2 84192 25536 84192 25536 0 digitalH.g\[28\].u.OUTN
rlabel metal2 83904 25578 83904 25578 0 digitalH.g\[28\].u.OUTP
rlabel metal2 84576 25998 84576 25998 0 digitalH.g\[29\].u.OUTN
rlabel metal2 84480 25116 84480 25116 0 digitalH.g\[29\].u.OUTP
rlabel metal2 73635 26702 73635 26702 0 digitalH.g\[2\].u.OUTN
rlabel metal2 70896 26628 70896 26628 0 digitalH.g\[2\].u.OUTP
rlabel metal2 84864 25956 84864 25956 0 digitalH.g\[30\].u.OUTN
rlabel metal2 84816 24780 84816 24780 0 digitalH.g\[30\].u.OUTP
rlabel metal2 85248 25956 85248 25956 0 digitalH.g\[31\].u.OUTN
rlabel metal2 85152 24528 85152 24528 0 digitalH.g\[31\].u.OUTP
rlabel metal2 85632 25956 85632 25956 0 digitalH.g\[32\].u.OUTN
rlabel metal2 85488 24780 85488 24780 0 digitalH.g\[32\].u.OUTP
rlabel metal2 86016 25956 86016 25956 0 digitalH.g\[33\].u.OUTN
rlabel metal2 85872 23940 85872 23940 0 digitalH.g\[33\].u.OUTP
rlabel metal2 86400 25914 86400 25914 0 digitalH.g\[34\].u.OUTN
rlabel metal2 86304 25578 86304 25578 0 digitalH.g\[34\].u.OUTP
rlabel metal3 87216 25536 87216 25536 0 digitalH.g\[35\].u.OUTN
rlabel metal2 86688 25158 86688 25158 0 digitalH.g\[35\].u.OUTP
rlabel metal2 87600 24612 87600 24612 0 digitalH.g\[36\].u.OUTN
rlabel metal2 87120 24780 87120 24780 0 digitalH.g\[36\].u.OUTP
rlabel metal2 87840 25956 87840 25956 0 digitalH.g\[37\].u.OUTN
rlabel metal2 87504 24780 87504 24780 0 digitalH.g\[37\].u.OUTP
rlabel metal2 88128 25956 88128 25956 0 digitalH.g\[38\].u.OUTN
rlabel metal2 87984 23940 87984 23940 0 digitalH.g\[38\].u.OUTP
rlabel metal2 88416 25956 88416 25956 0 digitalH.g\[39\].u.OUTN
rlabel metal2 88320 25578 88320 25578 0 digitalH.g\[39\].u.OUTP
rlabel metal2 73344 24864 73344 24864 0 digitalH.g\[3\].u.OUTN
rlabel metal2 73632 25536 73632 25536 0 digitalH.g\[3\].u.OUTP
rlabel metal2 88800 25956 88800 25956 0 digitalH.g\[40\].u.OUTN
rlabel metal2 88656 24780 88656 24780 0 digitalH.g\[40\].u.OUTP
rlabel metal2 89184 25956 89184 25956 0 digitalH.g\[41\].u.OUTN
rlabel metal2 89040 23940 89040 23940 0 digitalH.g\[41\].u.OUTP
rlabel metal3 89808 25536 89808 25536 0 digitalH.g\[42\].u.OUTN
rlabel metal2 89472 25578 89472 25578 0 digitalH.g\[42\].u.OUTP
rlabel metal2 90240 25956 90240 25956 0 digitalH.g\[43\].u.OUTN
rlabel metal2 89904 24780 89904 24780 0 digitalH.g\[43\].u.OUTP
rlabel metal2 90528 25956 90528 25956 0 digitalH.g\[44\].u.OUTN
rlabel metal2 90384 24780 90384 24780 0 digitalH.g\[44\].u.OUTP
rlabel metal2 90816 25956 90816 25956 0 digitalH.g\[45\].u.OUTN
rlabel metal2 90725 26576 90725 26576 0 digitalH.g\[45\].u.OUTP
rlabel metal2 91200 25956 91200 25956 0 digitalH.g\[46\].u.OUTN
rlabel metal2 91152 24780 91152 24780 0 digitalH.g\[46\].u.OUTP
rlabel metal2 91584 25956 91584 25956 0 digitalH.g\[47\].u.OUTN
rlabel metal2 91536 23940 91536 23940 0 digitalH.g\[47\].u.OUTP
rlabel metal2 92064 25956 92064 25956 0 digitalH.g\[48\].u.OUTN
rlabel metal2 91872 25578 91872 25578 0 digitalH.g\[48\].u.OUTP
rlabel metal2 92448 25158 92448 25158 0 digitalH.g\[49\].u.OUTN
rlabel metal2 92160 25578 92160 25578 0 digitalH.g\[49\].u.OUTP
rlabel metal3 73968 24780 73968 24780 0 digitalH.g\[4\].u.OUTN
rlabel metal2 74112 25956 74112 25956 0 digitalH.g\[4\].u.OUTP
rlabel metal2 92832 25956 92832 25956 0 digitalH.g\[50\].u.OUTN
rlabel metal2 92832 24780 92832 24780 0 digitalH.g\[50\].u.OUTP
rlabel metal2 93216 25956 93216 25956 0 digitalH.g\[51\].u.OUTN
rlabel metal2 93264 24780 93264 24780 0 digitalH.g\[51\].u.OUTP
rlabel metal2 93600 25956 93600 25956 0 digitalH.g\[52\].u.OUTN
rlabel metal2 93600 24654 93600 24654 0 digitalH.g\[52\].u.OUTP
rlabel metal2 94080 25956 94080 25956 0 digitalH.g\[53\].u.OUTN
rlabel metal2 93936 24780 93936 24780 0 digitalH.g\[53\].u.OUTP
rlabel metal2 94368 25956 94368 25956 0 digitalH.g\[54\].u.OUTN
rlabel metal2 94368 25074 94368 25074 0 digitalH.g\[54\].u.OUTP
rlabel metal2 94848 25956 94848 25956 0 digitalH.g\[55\].u.OUTN
rlabel metal2 94752 25578 94752 25578 0 digitalH.g\[55\].u.OUTP
rlabel metal2 95232 25956 95232 25956 0 digitalH.g\[56\].u.OUTN
rlabel metal2 95136 25578 95136 25578 0 digitalH.g\[56\].u.OUTP
rlabel metal3 95904 25536 95904 25536 0 digitalH.g\[57\].u.OUTN
rlabel metal2 95616 25578 95616 25578 0 digitalH.g\[57\].u.OUTP
rlabel metal2 96384 25956 96384 25956 0 digitalH.g\[58\].u.OUTN
rlabel metal2 96192 24864 96192 24864 0 digitalH.g\[58\].u.OUTP
rlabel metal3 96960 25536 96960 25536 0 digitalH.g\[59\].u.OUTN
rlabel metal2 96576 25662 96576 25662 0 digitalH.g\[59\].u.OUTP
rlabel metal3 75408 25536 75408 25536 0 digitalH.g\[5\].u.OUTN
rlabel metal2 69984 26670 69984 26670 0 digitalH.g\[5\].u.OUTP
rlabel metal2 96864 25956 96864 25956 0 digitalH.g\[60\].u.OUTN
rlabel metal2 96960 24948 96960 24948 0 digitalH.g\[60\].u.OUTP
rlabel metal2 97248 25956 97248 25956 0 digitalH.g\[61\].u.OUTN
rlabel metal2 97344 25074 97344 25074 0 digitalH.g\[61\].u.OUTP
rlabel metal2 97728 25956 97728 25956 0 digitalH.g\[62\].u.OUTN
rlabel metal2 97680 24780 97680 24780 0 digitalH.g\[62\].u.OUTP
rlabel metal2 98112 25956 98112 25956 0 digitalH.g\[63\].u.OUTN
rlabel metal2 98016 24780 98016 24780 0 digitalH.g\[63\].u.OUTP
rlabel metal2 97925 32014 97925 32014 0 digitalH.g\[64\].u.OUTN
rlabel metal2 98035 32140 98035 32140 0 digitalH.g\[64\].u.OUTP
rlabel metal2 97525 32014 97525 32014 0 digitalH.g\[65\].u.OUTN
rlabel metal2 97635 32140 97635 32140 0 digitalH.g\[65\].u.OUTP
rlabel metal2 97125 32014 97125 32014 0 digitalH.g\[66\].u.OUTN
rlabel metal2 97235 32140 97235 32140 0 digitalH.g\[66\].u.OUTP
rlabel metal2 96725 32056 96725 32056 0 digitalH.g\[67\].u.OUTN
rlabel metal2 96835 32140 96835 32140 0 digitalH.g\[67\].u.OUTP
rlabel metal2 96325 32014 96325 32014 0 digitalH.g\[68\].u.OUTN
rlabel metal2 96435 32140 96435 32140 0 digitalH.g\[68\].u.OUTP
rlabel metal2 95925 32098 95925 32098 0 digitalH.g\[69\].u.OUTN
rlabel metal2 96035 32056 96035 32056 0 digitalH.g\[69\].u.OUTP
rlabel metal2 76224 25998 76224 25998 0 digitalH.g\[6\].u.OUTN
rlabel metal2 74928 24780 74928 24780 0 digitalH.g\[6\].u.OUTP
rlabel metal2 95525 32014 95525 32014 0 digitalH.g\[70\].u.OUTN
rlabel metal2 95635 32140 95635 32140 0 digitalH.g\[70\].u.OUTP
rlabel metal2 95125 32014 95125 32014 0 digitalH.g\[71\].u.OUTN
rlabel metal2 95235 32140 95235 32140 0 digitalH.g\[71\].u.OUTP
rlabel metal2 94725 32014 94725 32014 0 digitalH.g\[72\].u.OUTN
rlabel metal2 94835 32140 94835 32140 0 digitalH.g\[72\].u.OUTP
rlabel metal2 94325 32014 94325 32014 0 digitalH.g\[73\].u.OUTN
rlabel metal2 94435 32140 94435 32140 0 digitalH.g\[73\].u.OUTP
rlabel metal2 93925 32014 93925 32014 0 digitalH.g\[74\].u.OUTN
rlabel metal2 94035 32140 94035 32140 0 digitalH.g\[74\].u.OUTP
rlabel metal2 93525 32014 93525 32014 0 digitalH.g\[75\].u.OUTN
rlabel metal2 93635 32140 93635 32140 0 digitalH.g\[75\].u.OUTP
rlabel metal2 93125 32014 93125 32014 0 digitalH.g\[76\].u.OUTN
rlabel metal2 93235 32140 93235 32140 0 digitalH.g\[76\].u.OUTP
rlabel metal2 92725 32014 92725 32014 0 digitalH.g\[77\].u.OUTN
rlabel metal2 92835 32140 92835 32140 0 digitalH.g\[77\].u.OUTP
rlabel metal2 92325 32056 92325 32056 0 digitalH.g\[78\].u.OUTN
rlabel metal2 92435 32140 92435 32140 0 digitalH.g\[78\].u.OUTP
rlabel metal2 91925 32014 91925 32014 0 digitalH.g\[79\].u.OUTN
rlabel metal2 92035 32140 92035 32140 0 digitalH.g\[79\].u.OUTP
rlabel metal2 75648 25578 75648 25578 0 digitalH.g\[7\].u.OUTN
rlabel metal2 75456 25578 75456 25578 0 digitalH.g\[7\].u.OUTP
rlabel metal2 91525 32014 91525 32014 0 digitalH.g\[80\].u.OUTN
rlabel metal2 91635 32140 91635 32140 0 digitalH.g\[80\].u.OUTP
rlabel metal2 91125 32098 91125 32098 0 digitalH.g\[81\].u.OUTN
rlabel metal2 91235 32140 91235 32140 0 digitalH.g\[81\].u.OUTP
rlabel metal2 90725 32182 90725 32182 0 digitalH.g\[82\].u.OUTN
rlabel metal2 90835 32140 90835 32140 0 digitalH.g\[82\].u.OUTP
rlabel metal2 90325 32056 90325 32056 0 digitalH.g\[83\].u.OUTN
rlabel metal2 90435 32014 90435 32014 0 digitalH.g\[83\].u.OUTP
rlabel metal3 90048 32844 90048 32844 0 digitalH.g\[84\].u.OUTN
rlabel metal2 90240 33432 90240 33432 0 digitalH.g\[84\].u.OUTP
rlabel metal2 89525 32014 89525 32014 0 digitalH.g\[85\].u.OUTN
rlabel metal2 89904 33432 89904 33432 0 digitalH.g\[85\].u.OUTP
rlabel metal3 89568 32928 89568 32928 0 digitalH.g\[86\].u.OUTN
rlabel metal2 89184 32466 89184 32466 0 digitalH.g\[86\].u.OUTP
rlabel metal3 89232 32844 89232 32844 0 digitalH.g\[87\].u.OUTN
rlabel metal2 89040 33432 89040 33432 0 digitalH.g\[87\].u.OUTP
rlabel metal2 88325 32014 88325 32014 0 digitalH.g\[88\].u.OUTN
rlabel metal2 88656 33432 88656 33432 0 digitalH.g\[88\].u.OUTP
rlabel metal3 88272 32844 88272 32844 0 digitalH.g\[89\].u.OUTN
rlabel metal3 88224 33096 88224 33096 0 digitalH.g\[89\].u.OUTP
rlabel metal3 76272 25452 76272 25452 0 digitalH.g\[8\].u.OUTN
rlabel metal2 75744 25956 75744 25956 0 digitalH.g\[8\].u.OUTP
rlabel metal3 88032 32928 88032 32928 0 digitalH.g\[90\].u.OUTN
rlabel metal2 87888 33432 87888 33432 0 digitalH.g\[90\].u.OUTP
rlabel metal2 87125 32140 87125 32140 0 digitalH.g\[91\].u.OUTN
rlabel metal2 87552 33432 87552 33432 0 digitalH.g\[91\].u.OUTP
rlabel metal3 86976 32844 86976 32844 0 digitalH.g\[92\].u.OUTN
rlabel metal3 87072 33096 87072 33096 0 digitalH.g\[92\].u.OUTP
rlabel metal3 86352 32844 86352 32844 0 digitalH.g\[93\].u.OUTN
rlabel metal2 86448 33432 86448 33432 0 digitalH.g\[93\].u.OUTP
rlabel metal2 85925 32140 85925 32140 0 digitalH.g\[94\].u.OUTN
rlabel metal2 86035 32014 86035 32014 0 digitalH.g\[94\].u.OUTP
rlabel metal3 85800 32760 85800 32760 0 digitalH.g\[95\].u.OUTN
rlabel metal2 85632 33432 85632 33432 0 digitalH.g\[95\].u.OUTP
rlabel metal2 85125 32140 85125 32140 0 digitalH.g\[96\].u.OUTN
rlabel metal2 85296 33432 85296 33432 0 digitalH.g\[96\].u.OUTP
rlabel metal2 84725 32014 84725 32014 0 digitalH.g\[97\].u.OUTN
rlabel metal2 84960 33096 84960 33096 0 digitalH.g\[97\].u.OUTP
rlabel metal3 84672 32844 84672 32844 0 digitalH.g\[98\].u.OUTN
rlabel metal2 84435 32014 84435 32014 0 digitalH.g\[98\].u.OUTP
rlabel metal2 83925 32014 83925 32014 0 digitalH.g\[99\].u.OUTN
rlabel metal2 84096 33432 84096 33432 0 digitalH.g\[99\].u.OUTP
rlabel metal2 76512 26040 76512 26040 0 digitalH.g\[9\].u.OUTN
rlabel metal2 76320 24780 76320 24780 0 digitalH.g\[9\].u.OUTP
rlabel metal2 72192 7518 72192 7518 0 digitalL.g\[0\].u.OUTN
rlabel metal2 71040 7854 71040 7854 0 digitalL.g\[0\].u.OUTP
rlabel metal2 83525 13324 83525 13324 0 digitalL.g\[100\].u.OUTN
rlabel metal2 83635 13366 83635 13366 0 digitalL.g\[100\].u.OUTP
rlabel metal2 83125 13324 83125 13324 0 digitalL.g\[101\].u.OUTN
rlabel metal2 83235 13366 83235 13366 0 digitalL.g\[101\].u.OUTP
rlabel metal2 82725 13324 82725 13324 0 digitalL.g\[102\].u.OUTN
rlabel metal2 82835 13366 82835 13366 0 digitalL.g\[102\].u.OUTP
rlabel metal2 82325 13324 82325 13324 0 digitalL.g\[103\].u.OUTN
rlabel metal2 82435 13366 82435 13366 0 digitalL.g\[103\].u.OUTP
rlabel metal2 81984 14028 81984 14028 0 digitalL.g\[104\].u.OUTN
rlabel metal2 82035 13324 82035 13324 0 digitalL.g\[104\].u.OUTP
rlabel metal2 81525 13324 81525 13324 0 digitalL.g\[105\].u.OUTN
rlabel metal2 81635 13366 81635 13366 0 digitalL.g\[105\].u.OUTP
rlabel metal2 81125 13324 81125 13324 0 digitalL.g\[106\].u.OUTN
rlabel metal2 81235 13240 81235 13240 0 digitalL.g\[106\].u.OUTP
rlabel metal2 80725 13366 80725 13366 0 digitalL.g\[107\].u.OUTN
rlabel metal2 80835 13366 80835 13366 0 digitalL.g\[107\].u.OUTP
rlabel metal2 80325 13282 80325 13282 0 digitalL.g\[108\].u.OUTN
rlabel metal2 80435 13366 80435 13366 0 digitalL.g\[108\].u.OUTP
rlabel metal2 79925 13324 79925 13324 0 digitalL.g\[109\].u.OUTN
rlabel metal2 80035 13366 80035 13366 0 digitalL.g\[109\].u.OUTP
rlabel metal2 76835 7802 76835 7802 0 digitalL.g\[10\].u.OUTN
rlabel metal2 76704 7140 76704 7140 0 digitalL.g\[10\].u.OUTP
rlabel metal2 79525 13324 79525 13324 0 digitalL.g\[110\].u.OUTN
rlabel metal2 79635 13324 79635 13324 0 digitalL.g\[110\].u.OUTP
rlabel metal2 79125 13324 79125 13324 0 digitalL.g\[111\].u.OUTN
rlabel metal2 79235 13366 79235 13366 0 digitalL.g\[111\].u.OUTP
rlabel metal2 78725 13366 78725 13366 0 digitalL.g\[112\].u.OUTN
rlabel metal2 78835 13366 78835 13366 0 digitalL.g\[112\].u.OUTP
rlabel metal2 78325 13366 78325 13366 0 digitalL.g\[113\].u.OUTN
rlabel metal2 78435 13324 78435 13324 0 digitalL.g\[113\].u.OUTP
rlabel metal2 77925 13324 77925 13324 0 digitalL.g\[114\].u.OUTN
rlabel metal2 78035 13366 78035 13366 0 digitalL.g\[114\].u.OUTP
rlabel metal2 77525 13282 77525 13282 0 digitalL.g\[115\].u.OUTN
rlabel metal2 77635 13282 77635 13282 0 digitalL.g\[115\].u.OUTP
rlabel metal2 77125 13324 77125 13324 0 digitalL.g\[116\].u.OUTN
rlabel metal2 77235 13324 77235 13324 0 digitalL.g\[116\].u.OUTP
rlabel metal2 76725 13324 76725 13324 0 digitalL.g\[117\].u.OUTN
rlabel metal2 76835 13366 76835 13366 0 digitalL.g\[117\].u.OUTP
rlabel metal2 76325 13366 76325 13366 0 digitalL.g\[118\].u.OUTN
rlabel metal2 76435 13366 76435 13366 0 digitalL.g\[118\].u.OUTP
rlabel metal2 75925 13324 75925 13324 0 digitalL.g\[119\].u.OUTN
rlabel metal2 76035 13366 76035 13366 0 digitalL.g\[119\].u.OUTP
rlabel metal3 77568 7392 77568 7392 0 digitalL.g\[11\].u.OUTN
rlabel metal2 77088 7140 77088 7140 0 digitalL.g\[11\].u.OUTP
rlabel metal2 75525 13282 75525 13282 0 digitalL.g\[120\].u.OUTN
rlabel metal2 75635 13366 75635 13366 0 digitalL.g\[120\].u.OUTP
rlabel metal2 75125 13366 75125 13366 0 digitalL.g\[121\].u.OUTN
rlabel metal2 75235 13408 75235 13408 0 digitalL.g\[121\].u.OUTP
rlabel metal2 74725 13324 74725 13324 0 digitalL.g\[122\].u.OUTN
rlabel metal2 74835 13366 74835 13366 0 digitalL.g\[122\].u.OUTP
rlabel metal3 72972 14532 72972 14532 0 digitalL.g\[123\].u.OUTN
rlabel metal2 74435 13366 74435 13366 0 digitalL.g\[123\].u.OUTP
rlabel metal2 73925 13366 73925 13366 0 digitalL.g\[124\].u.OUTN
rlabel metal2 74035 13324 74035 13324 0 digitalL.g\[124\].u.OUTP
rlabel metal2 73536 13692 73536 13692 0 digitalL.g\[125\].u.OUTN
rlabel metal2 73635 13366 73635 13366 0 digitalL.g\[125\].u.OUTP
rlabel metal2 70608 12600 70608 12600 0 digitalL.g\[126\].u.OUTN
rlabel metal2 70080 13524 70080 13524 0 digitalL.g\[126\].u.OUTP
rlabel metal2 70992 12600 70992 12600 0 digitalL.g\[127\].u.OUTN
rlabel metal2 72835 13366 72835 13366 0 digitalL.g\[127\].u.OUTP
rlabel metal2 78144 7434 78144 7434 0 digitalL.g\[12\].u.OUTN
rlabel metal2 77472 7140 77472 7140 0 digitalL.g\[12\].u.OUTP
rlabel metal3 78240 7392 78240 7392 0 digitalL.g\[13\].u.OUTN
rlabel metal2 77808 6636 77808 6636 0 digitalL.g\[13\].u.OUTP
rlabel metal2 79296 7518 79296 7518 0 digitalL.g\[14\].u.OUTN
rlabel metal2 78336 7140 78336 7140 0 digitalL.g\[14\].u.OUTP
rlabel metal3 79152 7392 79152 7392 0 digitalL.g\[15\].u.OUTN
rlabel metal2 78720 7140 78720 7140 0 digitalL.g\[15\].u.OUTP
rlabel metal3 79872 7308 79872 7308 0 digitalL.g\[16\].u.OUTN
rlabel metal2 79104 7140 79104 7140 0 digitalL.g\[16\].u.OUTP
rlabel metal2 80928 6930 80928 6930 0 digitalL.g\[17\].u.OUTN
rlabel metal2 79440 6636 79440 6636 0 digitalL.g\[17\].u.OUTP
rlabel metal3 80592 7392 80592 7392 0 digitalL.g\[18\].u.OUTN
rlabel metal2 79920 6636 79920 6636 0 digitalL.g\[18\].u.OUTP
rlabel metal3 80688 6636 80688 6636 0 digitalL.g\[19\].u.OUTN
rlabel metal2 80304 6636 80304 6636 0 digitalL.g\[19\].u.OUTP
rlabel metal2 73344 7518 73344 7518 0 digitalL.g\[1\].u.OUTN
rlabel metal2 72576 7434 72576 7434 0 digitalL.g\[1\].u.OUTP
rlabel metal3 81456 6972 81456 6972 0 digitalL.g\[20\].u.OUTN
rlabel metal2 80736 7140 80736 7140 0 digitalL.g\[20\].u.OUTP
rlabel metal2 82368 7434 82368 7434 0 digitalL.g\[21\].u.OUTN
rlabel metal2 81072 6804 81072 6804 0 digitalL.g\[21\].u.OUTP
rlabel metal3 82128 7392 82128 7392 0 digitalL.g\[22\].u.OUTN
rlabel metal2 81504 7140 81504 7140 0 digitalL.g\[22\].u.OUTP
rlabel metal2 82848 7476 82848 7476 0 digitalL.g\[23\].u.OUTN
rlabel metal2 81888 6888 81888 6888 0 digitalL.g\[23\].u.OUTP
rlabel metal3 83040 7308 83040 7308 0 digitalL.g\[24\].u.OUTN
rlabel metal2 82224 6636 82224 6636 0 digitalL.g\[24\].u.OUTP
rlabel metal2 84000 7434 84000 7434 0 digitalL.g\[25\].u.OUTN
rlabel metal2 82752 7140 82752 7140 0 digitalL.g\[25\].u.OUTP
rlabel metal2 83328 7140 83328 7140 0 digitalL.g\[26\].u.OUTN
rlabel metal2 83136 7140 83136 7140 0 digitalL.g\[26\].u.OUTP
rlabel metal2 84192 7518 84192 7518 0 digitalL.g\[27\].u.OUTN
rlabel metal2 83522 7644 83522 7644 0 digitalL.g\[27\].u.OUTP
rlabel metal3 84288 7392 84288 7392 0 digitalL.g\[28\].u.OUTN
rlabel metal2 83856 6636 83856 6636 0 digitalL.g\[28\].u.OUTP
rlabel metal2 85344 7602 85344 7602 0 digitalL.g\[29\].u.OUTN
rlabel metal2 84336 6636 84336 6636 0 digitalL.g\[29\].u.OUTP
rlabel metal2 73728 7518 73728 7518 0 digitalL.g\[2\].u.OUTN
rlabel metal2 73152 7266 73152 7266 0 digitalL.g\[2\].u.OUTP
rlabel metal2 85536 7434 85536 7434 0 digitalL.g\[30\].u.OUTN
rlabel metal2 84672 7140 84672 7140 0 digitalL.g\[30\].u.OUTP
rlabel metal2 85248 7560 85248 7560 0 digitalL.g\[31\].u.OUTN
rlabel metal2 85104 6636 85104 6636 0 digitalL.g\[31\].u.OUTP
rlabel metal3 86304 7308 86304 7308 0 digitalL.g\[32\].u.OUTN
rlabel metal2 85488 6636 85488 6636 0 digitalL.g\[32\].u.OUTP
rlabel metal3 86736 7056 86736 7056 0 digitalL.g\[33\].u.OUTN
rlabel metal2 85968 6636 85968 6636 0 digitalL.g\[33\].u.OUTP
rlabel metal3 86976 7392 86976 7392 0 digitalL.g\[34\].u.OUTN
rlabel metal2 86352 6636 86352 6636 0 digitalL.g\[34\].u.OUTP
rlabel metal2 87744 7434 87744 7434 0 digitalL.g\[35\].u.OUTN
rlabel metal2 86736 6636 86736 6636 0 digitalL.g\[35\].u.OUTP
rlabel metal3 87840 7308 87840 7308 0 digitalL.g\[36\].u.OUTN
rlabel metal2 87072 7140 87072 7140 0 digitalL.g\[36\].u.OUTP
rlabel metal2 88800 7476 88800 7476 0 digitalL.g\[37\].u.OUTN
rlabel metal2 87600 6636 87600 6636 0 digitalL.g\[37\].u.OUTP
rlabel metal3 88512 7392 88512 7392 0 digitalL.g\[38\].u.OUTN
rlabel metal2 87840 6636 87840 6636 0 digitalL.g\[38\].u.OUTP
rlabel metal2 89664 7434 89664 7434 0 digitalL.g\[39\].u.OUTN
rlabel metal2 88320 7140 88320 7140 0 digitalL.g\[39\].u.OUTP
rlabel metal2 73488 6552 73488 6552 0 digitalL.g\[3\].u.OUTN
rlabel metal2 73776 6636 73776 6636 0 digitalL.g\[3\].u.OUTP
rlabel metal3 89472 7308 89472 7308 0 digitalL.g\[40\].u.OUTN
rlabel metal2 88656 6636 88656 6636 0 digitalL.g\[40\].u.OUTP
rlabel metal3 89760 7392 89760 7392 0 digitalL.g\[41\].u.OUTN
rlabel metal2 89136 6636 89136 6636 0 digitalL.g\[41\].u.OUTP
rlabel metal2 90528 7560 90528 7560 0 digitalL.g\[42\].u.OUTN
rlabel metal2 89520 6636 89520 6636 0 digitalL.g\[42\].u.OUTP
rlabel metal2 90048 7560 90048 7560 0 digitalL.g\[43\].u.OUTN
rlabel metal2 89904 6636 89904 6636 0 digitalL.g\[43\].u.OUTP
rlabel metal2 90624 7644 90624 7644 0 digitalL.g\[44\].u.OUTN
rlabel metal2 90384 6636 90384 6636 0 digitalL.g\[44\].u.OUTP
rlabel metal2 91776 7518 91776 7518 0 digitalL.g\[45\].u.OUTN
rlabel metal2 90720 7014 90720 7014 0 digitalL.g\[45\].u.OUTP
rlabel metal2 91200 6552 91200 6552 0 digitalL.g\[46\].u.OUTN
rlabel metal2 91104 7140 91104 7140 0 digitalL.g\[46\].u.OUTP
rlabel metal3 92304 7224 92304 7224 0 digitalL.g\[47\].u.OUTN
rlabel metal2 91440 6636 91440 6636 0 digitalL.g\[47\].u.OUTP
rlabel metal3 92688 6972 92688 6972 0 digitalL.g\[48\].u.OUTN
rlabel metal2 91968 6972 91968 6972 0 digitalL.g\[48\].u.OUTP
rlabel metal2 93504 7434 93504 7434 0 digitalL.g\[49\].u.OUTN
rlabel metal2 92304 6636 92304 6636 0 digitalL.g\[49\].u.OUTP
rlabel metal3 74688 7224 74688 7224 0 digitalL.g\[4\].u.OUTN
rlabel metal2 74208 7140 74208 7140 0 digitalL.g\[4\].u.OUTP
rlabel metal3 93312 7392 93312 7392 0 digitalL.g\[50\].u.OUTN
rlabel metal2 92688 6636 92688 6636 0 digitalL.g\[50\].u.OUTP
rlabel metal3 94464 7098 94464 7098 0 digitalL.g\[51\].u.OUTN
rlabel metal2 93120 7140 93120 7140 0 digitalL.g\[51\].u.OUTP
rlabel metal2 94896 7140 94896 7140 0 digitalL.g\[52\].u.OUTN
rlabel metal2 93648 6636 93648 6636 0 digitalL.g\[52\].u.OUTP
rlabel metal2 94080 6300 94080 6300 0 digitalL.g\[53\].u.OUTN
rlabel metal4 93792 7224 93792 7224 0 digitalL.g\[53\].u.OUTP
rlabel metal3 95040 7224 95040 7224 0 digitalL.g\[54\].u.OUTN
rlabel metal2 94368 7140 94368 7140 0 digitalL.g\[54\].u.OUTP
rlabel metal3 95424 7308 95424 7308 0 digitalL.g\[55\].u.OUTN
rlabel metal2 94704 6636 94704 6636 0 digitalL.g\[55\].u.OUTP
rlabel metal3 96192 7182 96192 7182 0 digitalL.g\[56\].u.OUTN
rlabel metal2 95136 7140 95136 7140 0 digitalL.g\[56\].u.OUTP
rlabel metal3 96048 7392 96048 7392 0 digitalL.g\[57\].u.OUTN
rlabel metal2 95568 6636 95568 6636 0 digitalL.g\[57\].u.OUTP
rlabel metal3 96768 7140 96768 7140 0 digitalL.g\[58\].u.OUTN
rlabel metal2 96048 6636 96048 6636 0 digitalL.g\[58\].u.OUTP
rlabel metal3 97152 6972 97152 6972 0 digitalL.g\[59\].u.OUTN
rlabel metal2 96384 7140 96384 7140 0 digitalL.g\[59\].u.OUTP
rlabel metal3 75024 7392 75024 7392 0 digitalL.g\[5\].u.OUTN
rlabel metal2 74592 7140 74592 7140 0 digitalL.g\[5\].u.OUTP
rlabel metal3 97344 7392 97344 7392 0 digitalL.g\[60\].u.OUTN
rlabel metal2 96768 7140 96768 7140 0 digitalL.g\[60\].u.OUTP
rlabel metal3 97680 7308 97680 7308 0 digitalL.g\[61\].u.OUTN
rlabel metal2 97104 6636 97104 6636 0 digitalL.g\[61\].u.OUTP
rlabel metal3 98880 7098 98880 7098 0 digitalL.g\[62\].u.OUTN
rlabel metal2 97632 6636 97632 6636 0 digitalL.g\[62\].u.OUTP
rlabel metal2 99264 7434 99264 7434 0 digitalL.g\[63\].u.OUTN
rlabel metal2 97968 6636 97968 6636 0 digitalL.g\[63\].u.OUTP
rlabel metal2 97925 13324 97925 13324 0 digitalL.g\[64\].u.OUTN
rlabel metal2 98035 13366 98035 13366 0 digitalL.g\[64\].u.OUTP
rlabel metal2 97525 13324 97525 13324 0 digitalL.g\[65\].u.OUTN
rlabel metal2 97635 13366 97635 13366 0 digitalL.g\[65\].u.OUTP
rlabel metal2 97125 13282 97125 13282 0 digitalL.g\[66\].u.OUTN
rlabel metal2 97235 13366 97235 13366 0 digitalL.g\[66\].u.OUTP
rlabel metal2 96725 13282 96725 13282 0 digitalL.g\[67\].u.OUTN
rlabel metal2 96835 13366 96835 13366 0 digitalL.g\[67\].u.OUTP
rlabel metal2 96325 13324 96325 13324 0 digitalL.g\[68\].u.OUTN
rlabel metal2 96435 13366 96435 13366 0 digitalL.g\[68\].u.OUTP
rlabel metal2 95925 13324 95925 13324 0 digitalL.g\[69\].u.OUTN
rlabel metal2 96035 13366 96035 13366 0 digitalL.g\[69\].u.OUTP
rlabel metal2 75936 7434 75936 7434 0 digitalL.g\[6\].u.OUTN
rlabel metal2 75072 7140 75072 7140 0 digitalL.g\[6\].u.OUTP
rlabel metal2 95525 13366 95525 13366 0 digitalL.g\[70\].u.OUTN
rlabel metal2 95635 13366 95635 13366 0 digitalL.g\[70\].u.OUTP
rlabel metal2 95125 13324 95125 13324 0 digitalL.g\[71\].u.OUTN
rlabel metal2 95235 13366 95235 13366 0 digitalL.g\[71\].u.OUTP
rlabel metal2 94725 13324 94725 13324 0 digitalL.g\[72\].u.OUTN
rlabel metal2 94835 13366 94835 13366 0 digitalL.g\[72\].u.OUTP
rlabel metal2 94325 13366 94325 13366 0 digitalL.g\[73\].u.OUTN
rlabel metal2 94435 13366 94435 13366 0 digitalL.g\[73\].u.OUTP
rlabel metal2 93925 13324 93925 13324 0 digitalL.g\[74\].u.OUTN
rlabel metal2 94035 13366 94035 13366 0 digitalL.g\[74\].u.OUTP
rlabel metal2 93525 13324 93525 13324 0 digitalL.g\[75\].u.OUTN
rlabel metal2 93635 13366 93635 13366 0 digitalL.g\[75\].u.OUTP
rlabel metal2 93125 13366 93125 13366 0 digitalL.g\[76\].u.OUTN
rlabel metal2 93235 13366 93235 13366 0 digitalL.g\[76\].u.OUTP
rlabel metal2 92725 13366 92725 13366 0 digitalL.g\[77\].u.OUTN
rlabel metal2 92835 13366 92835 13366 0 digitalL.g\[77\].u.OUTP
rlabel metal2 92325 13282 92325 13282 0 digitalL.g\[78\].u.OUTN
rlabel metal2 92435 13366 92435 13366 0 digitalL.g\[78\].u.OUTP
rlabel metal2 91925 13282 91925 13282 0 digitalL.g\[79\].u.OUTN
rlabel metal2 92035 13366 92035 13366 0 digitalL.g\[79\].u.OUTP
rlabel metal2 76224 7518 76224 7518 0 digitalL.g\[7\].u.OUTN
rlabel metal2 75456 7140 75456 7140 0 digitalL.g\[7\].u.OUTP
rlabel metal2 91525 13282 91525 13282 0 digitalL.g\[80\].u.OUTN
rlabel metal2 91635 13324 91635 13324 0 digitalL.g\[80\].u.OUTP
rlabel metal2 91125 13282 91125 13282 0 digitalL.g\[81\].u.OUTN
rlabel metal2 91235 13324 91235 13324 0 digitalL.g\[81\].u.OUTP
rlabel metal2 90725 13366 90725 13366 0 digitalL.g\[82\].u.OUTN
rlabel metal2 90835 13324 90835 13324 0 digitalL.g\[82\].u.OUTP
rlabel metal2 90325 13324 90325 13324 0 digitalL.g\[83\].u.OUTN
rlabel metal2 90435 13324 90435 13324 0 digitalL.g\[83\].u.OUTP
rlabel metal2 89925 13324 89925 13324 0 digitalL.g\[84\].u.OUTN
rlabel metal2 90035 13366 90035 13366 0 digitalL.g\[84\].u.OUTP
rlabel metal2 89525 13366 89525 13366 0 digitalL.g\[85\].u.OUTN
rlabel metal2 89635 13366 89635 13366 0 digitalL.g\[85\].u.OUTP
rlabel metal2 89125 13366 89125 13366 0 digitalL.g\[86\].u.OUTN
rlabel metal2 89235 13282 89235 13282 0 digitalL.g\[86\].u.OUTP
rlabel metal2 88725 13282 88725 13282 0 digitalL.g\[87\].u.OUTN
rlabel metal2 88835 13324 88835 13324 0 digitalL.g\[87\].u.OUTP
rlabel metal2 88325 13324 88325 13324 0 digitalL.g\[88\].u.OUTN
rlabel metal2 88435 13240 88435 13240 0 digitalL.g\[88\].u.OUTP
rlabel metal2 87925 13366 87925 13366 0 digitalL.g\[89\].u.OUTN
rlabel metal2 88035 13366 88035 13366 0 digitalL.g\[89\].u.OUTP
rlabel metal3 76320 7224 76320 7224 0 digitalL.g\[8\].u.OUTN
rlabel metal2 75840 7140 75840 7140 0 digitalL.g\[8\].u.OUTP
rlabel metal2 87525 13366 87525 13366 0 digitalL.g\[90\].u.OUTN
rlabel metal2 87635 13366 87635 13366 0 digitalL.g\[90\].u.OUTP
rlabel metal2 87125 13366 87125 13366 0 digitalL.g\[91\].u.OUTN
rlabel metal2 87235 13366 87235 13366 0 digitalL.g\[91\].u.OUTP
rlabel metal2 86725 13324 86725 13324 0 digitalL.g\[92\].u.OUTN
rlabel metal2 86835 13366 86835 13366 0 digitalL.g\[92\].u.OUTP
rlabel metal2 86325 13324 86325 13324 0 digitalL.g\[93\].u.OUTN
rlabel metal2 86435 13366 86435 13366 0 digitalL.g\[93\].u.OUTP
rlabel metal2 85925 13324 85925 13324 0 digitalL.g\[94\].u.OUTN
rlabel metal2 86035 13366 86035 13366 0 digitalL.g\[94\].u.OUTP
rlabel metal2 85525 13324 85525 13324 0 digitalL.g\[95\].u.OUTN
rlabel metal2 85635 13366 85635 13366 0 digitalL.g\[95\].u.OUTP
rlabel metal2 85125 13324 85125 13324 0 digitalL.g\[96\].u.OUTN
rlabel metal2 85235 13366 85235 13366 0 digitalL.g\[96\].u.OUTP
rlabel metal2 84725 13282 84725 13282 0 digitalL.g\[97\].u.OUTN
rlabel metal2 84835 13282 84835 13282 0 digitalL.g\[97\].u.OUTP
rlabel metal2 84325 13366 84325 13366 0 digitalL.g\[98\].u.OUTN
rlabel metal2 84435 13366 84435 13366 0 digitalL.g\[98\].u.OUTP
rlabel metal2 83925 13366 83925 13366 0 digitalL.g\[99\].u.OUTN
rlabel metal2 84035 13366 84035 13366 0 digitalL.g\[99\].u.OUTP
rlabel metal3 76656 7392 76656 7392 0 digitalL.g\[9\].u.OUTN
rlabel metal2 76320 6636 76320 6636 0 digitalL.g\[9\].u.OUTP
rlabel metal2 71424 26376 71424 26376 0 digitalenH.g\[0\].u.OUTN
rlabel metal2 72325 26702 72325 26702 0 digitalenH.g\[0\].u.OUTP
rlabel metal2 98784 25998 98784 25998 0 digitalenH.g\[1\].u.OUTN
rlabel metal2 98400 25956 98400 25956 0 digitalenH.g\[1\].u.OUTP
rlabel metal2 98325 32056 98325 32056 0 digitalenH.g\[2\].u.OUTN
rlabel metal2 98435 32014 98435 32014 0 digitalenH.g\[2\].u.OUTP
rlabel metal3 71952 32844 71952 32844 0 digitalenH.g\[3\].u.OUTN
rlabel metal2 72435 32140 72435 32140 0 digitalenH.g\[3\].u.OUTP
rlabel metal2 71472 7392 71472 7392 0 digitalenL.g\[0\].u.OUTN
rlabel metal3 71874 7812 71874 7812 0 digitalenL.g\[0\].u.OUTP
rlabel metal2 98400 7140 98400 7140 0 digitalenL.g\[1\].u.OUTN
rlabel metal3 98400 7392 98400 7392 0 digitalenL.g\[1\].u.OUTP
rlabel metal2 98325 13324 98325 13324 0 digitalenL.g\[2\].u.OUTN
rlabel metal2 98435 13366 98435 13366 0 digitalenL.g\[2\].u.OUTP
rlabel metal2 71232 12978 71232 12978 0 digitalenL.g\[3\].u.OUTN
rlabel metal2 72435 13324 72435 13324 0 digitalenL.g\[3\].u.OUTP
rlabel metal3 1440 23100 1440 23100 0 net1
rlabel metal2 864 13314 864 13314 0 net10
rlabel metal2 95808 7140 95808 7140 0 net100
rlabel metal2 97344 7188 97344 7188 0 net101
rlabel metal2 97248 6594 97248 6594 0 net102
rlabel metal2 95232 7056 95232 7056 0 net103
rlabel metal2 93408 15372 93408 15372 0 net104
rlabel metal2 93840 15456 93840 15456 0 net105
rlabel metal2 94128 16296 94128 16296 0 net106
rlabel metal2 98448 15456 98448 15456 0 net107
rlabel metal2 97056 15204 97056 15204 0 net108
rlabel metal2 95760 15456 95760 15456 0 net109
rlabel metal2 1056 14490 1056 14490 0 net11
rlabel metal2 86688 7350 86688 7350 0 net110
rlabel metal2 70560 13608 70560 13608 0 net111
rlabel metal2 1680 10248 1680 10248 0 net112
rlabel metal3 366 15708 366 15708 0 net113
rlabel metal3 366 16548 366 16548 0 net114
rlabel metal3 366 17388 366 17388 0 net115
rlabel metal3 366 18228 366 18228 0 net116
rlabel metal3 366 19068 366 19068 0 net117
rlabel metal3 366 19908 366 19908 0 net118
rlabel metal3 366 20748 366 20748 0 net119
rlabel metal3 1152 14952 1152 14952 0 net12
rlabel metal3 366 21588 366 21588 0 net120
rlabel metal2 816 2688 816 2688 0 net13
rlabel metal2 912 3360 912 3360 0 net14
rlabel metal2 1248 4452 1248 4452 0 net15
rlabel metal3 1248 4200 1248 4200 0 net16
rlabel metal2 864 6006 864 6006 0 net17
rlabel metal3 1296 6636 1296 6636 0 net18
rlabel metal3 1200 7392 1200 7392 0 net19
rlabel metal3 1488 23772 1488 23772 0 net2
rlabel metal2 864 8778 864 8778 0 net20
rlabel metal5 73460 32844 73460 32844 0 net21
rlabel metal2 72384 32886 72384 32886 0 net22
rlabel metal2 70368 27594 70368 27594 0 net23
rlabel metal3 76224 24528 76224 24528 0 net24
rlabel metal2 75552 25410 75552 25410 0 net25
rlabel metal2 77856 24486 77856 24486 0 net26
rlabel metal3 77904 25284 77904 25284 0 net27
rlabel metal2 74688 25410 74688 25410 0 net28
rlabel metal3 80592 23856 80592 23856 0 net29
rlabel metal3 71520 13272 71520 13272 0 net3
rlabel metal2 81504 25242 81504 25242 0 net30
rlabel metal2 83280 24528 83280 24528 0 net31
rlabel metal3 83952 25284 83952 25284 0 net32
rlabel metal2 74832 25368 74832 25368 0 net33
rlabel metal2 76320 33222 76320 33222 0 net34
rlabel metal3 76320 33012 76320 33012 0 net35
rlabel metal2 78432 32928 78432 32928 0 net36
rlabel metal3 78816 33600 78816 33600 0 net37
rlabel metal2 75168 32886 75168 32886 0 net38
rlabel metal2 80928 33558 80928 33558 0 net39
rlabel metal2 71520 32802 71520 32802 0 net4
rlabel metal2 82848 33558 82848 33558 0 net40
rlabel metal2 84480 32928 84480 32928 0 net41
rlabel metal3 85872 32844 85872 32844 0 net42
rlabel metal2 83136 33054 83136 33054 0 net43
rlabel metal2 74688 33096 74688 33096 0 net44
rlabel metal2 86784 24486 86784 24486 0 net45
rlabel metal2 88752 25284 88752 25284 0 net46
rlabel metal2 91296 23898 91296 23898 0 net47
rlabel metal3 91104 25284 91104 25284 0 net48
rlabel metal2 93408 23898 93408 23898 0 net49
rlabel metal3 1152 8820 1152 8820 0 net5
rlabel metal3 93840 25284 93840 25284 0 net50
rlabel metal2 95424 24906 95424 24906 0 net51
rlabel metal2 96192 25242 96192 25242 0 net52
rlabel metal2 92352 25326 92352 25326 0 net53
rlabel metal2 87648 33012 87648 33012 0 net54
rlabel metal2 89760 32928 89760 32928 0 net55
rlabel metal2 89568 33348 89568 33348 0 net56
rlabel metal2 91296 34020 91296 34020 0 net57
rlabel metal2 89760 33390 89760 33390 0 net58
rlabel metal2 94368 33012 94368 33012 0 net59
rlabel metal2 864 10290 864 10290 0 net6
rlabel metal2 94176 33600 94176 33600 0 net60
rlabel metal2 96912 33600 96912 33600 0 net61
rlabel metal3 98640 32844 98640 32844 0 net62
rlabel metal3 96240 33600 96240 33600 0 net63
rlabel metal2 87072 33516 87072 33516 0 net64
rlabel metal3 1632 4872 1632 4872 0 net65
rlabel metal2 73056 14742 73056 14742 0 net66
rlabel metal2 70848 7980 70848 7980 0 net67
rlabel metal2 76032 7056 76032 7056 0 net68
rlabel metal3 76464 7140 76464 7140 0 net69
rlabel metal2 1440 10458 1440 10458 0 net7
rlabel metal3 78864 7140 78864 7140 0 net70
rlabel metal2 80640 7056 80640 7056 0 net71
rlabel metal2 75552 7266 75552 7266 0 net72
rlabel metal2 74112 15414 74112 15414 0 net73
rlabel metal2 74304 15750 74304 15750 0 net74
rlabel metal2 79776 15330 79776 15330 0 net75
rlabel metal2 79392 15414 79392 15414 0 net76
rlabel metal3 77088 16044 77088 16044 0 net77
rlabel metal2 80976 5712 80976 5712 0 net78
rlabel metal3 83808 7140 83808 7140 0 net79
rlabel metal2 1248 11466 1248 11466 0 net8
rlabel metal2 84576 7056 84576 7056 0 net80
rlabel metal3 86448 7140 86448 7140 0 net81
rlabel metal3 84048 7224 84048 7224 0 net82
rlabel metal2 82560 15876 82560 15876 0 net83
rlabel metal2 82224 16296 82224 16296 0 net84
rlabel metal2 83808 16338 83808 16338 0 net85
rlabel metal2 85056 15750 85056 15750 0 net86
rlabel metal3 84000 16296 84000 16296 0 net87
rlabel metal2 74688 7308 74688 7308 0 net88
rlabel metal3 88608 7140 88608 7140 0 net89
rlabel metal2 864 12390 864 12390 0 net9
rlabel metal3 89856 7140 89856 7140 0 net90
rlabel metal3 90480 7140 90480 7140 0 net91
rlabel metal2 93024 7224 93024 7224 0 net92
rlabel metal3 88752 7224 88752 7224 0 net93
rlabel metal2 87456 15918 87456 15918 0 net94
rlabel metal2 87984 15456 87984 15456 0 net95
rlabel metal3 89664 15456 89664 15456 0 net96
rlabel metal2 90528 15078 90528 15078 0 net97
rlabel metal3 86496 16296 86496 16296 0 net98
rlabel metal3 94656 7140 94656 7140 0 net99
rlabel metal3 318 22428 318 22428 0 ui_in[0]
rlabel metal3 366 23268 366 23268 0 ui_in[1]
rlabel metal3 366 24108 366 24108 0 ui_in[2]
rlabel metal3 366 24948 366 24948 0 ui_in[3]
rlabel metal3 366 8988 366 8988 0 uio_out[0]
rlabel metal3 366 9828 366 9828 0 uio_out[1]
rlabel metal3 366 10668 366 10668 0 uio_out[2]
rlabel metal3 366 11508 366 11508 0 uio_out[3]
rlabel metal3 366 12348 366 12348 0 uio_out[4]
rlabel metal3 366 13188 366 13188 0 uio_out[5]
rlabel metal3 366 14028 366 14028 0 uio_out[6]
rlabel metal3 366 14868 366 14868 0 uio_out[7]
rlabel metal3 366 2268 366 2268 0 uo_out[0]
rlabel metal3 366 3108 366 3108 0 uo_out[1]
rlabel metal3 558 3948 558 3948 0 uo_out[2]
rlabel metal2 672 4578 672 4578 0 uo_out[3]
rlabel metal3 366 5628 366 5628 0 uo_out[4]
rlabel metal3 366 6468 366 6468 0 uo_out[5]
rlabel metal3 366 7308 366 7308 0 uo_out[6]
rlabel metal3 366 8148 366 8148 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 100000 40000
<< end >>
