VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dac2u128out4in
  CLASS BLOCK ;
  FOREIGN dac2u128out4in ;
  ORIGIN 0 0 ;
  SIZE 133.800 BY 26.190 ;
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 73 0 133.8 26.19 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 0 0 60 26.19 ;
    END
  END VDD
#  PIN VbiasP[1]
#    PORT
#      LAYER Metal1 ;
#        RECT 0.9 14.95 132.9 19.88 ;
#    END
#  END VbiasP[1]
#  PIN Iout
#    PORT
#      LAYER Metal1 ;
#        RECT 0 12.745 133.8 13.445 ;
#    END
#  END Iout
#  PIN VbiasP[0]
#    PORT
#      LAYER Metal1 ;
#        RECT 0.9 6.31 132.9 11.24 ;
#    END
#  END VbiasP[0]
  PIN ON[64]
    PORT
      LAYER Metal2 ;
        RECT 130.03 25.9 130.32 26.19 ;
    END
  END ON[64]
  PIN ONB[64]
    PORT
      LAYER Metal2 ;
        RECT 129.48 25.9 129.77 26.19 ;
    END
  END ONB[64]
  PIN ON[65]
    PORT
      LAYER Metal2 ;
        RECT 128.03 25.9 128.32 26.19 ;
    END
  END ON[65]
  PIN ONB[65]
    PORT
      LAYER Metal2 ;
        RECT 127.48 25.9 127.77 26.19 ;
    END
  END ONB[65]
  PIN ON[66]
    PORT
      LAYER Metal2 ;
        RECT 126.03 25.9 126.32 26.19 ;
    END
  END ON[66]
  PIN ONB[66]
    PORT
      LAYER Metal2 ;
        RECT 125.48 25.9 125.77 26.19 ;
    END
  END ONB[66]
  PIN ON[67]
    PORT
      LAYER Metal2 ;
        RECT 124.03 25.9 124.32 26.19 ;
    END
  END ON[67]
  PIN ONB[67]
    PORT
      LAYER Metal2 ;
        RECT 123.48 25.9 123.77 26.19 ;
    END
  END ONB[67]
  PIN ON[68]
    PORT
      LAYER Metal2 ;
        RECT 122.03 25.9 122.32 26.19 ;
    END
  END ON[68]
  PIN ONB[68]
    PORT
      LAYER Metal2 ;
        RECT 121.48 25.9 121.77 26.19 ;
    END
  END ONB[68]
  PIN ON[69]
    PORT
      LAYER Metal2 ;
        RECT 120.03 25.9 120.32 26.19 ;
    END
  END ON[69]
  PIN ONB[69]
    PORT
      LAYER Metal2 ;
        RECT 119.48 25.9 119.77 26.19 ;
    END
  END ONB[69]
  PIN ON[70]
    PORT
      LAYER Metal2 ;
        RECT 118.03 25.9 118.32 26.19 ;
    END
  END ON[70]
  PIN ONB[70]
    PORT
      LAYER Metal2 ;
        RECT 117.48 25.9 117.77 26.19 ;
    END
  END ONB[70]
  PIN ON[71]
    PORT
      LAYER Metal2 ;
        RECT 116.03 25.9 116.32 26.19 ;
    END
  END ON[71]
  PIN ONB[71]
    PORT
      LAYER Metal2 ;
        RECT 115.48 25.9 115.77 26.19 ;
    END
  END ONB[71]
  PIN ON[72]
    PORT
      LAYER Metal2 ;
        RECT 114.03 25.9 114.32 26.19 ;
    END
  END ON[72]
  PIN ONB[72]
    PORT
      LAYER Metal2 ;
        RECT 113.48 25.9 113.77 26.19 ;
    END
  END ONB[72]
  PIN ON[73]
    PORT
      LAYER Metal2 ;
        RECT 112.03 25.9 112.32 26.19 ;
    END
  END ON[73]
  PIN ONB[73]
    PORT
      LAYER Metal2 ;
        RECT 111.48 25.9 111.77 26.19 ;
    END
  END ONB[73]
  PIN ON[74]
    PORT
      LAYER Metal2 ;
        RECT 110.03 25.9 110.32 26.19 ;
    END
  END ON[74]
  PIN ONB[74]
    PORT
      LAYER Metal2 ;
        RECT 109.48 25.9 109.77 26.19 ;
    END
  END ONB[74]
  PIN ON[75]
    PORT
      LAYER Metal2 ;
        RECT 108.03 25.9 108.32 26.19 ;
    END
  END ON[75]
  PIN ONB[75]
    PORT
      LAYER Metal2 ;
        RECT 107.48 25.9 107.77 26.19 ;
    END
  END ONB[75]
  PIN ON[76]
    PORT
      LAYER Metal2 ;
        RECT 106.03 25.9 106.32 26.19 ;
    END
  END ON[76]
  PIN ONB[76]
    PORT
      LAYER Metal2 ;
        RECT 105.48 25.9 105.77 26.19 ;
    END
  END ONB[76]
  PIN ON[77]
    PORT
      LAYER Metal2 ;
        RECT 104.03 25.9 104.32 26.19 ;
    END
  END ON[77]
  PIN ONB[77]
    PORT
      LAYER Metal2 ;
        RECT 103.48 25.9 103.77 26.19 ;
    END
  END ONB[77]
  PIN ON[78]
    PORT
      LAYER Metal2 ;
        RECT 102.03 25.9 102.32 26.19 ;
    END
  END ON[78]
  PIN ONB[78]
    PORT
      LAYER Metal2 ;
        RECT 101.48 25.9 101.77 26.19 ;
    END
  END ONB[78]
  PIN ON[79]
    PORT
      LAYER Metal2 ;
        RECT 100.03 25.9 100.32 26.19 ;
    END
  END ON[79]
  PIN ONB[79]
    PORT
      LAYER Metal2 ;
        RECT 99.48 25.9 99.77 26.19 ;
    END
  END ONB[79]
  PIN ON[80]
    PORT
      LAYER Metal2 ;
        RECT 98.03 25.9 98.32 26.19 ;
    END
  END ON[80]
  PIN ONB[80]
    PORT
      LAYER Metal2 ;
        RECT 97.48 25.9 97.77 26.19 ;
    END
  END ONB[80]
  PIN ON[81]
    PORT
      LAYER Metal2 ;
        RECT 96.03 25.9 96.32 26.19 ;
    END
  END ON[81]
  PIN ONB[81]
    PORT
      LAYER Metal2 ;
        RECT 95.48 25.9 95.77 26.19 ;
    END
  END ONB[81]
  PIN ON[82]
    PORT
      LAYER Metal2 ;
        RECT 94.03 25.9 94.32 26.19 ;
    END
  END ON[82]
  PIN ONB[82]
    PORT
      LAYER Metal2 ;
        RECT 93.48 25.9 93.77 26.19 ;
    END
  END ONB[82]
  PIN ON[83]
    PORT
      LAYER Metal2 ;
        RECT 92.03 25.9 92.32 26.19 ;
    END
  END ON[83]
  PIN ONB[83]
    PORT
      LAYER Metal2 ;
        RECT 91.48 25.9 91.77 26.19 ;
    END
  END ONB[83]
  PIN ON[84]
    PORT
      LAYER Metal2 ;
        RECT 90.03 25.9 90.32 26.19 ;
    END
  END ON[84]
  PIN ONB[84]
    PORT
      LAYER Metal2 ;
        RECT 89.48 25.9 89.77 26.19 ;
    END
  END ONB[84]
  PIN ON[85]
    PORT
      LAYER Metal2 ;
        RECT 88.03 25.9 88.32 26.19 ;
    END
  END ON[85]
  PIN ONB[85]
    PORT
      LAYER Metal2 ;
        RECT 87.48 25.9 87.77 26.19 ;
    END
  END ONB[85]
  PIN ON[86]
    PORT
      LAYER Metal2 ;
        RECT 86.03 25.9 86.32 26.19 ;
    END
  END ON[86]
  PIN ONB[86]
    PORT
      LAYER Metal2 ;
        RECT 85.48 25.9 85.77 26.19 ;
    END
  END ONB[86]
  PIN ON[87]
    PORT
      LAYER Metal2 ;
        RECT 84.03 25.9 84.32 26.19 ;
    END
  END ON[87]
  PIN ONB[87]
    PORT
      LAYER Metal2 ;
        RECT 83.48 25.9 83.77 26.19 ;
    END
  END ONB[87]
  PIN ON[88]
    PORT
      LAYER Metal2 ;
        RECT 82.03 25.9 82.32 26.19 ;
    END
  END ON[88]
  PIN ONB[88]
    PORT
      LAYER Metal2 ;
        RECT 81.48 25.9 81.77 26.19 ;
    END
  END ONB[88]
  PIN ON[89]
    PORT
      LAYER Metal2 ;
        RECT 80.03 25.9 80.32 26.19 ;
    END
  END ON[89]
  PIN ONB[89]
    PORT
      LAYER Metal2 ;
        RECT 79.48 25.9 79.77 26.19 ;
    END
  END ONB[89]
  PIN ON[90]
    PORT
      LAYER Metal2 ;
        RECT 78.03 25.9 78.32 26.19 ;
    END
  END ON[90]
  PIN ONB[90]
    PORT
      LAYER Metal2 ;
        RECT 77.48 25.9 77.77 26.19 ;
    END
  END ONB[90]
  PIN ON[91]
    PORT
      LAYER Metal2 ;
        RECT 76.03 25.9 76.32 26.19 ;
    END
  END ON[91]
  PIN ONB[91]
    PORT
      LAYER Metal2 ;
        RECT 75.48 25.9 75.77 26.19 ;
    END
  END ONB[91]
  PIN ON[92]
    PORT
      LAYER Metal2 ;
        RECT 74.03 25.9 74.32 26.19 ;
    END
  END ON[92]
  PIN ONB[92]
    PORT
      LAYER Metal2 ;
        RECT 73.48 25.9 73.77 26.19 ;
    END
  END ONB[92]
  PIN ON[93]
    PORT
      LAYER Metal2 ;
        RECT 72.03 25.9 72.32 26.19 ;
    END
  END ON[93]
  PIN ONB[93]
    PORT
      LAYER Metal2 ;
        RECT 71.48 25.9 71.77 26.19 ;
    END
  END ONB[93]
  PIN ON[94]
    PORT
      LAYER Metal2 ;
        RECT 70.03 25.9 70.32 26.19 ;
    END
  END ON[94]
  PIN ONB[94]
    PORT
      LAYER Metal2 ;
        RECT 69.48 25.9 69.77 26.19 ;
    END
  END ONB[94]
  PIN ON[95]
    PORT
      LAYER Metal2 ;
        RECT 68.03 25.9 68.32 26.19 ;
    END
  END ON[95]
  PIN ONB[95]
    PORT
      LAYER Metal2 ;
        RECT 67.48 25.9 67.77 26.19 ;
    END
  END ONB[95]
  PIN EN[2]
    PORT
      LAYER Metal2 ;
        RECT 132.03 25.9 132.32 26.19 ;
    END
  END EN[2]
  PIN ENB[2]
    PORT
      LAYER Metal2 ;
        RECT 131.48 25.9 131.77 26.19 ;
    END
  END ENB[2]
  PIN ON[97]
    PORT
      LAYER Metal2 ;
        RECT 64.03 25.9 64.32 26.19 ;
    END
  END ON[97]
  PIN ONB[97]
    PORT
      LAYER Metal2 ;
        RECT 63.48 25.9 63.77 26.19 ;
    END
  END ONB[97]
  PIN ON[98]
    PORT
      LAYER Metal2 ;
        RECT 62.03 25.9 62.32 26.19 ;
    END
  END ON[98]
  PIN ONB[98]
    PORT
      LAYER Metal2 ;
        RECT 61.48 25.9 61.77 26.19 ;
    END
  END ONB[98]
  PIN ON[99]
    PORT
      LAYER Metal2 ;
        RECT 60.03 25.9 60.32 26.19 ;
    END
  END ON[99]
  PIN ONB[99]
    PORT
      LAYER Metal2 ;
        RECT 59.48 25.9 59.77 26.19 ;
    END
  END ONB[99]
  PIN ON[100]
    PORT
      LAYER Metal2 ;
        RECT 58.03 25.9 58.32 26.19 ;
    END
  END ON[100]
  PIN ONB[100]
    PORT
      LAYER Metal2 ;
        RECT 57.48 25.9 57.77 26.19 ;
    END
  END ONB[100]
  PIN ON[101]
    PORT
      LAYER Metal2 ;
        RECT 56.03 25.9 56.32 26.19 ;
    END
  END ON[101]
  PIN ONB[101]
    PORT
      LAYER Metal2 ;
        RECT 55.48 25.9 55.77 26.19 ;
    END
  END ONB[101]
  PIN ON[102]
    PORT
      LAYER Metal2 ;
        RECT 54.03 25.9 54.32 26.19 ;
    END
  END ON[102]
  PIN ONB[102]
    PORT
      LAYER Metal2 ;
        RECT 53.48 25.9 53.77 26.19 ;
    END
  END ONB[102]
  PIN ON[103]
    PORT
      LAYER Metal2 ;
        RECT 52.03 25.9 52.32 26.19 ;
    END
  END ON[103]
  PIN ONB[103]
    PORT
      LAYER Metal2 ;
        RECT 51.48 25.9 51.77 26.19 ;
    END
  END ONB[103]
  PIN ON[104]
    PORT
      LAYER Metal2 ;
        RECT 50.03 25.9 50.32 26.19 ;
    END
  END ON[104]
  PIN ONB[104]
    PORT
      LAYER Metal2 ;
        RECT 49.48 25.9 49.77 26.19 ;
    END
  END ONB[104]
  PIN ON[105]
    PORT
      LAYER Metal2 ;
        RECT 48.03 25.9 48.32 26.19 ;
    END
  END ON[105]
  PIN ONB[105]
    PORT
      LAYER Metal2 ;
        RECT 47.48 25.9 47.77 26.19 ;
    END
  END ONB[105]
  PIN ON[106]
    PORT
      LAYER Metal2 ;
        RECT 46.03 25.9 46.32 26.19 ;
    END
  END ON[106]
  PIN ONB[106]
    PORT
      LAYER Metal2 ;
        RECT 45.48 25.9 45.77 26.19 ;
    END
  END ONB[106]
  PIN ON[107]
    PORT
      LAYER Metal2 ;
        RECT 44.03 25.9 44.32 26.19 ;
    END
  END ON[107]
  PIN ONB[107]
    PORT
      LAYER Metal2 ;
        RECT 43.48 25.9 43.77 26.19 ;
    END
  END ONB[107]
  PIN ON[108]
    PORT
      LAYER Metal2 ;
        RECT 42.03 25.9 42.32 26.19 ;
    END
  END ON[108]
  PIN ONB[108]
    PORT
      LAYER Metal2 ;
        RECT 41.48 25.9 41.77 26.19 ;
    END
  END ONB[108]
  PIN ON[109]
    PORT
      LAYER Metal2 ;
        RECT 40.03 25.9 40.32 26.19 ;
    END
  END ON[109]
  PIN ONB[109]
    PORT
      LAYER Metal2 ;
        RECT 39.48 25.9 39.77 26.19 ;
    END
  END ONB[109]
  PIN ON[110]
    PORT
      LAYER Metal2 ;
        RECT 38.03 25.9 38.32 26.19 ;
    END
  END ON[110]
  PIN ONB[110]
    PORT
      LAYER Metal2 ;
        RECT 37.48 25.9 37.77 26.19 ;
    END
  END ONB[110]
  PIN ON[111]
    PORT
      LAYER Metal2 ;
        RECT 36.03 25.9 36.32 26.19 ;
    END
  END ON[111]
  PIN ONB[111]
    PORT
      LAYER Metal2 ;
        RECT 35.48 25.9 35.77 26.19 ;
    END
  END ONB[111]
  PIN ON[112]
    PORT
      LAYER Metal2 ;
        RECT 34.03 25.9 34.32 26.19 ;
    END
  END ON[112]
  PIN ONB[112]
    PORT
      LAYER Metal2 ;
        RECT 33.48 25.9 33.77 26.19 ;
    END
  END ONB[112]
  PIN ON[113]
    PORT
      LAYER Metal2 ;
        RECT 32.03 25.9 32.32 26.19 ;
    END
  END ON[113]
  PIN ONB[113]
    PORT
      LAYER Metal2 ;
        RECT 31.48 25.9 31.77 26.19 ;
    END
  END ONB[113]
  PIN ON[114]
    PORT
      LAYER Metal2 ;
        RECT 30.03 25.9 30.32 26.19 ;
    END
  END ON[114]
  PIN ONB[114]
    PORT
      LAYER Metal2 ;
        RECT 29.48 25.9 29.77 26.19 ;
    END
  END ONB[114]
  PIN ON[115]
    PORT
      LAYER Metal2 ;
        RECT 28.03 25.9 28.32 26.19 ;
    END
  END ON[115]
  PIN ONB[115]
    PORT
      LAYER Metal2 ;
        RECT 27.48 25.9 27.77 26.19 ;
    END
  END ONB[115]
  PIN ON[116]
    PORT
      LAYER Metal2 ;
        RECT 26.03 25.9 26.32 26.19 ;
    END
  END ON[116]
  PIN ONB[116]
    PORT
      LAYER Metal2 ;
        RECT 25.48 25.9 25.77 26.19 ;
    END
  END ONB[116]
  PIN ON[117]
    PORT
      LAYER Metal2 ;
        RECT 24.03 25.9 24.32 26.19 ;
    END
  END ON[117]
  PIN ONB[117]
    PORT
      LAYER Metal2 ;
        RECT 23.48 25.9 23.77 26.19 ;
    END
  END ONB[117]
  PIN ON[118]
    PORT
      LAYER Metal2 ;
        RECT 22.03 25.9 22.32 26.19 ;
    END
  END ON[118]
  PIN ONB[118]
    PORT
      LAYER Metal2 ;
        RECT 21.48 25.9 21.77 26.19 ;
    END
  END ONB[118]
  PIN ON[119]
    PORT
      LAYER Metal2 ;
        RECT 20.03 25.9 20.32 26.19 ;
    END
  END ON[119]
  PIN ONB[119]
    PORT
      LAYER Metal2 ;
        RECT 19.48 25.9 19.77 26.19 ;
    END
  END ONB[119]
  PIN ON[120]
    PORT
      LAYER Metal2 ;
        RECT 18.03 25.9 18.32 26.19 ;
    END
  END ON[120]
  PIN ONB[120]
    PORT
      LAYER Metal2 ;
        RECT 17.48 25.9 17.77 26.19 ;
    END
  END ONB[120]
  PIN ON[121]
    PORT
      LAYER Metal2 ;
        RECT 16.03 25.9 16.32 26.19 ;
    END
  END ON[121]
  PIN ONB[121]
    PORT
      LAYER Metal2 ;
        RECT 15.48 25.9 15.77 26.19 ;
    END
  END ONB[121]
  PIN ON[122]
    PORT
      LAYER Metal2 ;
        RECT 14.03 25.9 14.32 26.19 ;
    END
  END ON[122]
  PIN ONB[122]
    PORT
      LAYER Metal2 ;
        RECT 13.48 25.9 13.77 26.19 ;
    END
  END ONB[122]
  PIN ON[123]
    PORT
      LAYER Metal2 ;
        RECT 12.03 25.9 12.32 26.19 ;
    END
  END ON[123]
  PIN ONB[123]
    PORT
      LAYER Metal2 ;
        RECT 11.48 25.9 11.77 26.19 ;
    END
  END ONB[123]
  PIN ON[124]
    PORT
      LAYER Metal2 ;
        RECT 10.03 25.9 10.32 26.19 ;
    END
  END ON[124]
  PIN ONB[124]
    PORT
      LAYER Metal2 ;
        RECT 9.48 25.9 9.77 26.19 ;
    END
  END ONB[124]
  PIN ON[125]
    PORT
      LAYER Metal2 ;
        RECT 8.03 25.9 8.32 26.19 ;
    END
  END ON[125]
  PIN ONB[125]
    PORT
      LAYER Metal2 ;
        RECT 7.48 25.9 7.77 26.19 ;
    END
  END ONB[125]
  PIN ON[126]
    PORT
      LAYER Metal2 ;
        RECT 6.03 25.9 6.32 26.19 ;
    END
  END ON[126]
  PIN ONB[126]
    PORT
      LAYER Metal2 ;
        RECT 5.48 25.9 5.77 26.19 ;
    END
  END ONB[126]
  PIN ON[127]
    PORT
      LAYER Metal2 ;
        RECT 4.03 25.9 4.32 26.19 ;
    END
  END ON[127]
  PIN ONB[127]
    PORT
      LAYER Metal2 ;
        RECT 3.48 25.9 3.77 26.19 ;
    END
  END ONB[127]
  PIN ON[96]
    PORT
      LAYER Metal2 ;
        RECT 66.03 25.9 66.32 26.19 ;
    END
  END ON[96]
  PIN ONB[96]
    PORT
      LAYER Metal2 ;
        RECT 65.48 25.9 65.77 26.19 ;
    END
  END ONB[96]
  PIN EN[3]
    PORT
      LAYER Metal2 ;
        RECT 2.03 25.9 2.32 26.19 ;
    END
  END EN[3]
  PIN ENB[3]
    PORT
      LAYER Metal2 ;
        RECT 1.48 25.9 1.77 26.19 ;
    END
  END ENB[3]
  PIN ON[0]
    PORT
      LAYER Metal2 ;
        RECT 3.48 0 3.77 0.29 ;
    END
  END ON[0]
  PIN ONB[0]
    PORT
      LAYER Metal2 ;
        RECT 4.03 0 4.32 0.29 ;
    END
  END ONB[0]
  PIN ON[1]
    PORT
      LAYER Metal2 ;
        RECT 5.48 0 5.77 0.29 ;
    END
  END ON[1]
  PIN ONB[1]
    PORT
      LAYER Metal2 ;
        RECT 6.03 0 6.32 0.29 ;
    END
  END ONB[1]
  PIN ON[2]
    PORT
      LAYER Metal2 ;
        RECT 7.48 0 7.77 0.29 ;
    END
  END ON[2]
  PIN ONB[2]
    PORT
      LAYER Metal2 ;
        RECT 8.03 0 8.32 0.29 ;
    END
  END ONB[2]
  PIN ON[3]
    PORT
      LAYER Metal2 ;
        RECT 9.48 0 9.77 0.29 ;
    END
  END ON[3]
  PIN ONB[3]
    PORT
      LAYER Metal2 ;
        RECT 10.03 0 10.32 0.29 ;
    END
  END ONB[3]
  PIN ON[4]
    PORT
      LAYER Metal2 ;
        RECT 11.48 0 11.77 0.29 ;
    END
  END ON[4]
  PIN ONB[4]
    PORT
      LAYER Metal2 ;
        RECT 12.03 0 12.32 0.29 ;
    END
  END ONB[4]
  PIN ON[5]
    PORT
      LAYER Metal2 ;
        RECT 13.48 0 13.77 0.29 ;
    END
  END ON[5]
  PIN ONB[5]
    PORT
      LAYER Metal2 ;
        RECT 14.03 0 14.32 0.29 ;
    END
  END ONB[5]
  PIN ON[6]
    PORT
      LAYER Metal2 ;
        RECT 15.48 0 15.77 0.29 ;
    END
  END ON[6]
  PIN ONB[6]
    PORT
      LAYER Metal2 ;
        RECT 16.03 0 16.32 0.29 ;
    END
  END ONB[6]
  PIN ON[7]
    PORT
      LAYER Metal2 ;
        RECT 17.48 0 17.77 0.29 ;
    END
  END ON[7]
  PIN ONB[7]
    PORT
      LAYER Metal2 ;
        RECT 18.03 0 18.32 0.29 ;
    END
  END ONB[7]
  PIN ON[8]
    PORT
      LAYER Metal2 ;
        RECT 19.48 0 19.77 0.29 ;
    END
  END ON[8]
  PIN ONB[8]
    PORT
      LAYER Metal2 ;
        RECT 20.03 0 20.32 0.29 ;
    END
  END ONB[8]
  PIN ON[9]
    PORT
      LAYER Metal2 ;
        RECT 21.48 0 21.77 0.29 ;
    END
  END ON[9]
  PIN ONB[9]
    PORT
      LAYER Metal2 ;
        RECT 22.03 0 22.32 0.29 ;
    END
  END ONB[9]
  PIN ON[10]
    PORT
      LAYER Metal2 ;
        RECT 23.48 0 23.77 0.29 ;
    END
  END ON[10]
  PIN ONB[10]
    PORT
      LAYER Metal2 ;
        RECT 24.03 0 24.32 0.29 ;
    END
  END ONB[10]
  PIN ON[11]
    PORT
      LAYER Metal2 ;
        RECT 25.48 0 25.77 0.29 ;
    END
  END ON[11]
  PIN ONB[11]
    PORT
      LAYER Metal2 ;
        RECT 26.03 0 26.32 0.29 ;
    END
  END ONB[11]
  PIN ON[12]
    PORT
      LAYER Metal2 ;
        RECT 27.48 0 27.77 0.29 ;
    END
  END ON[12]
  PIN ONB[12]
    PORT
      LAYER Metal2 ;
        RECT 28.03 0 28.32 0.29 ;
    END
  END ONB[12]
  PIN ON[13]
    PORT
      LAYER Metal2 ;
        RECT 29.48 0 29.77 0.29 ;
    END
  END ON[13]
  PIN ONB[13]
    PORT
      LAYER Metal2 ;
        RECT 30.03 0 30.32 0.29 ;
    END
  END ONB[13]
  PIN ON[14]
    PORT
      LAYER Metal2 ;
        RECT 31.48 0 31.77 0.29 ;
    END
  END ON[14]
  PIN ONB[14]
    PORT
      LAYER Metal2 ;
        RECT 32.03 0 32.32 0.29 ;
    END
  END ONB[14]
  PIN ON[15]
    PORT
      LAYER Metal2 ;
        RECT 33.48 0 33.77 0.29 ;
    END
  END ON[15]
  PIN ONB[15]
    PORT
      LAYER Metal2 ;
        RECT 34.03 0 34.32 0.29 ;
    END
  END ONB[15]
  PIN ON[16]
    PORT
      LAYER Metal2 ;
        RECT 35.48 0 35.77 0.29 ;
    END
  END ON[16]
  PIN ONB[16]
    PORT
      LAYER Metal2 ;
        RECT 36.03 0 36.32 0.29 ;
    END
  END ONB[16]
  PIN ON[17]
    PORT
      LAYER Metal2 ;
        RECT 37.48 0 37.77 0.29 ;
    END
  END ON[17]
  PIN ONB[17]
    PORT
      LAYER Metal2 ;
        RECT 38.03 0 38.32 0.29 ;
    END
  END ONB[17]
  PIN ON[18]
    PORT
      LAYER Metal2 ;
        RECT 39.48 0 39.77 0.29 ;
    END
  END ON[18]
  PIN ONB[18]
    PORT
      LAYER Metal2 ;
        RECT 40.03 0 40.32 0.29 ;
    END
  END ONB[18]
  PIN ON[19]
    PORT
      LAYER Metal2 ;
        RECT 41.48 0 41.77 0.29 ;
    END
  END ON[19]
  PIN ONB[19]
    PORT
      LAYER Metal2 ;
        RECT 42.03 0 42.32 0.29 ;
    END
  END ONB[19]
  PIN ON[20]
    PORT
      LAYER Metal2 ;
        RECT 43.48 0 43.77 0.29 ;
    END
  END ON[20]
  PIN ONB[20]
    PORT
      LAYER Metal2 ;
        RECT 44.03 0 44.32 0.29 ;
    END
  END ONB[20]
  PIN ON[21]
    PORT
      LAYER Metal2 ;
        RECT 45.48 0 45.77 0.29 ;
    END
  END ON[21]
  PIN ONB[21]
    PORT
      LAYER Metal2 ;
        RECT 46.03 0 46.32 0.29 ;
    END
  END ONB[21]
  PIN ON[22]
    PORT
      LAYER Metal2 ;
        RECT 47.48 0 47.77 0.29 ;
    END
  END ON[22]
  PIN ONB[22]
    PORT
      LAYER Metal2 ;
        RECT 48.03 0 48.32 0.29 ;
    END
  END ONB[22]
  PIN ON[23]
    PORT
      LAYER Metal2 ;
        RECT 49.48 0 49.77 0.29 ;
    END
  END ON[23]
  PIN ONB[23]
    PORT
      LAYER Metal2 ;
        RECT 50.03 0 50.32 0.29 ;
    END
  END ONB[23]
  PIN ON[24]
    PORT
      LAYER Metal2 ;
        RECT 51.48 0 51.77 0.29 ;
    END
  END ON[24]
  PIN ONB[24]
    PORT
      LAYER Metal2 ;
        RECT 52.03 0 52.32 0.29 ;
    END
  END ONB[24]
  PIN ON[25]
    PORT
      LAYER Metal2 ;
        RECT 53.48 0 53.77 0.29 ;
    END
  END ON[25]
  PIN ONB[25]
    PORT
      LAYER Metal2 ;
        RECT 54.03 0 54.32 0.29 ;
    END
  END ONB[25]
  PIN ON[26]
    PORT
      LAYER Metal2 ;
        RECT 55.48 0 55.77 0.29 ;
    END
  END ON[26]
  PIN ONB[26]
    PORT
      LAYER Metal2 ;
        RECT 56.03 0 56.32 0.29 ;
    END
  END ONB[26]
  PIN ON[27]
    PORT
      LAYER Metal2 ;
        RECT 57.48 0 57.77 0.29 ;
    END
  END ON[27]
  PIN ONB[27]
    PORT
      LAYER Metal2 ;
        RECT 58.03 0 58.32 0.29 ;
    END
  END ONB[27]
  PIN ON[28]
    PORT
      LAYER Metal2 ;
        RECT 59.48 0 59.77 0.29 ;
    END
  END ON[28]
  PIN ONB[28]
    PORT
      LAYER Metal2 ;
        RECT 60.03 0 60.32 0.29 ;
    END
  END ONB[28]
  PIN ON[29]
    PORT
      LAYER Metal2 ;
        RECT 61.48 0 61.77 0.29 ;
    END
  END ON[29]
  PIN ONB[29]
    PORT
      LAYER Metal2 ;
        RECT 62.03 0 62.32 0.29 ;
    END
  END ONB[29]
  PIN ON[30]
    PORT
      LAYER Metal2 ;
        RECT 63.48 0 63.77 0.29 ;
    END
  END ON[30]
  PIN ONB[30]
    PORT
      LAYER Metal2 ;
        RECT 64.03 0 64.32 0.29 ;
    END
  END ONB[30]
  PIN ON[31]
    PORT
      LAYER Metal2 ;
        RECT 65.48 0 65.77 0.29 ;
    END
  END ON[31]
  PIN ONB[31]
    PORT
      LAYER Metal2 ;
        RECT 66.03 0 66.32 0.29 ;
    END
  END ONB[31]
  PIN EN[0]
    PORT
      LAYER Metal2 ;
        RECT 1.48 0 1.77 0.29 ;
    END
  END EN[0]
  PIN ENB[0]
    PORT
      LAYER Metal2 ;
        RECT 2.03 0 2.32 0.29 ;
    END
  END ENB[0]
  PIN ON[33]
    PORT
      LAYER Metal2 ;
        RECT 69.48 0 69.77 0.29 ;
    END
  END ON[33]
  PIN ONB[33]
    PORT
      LAYER Metal2 ;
        RECT 70.03 0 70.32 0.29 ;
    END
  END ONB[33]
  PIN ON[34]
    PORT
      LAYER Metal2 ;
        RECT 71.48 0 71.77 0.29 ;
    END
  END ON[34]
  PIN ONB[34]
    PORT
      LAYER Metal2 ;
        RECT 72.03 0 72.32 0.29 ;
    END
  END ONB[34]
  PIN ON[35]
    PORT
      LAYER Metal2 ;
        RECT 73.48 0 73.77 0.29 ;
    END
  END ON[35]
  PIN ONB[35]
    PORT
      LAYER Metal2 ;
        RECT 74.03 0 74.32 0.29 ;
    END
  END ONB[35]
  PIN ON[36]
    PORT
      LAYER Metal2 ;
        RECT 75.48 0 75.77 0.29 ;
    END
  END ON[36]
  PIN ONB[36]
    PORT
      LAYER Metal2 ;
        RECT 76.03 0 76.32 0.29 ;
    END
  END ONB[36]
  PIN ON[37]
    PORT
      LAYER Metal2 ;
        RECT 77.48 0 77.77 0.29 ;
    END
  END ON[37]
  PIN ONB[37]
    PORT
      LAYER Metal2 ;
        RECT 78.03 0 78.32 0.29 ;
    END
  END ONB[37]
  PIN ON[38]
    PORT
      LAYER Metal2 ;
        RECT 79.48 0 79.77 0.29 ;
    END
  END ON[38]
  PIN ONB[38]
    PORT
      LAYER Metal2 ;
        RECT 80.03 0 80.32 0.29 ;
    END
  END ONB[38]
  PIN ON[39]
    PORT
      LAYER Metal2 ;
        RECT 81.48 0 81.77 0.29 ;
    END
  END ON[39]
  PIN ONB[39]
    PORT
      LAYER Metal2 ;
        RECT 82.03 0 82.32 0.29 ;
    END
  END ONB[39]
  PIN ON[40]
    PORT
      LAYER Metal2 ;
        RECT 83.48 0 83.77 0.29 ;
    END
  END ON[40]
  PIN ONB[40]
    PORT
      LAYER Metal2 ;
        RECT 84.03 0 84.32 0.29 ;
    END
  END ONB[40]
  PIN ON[41]
    PORT
      LAYER Metal2 ;
        RECT 85.48 0 85.77 0.29 ;
    END
  END ON[41]
  PIN ONB[41]
    PORT
      LAYER Metal2 ;
        RECT 86.03 0 86.32 0.29 ;
    END
  END ONB[41]
  PIN ON[42]
    PORT
      LAYER Metal2 ;
        RECT 87.48 0 87.77 0.29 ;
    END
  END ON[42]
  PIN ONB[42]
    PORT
      LAYER Metal2 ;
        RECT 88.03 0 88.32 0.29 ;
    END
  END ONB[42]
  PIN ON[43]
    PORT
      LAYER Metal2 ;
        RECT 89.48 0 89.77 0.29 ;
    END
  END ON[43]
  PIN ONB[43]
    PORT
      LAYER Metal2 ;
        RECT 90.03 0 90.32 0.29 ;
    END
  END ONB[43]
  PIN ON[44]
    PORT
      LAYER Metal2 ;
        RECT 91.48 0 91.77 0.29 ;
    END
  END ON[44]
  PIN ONB[44]
    PORT
      LAYER Metal2 ;
        RECT 92.03 0 92.32 0.29 ;
    END
  END ONB[44]
  PIN ON[45]
    PORT
      LAYER Metal2 ;
        RECT 93.48 0 93.77 0.29 ;
    END
  END ON[45]
  PIN ONB[45]
    PORT
      LAYER Metal2 ;
        RECT 94.03 0 94.32 0.29 ;
    END
  END ONB[45]
  PIN ON[46]
    PORT
      LAYER Metal2 ;
        RECT 95.48 0 95.77 0.29 ;
    END
  END ON[46]
  PIN ONB[46]
    PORT
      LAYER Metal2 ;
        RECT 96.03 0 96.32 0.29 ;
    END
  END ONB[46]
  PIN ON[47]
    PORT
      LAYER Metal2 ;
        RECT 97.48 0 97.77 0.29 ;
    END
  END ON[47]
  PIN ONB[47]
    PORT
      LAYER Metal2 ;
        RECT 98.03 0 98.32 0.29 ;
    END
  END ONB[47]
  PIN ON[48]
    PORT
      LAYER Metal2 ;
        RECT 99.48 0 99.77 0.29 ;
    END
  END ON[48]
  PIN ONB[48]
    PORT
      LAYER Metal2 ;
        RECT 100.03 0 100.32 0.29 ;
    END
  END ONB[48]
  PIN ON[49]
    PORT
      LAYER Metal2 ;
        RECT 101.48 0 101.77 0.29 ;
    END
  END ON[49]
  PIN ONB[49]
    PORT
      LAYER Metal2 ;
        RECT 102.03 0 102.32 0.29 ;
    END
  END ONB[49]
  PIN ON[50]
    PORT
      LAYER Metal2 ;
        RECT 103.48 0 103.77 0.29 ;
    END
  END ON[50]
  PIN ONB[50]
    PORT
      LAYER Metal2 ;
        RECT 104.03 0 104.32 0.29 ;
    END
  END ONB[50]
  PIN ON[51]
    PORT
      LAYER Metal2 ;
        RECT 105.48 0 105.77 0.29 ;
    END
  END ON[51]
  PIN ONB[51]
    PORT
      LAYER Metal2 ;
        RECT 106.03 0 106.32 0.29 ;
    END
  END ONB[51]
  PIN ON[52]
    PORT
      LAYER Metal2 ;
        RECT 107.48 0 107.77 0.29 ;
    END
  END ON[52]
  PIN ONB[52]
    PORT
      LAYER Metal2 ;
        RECT 108.03 0 108.32 0.29 ;
    END
  END ONB[52]
  PIN ON[53]
    PORT
      LAYER Metal2 ;
        RECT 109.48 0 109.77 0.29 ;
    END
  END ON[53]
  PIN ONB[53]
    PORT
      LAYER Metal2 ;
        RECT 110.03 0 110.32 0.29 ;
    END
  END ONB[53]
  PIN ON[54]
    PORT
      LAYER Metal2 ;
        RECT 111.48 0 111.77 0.29 ;
    END
  END ON[54]
  PIN ONB[54]
    PORT
      LAYER Metal2 ;
        RECT 112.03 0 112.32 0.29 ;
    END
  END ONB[54]
  PIN ON[55]
    PORT
      LAYER Metal2 ;
        RECT 113.48 0 113.77 0.29 ;
    END
  END ON[55]
  PIN ONB[55]
    PORT
      LAYER Metal2 ;
        RECT 114.03 0 114.32 0.29 ;
    END
  END ONB[55]
  PIN ON[56]
    PORT
      LAYER Metal2 ;
        RECT 115.48 0 115.77 0.29 ;
    END
  END ON[56]
  PIN ONB[56]
    PORT
      LAYER Metal2 ;
        RECT 116.03 0 116.32 0.29 ;
    END
  END ONB[56]
  PIN ON[57]
    PORT
      LAYER Metal2 ;
        RECT 117.48 0 117.77 0.29 ;
    END
  END ON[57]
  PIN ONB[57]
    PORT
      LAYER Metal2 ;
        RECT 118.03 0 118.32 0.29 ;
    END
  END ONB[57]
  PIN ON[58]
    PORT
      LAYER Metal2 ;
        RECT 119.48 0 119.77 0.29 ;
    END
  END ON[58]
  PIN ONB[58]
    PORT
      LAYER Metal2 ;
        RECT 120.03 0 120.32 0.29 ;
    END
  END ONB[58]
  PIN ON[59]
    PORT
      LAYER Metal2 ;
        RECT 121.48 0 121.77 0.29 ;
    END
  END ON[59]
  PIN ONB[59]
    PORT
      LAYER Metal2 ;
        RECT 122.03 0 122.32 0.29 ;
    END
  END ONB[59]
  PIN ON[60]
    PORT
      LAYER Metal2 ;
        RECT 123.48 0 123.77 0.29 ;
    END
  END ON[60]
  PIN ONB[60]
    PORT
      LAYER Metal2 ;
        RECT 124.03 0 124.32 0.29 ;
    END
  END ONB[60]
  PIN ON[61]
    PORT
      LAYER Metal2 ;
        RECT 125.48 0 125.77 0.29 ;
    END
  END ON[61]
  PIN ONB[61]
    PORT
      LAYER Metal2 ;
        RECT 126.03 0 126.32 0.29 ;
    END
  END ONB[61]
  PIN ON[62]
    PORT
      LAYER Metal2 ;
        RECT 127.48 0 127.77 0.29 ;
    END
  END ON[62]
  PIN ONB[62]
    PORT
      LAYER Metal2 ;
        RECT 128.03 0 128.32 0.29 ;
    END
  END ONB[62]
  PIN ON[63]
    PORT
      LAYER Metal2 ;
        RECT 129.48 0 129.77 0.29 ;
    END
  END ON[63]
  PIN ONB[63]
    PORT
      LAYER Metal2 ;
        RECT 130.03 0 130.32 0.29 ;
    END
  END ONB[63]
  PIN ON[32]
    PORT
      LAYER Metal2 ;
        RECT 67.48 0 67.77 0.29 ;
    END
  END ON[32]
  PIN ONB[32]
    PORT
      LAYER Metal2 ;
        RECT 68.03 0 68.32 0.29 ;
    END
  END ONB[32]
  PIN EN[1]
    PORT
      LAYER Metal2 ;
        RECT 131.48 0 131.77 0.29 ;
    END
  END EN[1]
  PIN ENB[1]
    PORT
      LAYER Metal2 ;
        RECT 132.03 0 132.32 0.29 ;
    END
  END ENB[1]
#  PIN VcascP[1]
#    PORT
#      LAYER Metal3 ;
#        RECT 0 20.93 133.8 21.63 ;
#    END
#  END VcascP[1]
#  PIN VcascP[0]
#    PORT
#      LAYER Metal3 ;
#        RECT 0 4.56 133.8 5.26 ;
#    END
#  END VcascP[0]
END dac2u128out4in
END LIBRARY

