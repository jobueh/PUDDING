** sch_path: /home/cmaier/EDA/PUDDING/xschem/pcascsrc16.sch
.subckt pcascsrc16 Vcp[15] Vcp[14] Vcp[13] Vcp[12] Vcp[11] Vcp[10] Vcp[9] Vcp[8] Vcp[7] Vcp[6] Vcp[5] Vcp[4] Vcp[3] Vcp[2] Vcp[1]
+ Vcp[0] Vbp Iout VDD
*.PININFO Vcp[15:0]:I Vbp:I Iout:O VDD:I
xsrc[15] VDD Vbp Vcp[15] Iout VDD pcascsrc
xsrc[14] VDD Vbp Vcp[14] Iout VDD pcascsrc
xsrc[13] VDD Vbp Vcp[13] Iout VDD pcascsrc
xsrc[12] VDD Vbp Vcp[12] Iout VDD pcascsrc
xsrc[11] VDD Vbp Vcp[11] Iout VDD pcascsrc
xsrc[10] VDD Vbp Vcp[10] Iout VDD pcascsrc
xsrc[9] VDD Vbp Vcp[9] Iout VDD pcascsrc
xsrc[8] VDD Vbp Vcp[8] Iout VDD pcascsrc
xsrc[7] VDD Vbp Vcp[7] Iout VDD pcascsrc
xsrc[6] VDD Vbp Vcp[6] Iout VDD pcascsrc
xsrc[5] VDD Vbp Vcp[5] Iout VDD pcascsrc
xsrc[4] VDD Vbp Vcp[4] Iout VDD pcascsrc
xsrc[3] VDD Vbp Vcp[3] Iout VDD pcascsrc
xsrc[2] VDD Vbp Vcp[2] Iout VDD pcascsrc
xsrc[1] VDD Vbp Vcp[1] Iout VDD pcascsrc
xsrc[0] VDD Vbp Vcp[0] Iout VDD pcascsrc
.ends

* expanding   symbol:  pcascsrc.sym # of pins=5
** sym_path: /home/cmaier/EDA/PUDDING/xschem/pcascsrc.sym
** sch_path: /home/cmaier/EDA/PUDDING/xschem/pcascsrc.sch
.subckt pcascsrc VDD VbiasP VcascodeP Iout NWELL
*.PININFO VcascodeP:I VbiasP:I Iout:O VDD:I NWELL:B
Msrc drain VbiasP VDD NWELL sg13_lv_pmos w=0.74u l=2u ng=1 m=1
Mcasc Iout VcascodeP drain NWELL sg13_lv_pmos w=0.3u l=0.3u ng=1 m=1
.ends

