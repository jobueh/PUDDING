module heichips25_pudding (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire \daisychain[0] ;
 wire \daisychain[100] ;
 wire \daisychain[101] ;
 wire \daisychain[102] ;
 wire \daisychain[103] ;
 wire \daisychain[104] ;
 wire \daisychain[105] ;
 wire \daisychain[106] ;
 wire \daisychain[107] ;
 wire \daisychain[108] ;
 wire \daisychain[109] ;
 wire \daisychain[10] ;
 wire \daisychain[110] ;
 wire \daisychain[111] ;
 wire \daisychain[112] ;
 wire \daisychain[113] ;
 wire \daisychain[114] ;
 wire \daisychain[115] ;
 wire \daisychain[116] ;
 wire \daisychain[117] ;
 wire \daisychain[118] ;
 wire \daisychain[119] ;
 wire \daisychain[11] ;
 wire \daisychain[120] ;
 wire \daisychain[121] ;
 wire \daisychain[122] ;
 wire \daisychain[123] ;
 wire \daisychain[124] ;
 wire \daisychain[125] ;
 wire \daisychain[126] ;
 wire \daisychain[127] ;
 wire \daisychain[12] ;
 wire \daisychain[13] ;
 wire \daisychain[14] ;
 wire \daisychain[15] ;
 wire \daisychain[16] ;
 wire \daisychain[17] ;
 wire \daisychain[18] ;
 wire \daisychain[19] ;
 wire \daisychain[1] ;
 wire \daisychain[20] ;
 wire \daisychain[21] ;
 wire \daisychain[22] ;
 wire \daisychain[23] ;
 wire \daisychain[24] ;
 wire \daisychain[25] ;
 wire \daisychain[26] ;
 wire \daisychain[27] ;
 wire \daisychain[28] ;
 wire \daisychain[29] ;
 wire \daisychain[2] ;
 wire \daisychain[30] ;
 wire \daisychain[31] ;
 wire \daisychain[32] ;
 wire \daisychain[33] ;
 wire \daisychain[34] ;
 wire \daisychain[35] ;
 wire \daisychain[36] ;
 wire \daisychain[37] ;
 wire \daisychain[38] ;
 wire \daisychain[39] ;
 wire \daisychain[3] ;
 wire \daisychain[40] ;
 wire \daisychain[41] ;
 wire \daisychain[42] ;
 wire \daisychain[43] ;
 wire \daisychain[44] ;
 wire \daisychain[45] ;
 wire \daisychain[46] ;
 wire \daisychain[47] ;
 wire \daisychain[48] ;
 wire \daisychain[49] ;
 wire \daisychain[4] ;
 wire \daisychain[50] ;
 wire \daisychain[51] ;
 wire \daisychain[52] ;
 wire \daisychain[53] ;
 wire \daisychain[54] ;
 wire \daisychain[55] ;
 wire \daisychain[56] ;
 wire \daisychain[57] ;
 wire \daisychain[58] ;
 wire \daisychain[59] ;
 wire \daisychain[5] ;
 wire \daisychain[60] ;
 wire \daisychain[61] ;
 wire \daisychain[62] ;
 wire \daisychain[63] ;
 wire \daisychain[64] ;
 wire \daisychain[65] ;
 wire \daisychain[66] ;
 wire \daisychain[67] ;
 wire \daisychain[68] ;
 wire \daisychain[69] ;
 wire \daisychain[6] ;
 wire \daisychain[70] ;
 wire \daisychain[71] ;
 wire \daisychain[72] ;
 wire \daisychain[73] ;
 wire \daisychain[74] ;
 wire \daisychain[75] ;
 wire \daisychain[76] ;
 wire \daisychain[77] ;
 wire \daisychain[78] ;
 wire \daisychain[79] ;
 wire \daisychain[7] ;
 wire \daisychain[80] ;
 wire \daisychain[81] ;
 wire \daisychain[82] ;
 wire \daisychain[83] ;
 wire \daisychain[84] ;
 wire \daisychain[85] ;
 wire \daisychain[86] ;
 wire \daisychain[87] ;
 wire \daisychain[88] ;
 wire \daisychain[89] ;
 wire \daisychain[8] ;
 wire \daisychain[90] ;
 wire \daisychain[91] ;
 wire \daisychain[92] ;
 wire \daisychain[93] ;
 wire \daisychain[94] ;
 wire \daisychain[95] ;
 wire \daisychain[96] ;
 wire \daisychain[97] ;
 wire \daisychain[98] ;
 wire \daisychain[99] ;
 wire \daisychain[9] ;
 wire \digitalenH.g[0].u.OUTN ;
 wire \digitalenH.g[0].u.OUTP ;
 wire \digitalenH.g[1].u.OUTN ;
 wire \digitalenH.g[1].u.OUTP ;
 wire \digitalenH.g[2].u.OUTN ;
 wire \digitalenH.g[2].u.OUTP ;
 wire \digitalenH.g[3].u.OUTN ;
 wire \digitalenH.g[3].u.OUTP ;
 wire \digitalenL.g[0].u.OUTN ;
 wire \digitalenL.g[0].u.OUTP ;
 wire \digitalenL.g[1].u.OUTN ;
 wire \digitalenL.g[1].u.OUTP ;
 wire \digitalenL.g[2].u.OUTN ;
 wire \digitalenL.g[2].u.OUTP ;
 wire \digitalenL.g[3].u.OUTN ;
 wire \digitalenL.g[3].u.OUTP ;
 wire net1;
 wire \state[0] ;
 wire \state[100] ;
 wire \state[101] ;
 wire \state[102] ;
 wire \state[103] ;
 wire \state[104] ;
 wire \state[105] ;
 wire \state[106] ;
 wire \state[107] ;
 wire \state[108] ;
 wire \state[109] ;
 wire \state[10] ;
 wire \state[110] ;
 wire \state[111] ;
 wire \state[112] ;
 wire \state[113] ;
 wire \state[114] ;
 wire \state[115] ;
 wire \state[116] ;
 wire \state[117] ;
 wire \state[118] ;
 wire \state[119] ;
 wire \state[11] ;
 wire \state[120] ;
 wire \state[121] ;
 wire \state[122] ;
 wire \state[123] ;
 wire \state[124] ;
 wire \state[125] ;
 wire \state[126] ;
 wire \state[127] ;
 wire \state[12] ;
 wire \state[13] ;
 wire \state[14] ;
 wire \state[15] ;
 wire \state[16] ;
 wire \state[17] ;
 wire \state[18] ;
 wire \state[19] ;
 wire \state[1] ;
 wire \state[20] ;
 wire \state[21] ;
 wire \state[22] ;
 wire \state[23] ;
 wire \state[24] ;
 wire \state[25] ;
 wire \state[26] ;
 wire \state[27] ;
 wire \state[28] ;
 wire \state[29] ;
 wire \state[2] ;
 wire \state[30] ;
 wire \state[31] ;
 wire \state[32] ;
 wire \state[33] ;
 wire \state[34] ;
 wire \state[35] ;
 wire \state[36] ;
 wire \state[37] ;
 wire \state[38] ;
 wire \state[39] ;
 wire \state[3] ;
 wire \state[40] ;
 wire \state[41] ;
 wire \state[42] ;
 wire \state[43] ;
 wire \state[44] ;
 wire \state[45] ;
 wire \state[46] ;
 wire \state[47] ;
 wire \state[48] ;
 wire \state[49] ;
 wire \state[4] ;
 wire \state[50] ;
 wire \state[51] ;
 wire \state[52] ;
 wire \state[53] ;
 wire \state[54] ;
 wire \state[55] ;
 wire \state[56] ;
 wire \state[57] ;
 wire \state[58] ;
 wire \state[59] ;
 wire \state[5] ;
 wire \state[60] ;
 wire \state[61] ;
 wire \state[62] ;
 wire \state[63] ;
 wire \state[64] ;
 wire \state[65] ;
 wire \state[66] ;
 wire \state[67] ;
 wire \state[68] ;
 wire \state[69] ;
 wire \state[6] ;
 wire \state[70] ;
 wire \state[71] ;
 wire \state[72] ;
 wire \state[73] ;
 wire \state[74] ;
 wire \state[75] ;
 wire \state[76] ;
 wire \state[77] ;
 wire \state[78] ;
 wire \state[79] ;
 wire \state[7] ;
 wire \state[80] ;
 wire \state[81] ;
 wire \state[82] ;
 wire \state[83] ;
 wire \state[84] ;
 wire \state[85] ;
 wire \state[86] ;
 wire \state[87] ;
 wire \state[88] ;
 wire \state[89] ;
 wire \state[8] ;
 wire \state[90] ;
 wire \state[91] ;
 wire \state[92] ;
 wire \state[93] ;
 wire \state[94] ;
 wire \state[95] ;
 wire \state[96] ;
 wire \state[97] ;
 wire \state[98] ;
 wire \state[99] ;
 wire \state[9] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire clknet_leaf_0_clk;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_inv_1 _1283_ (.Y(_0030_),
    .A(\state[127] ));
 sg13g2_inv_1 _1284_ (.Y(_1026_),
    .A(net211));
 sg13g2_inv_1 _1285_ (.Y(_0029_),
    .A(\state[126] ));
 sg13g2_inv_1 _1286_ (.Y(_0028_),
    .A(\state[125] ));
 sg13g2_inv_1 _1287_ (.Y(_0027_),
    .A(\state[124] ));
 sg13g2_inv_1 _1288_ (.Y(_0026_),
    .A(\state[123] ));
 sg13g2_inv_1 _1289_ (.Y(_0025_),
    .A(\state[122] ));
 sg13g2_inv_1 _1290_ (.Y(_0024_),
    .A(\state[121] ));
 sg13g2_inv_1 _1291_ (.Y(_0023_),
    .A(\state[120] ));
 sg13g2_inv_1 _1292_ (.Y(_0021_),
    .A(\state[119] ));
 sg13g2_inv_1 _1293_ (.Y(_0020_),
    .A(\state[118] ));
 sg13g2_inv_1 _1294_ (.Y(_0019_),
    .A(\state[117] ));
 sg13g2_inv_1 _1295_ (.Y(_0018_),
    .A(\state[116] ));
 sg13g2_inv_1 _1296_ (.Y(_0017_),
    .A(\state[115] ));
 sg13g2_inv_1 _1297_ (.Y(_0016_),
    .A(\state[114] ));
 sg13g2_inv_1 _1298_ (.Y(_0015_),
    .A(\state[113] ));
 sg13g2_inv_1 _1299_ (.Y(_0014_),
    .A(\state[112] ));
 sg13g2_inv_1 _1300_ (.Y(_0013_),
    .A(\state[111] ));
 sg13g2_inv_1 _1301_ (.Y(_0012_),
    .A(\state[110] ));
 sg13g2_inv_1 _1302_ (.Y(_0010_),
    .A(\state[109] ));
 sg13g2_inv_1 _1303_ (.Y(_0009_),
    .A(\state[108] ));
 sg13g2_inv_1 _1304_ (.Y(_0008_),
    .A(\state[107] ));
 sg13g2_inv_1 _1305_ (.Y(_0007_),
    .A(\state[106] ));
 sg13g2_inv_1 _1306_ (.Y(_0006_),
    .A(\state[105] ));
 sg13g2_inv_1 _1307_ (.Y(_0005_),
    .A(\state[104] ));
 sg13g2_inv_1 _1308_ (.Y(_0004_),
    .A(\state[103] ));
 sg13g2_inv_1 _1309_ (.Y(_0003_),
    .A(\state[102] ));
 sg13g2_inv_1 _1310_ (.Y(_0002_),
    .A(\state[101] ));
 sg13g2_inv_1 _1311_ (.Y(_0001_),
    .A(\state[100] ));
 sg13g2_inv_1 _1312_ (.Y(_0126_),
    .A(\state[99] ));
 sg13g2_inv_1 _1313_ (.Y(_0125_),
    .A(\state[98] ));
 sg13g2_inv_1 _1314_ (.Y(_0124_),
    .A(\state[97] ));
 sg13g2_inv_1 _1315_ (.Y(_0123_),
    .A(\state[96] ));
 sg13g2_inv_1 _1316_ (.Y(_0122_),
    .A(\state[95] ));
 sg13g2_inv_1 _1317_ (.Y(_0121_),
    .A(\state[94] ));
 sg13g2_inv_1 _1318_ (.Y(_0120_),
    .A(\state[93] ));
 sg13g2_inv_1 _1319_ (.Y(_0119_),
    .A(\state[92] ));
 sg13g2_inv_1 _1320_ (.Y(_0118_),
    .A(\state[91] ));
 sg13g2_inv_1 _1321_ (.Y(_0117_),
    .A(\state[90] ));
 sg13g2_inv_1 _1322_ (.Y(_0115_),
    .A(\state[89] ));
 sg13g2_inv_1 _1323_ (.Y(_0114_),
    .A(\state[88] ));
 sg13g2_inv_1 _1324_ (.Y(_0113_),
    .A(\state[87] ));
 sg13g2_inv_1 _1325_ (.Y(_0112_),
    .A(\state[86] ));
 sg13g2_inv_1 _1326_ (.Y(_0111_),
    .A(\state[85] ));
 sg13g2_inv_1 _1327_ (.Y(_0110_),
    .A(\state[84] ));
 sg13g2_inv_1 _1328_ (.Y(_0109_),
    .A(\state[83] ));
 sg13g2_inv_1 _1329_ (.Y(_0108_),
    .A(\state[82] ));
 sg13g2_inv_1 _1330_ (.Y(_0107_),
    .A(\state[81] ));
 sg13g2_inv_1 _1331_ (.Y(_0106_),
    .A(\state[80] ));
 sg13g2_inv_1 _1332_ (.Y(_0104_),
    .A(\state[79] ));
 sg13g2_inv_1 _1333_ (.Y(_0103_),
    .A(\state[78] ));
 sg13g2_inv_1 _1334_ (.Y(_0102_),
    .A(\state[77] ));
 sg13g2_inv_1 _1335_ (.Y(_0101_),
    .A(\state[76] ));
 sg13g2_inv_1 _1336_ (.Y(_0100_),
    .A(\state[75] ));
 sg13g2_inv_1 _1337_ (.Y(_0099_),
    .A(\state[74] ));
 sg13g2_inv_1 _1338_ (.Y(_0098_),
    .A(\state[73] ));
 sg13g2_inv_1 _1339_ (.Y(_0097_),
    .A(\state[72] ));
 sg13g2_inv_1 _1340_ (.Y(_0096_),
    .A(\state[71] ));
 sg13g2_inv_1 _1341_ (.Y(_0095_),
    .A(\state[70] ));
 sg13g2_inv_1 _1342_ (.Y(_0093_),
    .A(\state[69] ));
 sg13g2_inv_1 _1343_ (.Y(_0092_),
    .A(\state[68] ));
 sg13g2_inv_1 _1344_ (.Y(_0091_),
    .A(\state[67] ));
 sg13g2_inv_1 _1345_ (.Y(_0090_),
    .A(\state[66] ));
 sg13g2_inv_1 _1346_ (.Y(_0089_),
    .A(\state[65] ));
 sg13g2_inv_1 _1347_ (.Y(_0088_),
    .A(\state[64] ));
 sg13g2_inv_1 _1348_ (.Y(_0087_),
    .A(\state[63] ));
 sg13g2_inv_1 _1349_ (.Y(_0086_),
    .A(\state[62] ));
 sg13g2_inv_1 _1350_ (.Y(_0085_),
    .A(\state[61] ));
 sg13g2_inv_1 _1351_ (.Y(_0084_),
    .A(\state[60] ));
 sg13g2_inv_1 _1352_ (.Y(_0082_),
    .A(\state[59] ));
 sg13g2_inv_1 _1353_ (.Y(_0081_),
    .A(\state[58] ));
 sg13g2_inv_1 _1354_ (.Y(_0080_),
    .A(\state[57] ));
 sg13g2_inv_1 _1355_ (.Y(_0079_),
    .A(\state[56] ));
 sg13g2_inv_1 _1356_ (.Y(_0078_),
    .A(\state[55] ));
 sg13g2_inv_1 _1357_ (.Y(_0077_),
    .A(\state[54] ));
 sg13g2_inv_1 _1358_ (.Y(_0076_),
    .A(\state[53] ));
 sg13g2_inv_1 _1359_ (.Y(_0075_),
    .A(\state[52] ));
 sg13g2_inv_1 _1360_ (.Y(_0074_),
    .A(\state[51] ));
 sg13g2_inv_1 _1361_ (.Y(_0073_),
    .A(\state[50] ));
 sg13g2_inv_1 _1362_ (.Y(_0071_),
    .A(\state[49] ));
 sg13g2_inv_1 _1363_ (.Y(_0070_),
    .A(\state[48] ));
 sg13g2_inv_1 _1364_ (.Y(_0069_),
    .A(\state[47] ));
 sg13g2_inv_1 _1365_ (.Y(_0068_),
    .A(\state[46] ));
 sg13g2_inv_1 _1366_ (.Y(_0067_),
    .A(\state[45] ));
 sg13g2_inv_1 _1367_ (.Y(_0066_),
    .A(\state[44] ));
 sg13g2_inv_1 _1368_ (.Y(_0065_),
    .A(\state[43] ));
 sg13g2_inv_1 _1369_ (.Y(_0064_),
    .A(\state[42] ));
 sg13g2_inv_1 _1370_ (.Y(_0063_),
    .A(\state[41] ));
 sg13g2_inv_1 _1371_ (.Y(_0062_),
    .A(\state[40] ));
 sg13g2_inv_1 _1372_ (.Y(_0060_),
    .A(\state[39] ));
 sg13g2_inv_1 _1373_ (.Y(_0059_),
    .A(\state[38] ));
 sg13g2_inv_1 _1374_ (.Y(_0058_),
    .A(\state[37] ));
 sg13g2_inv_1 _1375_ (.Y(_0057_),
    .A(\state[36] ));
 sg13g2_inv_1 _1376_ (.Y(_0056_),
    .A(\state[35] ));
 sg13g2_inv_1 _1377_ (.Y(_0055_),
    .A(\state[34] ));
 sg13g2_inv_1 _1378_ (.Y(_0054_),
    .A(\state[33] ));
 sg13g2_inv_1 _1379_ (.Y(_0053_),
    .A(\state[32] ));
 sg13g2_inv_1 _1380_ (.Y(_0052_),
    .A(\state[31] ));
 sg13g2_inv_1 _1381_ (.Y(_0051_),
    .A(\state[30] ));
 sg13g2_inv_1 _1382_ (.Y(_0049_),
    .A(\state[29] ));
 sg13g2_inv_1 _1383_ (.Y(_0048_),
    .A(\state[28] ));
 sg13g2_inv_1 _1384_ (.Y(_0047_),
    .A(\state[27] ));
 sg13g2_inv_1 _1385_ (.Y(_0046_),
    .A(\state[26] ));
 sg13g2_inv_1 _1386_ (.Y(_0045_),
    .A(\state[25] ));
 sg13g2_inv_1 _1387_ (.Y(_0044_),
    .A(\state[24] ));
 sg13g2_inv_1 _1388_ (.Y(_0043_),
    .A(\state[23] ));
 sg13g2_inv_1 _1389_ (.Y(_0042_),
    .A(\state[22] ));
 sg13g2_inv_1 _1390_ (.Y(_0041_),
    .A(\state[21] ));
 sg13g2_inv_1 _1391_ (.Y(_0040_),
    .A(\state[20] ));
 sg13g2_inv_1 _1392_ (.Y(_0038_),
    .A(\state[19] ));
 sg13g2_inv_1 _1393_ (.Y(_0037_),
    .A(\state[18] ));
 sg13g2_inv_1 _1394_ (.Y(_0036_),
    .A(\state[17] ));
 sg13g2_inv_1 _1395_ (.Y(_0035_),
    .A(\state[16] ));
 sg13g2_inv_1 _1396_ (.Y(_0034_),
    .A(\state[15] ));
 sg13g2_inv_1 _1397_ (.Y(_0033_),
    .A(\state[14] ));
 sg13g2_inv_1 _1398_ (.Y(_0032_),
    .A(\state[13] ));
 sg13g2_inv_1 _1399_ (.Y(_0031_),
    .A(\state[12] ));
 sg13g2_inv_1 _1400_ (.Y(_0022_),
    .A(\state[11] ));
 sg13g2_inv_1 _1401_ (.Y(_0011_),
    .A(\state[10] ));
 sg13g2_inv_1 _1402_ (.Y(_0127_),
    .A(\state[9] ));
 sg13g2_inv_1 _1403_ (.Y(_0116_),
    .A(\state[8] ));
 sg13g2_inv_1 _1404_ (.Y(_0105_),
    .A(\state[7] ));
 sg13g2_inv_1 _1405_ (.Y(_0094_),
    .A(\state[6] ));
 sg13g2_inv_1 _1406_ (.Y(_0083_),
    .A(\state[5] ));
 sg13g2_inv_1 _1407_ (.Y(_0072_),
    .A(\state[4] ));
 sg13g2_inv_1 _1408_ (.Y(_0061_),
    .A(\state[3] ));
 sg13g2_inv_1 _1409_ (.Y(_0050_),
    .A(\state[2] ));
 sg13g2_inv_1 _1410_ (.Y(_0039_),
    .A(\state[1] ));
 sg13g2_inv_1 _1411_ (.Y(_0000_),
    .A(\state[0] ));
 sg13g2_inv_1 _1412_ (.Y(_0158_),
    .A(\daisychain[127] ));
 sg13g2_inv_1 _1413_ (.Y(_0157_),
    .A(\daisychain[126] ));
 sg13g2_inv_1 _1414_ (.Y(_0156_),
    .A(\daisychain[125] ));
 sg13g2_inv_1 _1415_ (.Y(_0155_),
    .A(\daisychain[124] ));
 sg13g2_inv_1 _1416_ (.Y(_0154_),
    .A(\daisychain[123] ));
 sg13g2_inv_1 _1417_ (.Y(_0153_),
    .A(\daisychain[122] ));
 sg13g2_inv_1 _1418_ (.Y(_0152_),
    .A(\daisychain[121] ));
 sg13g2_inv_1 _1419_ (.Y(_0151_),
    .A(\daisychain[120] ));
 sg13g2_inv_1 _1420_ (.Y(_0149_),
    .A(\daisychain[119] ));
 sg13g2_inv_1 _1421_ (.Y(_0148_),
    .A(\daisychain[118] ));
 sg13g2_inv_1 _1422_ (.Y(_0147_),
    .A(\daisychain[117] ));
 sg13g2_inv_1 _1423_ (.Y(_0146_),
    .A(\daisychain[116] ));
 sg13g2_inv_1 _1424_ (.Y(_0145_),
    .A(\daisychain[115] ));
 sg13g2_inv_1 _1425_ (.Y(_0144_),
    .A(\daisychain[114] ));
 sg13g2_inv_1 _1426_ (.Y(_0143_),
    .A(\daisychain[113] ));
 sg13g2_inv_1 _1427_ (.Y(_0142_),
    .A(\daisychain[112] ));
 sg13g2_inv_1 _1428_ (.Y(_0141_),
    .A(\daisychain[111] ));
 sg13g2_inv_1 _1429_ (.Y(_0140_),
    .A(\daisychain[110] ));
 sg13g2_inv_1 _1430_ (.Y(_0138_),
    .A(\daisychain[109] ));
 sg13g2_inv_1 _1431_ (.Y(_0137_),
    .A(\daisychain[108] ));
 sg13g2_inv_1 _1432_ (.Y(_0136_),
    .A(\daisychain[107] ));
 sg13g2_inv_1 _1433_ (.Y(_0135_),
    .A(\daisychain[106] ));
 sg13g2_inv_1 _1434_ (.Y(_0134_),
    .A(\daisychain[105] ));
 sg13g2_inv_1 _1435_ (.Y(_0133_),
    .A(\daisychain[104] ));
 sg13g2_inv_1 _1436_ (.Y(_0132_),
    .A(\daisychain[103] ));
 sg13g2_inv_1 _1437_ (.Y(_0131_),
    .A(\daisychain[102] ));
 sg13g2_inv_1 _1438_ (.Y(_0130_),
    .A(\daisychain[101] ));
 sg13g2_inv_1 _1439_ (.Y(_0129_),
    .A(\daisychain[100] ));
 sg13g2_inv_1 _1440_ (.Y(_0254_),
    .A(\daisychain[99] ));
 sg13g2_inv_1 _1441_ (.Y(_0253_),
    .A(\daisychain[98] ));
 sg13g2_inv_1 _1442_ (.Y(_0252_),
    .A(\daisychain[97] ));
 sg13g2_inv_1 _1443_ (.Y(_0251_),
    .A(\daisychain[96] ));
 sg13g2_inv_1 _1444_ (.Y(_0250_),
    .A(\daisychain[95] ));
 sg13g2_inv_1 _1445_ (.Y(_0249_),
    .A(\daisychain[94] ));
 sg13g2_inv_1 _1446_ (.Y(_0248_),
    .A(\daisychain[93] ));
 sg13g2_inv_1 _1447_ (.Y(_0247_),
    .A(\daisychain[92] ));
 sg13g2_inv_1 _1448_ (.Y(_0246_),
    .A(\daisychain[91] ));
 sg13g2_inv_1 _1449_ (.Y(_0245_),
    .A(\daisychain[90] ));
 sg13g2_inv_1 _1450_ (.Y(_0243_),
    .A(\daisychain[89] ));
 sg13g2_inv_1 _1451_ (.Y(_0242_),
    .A(\daisychain[88] ));
 sg13g2_inv_1 _1452_ (.Y(_0241_),
    .A(\daisychain[87] ));
 sg13g2_inv_1 _1453_ (.Y(_0240_),
    .A(\daisychain[86] ));
 sg13g2_inv_1 _1454_ (.Y(_0239_),
    .A(\daisychain[85] ));
 sg13g2_inv_1 _1455_ (.Y(_0238_),
    .A(\daisychain[84] ));
 sg13g2_inv_1 _1456_ (.Y(_0237_),
    .A(\daisychain[83] ));
 sg13g2_inv_1 _1457_ (.Y(_0236_),
    .A(\daisychain[82] ));
 sg13g2_inv_1 _1458_ (.Y(_0235_),
    .A(\daisychain[81] ));
 sg13g2_inv_1 _1459_ (.Y(_0234_),
    .A(\daisychain[80] ));
 sg13g2_inv_1 _1460_ (.Y(_0232_),
    .A(\daisychain[79] ));
 sg13g2_inv_1 _1461_ (.Y(_0231_),
    .A(\daisychain[78] ));
 sg13g2_inv_1 _1462_ (.Y(_0230_),
    .A(\daisychain[77] ));
 sg13g2_inv_1 _1463_ (.Y(_0229_),
    .A(\daisychain[76] ));
 sg13g2_inv_1 _1464_ (.Y(_0228_),
    .A(\daisychain[75] ));
 sg13g2_inv_1 _1465_ (.Y(_0227_),
    .A(\daisychain[74] ));
 sg13g2_inv_1 _1466_ (.Y(_0226_),
    .A(\daisychain[73] ));
 sg13g2_inv_1 _1467_ (.Y(_0225_),
    .A(\daisychain[72] ));
 sg13g2_inv_1 _1468_ (.Y(_0224_),
    .A(\daisychain[71] ));
 sg13g2_inv_1 _1469_ (.Y(_0223_),
    .A(\daisychain[70] ));
 sg13g2_inv_1 _1470_ (.Y(_0221_),
    .A(\daisychain[69] ));
 sg13g2_inv_1 _1471_ (.Y(_0220_),
    .A(\daisychain[68] ));
 sg13g2_inv_1 _1472_ (.Y(_0219_),
    .A(\daisychain[67] ));
 sg13g2_inv_1 _1473_ (.Y(_0218_),
    .A(\daisychain[66] ));
 sg13g2_inv_1 _1474_ (.Y(_0217_),
    .A(\daisychain[65] ));
 sg13g2_inv_1 _1475_ (.Y(_0216_),
    .A(\daisychain[64] ));
 sg13g2_inv_1 _1476_ (.Y(_0215_),
    .A(\daisychain[63] ));
 sg13g2_inv_1 _1477_ (.Y(_0214_),
    .A(\daisychain[62] ));
 sg13g2_inv_1 _1478_ (.Y(_0213_),
    .A(\daisychain[61] ));
 sg13g2_inv_1 _1479_ (.Y(_0212_),
    .A(\daisychain[60] ));
 sg13g2_inv_1 _1480_ (.Y(_0210_),
    .A(\daisychain[59] ));
 sg13g2_inv_1 _1481_ (.Y(_0209_),
    .A(\daisychain[58] ));
 sg13g2_inv_1 _1482_ (.Y(_0208_),
    .A(\daisychain[57] ));
 sg13g2_inv_1 _1483_ (.Y(_0207_),
    .A(\daisychain[56] ));
 sg13g2_inv_1 _1484_ (.Y(_0206_),
    .A(\daisychain[55] ));
 sg13g2_inv_1 _1485_ (.Y(_0205_),
    .A(\daisychain[54] ));
 sg13g2_inv_1 _1486_ (.Y(_0204_),
    .A(\daisychain[53] ));
 sg13g2_inv_1 _1487_ (.Y(_0203_),
    .A(\daisychain[52] ));
 sg13g2_inv_1 _1488_ (.Y(_0202_),
    .A(\daisychain[51] ));
 sg13g2_inv_1 _1489_ (.Y(_0201_),
    .A(\daisychain[50] ));
 sg13g2_inv_1 _1490_ (.Y(_0199_),
    .A(\daisychain[49] ));
 sg13g2_inv_1 _1491_ (.Y(_0198_),
    .A(\daisychain[48] ));
 sg13g2_inv_1 _1492_ (.Y(_0197_),
    .A(\daisychain[47] ));
 sg13g2_inv_1 _1493_ (.Y(_0196_),
    .A(\daisychain[46] ));
 sg13g2_inv_1 _1494_ (.Y(_0195_),
    .A(\daisychain[45] ));
 sg13g2_inv_1 _1495_ (.Y(_0194_),
    .A(\daisychain[44] ));
 sg13g2_inv_1 _1496_ (.Y(_0193_),
    .A(\daisychain[43] ));
 sg13g2_inv_1 _1497_ (.Y(_0192_),
    .A(\daisychain[42] ));
 sg13g2_inv_1 _1498_ (.Y(_0191_),
    .A(\daisychain[41] ));
 sg13g2_inv_1 _1499_ (.Y(_0190_),
    .A(\daisychain[40] ));
 sg13g2_inv_1 _1500_ (.Y(_0188_),
    .A(\daisychain[39] ));
 sg13g2_inv_1 _1501_ (.Y(_0187_),
    .A(\daisychain[38] ));
 sg13g2_inv_1 _1502_ (.Y(_0186_),
    .A(\daisychain[37] ));
 sg13g2_inv_1 _1503_ (.Y(_0185_),
    .A(\daisychain[36] ));
 sg13g2_inv_1 _1504_ (.Y(_0184_),
    .A(\daisychain[35] ));
 sg13g2_inv_1 _1505_ (.Y(_0183_),
    .A(\daisychain[34] ));
 sg13g2_inv_1 _1506_ (.Y(_0182_),
    .A(\daisychain[33] ));
 sg13g2_inv_1 _1507_ (.Y(_0181_),
    .A(\daisychain[32] ));
 sg13g2_inv_1 _1508_ (.Y(_0180_),
    .A(\daisychain[31] ));
 sg13g2_inv_1 _1509_ (.Y(_0179_),
    .A(\daisychain[30] ));
 sg13g2_inv_1 _1510_ (.Y(_0177_),
    .A(\daisychain[29] ));
 sg13g2_inv_1 _1511_ (.Y(_0176_),
    .A(\daisychain[28] ));
 sg13g2_inv_1 _1512_ (.Y(_0175_),
    .A(\daisychain[27] ));
 sg13g2_inv_1 _1513_ (.Y(_0174_),
    .A(\daisychain[26] ));
 sg13g2_inv_1 _1514_ (.Y(_0173_),
    .A(\daisychain[25] ));
 sg13g2_inv_1 _1515_ (.Y(_0172_),
    .A(\daisychain[24] ));
 sg13g2_inv_1 _1516_ (.Y(_0171_),
    .A(\daisychain[23] ));
 sg13g2_inv_1 _1517_ (.Y(_0170_),
    .A(\daisychain[22] ));
 sg13g2_inv_1 _1518_ (.Y(_0169_),
    .A(\daisychain[21] ));
 sg13g2_inv_1 _1519_ (.Y(_0168_),
    .A(\daisychain[20] ));
 sg13g2_inv_1 _1520_ (.Y(_0166_),
    .A(\daisychain[19] ));
 sg13g2_inv_1 _1521_ (.Y(_0165_),
    .A(\daisychain[18] ));
 sg13g2_inv_1 _1522_ (.Y(_0164_),
    .A(\daisychain[17] ));
 sg13g2_inv_1 _1523_ (.Y(_0163_),
    .A(\daisychain[16] ));
 sg13g2_inv_1 _1524_ (.Y(_0162_),
    .A(\daisychain[15] ));
 sg13g2_inv_1 _1525_ (.Y(_0161_),
    .A(\daisychain[14] ));
 sg13g2_inv_1 _1526_ (.Y(_0160_),
    .A(\daisychain[13] ));
 sg13g2_inv_1 _1527_ (.Y(_0159_),
    .A(\daisychain[12] ));
 sg13g2_inv_1 _1528_ (.Y(_0150_),
    .A(\daisychain[11] ));
 sg13g2_inv_1 _1529_ (.Y(_0139_),
    .A(\daisychain[10] ));
 sg13g2_inv_1 _1530_ (.Y(_0255_),
    .A(\daisychain[9] ));
 sg13g2_inv_1 _1531_ (.Y(_0244_),
    .A(\daisychain[8] ));
 sg13g2_inv_1 _1532_ (.Y(_0233_),
    .A(\daisychain[7] ));
 sg13g2_inv_1 _1533_ (.Y(_0222_),
    .A(\daisychain[6] ));
 sg13g2_inv_1 _1534_ (.Y(_0211_),
    .A(\daisychain[5] ));
 sg13g2_inv_1 _1535_ (.Y(_0200_),
    .A(\daisychain[4] ));
 sg13g2_inv_1 _1536_ (.Y(_0189_),
    .A(\daisychain[3] ));
 sg13g2_inv_1 _1537_ (.Y(_0178_),
    .A(\daisychain[2] ));
 sg13g2_inv_1 _1538_ (.Y(_0167_),
    .A(\daisychain[1] ));
 sg13g2_inv_1 _1539_ (.Y(_0128_),
    .A(\daisychain[0] ));
 sg13g2_inv_1 _1540_ (.Y(_0512_),
    .A(net1));
 sg13g2_o21ai_1 _1541_ (.B1(net211),
    .Y(_0513_),
    .A1(\state[0] ),
    .A2(net170));
 sg13g2_a21o_1 _1542_ (.A2(net170),
    .A1(_0128_),
    .B1(_0513_),
    .X(_0514_));
 sg13g2_nor2_1 _1543_ (.A(net211),
    .B(net3),
    .Y(_0515_));
 sg13g2_a21oi_1 _1544_ (.A1(net123),
    .A2(net2),
    .Y(_0516_),
    .B1(net35));
 sg13g2_a221oi_1 _1545_ (.B2(_0514_),
    .C1(net79),
    .B1(_0516_),
    .A1(_0128_),
    .Y(_0256_),
    .A2(net35));
 sg13g2_o21ai_1 _1546_ (.B1(net211),
    .Y(_0517_),
    .A1(\state[1] ),
    .A2(net170));
 sg13g2_a21o_1 _1547_ (.A2(net170),
    .A1(_0167_),
    .B1(_0517_),
    .X(_0518_));
 sg13g2_a21oi_1 _1548_ (.A1(net124),
    .A2(\daisychain[0] ),
    .Y(_0519_),
    .B1(net34));
 sg13g2_a221oi_1 _1549_ (.B2(_0519_),
    .C1(net80),
    .B1(_0518_),
    .A1(_0167_),
    .Y(_0257_),
    .A2(net34));
 sg13g2_o21ai_1 _1550_ (.B1(net205),
    .Y(_0520_),
    .A1(\state[2] ),
    .A2(net160));
 sg13g2_a21o_1 _1551_ (.A2(net160),
    .A1(_0178_),
    .B1(_0520_),
    .X(_0521_));
 sg13g2_a21oi_1 _1552_ (.A1(net124),
    .A2(\daisychain[1] ),
    .Y(_0522_),
    .B1(net34));
 sg13g2_a221oi_1 _1553_ (.B2(_0522_),
    .C1(net80),
    .B1(_0521_),
    .A1(_0178_),
    .Y(_0258_),
    .A2(net34));
 sg13g2_o21ai_1 _1554_ (.B1(net205),
    .Y(_0523_),
    .A1(\state[3] ),
    .A2(net161));
 sg13g2_a21o_1 _1555_ (.A2(net161),
    .A1(_0189_),
    .B1(_0523_),
    .X(_0524_));
 sg13g2_a21oi_1 _1556_ (.A1(net124),
    .A2(\daisychain[2] ),
    .Y(_0525_),
    .B1(net34));
 sg13g2_a221oi_1 _1557_ (.B2(_0525_),
    .C1(net80),
    .B1(_0524_),
    .A1(_0189_),
    .Y(_0259_),
    .A2(net34));
 sg13g2_o21ai_1 _1558_ (.B1(net207),
    .Y(_0526_),
    .A1(\state[4] ),
    .A2(net165));
 sg13g2_a21o_1 _1559_ (.A2(net175),
    .A1(_0200_),
    .B1(_0526_),
    .X(_0527_));
 sg13g2_a21oi_1 _1560_ (.A1(net128),
    .A2(\daisychain[3] ),
    .Y(_0528_),
    .B1(net41));
 sg13g2_a221oi_1 _1561_ (.B2(_0528_),
    .C1(net84),
    .B1(_0527_),
    .A1(_0200_),
    .Y(_0260_),
    .A2(net41));
 sg13g2_o21ai_1 _1562_ (.B1(net207),
    .Y(_0529_),
    .A1(\state[5] ),
    .A2(net165));
 sg13g2_a21o_1 _1563_ (.A2(net166),
    .A1(_0211_),
    .B1(_0529_),
    .X(_0530_));
 sg13g2_a21oi_1 _1564_ (.A1(net128),
    .A2(\daisychain[4] ),
    .Y(_0531_),
    .B1(net41));
 sg13g2_a221oi_1 _1565_ (.B2(_0531_),
    .C1(net75),
    .B1(_0530_),
    .A1(_0211_),
    .Y(_0261_),
    .A2(net29));
 sg13g2_o21ai_1 _1566_ (.B1(net207),
    .Y(_0532_),
    .A1(\state[6] ),
    .A2(net166));
 sg13g2_a21o_1 _1567_ (.A2(net166),
    .A1(_0222_),
    .B1(_0532_),
    .X(_0533_));
 sg13g2_a21oi_1 _1568_ (.A1(net114),
    .A2(\daisychain[5] ),
    .Y(_0534_),
    .B1(net25));
 sg13g2_a221oi_1 _1569_ (.B2(_0534_),
    .C1(net70),
    .B1(_0533_),
    .A1(_0222_),
    .Y(_0262_),
    .A2(net25));
 sg13g2_o21ai_1 _1570_ (.B1(net205),
    .Y(_0535_),
    .A1(\state[7] ),
    .A2(net160));
 sg13g2_a21o_1 _1571_ (.A2(net160),
    .A1(_0233_),
    .B1(_0535_),
    .X(_0536_));
 sg13g2_a21oi_1 _1572_ (.A1(net114),
    .A2(\daisychain[6] ),
    .Y(_0537_),
    .B1(net25));
 sg13g2_a221oi_1 _1573_ (.B2(_0537_),
    .C1(net70),
    .B1(_0536_),
    .A1(_0233_),
    .Y(_0263_),
    .A2(net26));
 sg13g2_o21ai_1 _1574_ (.B1(net206),
    .Y(_0538_),
    .A1(\state[8] ),
    .A2(net169));
 sg13g2_a21o_1 _1575_ (.A2(net169),
    .A1(_0244_),
    .B1(_0538_),
    .X(_0539_));
 sg13g2_a21oi_1 _1576_ (.A1(net114),
    .A2(\daisychain[7] ),
    .Y(_0540_),
    .B1(net25));
 sg13g2_a221oi_1 _1577_ (.B2(_0540_),
    .C1(net70),
    .B1(_0539_),
    .A1(_0244_),
    .Y(_0264_),
    .A2(net33));
 sg13g2_o21ai_1 _1578_ (.B1(net206),
    .Y(_0541_),
    .A1(\state[9] ),
    .A2(net164));
 sg13g2_a21o_1 _1579_ (.A2(net164),
    .A1(_0255_),
    .B1(_0541_),
    .X(_0542_));
 sg13g2_a21oi_1 _1580_ (.A1(net117),
    .A2(\daisychain[8] ),
    .Y(_0543_),
    .B1(net28));
 sg13g2_a221oi_1 _1581_ (.B2(_0543_),
    .C1(net74),
    .B1(_0542_),
    .A1(_0255_),
    .Y(_0265_),
    .A2(net28));
 sg13g2_o21ai_1 _1582_ (.B1(net206),
    .Y(_0544_),
    .A1(\state[10] ),
    .A2(net164));
 sg13g2_a21o_1 _1583_ (.A2(net164),
    .A1(_0139_),
    .B1(_0544_),
    .X(_0545_));
 sg13g2_a21oi_1 _1584_ (.A1(net117),
    .A2(\daisychain[9] ),
    .Y(_0546_),
    .B1(net28));
 sg13g2_a221oi_1 _1585_ (.B2(_0546_),
    .C1(net74),
    .B1(_0545_),
    .A1(_0139_),
    .Y(_0266_),
    .A2(net28));
 sg13g2_o21ai_1 _1586_ (.B1(net206),
    .Y(_0547_),
    .A1(\state[11] ),
    .A2(net162));
 sg13g2_a21o_1 _1587_ (.A2(net162),
    .A1(_0150_),
    .B1(_0547_),
    .X(_0548_));
 sg13g2_a21oi_1 _1588_ (.A1(net116),
    .A2(\daisychain[10] ),
    .Y(_0549_),
    .B1(net27));
 sg13g2_a221oi_1 _1589_ (.B2(_0549_),
    .C1(net73),
    .B1(_0548_),
    .A1(_0150_),
    .Y(_0267_),
    .A2(net27));
 sg13g2_o21ai_1 _1590_ (.B1(net206),
    .Y(_0550_),
    .A1(\state[12] ),
    .A2(net162));
 sg13g2_a21o_1 _1591_ (.A2(net162),
    .A1(_0159_),
    .B1(_0550_),
    .X(_0551_));
 sg13g2_a21oi_1 _1592_ (.A1(net116),
    .A2(\daisychain[11] ),
    .Y(_0552_),
    .B1(net27));
 sg13g2_a221oi_1 _1593_ (.B2(_0552_),
    .C1(net73),
    .B1(_0551_),
    .A1(_0159_),
    .Y(_0268_),
    .A2(net27));
 sg13g2_o21ai_1 _1594_ (.B1(net218),
    .Y(_0553_),
    .A1(\state[13] ),
    .A2(net184));
 sg13g2_a21o_1 _1595_ (.A2(net184),
    .A1(_0160_),
    .B1(_0553_),
    .X(_0554_));
 sg13g2_a21oi_1 _1596_ (.A1(net138),
    .A2(\daisychain[12] ),
    .Y(_0555_),
    .B1(net52));
 sg13g2_a221oi_1 _1597_ (.B2(_0555_),
    .C1(net92),
    .B1(_0554_),
    .A1(_0160_),
    .Y(_0269_),
    .A2(net52));
 sg13g2_o21ai_1 _1598_ (.B1(net206),
    .Y(_0556_),
    .A1(\state[14] ),
    .A2(net162));
 sg13g2_a21o_1 _1599_ (.A2(net162),
    .A1(_0161_),
    .B1(_0556_),
    .X(_0557_));
 sg13g2_a21oi_1 _1600_ (.A1(net116),
    .A2(\daisychain[13] ),
    .Y(_0558_),
    .B1(net27));
 sg13g2_a221oi_1 _1601_ (.B2(_0558_),
    .C1(net73),
    .B1(_0557_),
    .A1(_0161_),
    .Y(_0270_),
    .A2(net27));
 sg13g2_o21ai_1 _1602_ (.B1(net207),
    .Y(_0559_),
    .A1(\state[15] ),
    .A2(net167));
 sg13g2_a21o_1 _1603_ (.A2(net167),
    .A1(_0162_),
    .B1(_0559_),
    .X(_0560_));
 sg13g2_a21oi_1 _1604_ (.A1(net119),
    .A2(\daisychain[14] ),
    .Y(_0561_),
    .B1(net30));
 sg13g2_a221oi_1 _1605_ (.B2(_0561_),
    .C1(net76),
    .B1(_0560_),
    .A1(_0162_),
    .Y(_0271_),
    .A2(net30));
 sg13g2_o21ai_1 _1606_ (.B1(net213),
    .Y(_0562_),
    .A1(\state[16] ),
    .A2(net177));
 sg13g2_a21o_1 _1607_ (.A2(net177),
    .A1(_0163_),
    .B1(_0562_),
    .X(_0563_));
 sg13g2_a21oi_1 _1608_ (.A1(net129),
    .A2(\daisychain[15] ),
    .Y(_0564_),
    .B1(net42));
 sg13g2_a221oi_1 _1609_ (.B2(_0564_),
    .C1(net85),
    .B1(_0563_),
    .A1(_0163_),
    .Y(_0272_),
    .A2(net42));
 sg13g2_o21ai_1 _1610_ (.B1(net220),
    .Y(_0565_),
    .A1(\state[17] ),
    .A2(net187));
 sg13g2_a21o_1 _1611_ (.A2(net187),
    .A1(_0164_),
    .B1(_0565_),
    .X(_0566_));
 sg13g2_a21oi_1 _1612_ (.A1(net148),
    .A2(\daisychain[16] ),
    .Y(_0567_),
    .B1(net57));
 sg13g2_a221oi_1 _1613_ (.B2(_0567_),
    .C1(net102),
    .B1(_0566_),
    .A1(_0164_),
    .Y(_0273_),
    .A2(net57));
 sg13g2_o21ai_1 _1614_ (.B1(net213),
    .Y(_0568_),
    .A1(\state[18] ),
    .A2(net177));
 sg13g2_a21o_1 _1615_ (.A2(net177),
    .A1(_0165_),
    .B1(_0568_),
    .X(_0569_));
 sg13g2_a21oi_1 _1616_ (.A1(net129),
    .A2(\daisychain[17] ),
    .Y(_0570_),
    .B1(net42));
 sg13g2_a221oi_1 _1617_ (.B2(_0570_),
    .C1(net85),
    .B1(_0569_),
    .A1(_0165_),
    .Y(_0274_),
    .A2(net42));
 sg13g2_o21ai_1 _1618_ (.B1(net213),
    .Y(_0571_),
    .A1(\state[19] ),
    .A2(net175));
 sg13g2_a21o_1 _1619_ (.A2(net175),
    .A1(_0166_),
    .B1(_0571_),
    .X(_0572_));
 sg13g2_a21oi_1 _1620_ (.A1(net129),
    .A2(\daisychain[18] ),
    .Y(_0573_),
    .B1(net42));
 sg13g2_a221oi_1 _1621_ (.B2(_0573_),
    .C1(net84),
    .B1(_0572_),
    .A1(_0166_),
    .Y(_0275_),
    .A2(net41));
 sg13g2_o21ai_1 _1622_ (.B1(net207),
    .Y(_0574_),
    .A1(\state[20] ),
    .A2(net165));
 sg13g2_a21o_1 _1623_ (.A2(net165),
    .A1(_0168_),
    .B1(_0574_),
    .X(_0575_));
 sg13g2_a21oi_1 _1624_ (.A1(net118),
    .A2(\daisychain[19] ),
    .Y(_0576_),
    .B1(net29));
 sg13g2_a221oi_1 _1625_ (.B2(_0576_),
    .C1(net75),
    .B1(_0575_),
    .A1(_0168_),
    .Y(_0276_),
    .A2(net29));
 sg13g2_o21ai_1 _1626_ (.B1(net207),
    .Y(_0577_),
    .A1(\state[21] ),
    .A2(net165));
 sg13g2_a21o_1 _1627_ (.A2(net165),
    .A1(_0169_),
    .B1(_0577_),
    .X(_0578_));
 sg13g2_a21oi_1 _1628_ (.A1(net118),
    .A2(\daisychain[20] ),
    .Y(_0579_),
    .B1(net29));
 sg13g2_a221oi_1 _1629_ (.B2(_0579_),
    .C1(net75),
    .B1(_0578_),
    .A1(_0169_),
    .Y(_0277_),
    .A2(net29));
 sg13g2_o21ai_1 _1630_ (.B1(net223),
    .Y(_0580_),
    .A1(\state[22] ),
    .A2(net194));
 sg13g2_a21o_1 _1631_ (.A2(net194),
    .A1(_0170_),
    .B1(_0580_),
    .X(_0581_));
 sg13g2_a21oi_1 _1632_ (.A1(net148),
    .A2(\daisychain[21] ),
    .Y(_0582_),
    .B1(net57));
 sg13g2_a221oi_1 _1633_ (.B2(_0582_),
    .C1(net102),
    .B1(_0581_),
    .A1(_0170_),
    .Y(_0278_),
    .A2(net57));
 sg13g2_o21ai_1 _1634_ (.B1(net223),
    .Y(_0583_),
    .A1(\state[23] ),
    .A2(net194));
 sg13g2_a21o_1 _1635_ (.A2(net194),
    .A1(_0171_),
    .B1(_0583_),
    .X(_0584_));
 sg13g2_a21oi_1 _1636_ (.A1(net148),
    .A2(\daisychain[22] ),
    .Y(_0585_),
    .B1(net57));
 sg13g2_a221oi_1 _1637_ (.B2(_0585_),
    .C1(net102),
    .B1(_0584_),
    .A1(_0171_),
    .Y(_0279_),
    .A2(net57));
 sg13g2_o21ai_1 _1638_ (.B1(net223),
    .Y(_0586_),
    .A1(\state[24] ),
    .A2(net195));
 sg13g2_a21o_1 _1639_ (.A2(net195),
    .A1(_0172_),
    .B1(_0586_),
    .X(_0587_));
 sg13g2_a21oi_1 _1640_ (.A1(net149),
    .A2(\daisychain[23] ),
    .Y(_0588_),
    .B1(net58));
 sg13g2_a221oi_1 _1641_ (.B2(_0588_),
    .C1(net103),
    .B1(_0587_),
    .A1(_0172_),
    .Y(_0280_),
    .A2(net58));
 sg13g2_o21ai_1 _1642_ (.B1(net223),
    .Y(_0589_),
    .A1(\state[25] ),
    .A2(net194));
 sg13g2_a21o_1 _1643_ (.A2(net194),
    .A1(_0173_),
    .B1(_0589_),
    .X(_0590_));
 sg13g2_a21oi_1 _1644_ (.A1(net148),
    .A2(\daisychain[24] ),
    .Y(_0591_),
    .B1(net57));
 sg13g2_a221oi_1 _1645_ (.B2(_0591_),
    .C1(net102),
    .B1(_0590_),
    .A1(_0173_),
    .Y(_0281_),
    .A2(net57));
 sg13g2_o21ai_1 _1646_ (.B1(net208),
    .Y(_0592_),
    .A1(\state[26] ),
    .A2(net167));
 sg13g2_a21o_1 _1647_ (.A2(net167),
    .A1(_0174_),
    .B1(_0592_),
    .X(_0593_));
 sg13g2_a21oi_1 _1648_ (.A1(net119),
    .A2(\daisychain[25] ),
    .Y(_0594_),
    .B1(net30));
 sg13g2_a221oi_1 _1649_ (.B2(_0594_),
    .C1(net76),
    .B1(_0593_),
    .A1(_0174_),
    .Y(_0282_),
    .A2(net30));
 sg13g2_o21ai_1 _1650_ (.B1(net208),
    .Y(_0595_),
    .A1(\state[27] ),
    .A2(net167));
 sg13g2_a21o_1 _1651_ (.A2(net167),
    .A1(_0175_),
    .B1(_0595_),
    .X(_0596_));
 sg13g2_a21oi_1 _1652_ (.A1(net119),
    .A2(\daisychain[26] ),
    .Y(_0597_),
    .B1(net30));
 sg13g2_a221oi_1 _1653_ (.B2(_0597_),
    .C1(net76),
    .B1(_0596_),
    .A1(_0175_),
    .Y(_0283_),
    .A2(net30));
 sg13g2_o21ai_1 _1654_ (.B1(net207),
    .Y(_0598_),
    .A1(\state[28] ),
    .A2(net165));
 sg13g2_a21o_1 _1655_ (.A2(net165),
    .A1(_0176_),
    .B1(_0598_),
    .X(_0599_));
 sg13g2_a21oi_1 _1656_ (.A1(net118),
    .A2(\daisychain[27] ),
    .Y(_0600_),
    .B1(net29));
 sg13g2_a221oi_1 _1657_ (.B2(_0600_),
    .C1(net75),
    .B1(_0599_),
    .A1(_0176_),
    .Y(_0284_),
    .A2(net29));
 sg13g2_o21ai_1 _1658_ (.B1(net207),
    .Y(_0601_),
    .A1(\state[29] ),
    .A2(net166));
 sg13g2_a21o_1 _1659_ (.A2(net166),
    .A1(_0177_),
    .B1(_0601_),
    .X(_0602_));
 sg13g2_a21oi_1 _1660_ (.A1(net118),
    .A2(\daisychain[28] ),
    .Y(_0603_),
    .B1(net29));
 sg13g2_a221oi_1 _1661_ (.B2(_0603_),
    .C1(net75),
    .B1(_0602_),
    .A1(_0177_),
    .Y(_0285_),
    .A2(net32));
 sg13g2_o21ai_1 _1662_ (.B1(net208),
    .Y(_0604_),
    .A1(\state[30] ),
    .A2(net168));
 sg13g2_a21o_1 _1663_ (.A2(net168),
    .A1(_0179_),
    .B1(_0604_),
    .X(_0605_));
 sg13g2_a21oi_1 _1664_ (.A1(net119),
    .A2(\daisychain[29] ),
    .Y(_0606_),
    .B1(net31));
 sg13g2_a221oi_1 _1665_ (.B2(_0606_),
    .C1(net76),
    .B1(_0605_),
    .A1(_0179_),
    .Y(_0286_),
    .A2(net31));
 sg13g2_o21ai_1 _1666_ (.B1(net206),
    .Y(_0607_),
    .A1(\state[31] ),
    .A2(net162));
 sg13g2_a21o_1 _1667_ (.A2(net163),
    .A1(_0180_),
    .B1(_0607_),
    .X(_0608_));
 sg13g2_a21oi_1 _1668_ (.A1(net120),
    .A2(\daisychain[30] ),
    .Y(_0609_),
    .B1(net31));
 sg13g2_a221oi_1 _1669_ (.B2(_0609_),
    .C1(net77),
    .B1(_0608_),
    .A1(_0180_),
    .Y(_0287_),
    .A2(net31));
 sg13g2_o21ai_1 _1670_ (.B1(net208),
    .Y(_0610_),
    .A1(\state[32] ),
    .A2(net167));
 sg13g2_a21o_1 _1671_ (.A2(net167),
    .A1(_0181_),
    .B1(_0610_),
    .X(_0611_));
 sg13g2_a21oi_1 _1672_ (.A1(net119),
    .A2(\daisychain[31] ),
    .Y(_0612_),
    .B1(net30));
 sg13g2_a221oi_1 _1673_ (.B2(_0612_),
    .C1(net76),
    .B1(_0611_),
    .A1(_0181_),
    .Y(_0288_),
    .A2(net30));
 sg13g2_o21ai_1 _1674_ (.B1(net209),
    .Y(_0613_),
    .A1(\state[33] ),
    .A2(net163));
 sg13g2_a21o_1 _1675_ (.A2(net163),
    .A1(_0182_),
    .B1(_0613_),
    .X(_0614_));
 sg13g2_a21oi_1 _1676_ (.A1(net116),
    .A2(\daisychain[32] ),
    .Y(_0615_),
    .B1(net27));
 sg13g2_a221oi_1 _1677_ (.B2(_0615_),
    .C1(net73),
    .B1(_0614_),
    .A1(_0182_),
    .Y(_0289_),
    .A2(net27));
 sg13g2_o21ai_1 _1678_ (.B1(net206),
    .Y(_0616_),
    .A1(\state[34] ),
    .A2(net164));
 sg13g2_a21o_1 _1679_ (.A2(net164),
    .A1(_0183_),
    .B1(_0616_),
    .X(_0617_));
 sg13g2_a21oi_1 _1680_ (.A1(net117),
    .A2(\daisychain[33] ),
    .Y(_0618_),
    .B1(net28));
 sg13g2_a221oi_1 _1681_ (.B2(_0618_),
    .C1(net74),
    .B1(_0617_),
    .A1(_0183_),
    .Y(_0290_),
    .A2(net28));
 sg13g2_o21ai_1 _1682_ (.B1(net218),
    .Y(_0619_),
    .A1(\state[35] ),
    .A2(net162));
 sg13g2_a21o_1 _1683_ (.A2(net184),
    .A1(_0184_),
    .B1(_0619_),
    .X(_0620_));
 sg13g2_a21oi_1 _1684_ (.A1(net116),
    .A2(\daisychain[34] ),
    .Y(_0621_),
    .B1(net28));
 sg13g2_a221oi_1 _1685_ (.B2(_0621_),
    .C1(net92),
    .B1(_0620_),
    .A1(_0184_),
    .Y(_0291_),
    .A2(net52));
 sg13g2_o21ai_1 _1686_ (.B1(net209),
    .Y(_0622_),
    .A1(\state[36] ),
    .A2(net163));
 sg13g2_a21o_1 _1687_ (.A2(net186),
    .A1(_0185_),
    .B1(_0622_),
    .X(_0623_));
 sg13g2_a21oi_1 _1688_ (.A1(net140),
    .A2(\daisychain[35] ),
    .Y(_0624_),
    .B1(net49));
 sg13g2_a221oi_1 _1689_ (.B2(_0624_),
    .C1(net94),
    .B1(_0623_),
    .A1(_0185_),
    .Y(_0292_),
    .A2(net49));
 sg13g2_o21ai_1 _1690_ (.B1(net218),
    .Y(_0625_),
    .A1(\state[37] ),
    .A2(net184));
 sg13g2_a21o_1 _1691_ (.A2(net184),
    .A1(_0186_),
    .B1(_0625_),
    .X(_0626_));
 sg13g2_a21oi_1 _1692_ (.A1(net140),
    .A2(\daisychain[36] ),
    .Y(_0627_),
    .B1(net49));
 sg13g2_a221oi_1 _1693_ (.B2(_0627_),
    .C1(net94),
    .B1(_0626_),
    .A1(_0186_),
    .Y(_0293_),
    .A2(net49));
 sg13g2_o21ai_1 _1694_ (.B1(net218),
    .Y(_0628_),
    .A1(\state[38] ),
    .A2(net184));
 sg13g2_a21o_1 _1695_ (.A2(net187),
    .A1(_0187_),
    .B1(_0628_),
    .X(_0629_));
 sg13g2_a21oi_1 _1696_ (.A1(net140),
    .A2(\daisychain[37] ),
    .Y(_0630_),
    .B1(net49));
 sg13g2_a221oi_1 _1697_ (.B2(_0630_),
    .C1(net94),
    .B1(_0629_),
    .A1(_0187_),
    .Y(_0294_),
    .A2(net49));
 sg13g2_o21ai_1 _1698_ (.B1(net223),
    .Y(_0631_),
    .A1(\state[39] ),
    .A2(net195));
 sg13g2_a21o_1 _1699_ (.A2(net195),
    .A1(_0188_),
    .B1(_0631_),
    .X(_0632_));
 sg13g2_a21oi_1 _1700_ (.A1(net149),
    .A2(\daisychain[38] ),
    .Y(_0633_),
    .B1(net58));
 sg13g2_a221oi_1 _1701_ (.B2(_0633_),
    .C1(net103),
    .B1(_0632_),
    .A1(_0188_),
    .Y(_0295_),
    .A2(net58));
 sg13g2_o21ai_1 _1702_ (.B1(net220),
    .Y(_0634_),
    .A1(\state[40] ),
    .A2(net187));
 sg13g2_a21o_1 _1703_ (.A2(net195),
    .A1(_0190_),
    .B1(_0634_),
    .X(_0635_));
 sg13g2_a21oi_1 _1704_ (.A1(net149),
    .A2(\daisychain[39] ),
    .Y(_0636_),
    .B1(net58));
 sg13g2_a221oi_1 _1705_ (.B2(_0636_),
    .C1(net103),
    .B1(_0635_),
    .A1(_0190_),
    .Y(_0296_),
    .A2(net58));
 sg13g2_o21ai_1 _1706_ (.B1(net218),
    .Y(_0637_),
    .A1(\state[41] ),
    .A2(net186));
 sg13g2_a21o_1 _1707_ (.A2(net187),
    .A1(_0191_),
    .B1(_0637_),
    .X(_0638_));
 sg13g2_a21oi_1 _1708_ (.A1(net140),
    .A2(\daisychain[40] ),
    .Y(_0639_),
    .B1(net49));
 sg13g2_a221oi_1 _1709_ (.B2(_0639_),
    .C1(net94),
    .B1(_0638_),
    .A1(_0191_),
    .Y(_0297_),
    .A2(net49));
 sg13g2_o21ai_1 _1710_ (.B1(net218),
    .Y(_0640_),
    .A1(\state[42] ),
    .A2(net184));
 sg13g2_a21o_1 _1711_ (.A2(net184),
    .A1(_0192_),
    .B1(_0640_),
    .X(_0641_));
 sg13g2_a21oi_1 _1712_ (.A1(net140),
    .A2(\daisychain[41] ),
    .Y(_0642_),
    .B1(net51));
 sg13g2_a221oi_1 _1713_ (.B2(_0642_),
    .C1(net94),
    .B1(_0641_),
    .A1(_0192_),
    .Y(_0298_),
    .A2(net51));
 sg13g2_o21ai_1 _1714_ (.B1(net218),
    .Y(_0643_),
    .A1(\state[43] ),
    .A2(net185));
 sg13g2_a21o_1 _1715_ (.A2(net185),
    .A1(_0193_),
    .B1(_0643_),
    .X(_0644_));
 sg13g2_a21oi_1 _1716_ (.A1(net140),
    .A2(\daisychain[42] ),
    .Y(_0645_),
    .B1(net50));
 sg13g2_a221oi_1 _1717_ (.B2(_0645_),
    .C1(net94),
    .B1(_0644_),
    .A1(_0193_),
    .Y(_0299_),
    .A2(net50));
 sg13g2_o21ai_1 _1718_ (.B1(net218),
    .Y(_0646_),
    .A1(\state[44] ),
    .A2(net185));
 sg13g2_a21o_1 _1719_ (.A2(net185),
    .A1(_0194_),
    .B1(_0646_),
    .X(_0647_));
 sg13g2_a21oi_1 _1720_ (.A1(net141),
    .A2(\daisychain[43] ),
    .Y(_0648_),
    .B1(net50));
 sg13g2_a221oi_1 _1721_ (.B2(_0648_),
    .C1(net94),
    .B1(_0647_),
    .A1(_0194_),
    .Y(_0300_),
    .A2(net50));
 sg13g2_o21ai_1 _1722_ (.B1(net219),
    .Y(_0649_),
    .A1(\state[45] ),
    .A2(net185));
 sg13g2_a21o_1 _1723_ (.A2(net185),
    .A1(_0195_),
    .B1(_0649_),
    .X(_0650_));
 sg13g2_a21oi_1 _1724_ (.A1(net141),
    .A2(\daisychain[44] ),
    .Y(_0651_),
    .B1(net50));
 sg13g2_a221oi_1 _1725_ (.B2(_0651_),
    .C1(net95),
    .B1(_0650_),
    .A1(_0195_),
    .Y(_0301_),
    .A2(net50));
 sg13g2_o21ai_1 _1726_ (.B1(net219),
    .Y(_0652_),
    .A1(\state[46] ),
    .A2(net185));
 sg13g2_a21o_1 _1727_ (.A2(net187),
    .A1(_0196_),
    .B1(_0652_),
    .X(_0653_));
 sg13g2_a21oi_1 _1728_ (.A1(net141),
    .A2(\daisychain[45] ),
    .Y(_0654_),
    .B1(net50));
 sg13g2_a221oi_1 _1729_ (.B2(_0654_),
    .C1(net95),
    .B1(_0653_),
    .A1(_0196_),
    .Y(_0302_),
    .A2(net50));
 sg13g2_o21ai_1 _1730_ (.B1(net219),
    .Y(_0655_),
    .A1(\state[47] ),
    .A2(net185));
 sg13g2_a21o_1 _1731_ (.A2(net187),
    .A1(_0197_),
    .B1(_0655_),
    .X(_0656_));
 sg13g2_a21oi_1 _1732_ (.A1(net154),
    .A2(\daisychain[46] ),
    .Y(_0657_),
    .B1(net62));
 sg13g2_a221oi_1 _1733_ (.B2(_0657_),
    .C1(net106),
    .B1(_0656_),
    .A1(_0197_),
    .Y(_0303_),
    .A2(net62));
 sg13g2_o21ai_1 _1734_ (.B1(net222),
    .Y(_0658_),
    .A1(\state[48] ),
    .A2(net192));
 sg13g2_a21o_1 _1735_ (.A2(net192),
    .A1(_0198_),
    .B1(_0658_),
    .X(_0659_));
 sg13g2_a21oi_1 _1736_ (.A1(net154),
    .A2(\daisychain[47] ),
    .Y(_0660_),
    .B1(net62));
 sg13g2_a221oi_1 _1737_ (.B2(_0660_),
    .C1(net106),
    .B1(_0659_),
    .A1(_0198_),
    .Y(_0304_),
    .A2(net62));
 sg13g2_o21ai_1 _1738_ (.B1(net221),
    .Y(_0661_),
    .A1(\state[49] ),
    .A2(net188));
 sg13g2_a21o_1 _1739_ (.A2(net192),
    .A1(_0199_),
    .B1(_0661_),
    .X(_0662_));
 sg13g2_a21oi_1 _1740_ (.A1(net145),
    .A2(\daisychain[48] ),
    .Y(_0663_),
    .B1(net55));
 sg13g2_a221oi_1 _1741_ (.B2(_0663_),
    .C1(net99),
    .B1(_0662_),
    .A1(_0199_),
    .Y(_0305_),
    .A2(net55));
 sg13g2_o21ai_1 _1742_ (.B1(net219),
    .Y(_0664_),
    .A1(\state[50] ),
    .A2(net186));
 sg13g2_a21o_1 _1743_ (.A2(net186),
    .A1(_0201_),
    .B1(_0664_),
    .X(_0665_));
 sg13g2_a21oi_1 _1744_ (.A1(net141),
    .A2(\daisychain[49] ),
    .Y(_0666_),
    .B1(net51));
 sg13g2_a221oi_1 _1745_ (.B2(_0666_),
    .C1(net95),
    .B1(_0665_),
    .A1(_0201_),
    .Y(_0306_),
    .A2(net51));
 sg13g2_o21ai_1 _1746_ (.B1(net221),
    .Y(_0667_),
    .A1(\state[51] ),
    .A2(net188));
 sg13g2_a21o_1 _1747_ (.A2(net188),
    .A1(_0202_),
    .B1(_0667_),
    .X(_0668_));
 sg13g2_a21oi_1 _1748_ (.A1(net145),
    .A2(\daisychain[50] ),
    .Y(_0669_),
    .B1(net55));
 sg13g2_a221oi_1 _1749_ (.B2(_0669_),
    .C1(net99),
    .B1(_0668_),
    .A1(_0202_),
    .Y(_0307_),
    .A2(net55));
 sg13g2_o21ai_1 _1750_ (.B1(net221),
    .Y(_0670_),
    .A1(\state[52] ),
    .A2(net188));
 sg13g2_a21o_1 _1751_ (.A2(net188),
    .A1(_0203_),
    .B1(_0670_),
    .X(_0671_));
 sg13g2_a21oi_1 _1752_ (.A1(net145),
    .A2(\daisychain[51] ),
    .Y(_0672_),
    .B1(net55));
 sg13g2_a221oi_1 _1753_ (.B2(_0672_),
    .C1(net99),
    .B1(_0671_),
    .A1(_0203_),
    .Y(_0308_),
    .A2(net55));
 sg13g2_o21ai_1 _1754_ (.B1(net221),
    .Y(_0673_),
    .A1(\state[53] ),
    .A2(net189));
 sg13g2_a21o_1 _1755_ (.A2(net189),
    .A1(_0204_),
    .B1(_0673_),
    .X(_0674_));
 sg13g2_a21oi_1 _1756_ (.A1(net145),
    .A2(\daisychain[52] ),
    .Y(_0675_),
    .B1(net53));
 sg13g2_a221oi_1 _1757_ (.B2(_0675_),
    .C1(net99),
    .B1(_0674_),
    .A1(_0204_),
    .Y(_0309_),
    .A2(net53));
 sg13g2_o21ai_1 _1758_ (.B1(net222),
    .Y(_0676_),
    .A1(\state[54] ),
    .A2(net192));
 sg13g2_a21o_1 _1759_ (.A2(net192),
    .A1(_0205_),
    .B1(_0676_),
    .X(_0677_));
 sg13g2_a21oi_1 _1760_ (.A1(net153),
    .A2(\daisychain[53] ),
    .Y(_0678_),
    .B1(net63));
 sg13g2_a221oi_1 _1761_ (.B2(_0678_),
    .C1(net107),
    .B1(_0677_),
    .A1(_0205_),
    .Y(_0310_),
    .A2(net53));
 sg13g2_o21ai_1 _1762_ (.B1(net222),
    .Y(_0679_),
    .A1(\state[55] ),
    .A2(net192));
 sg13g2_a21o_1 _1763_ (.A2(net192),
    .A1(_0206_),
    .B1(_0679_),
    .X(_0680_));
 sg13g2_a21oi_1 _1764_ (.A1(net153),
    .A2(\daisychain[54] ),
    .Y(_0681_),
    .B1(net53));
 sg13g2_a221oi_1 _1765_ (.B2(_0681_),
    .C1(net99),
    .B1(_0680_),
    .A1(_0206_),
    .Y(_0311_),
    .A2(net53));
 sg13g2_o21ai_1 _1766_ (.B1(net221),
    .Y(_0682_),
    .A1(\state[56] ),
    .A2(net189));
 sg13g2_a21o_1 _1767_ (.A2(net189),
    .A1(_0207_),
    .B1(_0682_),
    .X(_0683_));
 sg13g2_a21oi_1 _1768_ (.A1(net145),
    .A2(\daisychain[55] ),
    .Y(_0684_),
    .B1(net53));
 sg13g2_a221oi_1 _1769_ (.B2(_0684_),
    .C1(net99),
    .B1(_0683_),
    .A1(_0207_),
    .Y(_0312_),
    .A2(net53));
 sg13g2_o21ai_1 _1770_ (.B1(net221),
    .Y(_0685_),
    .A1(\state[57] ),
    .A2(net188));
 sg13g2_a21o_1 _1771_ (.A2(net191),
    .A1(_0208_),
    .B1(_0685_),
    .X(_0686_));
 sg13g2_a21oi_1 _1772_ (.A1(net145),
    .A2(\daisychain[56] ),
    .Y(_0687_),
    .B1(net53));
 sg13g2_a221oi_1 _1773_ (.B2(_0687_),
    .C1(net97),
    .B1(_0686_),
    .A1(_0208_),
    .Y(_0313_),
    .A2(net56));
 sg13g2_o21ai_1 _1774_ (.B1(net221),
    .Y(_0688_),
    .A1(\state[58] ),
    .A2(net188));
 sg13g2_a21o_1 _1775_ (.A2(net188),
    .A1(_0209_),
    .B1(_0688_),
    .X(_0689_));
 sg13g2_a21oi_1 _1776_ (.A1(net144),
    .A2(\daisychain[57] ),
    .Y(_0690_),
    .B1(net56));
 sg13g2_a221oi_1 _1777_ (.B2(_0690_),
    .C1(net97),
    .B1(_0689_),
    .A1(_0209_),
    .Y(_0314_),
    .A2(net56));
 sg13g2_o21ai_1 _1778_ (.B1(net221),
    .Y(_0691_),
    .A1(\state[59] ),
    .A2(net189));
 sg13g2_a21o_1 _1779_ (.A2(net189),
    .A1(_0210_),
    .B1(_0691_),
    .X(_0692_));
 sg13g2_a21oi_1 _1780_ (.A1(net143),
    .A2(\daisychain[58] ),
    .Y(_0693_),
    .B1(net56));
 sg13g2_a221oi_1 _1781_ (.B2(_0693_),
    .C1(net97),
    .B1(_0692_),
    .A1(_0210_),
    .Y(_0315_),
    .A2(net56));
 sg13g2_o21ai_1 _1782_ (.B1(net222),
    .Y(_0694_),
    .A1(\state[60] ),
    .A2(net189));
 sg13g2_a21o_1 _1783_ (.A2(net189),
    .A1(_0212_),
    .B1(_0694_),
    .X(_0695_));
 sg13g2_a21oi_1 _1784_ (.A1(net143),
    .A2(\daisychain[59] ),
    .Y(_0696_),
    .B1(net56));
 sg13g2_a221oi_1 _1785_ (.B2(_0696_),
    .C1(net98),
    .B1(_0695_),
    .A1(_0212_),
    .Y(_0316_),
    .A2(net56));
 sg13g2_o21ai_1 _1786_ (.B1(net222),
    .Y(_0697_),
    .A1(\state[61] ),
    .A2(net190));
 sg13g2_a21o_1 _1787_ (.A2(net190),
    .A1(_0213_),
    .B1(_0697_),
    .X(_0698_));
 sg13g2_a21oi_1 _1788_ (.A1(net146),
    .A2(\daisychain[60] ),
    .Y(_0699_),
    .B1(net54));
 sg13g2_a221oi_1 _1789_ (.B2(_0699_),
    .C1(net100),
    .B1(_0698_),
    .A1(_0213_),
    .Y(_0317_),
    .A2(net54));
 sg13g2_o21ai_1 _1790_ (.B1(net222),
    .Y(_0700_),
    .A1(\state[62] ),
    .A2(net190));
 sg13g2_a21o_1 _1791_ (.A2(net190),
    .A1(_0214_),
    .B1(_0700_),
    .X(_0701_));
 sg13g2_a21oi_1 _1792_ (.A1(net146),
    .A2(\daisychain[61] ),
    .Y(_0702_),
    .B1(net54));
 sg13g2_a221oi_1 _1793_ (.B2(_0702_),
    .C1(net100),
    .B1(_0701_),
    .A1(_0214_),
    .Y(_0318_),
    .A2(net54));
 sg13g2_o21ai_1 _1794_ (.B1(net222),
    .Y(_0703_),
    .A1(\state[63] ),
    .A2(net192));
 sg13g2_a21o_1 _1795_ (.A2(net193),
    .A1(_0215_),
    .B1(_0703_),
    .X(_0704_));
 sg13g2_a21oi_1 _1796_ (.A1(net153),
    .A2(\daisychain[62] ),
    .Y(_0705_),
    .B1(net63));
 sg13g2_a221oi_1 _1797_ (.B2(_0705_),
    .C1(net107),
    .B1(_0704_),
    .A1(_0215_),
    .Y(_0319_),
    .A2(net63));
 sg13g2_o21ai_1 _1798_ (.B1(net225),
    .Y(_0706_),
    .A1(\state[64] ),
    .A2(net199));
 sg13g2_a21o_1 _1799_ (.A2(net199),
    .A1(_0216_),
    .B1(_0706_),
    .X(_0707_));
 sg13g2_a21oi_1 _1800_ (.A1(net153),
    .A2(\daisychain[63] ),
    .Y(_0708_),
    .B1(net63));
 sg13g2_a221oi_1 _1801_ (.B2(_0708_),
    .C1(net107),
    .B1(_0707_),
    .A1(_0216_),
    .Y(_0320_),
    .A2(net63));
 sg13g2_o21ai_1 _1802_ (.B1(net225),
    .Y(_0709_),
    .A1(\state[65] ),
    .A2(net200));
 sg13g2_a21o_1 _1803_ (.A2(net200),
    .A1(_0217_),
    .B1(_0709_),
    .X(_0710_));
 sg13g2_a21oi_1 _1804_ (.A1(net153),
    .A2(\daisychain[64] ),
    .Y(_0711_),
    .B1(net63));
 sg13g2_a221oi_1 _1805_ (.B2(_0711_),
    .C1(net107),
    .B1(_0710_),
    .A1(_0217_),
    .Y(_0321_),
    .A2(net63));
 sg13g2_o21ai_1 _1806_ (.B1(net225),
    .Y(_0712_),
    .A1(\state[66] ),
    .A2(net200));
 sg13g2_a21o_1 _1807_ (.A2(net200),
    .A1(_0218_),
    .B1(_0712_),
    .X(_0713_));
 sg13g2_a21oi_1 _1808_ (.A1(net157),
    .A2(\daisychain[65] ),
    .Y(_0714_),
    .B1(net64));
 sg13g2_a221oi_1 _1809_ (.B2(_0714_),
    .C1(net107),
    .B1(_0713_),
    .A1(_0218_),
    .Y(_0322_),
    .A2(net63));
 sg13g2_o21ai_1 _1810_ (.B1(net225),
    .Y(_0715_),
    .A1(\state[67] ),
    .A2(net201));
 sg13g2_a21o_1 _1811_ (.A2(net201),
    .A1(_0219_),
    .B1(_0715_),
    .X(_0716_));
 sg13g2_a21oi_1 _1812_ (.A1(net155),
    .A2(\daisychain[66] ),
    .Y(_0717_),
    .B1(net65));
 sg13g2_a221oi_1 _1813_ (.B2(_0717_),
    .C1(net108),
    .B1(_0716_),
    .A1(_0219_),
    .Y(_0323_),
    .A2(net65));
 sg13g2_o21ai_1 _1814_ (.B1(net225),
    .Y(_0718_),
    .A1(\state[68] ),
    .A2(net202));
 sg13g2_a21o_1 _1815_ (.A2(net202),
    .A1(_0220_),
    .B1(_0718_),
    .X(_0719_));
 sg13g2_a21oi_1 _1816_ (.A1(net155),
    .A2(\daisychain[67] ),
    .Y(_0720_),
    .B1(net66));
 sg13g2_a221oi_1 _1817_ (.B2(_0720_),
    .C1(net108),
    .B1(_0719_),
    .A1(_0220_),
    .Y(_0324_),
    .A2(net66));
 sg13g2_o21ai_1 _1818_ (.B1(net226),
    .Y(_0721_),
    .A1(\state[69] ),
    .A2(net202));
 sg13g2_a21o_1 _1819_ (.A2(net202),
    .A1(_0221_),
    .B1(_0721_),
    .X(_0722_));
 sg13g2_a21oi_1 _1820_ (.A1(net156),
    .A2(\daisychain[68] ),
    .Y(_0723_),
    .B1(net66));
 sg13g2_a221oi_1 _1821_ (.B2(_0723_),
    .C1(net109),
    .B1(_0722_),
    .A1(_0221_),
    .Y(_0325_),
    .A2(net66));
 sg13g2_o21ai_1 _1822_ (.B1(net226),
    .Y(_0724_),
    .A1(\state[70] ),
    .A2(net201));
 sg13g2_a21o_1 _1823_ (.A2(net201),
    .A1(_0223_),
    .B1(_0724_),
    .X(_0725_));
 sg13g2_a21oi_1 _1824_ (.A1(net155),
    .A2(\daisychain[69] ),
    .Y(_0726_),
    .B1(net65));
 sg13g2_a221oi_1 _1825_ (.B2(_0726_),
    .C1(net108),
    .B1(_0725_),
    .A1(_0223_),
    .Y(_0326_),
    .A2(net65));
 sg13g2_o21ai_1 _1826_ (.B1(net224),
    .Y(_0727_),
    .A1(\state[71] ),
    .A2(net197));
 sg13g2_a21o_1 _1827_ (.A2(net197),
    .A1(_0224_),
    .B1(_0727_),
    .X(_0728_));
 sg13g2_a21oi_1 _1828_ (.A1(net151),
    .A2(\daisychain[70] ),
    .Y(_0729_),
    .B1(net60));
 sg13g2_a221oi_1 _1829_ (.B2(_0729_),
    .C1(net105),
    .B1(_0728_),
    .A1(_0224_),
    .Y(_0327_),
    .A2(net60));
 sg13g2_o21ai_1 _1830_ (.B1(net226),
    .Y(_0730_),
    .A1(\state[72] ),
    .A2(net201));
 sg13g2_a21o_1 _1831_ (.A2(net201),
    .A1(_0225_),
    .B1(_0730_),
    .X(_0731_));
 sg13g2_a21oi_1 _1832_ (.A1(net155),
    .A2(\daisychain[71] ),
    .Y(_0732_),
    .B1(net65));
 sg13g2_a221oi_1 _1833_ (.B2(_0732_),
    .C1(net108),
    .B1(_0731_),
    .A1(_0225_),
    .Y(_0328_),
    .A2(net65));
 sg13g2_o21ai_1 _1834_ (.B1(net226),
    .Y(_0733_),
    .A1(\state[73] ),
    .A2(net202));
 sg13g2_a21o_1 _1835_ (.A2(net202),
    .A1(_0226_),
    .B1(_0733_),
    .X(_0734_));
 sg13g2_a21oi_1 _1836_ (.A1(net156),
    .A2(\daisychain[72] ),
    .Y(_0735_),
    .B1(net66));
 sg13g2_a221oi_1 _1837_ (.B2(_0735_),
    .C1(net109),
    .B1(_0734_),
    .A1(_0226_),
    .Y(_0329_),
    .A2(net66));
 sg13g2_o21ai_1 _1838_ (.B1(net225),
    .Y(_0736_),
    .A1(\state[74] ),
    .A2(net199));
 sg13g2_a21o_1 _1839_ (.A2(net199),
    .A1(_0227_),
    .B1(_0736_),
    .X(_0737_));
 sg13g2_a21oi_1 _1840_ (.A1(net154),
    .A2(\daisychain[73] ),
    .Y(_0738_),
    .B1(net62));
 sg13g2_a221oi_1 _1841_ (.B2(_0738_),
    .C1(net106),
    .B1(_0737_),
    .A1(_0227_),
    .Y(_0330_),
    .A2(net62));
 sg13g2_o21ai_1 _1842_ (.B1(net225),
    .Y(_0739_),
    .A1(\state[75] ),
    .A2(net199));
 sg13g2_a21o_1 _1843_ (.A2(net199),
    .A1(_0228_),
    .B1(_0739_),
    .X(_0740_));
 sg13g2_a21oi_1 _1844_ (.A1(net154),
    .A2(\daisychain[74] ),
    .Y(_0741_),
    .B1(net64));
 sg13g2_a221oi_1 _1845_ (.B2(_0741_),
    .C1(net106),
    .B1(_0740_),
    .A1(_0228_),
    .Y(_0331_),
    .A2(net62));
 sg13g2_o21ai_1 _1846_ (.B1(net225),
    .Y(_0742_),
    .A1(\state[76] ),
    .A2(net199));
 sg13g2_a21o_1 _1847_ (.A2(net199),
    .A1(_0229_),
    .B1(_0742_),
    .X(_0743_));
 sg13g2_a21oi_1 _1848_ (.A1(net154),
    .A2(\daisychain[75] ),
    .Y(_0744_),
    .B1(net64));
 sg13g2_a221oi_1 _1849_ (.B2(_0744_),
    .C1(net106),
    .B1(_0743_),
    .A1(_0229_),
    .Y(_0332_),
    .A2(net62));
 sg13g2_o21ai_1 _1850_ (.B1(net226),
    .Y(_0745_),
    .A1(\state[77] ),
    .A2(net201));
 sg13g2_a21o_1 _1851_ (.A2(net201),
    .A1(_0230_),
    .B1(_0745_),
    .X(_0746_));
 sg13g2_a21oi_1 _1852_ (.A1(net155),
    .A2(\daisychain[76] ),
    .Y(_0747_),
    .B1(net65));
 sg13g2_a221oi_1 _1853_ (.B2(_0747_),
    .C1(net108),
    .B1(_0746_),
    .A1(_0230_),
    .Y(_0333_),
    .A2(net65));
 sg13g2_o21ai_1 _1854_ (.B1(net224),
    .Y(_0748_),
    .A1(\state[78] ),
    .A2(net196));
 sg13g2_a21o_1 _1855_ (.A2(net196),
    .A1(_0231_),
    .B1(_0748_),
    .X(_0749_));
 sg13g2_a21oi_1 _1856_ (.A1(net151),
    .A2(\daisychain[77] ),
    .Y(_0750_),
    .B1(net60));
 sg13g2_a221oi_1 _1857_ (.B2(_0750_),
    .C1(net105),
    .B1(_0749_),
    .A1(_0231_),
    .Y(_0334_),
    .A2(net60));
 sg13g2_o21ai_1 _1858_ (.B1(net224),
    .Y(_0751_),
    .A1(\state[79] ),
    .A2(net196));
 sg13g2_a21o_1 _1859_ (.A2(net196),
    .A1(_0232_),
    .B1(_0751_),
    .X(_0752_));
 sg13g2_a21oi_1 _1860_ (.A1(net150),
    .A2(\daisychain[78] ),
    .Y(_0753_),
    .B1(net59));
 sg13g2_a221oi_1 _1861_ (.B2(_0753_),
    .C1(net104),
    .B1(_0752_),
    .A1(_0232_),
    .Y(_0335_),
    .A2(net59));
 sg13g2_o21ai_1 _1862_ (.B1(net223),
    .Y(_0754_),
    .A1(\state[80] ),
    .A2(net194));
 sg13g2_a21o_1 _1863_ (.A2(net194),
    .A1(_0234_),
    .B1(_0754_),
    .X(_0755_));
 sg13g2_a21oi_1 _1864_ (.A1(net150),
    .A2(\daisychain[79] ),
    .Y(_0756_),
    .B1(net59));
 sg13g2_a221oi_1 _1865_ (.B2(_0756_),
    .C1(net104),
    .B1(_0755_),
    .A1(_0234_),
    .Y(_0336_),
    .A2(net59));
 sg13g2_o21ai_1 _1866_ (.B1(net224),
    .Y(_0757_),
    .A1(\state[81] ),
    .A2(net197));
 sg13g2_a21o_1 _1867_ (.A2(net197),
    .A1(_0235_),
    .B1(_0757_),
    .X(_0758_));
 sg13g2_a21oi_1 _1868_ (.A1(net151),
    .A2(\daisychain[80] ),
    .Y(_0759_),
    .B1(net60));
 sg13g2_a221oi_1 _1869_ (.B2(_0759_),
    .C1(net105),
    .B1(_0758_),
    .A1(_0235_),
    .Y(_0337_),
    .A2(net60));
 sg13g2_o21ai_1 _1870_ (.B1(net211),
    .Y(_0760_),
    .A1(\state[82] ),
    .A2(net172));
 sg13g2_a21o_1 _1871_ (.A2(net172),
    .A1(_0236_),
    .B1(_0760_),
    .X(_0761_));
 sg13g2_a21oi_1 _1872_ (.A1(net123),
    .A2(\daisychain[81] ),
    .Y(_0762_),
    .B1(net35));
 sg13g2_a221oi_1 _1873_ (.B2(_0762_),
    .C1(net79),
    .B1(_0761_),
    .A1(_0236_),
    .Y(_0338_),
    .A2(net35));
 sg13g2_o21ai_1 _1874_ (.B1(net211),
    .Y(_0763_),
    .A1(\state[83] ),
    .A2(net172));
 sg13g2_a21o_1 _1875_ (.A2(net172),
    .A1(_0237_),
    .B1(_0763_),
    .X(_0764_));
 sg13g2_a21oi_1 _1876_ (.A1(net123),
    .A2(\daisychain[82] ),
    .Y(_0765_),
    .B1(net35));
 sg13g2_a221oi_1 _1877_ (.B2(_0765_),
    .C1(net79),
    .B1(_0764_),
    .A1(_0237_),
    .Y(_0339_),
    .A2(net35));
 sg13g2_o21ai_1 _1878_ (.B1(net211),
    .Y(_0766_),
    .A1(\state[84] ),
    .A2(net172));
 sg13g2_a21o_1 _1879_ (.A2(net172),
    .A1(_0238_),
    .B1(_0766_),
    .X(_0767_));
 sg13g2_a21oi_1 _1880_ (.A1(net123),
    .A2(\daisychain[83] ),
    .Y(_0768_),
    .B1(net35));
 sg13g2_a221oi_1 _1881_ (.B2(_0768_),
    .C1(net79),
    .B1(_0767_),
    .A1(_0238_),
    .Y(_0340_),
    .A2(net35));
 sg13g2_o21ai_1 _1882_ (.B1(net212),
    .Y(_0769_),
    .A1(\state[85] ),
    .A2(net173));
 sg13g2_a21o_1 _1883_ (.A2(net173),
    .A1(_0239_),
    .B1(_0769_),
    .X(_0770_));
 sg13g2_a21oi_1 _1884_ (.A1(net126),
    .A2(\daisychain[84] ),
    .Y(_0771_),
    .B1(net37));
 sg13g2_a221oi_1 _1885_ (.B2(_0771_),
    .C1(net82),
    .B1(_0770_),
    .A1(_0239_),
    .Y(_0341_),
    .A2(net37));
 sg13g2_o21ai_1 _1886_ (.B1(net212),
    .Y(_0772_),
    .A1(\state[86] ),
    .A2(net174));
 sg13g2_a21o_1 _1887_ (.A2(net174),
    .A1(_0240_),
    .B1(_0772_),
    .X(_0773_));
 sg13g2_a21oi_1 _1888_ (.A1(net127),
    .A2(\daisychain[85] ),
    .Y(_0774_),
    .B1(net38));
 sg13g2_a221oi_1 _1889_ (.B2(_0774_),
    .C1(net83),
    .B1(_0773_),
    .A1(_0240_),
    .Y(_0342_),
    .A2(net38));
 sg13g2_o21ai_1 _1890_ (.B1(net212),
    .Y(_0775_),
    .A1(\state[87] ),
    .A2(net173));
 sg13g2_a21o_1 _1891_ (.A2(net173),
    .A1(_0241_),
    .B1(_0775_),
    .X(_0776_));
 sg13g2_a21oi_1 _1892_ (.A1(net127),
    .A2(\daisychain[86] ),
    .Y(_0777_),
    .B1(net38));
 sg13g2_a221oi_1 _1893_ (.B2(_0777_),
    .C1(net83),
    .B1(_0776_),
    .A1(_0241_),
    .Y(_0343_),
    .A2(net38));
 sg13g2_o21ai_1 _1894_ (.B1(net211),
    .Y(_0778_),
    .A1(\state[88] ),
    .A2(net170));
 sg13g2_a21o_1 _1895_ (.A2(net173),
    .A1(_0242_),
    .B1(_0778_),
    .X(_0779_));
 sg13g2_a21oi_1 _1896_ (.A1(net127),
    .A2(\daisychain[87] ),
    .Y(_0780_),
    .B1(net38));
 sg13g2_a221oi_1 _1897_ (.B2(_0780_),
    .C1(net83),
    .B1(_0779_),
    .A1(_0242_),
    .Y(_0344_),
    .A2(net38));
 sg13g2_o21ai_1 _1898_ (.B1(net214),
    .Y(_0781_),
    .A1(\state[89] ),
    .A2(net178));
 sg13g2_a21o_1 _1899_ (.A2(net178),
    .A1(_0243_),
    .B1(_0781_),
    .X(_0782_));
 sg13g2_a21oi_1 _1900_ (.A1(net133),
    .A2(\daisychain[88] ),
    .Y(_0783_),
    .B1(net46));
 sg13g2_a221oi_1 _1901_ (.B2(_0783_),
    .C1(net85),
    .B1(_0782_),
    .A1(_0243_),
    .Y(_0345_),
    .A2(net42));
 sg13g2_o21ai_1 _1902_ (.B1(net223),
    .Y(_0784_),
    .A1(\state[90] ),
    .A2(net195));
 sg13g2_a21o_1 _1903_ (.A2(net195),
    .A1(_0245_),
    .B1(_0784_),
    .X(_0785_));
 sg13g2_a21oi_1 _1904_ (.A1(net150),
    .A2(\daisychain[89] ),
    .Y(_0786_),
    .B1(net59));
 sg13g2_a221oi_1 _1905_ (.B2(_0786_),
    .C1(net104),
    .B1(_0785_),
    .A1(_0245_),
    .Y(_0346_),
    .A2(net59));
 sg13g2_o21ai_1 _1906_ (.B1(net223),
    .Y(_0787_),
    .A1(\state[91] ),
    .A2(net198));
 sg13g2_a21o_1 _1907_ (.A2(net198),
    .A1(_0246_),
    .B1(_0787_),
    .X(_0788_));
 sg13g2_a21oi_1 _1908_ (.A1(net151),
    .A2(\daisychain[90] ),
    .Y(_0789_),
    .B1(net60));
 sg13g2_a221oi_1 _1909_ (.B2(_0789_),
    .C1(net105),
    .B1(_0788_),
    .A1(_0246_),
    .Y(_0347_),
    .A2(net60));
 sg13g2_o21ai_1 _1910_ (.B1(net224),
    .Y(_0790_),
    .A1(\state[92] ),
    .A2(net197));
 sg13g2_a21o_1 _1911_ (.A2(net197),
    .A1(_0247_),
    .B1(_0790_),
    .X(_0791_));
 sg13g2_a21oi_1 _1912_ (.A1(net151),
    .A2(\daisychain[91] ),
    .Y(_0792_),
    .B1(net61));
 sg13g2_a221oi_1 _1913_ (.B2(_0792_),
    .C1(net105),
    .B1(_0791_),
    .A1(_0247_),
    .Y(_0348_),
    .A2(net61));
 sg13g2_o21ai_1 _1914_ (.B1(net224),
    .Y(_0793_),
    .A1(\state[93] ),
    .A2(net196));
 sg13g2_a21o_1 _1915_ (.A2(net196),
    .A1(_0248_),
    .B1(_0793_),
    .X(_0794_));
 sg13g2_a21oi_1 _1916_ (.A1(net150),
    .A2(\daisychain[92] ),
    .Y(_0795_),
    .B1(net59));
 sg13g2_a221oi_1 _1917_ (.B2(_0795_),
    .C1(net104),
    .B1(_0794_),
    .A1(_0248_),
    .Y(_0349_),
    .A2(net59));
 sg13g2_o21ai_1 _1918_ (.B1(net215),
    .Y(_0796_),
    .A1(\state[94] ),
    .A2(net180));
 sg13g2_a21o_1 _1919_ (.A2(net180),
    .A1(_0249_),
    .B1(_0796_),
    .X(_0797_));
 sg13g2_a21oi_1 _1920_ (.A1(net134),
    .A2(\daisychain[93] ),
    .Y(_0798_),
    .B1(net47));
 sg13g2_a221oi_1 _1921_ (.B2(_0798_),
    .C1(net89),
    .B1(_0797_),
    .A1(_0249_),
    .Y(_0350_),
    .A2(net47));
 sg13g2_o21ai_1 _1922_ (.B1(net214),
    .Y(_0799_),
    .A1(\state[95] ),
    .A2(net177));
 sg13g2_a21o_1 _1923_ (.A2(net177),
    .A1(_0250_),
    .B1(_0799_),
    .X(_0800_));
 sg13g2_a21oi_1 _1924_ (.A1(net129),
    .A2(\daisychain[94] ),
    .Y(_0801_),
    .B1(net42));
 sg13g2_a221oi_1 _1925_ (.B2(_0801_),
    .C1(net85),
    .B1(_0800_),
    .A1(_0250_),
    .Y(_0351_),
    .A2(net43));
 sg13g2_o21ai_1 _1926_ (.B1(net214),
    .Y(_0802_),
    .A1(\state[96] ),
    .A2(net177));
 sg13g2_a21o_1 _1927_ (.A2(net177),
    .A1(_0251_),
    .B1(_0802_),
    .X(_0803_));
 sg13g2_a21oi_1 _1928_ (.A1(net129),
    .A2(\daisychain[95] ),
    .Y(_0804_),
    .B1(net43));
 sg13g2_a221oi_1 _1929_ (.B2(_0804_),
    .C1(net86),
    .B1(_0803_),
    .A1(_0251_),
    .Y(_0352_),
    .A2(net42));
 sg13g2_o21ai_1 _1930_ (.B1(net213),
    .Y(_0805_),
    .A1(\state[97] ),
    .A2(net175));
 sg13g2_a21o_1 _1931_ (.A2(net175),
    .A1(_0252_),
    .B1(_0805_),
    .X(_0806_));
 sg13g2_a21oi_1 _1932_ (.A1(net128),
    .A2(\daisychain[96] ),
    .Y(_0807_),
    .B1(net41));
 sg13g2_a221oi_1 _1933_ (.B2(_0807_),
    .C1(net84),
    .B1(_0806_),
    .A1(_0252_),
    .Y(_0353_),
    .A2(net41));
 sg13g2_o21ai_1 _1934_ (.B1(net213),
    .Y(_0808_),
    .A1(\state[98] ),
    .A2(net175));
 sg13g2_a21o_1 _1935_ (.A2(net176),
    .A1(_0253_),
    .B1(_0808_),
    .X(_0809_));
 sg13g2_a21oi_1 _1936_ (.A1(net128),
    .A2(\daisychain[97] ),
    .Y(_0810_),
    .B1(net41));
 sg13g2_a221oi_1 _1937_ (.B2(_0810_),
    .C1(net84),
    .B1(_0809_),
    .A1(_0253_),
    .Y(_0354_),
    .A2(net41));
 sg13g2_o21ai_1 _1938_ (.B1(net214),
    .Y(_0811_),
    .A1(\state[99] ),
    .A2(net178));
 sg13g2_a21o_1 _1939_ (.A2(net180),
    .A1(_0254_),
    .B1(_0811_),
    .X(_0812_));
 sg13g2_a21oi_1 _1940_ (.A1(net133),
    .A2(\daisychain[98] ),
    .Y(_0813_),
    .B1(net46));
 sg13g2_a221oi_1 _1941_ (.B2(_0813_),
    .C1(net89),
    .B1(_0812_),
    .A1(_0254_),
    .Y(_0355_),
    .A2(net46));
 sg13g2_o21ai_1 _1942_ (.B1(net215),
    .Y(_0814_),
    .A1(\state[100] ),
    .A2(net180));
 sg13g2_a21o_1 _1943_ (.A2(net180),
    .A1(_0129_),
    .B1(_0814_),
    .X(_0815_));
 sg13g2_a21oi_1 _1944_ (.A1(net133),
    .A2(\daisychain[99] ),
    .Y(_0816_),
    .B1(net46));
 sg13g2_a221oi_1 _1945_ (.B2(_0816_),
    .C1(net89),
    .B1(_0815_),
    .A1(_0129_),
    .Y(_0356_),
    .A2(net46));
 sg13g2_o21ai_1 _1946_ (.B1(net215),
    .Y(_0817_),
    .A1(\state[101] ),
    .A2(net181));
 sg13g2_a21o_1 _1947_ (.A2(net180),
    .A1(_0130_),
    .B1(_0817_),
    .X(_0818_));
 sg13g2_a21oi_1 _1948_ (.A1(net133),
    .A2(\daisychain[100] ),
    .Y(_0819_),
    .B1(net47));
 sg13g2_a221oi_1 _1949_ (.B2(_0819_),
    .C1(net89),
    .B1(_0818_),
    .A1(_0130_),
    .Y(_0357_),
    .A2(net47));
 sg13g2_o21ai_1 _1950_ (.B1(net224),
    .Y(_0820_),
    .A1(\state[102] ),
    .A2(net196));
 sg13g2_a21o_1 _1951_ (.A2(net196),
    .A1(_0131_),
    .B1(_0820_),
    .X(_0821_));
 sg13g2_a21oi_1 _1952_ (.A1(net150),
    .A2(\daisychain[101] ),
    .Y(_0822_),
    .B1(net61));
 sg13g2_a221oi_1 _1953_ (.B2(_0822_),
    .C1(net104),
    .B1(_0821_),
    .A1(_0131_),
    .Y(_0358_),
    .A2(net61));
 sg13g2_o21ai_1 _1954_ (.B1(net216),
    .Y(_0823_),
    .A1(\state[103] ),
    .A2(net179));
 sg13g2_a21o_1 _1955_ (.A2(net181),
    .A1(_0132_),
    .B1(_0823_),
    .X(_0824_));
 sg13g2_a21oi_1 _1956_ (.A1(net134),
    .A2(\daisychain[102] ),
    .Y(_0825_),
    .B1(net47));
 sg13g2_a221oi_1 _1957_ (.B2(_0825_),
    .C1(net87),
    .B1(_0824_),
    .A1(_0132_),
    .Y(_0359_),
    .A2(net44));
 sg13g2_o21ai_1 _1958_ (.B1(net216),
    .Y(_0826_),
    .A1(\state[104] ),
    .A2(net180));
 sg13g2_a21o_1 _1959_ (.A2(net180),
    .A1(_0133_),
    .B1(_0826_),
    .X(_0827_));
 sg13g2_a21oi_1 _1960_ (.A1(net133),
    .A2(\daisychain[103] ),
    .Y(_0828_),
    .B1(net46));
 sg13g2_a221oi_1 _1961_ (.B2(_0828_),
    .C1(net89),
    .B1(_0827_),
    .A1(_0133_),
    .Y(_0360_),
    .A2(net46));
 sg13g2_o21ai_1 _1962_ (.B1(net216),
    .Y(_0829_),
    .A1(\state[105] ),
    .A2(net181));
 sg13g2_a21o_1 _1963_ (.A2(net181),
    .A1(_0134_),
    .B1(_0829_),
    .X(_0830_));
 sg13g2_a21oi_1 _1964_ (.A1(net133),
    .A2(\daisychain[104] ),
    .Y(_0831_),
    .B1(net46));
 sg13g2_a221oi_1 _1965_ (.B2(_0831_),
    .C1(net89),
    .B1(_0830_),
    .A1(_0134_),
    .Y(_0361_),
    .A2(net47));
 sg13g2_o21ai_1 _1966_ (.B1(net215),
    .Y(_0832_),
    .A1(\state[106] ),
    .A2(net179));
 sg13g2_a21o_1 _1967_ (.A2(net182),
    .A1(_0135_),
    .B1(_0832_),
    .X(_0833_));
 sg13g2_a21oi_1 _1968_ (.A1(net131),
    .A2(\daisychain[105] ),
    .Y(_0834_),
    .B1(net45));
 sg13g2_a221oi_1 _1969_ (.B2(_0834_),
    .C1(net87),
    .B1(_0833_),
    .A1(_0135_),
    .Y(_0362_),
    .A2(net45));
 sg13g2_o21ai_1 _1970_ (.B1(net215),
    .Y(_0835_),
    .A1(\state[107] ),
    .A2(net179));
 sg13g2_a21o_1 _1971_ (.A2(net179),
    .A1(_0136_),
    .B1(_0835_),
    .X(_0836_));
 sg13g2_a21oi_1 _1972_ (.A1(net131),
    .A2(\daisychain[106] ),
    .Y(_0837_),
    .B1(net44));
 sg13g2_a221oi_1 _1973_ (.B2(_0837_),
    .C1(net87),
    .B1(_0836_),
    .A1(_0136_),
    .Y(_0363_),
    .A2(net44));
 sg13g2_o21ai_1 _1974_ (.B1(net215),
    .Y(_0838_),
    .A1(\state[108] ),
    .A2(net179));
 sg13g2_a21o_1 _1975_ (.A2(net179),
    .A1(_0137_),
    .B1(_0838_),
    .X(_0839_));
 sg13g2_a21oi_1 _1976_ (.A1(net131),
    .A2(\daisychain[107] ),
    .Y(_0840_),
    .B1(net44));
 sg13g2_a221oi_1 _1977_ (.B2(_0840_),
    .C1(net87),
    .B1(_0839_),
    .A1(_0137_),
    .Y(_0364_),
    .A2(net44));
 sg13g2_o21ai_1 _1978_ (.B1(net213),
    .Y(_0841_),
    .A1(\state[109] ),
    .A2(net176));
 sg13g2_a21o_1 _1979_ (.A2(net176),
    .A1(_0138_),
    .B1(_0841_),
    .X(_0842_));
 sg13g2_a21oi_1 _1980_ (.A1(net131),
    .A2(\daisychain[108] ),
    .Y(_0843_),
    .B1(net44));
 sg13g2_a221oi_1 _1981_ (.B2(_0843_),
    .C1(net87),
    .B1(_0842_),
    .A1(_0138_),
    .Y(_0365_),
    .A2(net44));
 sg13g2_o21ai_1 _1982_ (.B1(net213),
    .Y(_0844_),
    .A1(\state[110] ),
    .A2(net175));
 sg13g2_a21o_1 _1983_ (.A2(net176),
    .A1(_0140_),
    .B1(_0844_),
    .X(_0845_));
 sg13g2_a21oi_1 _1984_ (.A1(net128),
    .A2(\daisychain[109] ),
    .Y(_0846_),
    .B1(net43));
 sg13g2_a221oi_1 _1985_ (.B2(_0846_),
    .C1(net84),
    .B1(_0845_),
    .A1(_0140_),
    .Y(_0366_),
    .A2(net43));
 sg13g2_o21ai_1 _1986_ (.B1(net213),
    .Y(_0847_),
    .A1(\state[111] ),
    .A2(net170));
 sg13g2_a21o_1 _1987_ (.A2(net175),
    .A1(_0141_),
    .B1(_0847_),
    .X(_0848_));
 sg13g2_a21oi_1 _1988_ (.A1(net128),
    .A2(\daisychain[110] ),
    .Y(_0849_),
    .B1(net43));
 sg13g2_a221oi_1 _1989_ (.B2(_0849_),
    .C1(net80),
    .B1(_0848_),
    .A1(_0141_),
    .Y(_0367_),
    .A2(net34));
 sg13g2_o21ai_1 _1990_ (.B1(net212),
    .Y(_0850_),
    .A1(\state[112] ),
    .A2(net170));
 sg13g2_a21o_1 _1991_ (.A2(net170),
    .A1(_0142_),
    .B1(_0850_),
    .X(_0851_));
 sg13g2_a21oi_1 _1992_ (.A1(net124),
    .A2(\daisychain[111] ),
    .Y(_0852_),
    .B1(net34));
 sg13g2_a221oi_1 _1993_ (.B2(_0852_),
    .C1(net80),
    .B1(_0851_),
    .A1(_0142_),
    .Y(_0368_),
    .A2(net36));
 sg13g2_o21ai_1 _1994_ (.B1(net212),
    .Y(_0853_),
    .A1(\state[113] ),
    .A2(net171));
 sg13g2_a21o_1 _1995_ (.A2(net171),
    .A1(_0143_),
    .B1(_0853_),
    .X(_0854_));
 sg13g2_a21oi_1 _1996_ (.A1(net124),
    .A2(\daisychain[112] ),
    .Y(_0855_),
    .B1(net36));
 sg13g2_a221oi_1 _1997_ (.B2(_0855_),
    .C1(net81),
    .B1(_0854_),
    .A1(_0143_),
    .Y(_0369_),
    .A2(net36));
 sg13g2_o21ai_1 _1998_ (.B1(net212),
    .Y(_0856_),
    .A1(\state[114] ),
    .A2(net171));
 sg13g2_a21o_1 _1999_ (.A2(net171),
    .A1(_0144_),
    .B1(_0856_),
    .X(_0857_));
 sg13g2_a21oi_1 _2000_ (.A1(net126),
    .A2(\daisychain[113] ),
    .Y(_0858_),
    .B1(net37));
 sg13g2_a221oi_1 _2001_ (.B2(_0858_),
    .C1(net82),
    .B1(_0857_),
    .A1(_0144_),
    .Y(_0370_),
    .A2(net37));
 sg13g2_o21ai_1 _2002_ (.B1(net215),
    .Y(_0859_),
    .A1(\state[115] ),
    .A2(net179));
 sg13g2_a21o_1 _2003_ (.A2(net179),
    .A1(_0145_),
    .B1(_0859_),
    .X(_0860_));
 sg13g2_a21oi_1 _2004_ (.A1(net131),
    .A2(\daisychain[114] ),
    .Y(_0861_),
    .B1(net37));
 sg13g2_a221oi_1 _2005_ (.B2(_0861_),
    .C1(net87),
    .B1(_0860_),
    .A1(_0145_),
    .Y(_0371_),
    .A2(net44));
 sg13g2_o21ai_1 _2006_ (.B1(net215),
    .Y(_0862_),
    .A1(\state[116] ),
    .A2(net182));
 sg13g2_a21o_1 _2007_ (.A2(net182),
    .A1(_0146_),
    .B1(_0862_),
    .X(_0863_));
 sg13g2_a21oi_1 _2008_ (.A1(net132),
    .A2(\daisychain[115] ),
    .Y(_0864_),
    .B1(net45));
 sg13g2_a221oi_1 _2009_ (.B2(_0864_),
    .C1(net88),
    .B1(_0863_),
    .A1(_0146_),
    .Y(_0372_),
    .A2(net45));
 sg13g2_o21ai_1 _2010_ (.B1(net212),
    .Y(_0865_),
    .A1(\state[117] ),
    .A2(net173));
 sg13g2_a21o_1 _2011_ (.A2(net174),
    .A1(_0147_),
    .B1(_0865_),
    .X(_0866_));
 sg13g2_a21oi_1 _2012_ (.A1(net126),
    .A2(\daisychain[116] ),
    .Y(_0867_),
    .B1(net37));
 sg13g2_a221oi_1 _2013_ (.B2(_0867_),
    .C1(net82),
    .B1(_0866_),
    .A1(_0147_),
    .Y(_0373_),
    .A2(net39));
 sg13g2_o21ai_1 _2014_ (.B1(net217),
    .Y(_0868_),
    .A1(\state[118] ),
    .A2(net174));
 sg13g2_a21o_1 _2015_ (.A2(net174),
    .A1(_0148_),
    .B1(_0868_),
    .X(_0869_));
 sg13g2_a21oi_1 _2016_ (.A1(net126),
    .A2(\daisychain[117] ),
    .Y(_0870_),
    .B1(net39));
 sg13g2_a221oi_1 _2017_ (.B2(_0870_),
    .C1(net82),
    .B1(_0869_),
    .A1(_0148_),
    .Y(_0374_),
    .A2(net39));
 sg13g2_o21ai_1 _2018_ (.B1(net217),
    .Y(_0871_),
    .A1(\state[119] ),
    .A2(net173));
 sg13g2_a21o_1 _2019_ (.A2(net173),
    .A1(_0149_),
    .B1(_0871_),
    .X(_0872_));
 sg13g2_a21oi_1 _2020_ (.A1(net126),
    .A2(\daisychain[118] ),
    .Y(_0873_),
    .B1(net37));
 sg13g2_a221oi_1 _2021_ (.B2(_0873_),
    .C1(net82),
    .B1(_0872_),
    .A1(_0149_),
    .Y(_0375_),
    .A2(net37));
 sg13g2_o21ai_1 _2022_ (.B1(net217),
    .Y(_0874_),
    .A1(\state[120] ),
    .A2(net174));
 sg13g2_a21o_1 _2023_ (.A2(net174),
    .A1(_0151_),
    .B1(_0874_),
    .X(_0875_));
 sg13g2_a21oi_1 _2024_ (.A1(net127),
    .A2(\daisychain[119] ),
    .Y(_0876_),
    .B1(net38));
 sg13g2_a221oi_1 _2025_ (.B2(_0876_),
    .C1(net83),
    .B1(_0875_),
    .A1(_0151_),
    .Y(_0376_),
    .A2(net38));
 sg13g2_o21ai_1 _2026_ (.B1(net205),
    .Y(_0877_),
    .A1(\state[121] ),
    .A2(net159));
 sg13g2_a21o_1 _2027_ (.A2(net159),
    .A1(_0152_),
    .B1(_0877_),
    .X(_0878_));
 sg13g2_a21oi_1 _2028_ (.A1(net113),
    .A2(\daisychain[120] ),
    .Y(_0879_),
    .B1(net24));
 sg13g2_a221oi_1 _2029_ (.B2(_0879_),
    .C1(net69),
    .B1(_0878_),
    .A1(_0152_),
    .Y(_0377_),
    .A2(net24));
 sg13g2_o21ai_1 _2030_ (.B1(net205),
    .Y(_0880_),
    .A1(\state[122] ),
    .A2(net160));
 sg13g2_a21o_1 _2031_ (.A2(net160),
    .A1(_0153_),
    .B1(_0880_),
    .X(_0881_));
 sg13g2_a21oi_1 _2032_ (.A1(net114),
    .A2(\daisychain[121] ),
    .Y(_0882_),
    .B1(net25));
 sg13g2_a221oi_1 _2033_ (.B2(_0882_),
    .C1(net70),
    .B1(_0881_),
    .A1(_0153_),
    .Y(_0378_),
    .A2(net25));
 sg13g2_o21ai_1 _2034_ (.B1(net210),
    .Y(_0883_),
    .A1(\state[123] ),
    .A2(net160));
 sg13g2_a21o_1 _2035_ (.A2(net160),
    .A1(_0154_),
    .B1(_0883_),
    .X(_0884_));
 sg13g2_a21oi_1 _2036_ (.A1(net115),
    .A2(\daisychain[122] ),
    .Y(_0885_),
    .B1(net25));
 sg13g2_a221oi_1 _2037_ (.B2(_0885_),
    .C1(net71),
    .B1(_0884_),
    .A1(_0154_),
    .Y(_0379_),
    .A2(net25));
 sg13g2_o21ai_1 _2038_ (.B1(net210),
    .Y(_0886_),
    .A1(\state[124] ),
    .A2(net159));
 sg13g2_a21o_1 _2039_ (.A2(net161),
    .A1(_0155_),
    .B1(_0886_),
    .X(_0887_));
 sg13g2_a21oi_1 _2040_ (.A1(net113),
    .A2(\daisychain[123] ),
    .Y(_0888_),
    .B1(net24));
 sg13g2_a221oi_1 _2041_ (.B2(_0888_),
    .C1(net71),
    .B1(_0887_),
    .A1(_0155_),
    .Y(_0380_),
    .A2(net24));
 sg13g2_o21ai_1 _2042_ (.B1(net205),
    .Y(_0889_),
    .A1(\state[125] ),
    .A2(net159));
 sg13g2_a21o_1 _2043_ (.A2(net159),
    .A1(_0156_),
    .B1(_0889_),
    .X(_0890_));
 sg13g2_a21oi_1 _2044_ (.A1(net113),
    .A2(\daisychain[124] ),
    .Y(_0891_),
    .B1(net24));
 sg13g2_a221oi_1 _2045_ (.B2(_0891_),
    .C1(net69),
    .B1(_0890_),
    .A1(_0156_),
    .Y(_0381_),
    .A2(net24));
 sg13g2_o21ai_1 _2046_ (.B1(net205),
    .Y(_0892_),
    .A1(\state[126] ),
    .A2(net159));
 sg13g2_a21o_1 _2047_ (.A2(net159),
    .A1(_0157_),
    .B1(_0892_),
    .X(_0893_));
 sg13g2_a21oi_1 _2048_ (.A1(net113),
    .A2(\daisychain[125] ),
    .Y(_0894_),
    .B1(net24));
 sg13g2_a221oi_1 _2049_ (.B2(_0894_),
    .C1(net69),
    .B1(_0893_),
    .A1(_0157_),
    .Y(_0382_),
    .A2(net24));
 sg13g2_o21ai_1 _2050_ (.B1(net205),
    .Y(_0895_),
    .A1(\state[127] ),
    .A2(net159));
 sg13g2_a21o_1 _2051_ (.A2(net161),
    .A1(_0158_),
    .B1(_0895_),
    .X(_0896_));
 sg13g2_a21oi_1 _2052_ (.A1(net113),
    .A2(\daisychain[126] ),
    .Y(_0897_),
    .B1(net26));
 sg13g2_a221oi_1 _2053_ (.B2(_0897_),
    .C1(net69),
    .B1(_0896_),
    .A1(_0158_),
    .Y(_0383_),
    .A2(net26));
 sg13g2_nand2_1 _2054_ (.Y(_0898_),
    .A(net123),
    .B(\state[0] ));
 sg13g2_a21oi_1 _2055_ (.A1(_0514_),
    .A2(_0898_),
    .Y(_0384_),
    .B1(net79));
 sg13g2_nand2_1 _2056_ (.Y(_0899_),
    .A(net124),
    .B(\state[1] ));
 sg13g2_a21oi_1 _2057_ (.A1(_0518_),
    .A2(_0899_),
    .Y(_0385_),
    .B1(net80));
 sg13g2_nand2_1 _2058_ (.Y(_0900_),
    .A(net115),
    .B(\state[2] ));
 sg13g2_a21oi_1 _2059_ (.A1(_0521_),
    .A2(_0900_),
    .Y(_0386_),
    .B1(net71));
 sg13g2_nand2_1 _2060_ (.Y(_0901_),
    .A(net115),
    .B(\state[3] ));
 sg13g2_a21oi_1 _2061_ (.A1(_0524_),
    .A2(_0901_),
    .Y(_0387_),
    .B1(net71));
 sg13g2_nand2_1 _2062_ (.Y(_0902_),
    .A(net118),
    .B(\state[4] ));
 sg13g2_a21oi_1 _2063_ (.A1(_0527_),
    .A2(_0902_),
    .Y(_0388_),
    .B1(net77));
 sg13g2_nand2_1 _2064_ (.Y(_0903_),
    .A(net121),
    .B(\state[5] ));
 sg13g2_a21oi_1 _2065_ (.A1(_0530_),
    .A2(_0903_),
    .Y(_0389_),
    .B1(net77));
 sg13g2_nand2_1 _2066_ (.Y(_0904_),
    .A(net114),
    .B(\state[6] ));
 sg13g2_a21oi_1 _2067_ (.A1(_0533_),
    .A2(_0904_),
    .Y(_0390_),
    .B1(net70));
 sg13g2_nand2_1 _2068_ (.Y(_0905_),
    .A(net114),
    .B(\state[7] ));
 sg13g2_a21oi_1 _2069_ (.A1(_0536_),
    .A2(_0905_),
    .Y(_0391_),
    .B1(net70));
 sg13g2_nand2_1 _2070_ (.Y(_0906_),
    .A(net137),
    .B(\state[8] ));
 sg13g2_a21oi_1 _2071_ (.A1(_0539_),
    .A2(_0906_),
    .Y(_0392_),
    .B1(net78));
 sg13g2_nand2_1 _2072_ (.Y(_0907_),
    .A(net117),
    .B(\state[9] ));
 sg13g2_a21oi_1 _2073_ (.A1(_0542_),
    .A2(_0907_),
    .Y(_0393_),
    .B1(net74));
 sg13g2_nand2_1 _2074_ (.Y(_0908_),
    .A(net117),
    .B(\state[10] ));
 sg13g2_a21oi_1 _2075_ (.A1(_0545_),
    .A2(_0908_),
    .Y(_0394_),
    .B1(net74));
 sg13g2_nand2_1 _2076_ (.Y(_0909_),
    .A(net116),
    .B(\state[11] ));
 sg13g2_a21oi_1 _2077_ (.A1(_0548_),
    .A2(_0909_),
    .Y(_0395_),
    .B1(net73));
 sg13g2_nand2_1 _2078_ (.Y(_0910_),
    .A(net116),
    .B(\state[12] ));
 sg13g2_a21oi_1 _2079_ (.A1(_0551_),
    .A2(_0910_),
    .Y(_0396_),
    .B1(net73));
 sg13g2_nand2_1 _2080_ (.Y(_0911_),
    .A(net138),
    .B(\state[13] ));
 sg13g2_a21oi_1 _2081_ (.A1(_0554_),
    .A2(_0911_),
    .Y(_0397_),
    .B1(net92));
 sg13g2_nand2_1 _2082_ (.Y(_0912_),
    .A(net116),
    .B(\state[14] ));
 sg13g2_a21oi_1 _2083_ (.A1(_0557_),
    .A2(_0912_),
    .Y(_0398_),
    .B1(net73));
 sg13g2_nand2_1 _2084_ (.Y(_0913_),
    .A(net120),
    .B(\state[15] ));
 sg13g2_a21oi_1 _2085_ (.A1(_0560_),
    .A2(_0913_),
    .Y(_0399_),
    .B1(net77));
 sg13g2_nand2_1 _2086_ (.Y(_0914_),
    .A(net120),
    .B(\state[16] ));
 sg13g2_a21oi_1 _2087_ (.A1(_0563_),
    .A2(_0914_),
    .Y(_0400_),
    .B1(net85));
 sg13g2_nand2_1 _2088_ (.Y(_0915_),
    .A(net140),
    .B(\state[17] ));
 sg13g2_a21oi_1 _2089_ (.A1(_0566_),
    .A2(_0915_),
    .Y(_0401_),
    .B1(net94));
 sg13g2_nand2_1 _2090_ (.Y(_0916_),
    .A(net129),
    .B(\state[18] ));
 sg13g2_a21oi_1 _2091_ (.A1(_0569_),
    .A2(_0916_),
    .Y(_0402_),
    .B1(net85));
 sg13g2_nand2_1 _2092_ (.Y(_0917_),
    .A(net121),
    .B(\state[19] ));
 sg13g2_a21oi_1 _2093_ (.A1(_0572_),
    .A2(_0917_),
    .Y(_0403_),
    .B1(net84));
 sg13g2_nand2_1 _2094_ (.Y(_0918_),
    .A(net118),
    .B(\state[20] ));
 sg13g2_a21oi_1 _2095_ (.A1(_0575_),
    .A2(_0918_),
    .Y(_0404_),
    .B1(net75));
 sg13g2_nand2_1 _2096_ (.Y(_0919_),
    .A(net118),
    .B(\state[21] ));
 sg13g2_a21oi_1 _2097_ (.A1(_0578_),
    .A2(_0919_),
    .Y(_0405_),
    .B1(net75));
 sg13g2_nand2_1 _2098_ (.Y(_0920_),
    .A(net148),
    .B(\state[22] ));
 sg13g2_a21oi_1 _2099_ (.A1(_0581_),
    .A2(_0920_),
    .Y(_0406_),
    .B1(net102));
 sg13g2_nand2_1 _2100_ (.Y(_0921_),
    .A(net148),
    .B(\state[23] ));
 sg13g2_a21oi_1 _2101_ (.A1(_0584_),
    .A2(_0921_),
    .Y(_0407_),
    .B1(net102));
 sg13g2_nand2_1 _2102_ (.Y(_0922_),
    .A(net149),
    .B(\state[24] ));
 sg13g2_a21oi_1 _2103_ (.A1(_0587_),
    .A2(_0922_),
    .Y(_0408_),
    .B1(net103));
 sg13g2_nand2_1 _2104_ (.Y(_0923_),
    .A(net140),
    .B(\state[25] ));
 sg13g2_a21oi_1 _2105_ (.A1(_0590_),
    .A2(_0923_),
    .Y(_0409_),
    .B1(net102));
 sg13g2_nand2_1 _2106_ (.Y(_0924_),
    .A(net119),
    .B(\state[26] ));
 sg13g2_a21oi_1 _2107_ (.A1(_0593_),
    .A2(_0924_),
    .Y(_0410_),
    .B1(net76));
 sg13g2_nand2_1 _2108_ (.Y(_0925_),
    .A(net119),
    .B(\state[27] ));
 sg13g2_a21oi_1 _2109_ (.A1(_0596_),
    .A2(_0925_),
    .Y(_0411_),
    .B1(net76));
 sg13g2_nand2_1 _2110_ (.Y(_0926_),
    .A(net118),
    .B(\state[28] ));
 sg13g2_a21oi_1 _2111_ (.A1(_0599_),
    .A2(_0926_),
    .Y(_0412_),
    .B1(net75));
 sg13g2_nand2_1 _2112_ (.Y(_0927_),
    .A(net121),
    .B(\state[29] ));
 sg13g2_a21oi_1 _2113_ (.A1(_0602_),
    .A2(_0927_),
    .Y(_0413_),
    .B1(net77));
 sg13g2_nand2_1 _2114_ (.Y(_0928_),
    .A(net120),
    .B(\state[30] ));
 sg13g2_a21oi_1 _2115_ (.A1(_0605_),
    .A2(_0928_),
    .Y(_0414_),
    .B1(net77));
 sg13g2_nand2_1 _2116_ (.Y(_0929_),
    .A(net122),
    .B(\state[31] ));
 sg13g2_a21oi_1 _2117_ (.A1(_0608_),
    .A2(_0929_),
    .Y(_0415_),
    .B1(net73));
 sg13g2_nand2_1 _2118_ (.Y(_0930_),
    .A(net119),
    .B(\state[32] ));
 sg13g2_a21oi_1 _2119_ (.A1(_0611_),
    .A2(_0930_),
    .Y(_0416_),
    .B1(net76));
 sg13g2_nand2_1 _2120_ (.Y(_0931_),
    .A(net122),
    .B(\state[33] ));
 sg13g2_a21oi_1 _2121_ (.A1(_0614_),
    .A2(_0931_),
    .Y(_0417_),
    .B1(net78));
 sg13g2_nand2_1 _2122_ (.Y(_0932_),
    .A(net117),
    .B(\state[34] ));
 sg13g2_a21oi_1 _2123_ (.A1(_0617_),
    .A2(_0932_),
    .Y(_0418_),
    .B1(net74));
 sg13g2_nand2_1 _2124_ (.Y(_0933_),
    .A(net138),
    .B(\state[35] ));
 sg13g2_a21oi_1 _2125_ (.A1(_0620_),
    .A2(_0933_),
    .Y(_0419_),
    .B1(net92));
 sg13g2_nand2_1 _2126_ (.Y(_0934_),
    .A(net117),
    .B(\state[36] ));
 sg13g2_a21oi_1 _2127_ (.A1(_0623_),
    .A2(_0934_),
    .Y(_0420_),
    .B1(net74));
 sg13g2_nand2_1 _2128_ (.Y(_0935_),
    .A(net138),
    .B(\state[37] ));
 sg13g2_a21oi_1 _2129_ (.A1(_0626_),
    .A2(_0935_),
    .Y(_0421_),
    .B1(net92));
 sg13g2_nand2_1 _2130_ (.Y(_0936_),
    .A(net138),
    .B(\state[38] ));
 sg13g2_a21oi_1 _2131_ (.A1(_0629_),
    .A2(_0936_),
    .Y(_0422_),
    .B1(net92));
 sg13g2_nand2_1 _2132_ (.Y(_0937_),
    .A(net149),
    .B(\state[39] ));
 sg13g2_a21oi_1 _2133_ (.A1(_0632_),
    .A2(_0937_),
    .Y(_0423_),
    .B1(net103));
 sg13g2_nand2_1 _2134_ (.Y(_0938_),
    .A(net141),
    .B(\state[40] ));
 sg13g2_a21oi_1 _2135_ (.A1(_0635_),
    .A2(_0938_),
    .Y(_0424_),
    .B1(net95));
 sg13g2_nand2_1 _2136_ (.Y(_0939_),
    .A(net138),
    .B(\state[41] ));
 sg13g2_a21oi_1 _2137_ (.A1(_0638_),
    .A2(_0939_),
    .Y(_0425_),
    .B1(net92));
 sg13g2_nand2_1 _2138_ (.Y(_0940_),
    .A(net138),
    .B(\state[42] ));
 sg13g2_a21oi_1 _2139_ (.A1(_0641_),
    .A2(_0940_),
    .Y(_0426_),
    .B1(net92));
 sg13g2_nand2_1 _2140_ (.Y(_0941_),
    .A(net138),
    .B(\state[43] ));
 sg13g2_a21oi_1 _2141_ (.A1(_0644_),
    .A2(_0941_),
    .Y(_0427_),
    .B1(net93));
 sg13g2_nand2_1 _2142_ (.Y(_0942_),
    .A(net139),
    .B(\state[44] ));
 sg13g2_a21oi_1 _2143_ (.A1(_0647_),
    .A2(_0942_),
    .Y(_0428_),
    .B1(net93));
 sg13g2_nand2_1 _2144_ (.Y(_0943_),
    .A(net139),
    .B(\state[45] ));
 sg13g2_a21oi_1 _2145_ (.A1(_0650_),
    .A2(_0943_),
    .Y(_0429_),
    .B1(net93));
 sg13g2_nand2_1 _2146_ (.Y(_0944_),
    .A(net139),
    .B(\state[46] ));
 sg13g2_a21oi_1 _2147_ (.A1(_0653_),
    .A2(_0944_),
    .Y(_0430_),
    .B1(net93));
 sg13g2_nand2_1 _2148_ (.Y(_0945_),
    .A(net139),
    .B(\state[47] ));
 sg13g2_a21oi_1 _2149_ (.A1(_0656_),
    .A2(_0945_),
    .Y(_0431_),
    .B1(net93));
 sg13g2_nand2_1 _2150_ (.Y(_0946_),
    .A(net145),
    .B(\state[48] ));
 sg13g2_a21oi_1 _2151_ (.A1(_0659_),
    .A2(_0946_),
    .Y(_0432_),
    .B1(net99));
 sg13g2_nand2_1 _2152_ (.Y(_0947_),
    .A(net144),
    .B(\state[49] ));
 sg13g2_a21oi_1 _2153_ (.A1(_0662_),
    .A2(_0947_),
    .Y(_0433_),
    .B1(net97));
 sg13g2_nand2_1 _2154_ (.Y(_0948_),
    .A(net139),
    .B(\state[50] ));
 sg13g2_a21oi_1 _2155_ (.A1(_0665_),
    .A2(_0948_),
    .Y(_0434_),
    .B1(net93));
 sg13g2_nand2_1 _2156_ (.Y(_0949_),
    .A(net144),
    .B(\state[51] ));
 sg13g2_a21oi_1 _2157_ (.A1(_0668_),
    .A2(_0949_),
    .Y(_0435_),
    .B1(net97));
 sg13g2_nand2_1 _2158_ (.Y(_0950_),
    .A(net144),
    .B(\state[52] ));
 sg13g2_a21oi_1 _2159_ (.A1(_0671_),
    .A2(_0950_),
    .Y(_0436_),
    .B1(net97));
 sg13g2_nand2_1 _2160_ (.Y(_0951_),
    .A(net143),
    .B(\state[53] ));
 sg13g2_a21oi_1 _2161_ (.A1(_0674_),
    .A2(_0951_),
    .Y(_0437_),
    .B1(net98));
 sg13g2_nand2_1 _2162_ (.Y(_0952_),
    .A(net145),
    .B(\state[54] ));
 sg13g2_a21oi_1 _2163_ (.A1(_0677_),
    .A2(_0952_),
    .Y(_0438_),
    .B1(net99));
 sg13g2_nand2_1 _2164_ (.Y(_0953_),
    .A(net146),
    .B(\state[55] ));
 sg13g2_a21oi_1 _2165_ (.A1(_0680_),
    .A2(_0953_),
    .Y(_0439_),
    .B1(net100));
 sg13g2_nand2_1 _2166_ (.Y(_0954_),
    .A(net143),
    .B(\state[56] ));
 sg13g2_a21oi_1 _2167_ (.A1(_0683_),
    .A2(_0954_),
    .Y(_0440_),
    .B1(net98));
 sg13g2_nand2_1 _2168_ (.Y(_0955_),
    .A(net143),
    .B(\state[57] ));
 sg13g2_a21oi_1 _2169_ (.A1(_0686_),
    .A2(_0955_),
    .Y(_0441_),
    .B1(net97));
 sg13g2_nand2_1 _2170_ (.Y(_0956_),
    .A(net144),
    .B(\state[58] ));
 sg13g2_a21oi_1 _2171_ (.A1(_0689_),
    .A2(_0956_),
    .Y(_0442_),
    .B1(net97));
 sg13g2_nand2_1 _2172_ (.Y(_0957_),
    .A(net143),
    .B(\state[59] ));
 sg13g2_a21oi_1 _2173_ (.A1(_0692_),
    .A2(_0957_),
    .Y(_0443_),
    .B1(net98));
 sg13g2_nand2_1 _2174_ (.Y(_0958_),
    .A(net143),
    .B(\state[60] ));
 sg13g2_a21oi_1 _2175_ (.A1(_0695_),
    .A2(_0958_),
    .Y(_0444_),
    .B1(net98));
 sg13g2_nand2_1 _2176_ (.Y(_0959_),
    .A(net143),
    .B(\state[61] ));
 sg13g2_a21oi_1 _2177_ (.A1(_0698_),
    .A2(_0959_),
    .Y(_0445_),
    .B1(net98));
 sg13g2_nand2_1 _2178_ (.Y(_0960_),
    .A(net144),
    .B(\state[62] ));
 sg13g2_a21oi_1 _2179_ (.A1(_0701_),
    .A2(_0960_),
    .Y(_0446_),
    .B1(net98));
 sg13g2_nand2_1 _2180_ (.Y(_0961_),
    .A(net146),
    .B(\state[63] ));
 sg13g2_a21oi_1 _2181_ (.A1(_0704_),
    .A2(_0961_),
    .Y(_0447_),
    .B1(net100));
 sg13g2_nand2_1 _2182_ (.Y(_0962_),
    .A(net153),
    .B(\state[64] ));
 sg13g2_a21oi_1 _2183_ (.A1(_0707_),
    .A2(_0962_),
    .Y(_0448_),
    .B1(net107));
 sg13g2_nand2_1 _2184_ (.Y(_0963_),
    .A(net153),
    .B(\state[65] ));
 sg13g2_a21oi_1 _2185_ (.A1(_0710_),
    .A2(_0963_),
    .Y(_0449_),
    .B1(net107));
 sg13g2_nand2_1 _2186_ (.Y(_0964_),
    .A(net153),
    .B(\state[66] ));
 sg13g2_a21oi_1 _2187_ (.A1(_0713_),
    .A2(_0964_),
    .Y(_0450_),
    .B1(net107));
 sg13g2_nand2_1 _2188_ (.Y(_0965_),
    .A(net156),
    .B(\state[67] ));
 sg13g2_a21oi_1 _2189_ (.A1(_0716_),
    .A2(_0965_),
    .Y(_0451_),
    .B1(net109));
 sg13g2_nand2_1 _2190_ (.Y(_0966_),
    .A(net156),
    .B(\state[68] ));
 sg13g2_a21oi_1 _2191_ (.A1(_0719_),
    .A2(_0966_),
    .Y(_0452_),
    .B1(net109));
 sg13g2_nand2_1 _2192_ (.Y(_0967_),
    .A(net156),
    .B(\state[69] ));
 sg13g2_a21oi_1 _2193_ (.A1(_0722_),
    .A2(_0967_),
    .Y(_0453_),
    .B1(net109));
 sg13g2_nand2_1 _2194_ (.Y(_0968_),
    .A(net155),
    .B(\state[70] ));
 sg13g2_a21oi_1 _2195_ (.A1(_0725_),
    .A2(_0968_),
    .Y(_0454_),
    .B1(net108));
 sg13g2_nand2_1 _2196_ (.Y(_0969_),
    .A(net151),
    .B(\state[71] ));
 sg13g2_a21oi_1 _2197_ (.A1(_0728_),
    .A2(_0969_),
    .Y(_0455_),
    .B1(net105));
 sg13g2_nand2_1 _2198_ (.Y(_0970_),
    .A(net155),
    .B(\state[72] ));
 sg13g2_a21oi_1 _2199_ (.A1(_0731_),
    .A2(_0970_),
    .Y(_0456_),
    .B1(net108));
 sg13g2_nand2_1 _2200_ (.Y(_0971_),
    .A(net156),
    .B(\state[73] ));
 sg13g2_a21oi_1 _2201_ (.A1(_0734_),
    .A2(_0971_),
    .Y(_0457_),
    .B1(net109));
 sg13g2_nand2_1 _2202_ (.Y(_0972_),
    .A(net154),
    .B(\state[74] ));
 sg13g2_a21oi_1 _2203_ (.A1(_0737_),
    .A2(_0972_),
    .Y(_0458_),
    .B1(net106));
 sg13g2_nand2_1 _2204_ (.Y(_0973_),
    .A(net154),
    .B(\state[75] ));
 sg13g2_a21oi_1 _2205_ (.A1(_0740_),
    .A2(_0973_),
    .Y(_0459_),
    .B1(net106));
 sg13g2_nand2_1 _2206_ (.Y(_0974_),
    .A(net154),
    .B(\state[76] ));
 sg13g2_a21oi_1 _2207_ (.A1(_0743_),
    .A2(_0974_),
    .Y(_0460_),
    .B1(net106));
 sg13g2_nand2_1 _2208_ (.Y(_0975_),
    .A(net155),
    .B(\state[77] ));
 sg13g2_a21oi_1 _2209_ (.A1(_0746_),
    .A2(_0975_),
    .Y(_0461_),
    .B1(net108));
 sg13g2_nand2_1 _2210_ (.Y(_0976_),
    .A(net150),
    .B(\state[78] ));
 sg13g2_a21oi_1 _2211_ (.A1(_0749_),
    .A2(_0976_),
    .Y(_0462_),
    .B1(net104));
 sg13g2_nand2_1 _2212_ (.Y(_0977_),
    .A(net150),
    .B(\state[79] ));
 sg13g2_a21oi_1 _2213_ (.A1(_0752_),
    .A2(_0977_),
    .Y(_0463_),
    .B1(net104));
 sg13g2_nand2_1 _2214_ (.Y(_0978_),
    .A(net148),
    .B(\state[80] ));
 sg13g2_a21oi_1 _2215_ (.A1(_0755_),
    .A2(_0978_),
    .Y(_0464_),
    .B1(net102));
 sg13g2_nand2_1 _2216_ (.Y(_0979_),
    .A(net151),
    .B(\state[81] ));
 sg13g2_a21oi_1 _2217_ (.A1(_0758_),
    .A2(_0979_),
    .Y(_0465_),
    .B1(net105));
 sg13g2_nand2_1 _2218_ (.Y(_0980_),
    .A(net123),
    .B(\state[82] ));
 sg13g2_a21oi_1 _2219_ (.A1(_0761_),
    .A2(_0980_),
    .Y(_0466_),
    .B1(net79));
 sg13g2_nand2_1 _2220_ (.Y(_0981_),
    .A(net123),
    .B(\state[83] ));
 sg13g2_a21oi_1 _2221_ (.A1(_0764_),
    .A2(_0981_),
    .Y(_0467_),
    .B1(net79));
 sg13g2_nand2_1 _2222_ (.Y(_0982_),
    .A(net123),
    .B(\state[84] ));
 sg13g2_a21oi_1 _2223_ (.A1(_0767_),
    .A2(_0982_),
    .Y(_0468_),
    .B1(net79));
 sg13g2_nand2_1 _2224_ (.Y(_0983_),
    .A(net126),
    .B(\state[85] ));
 sg13g2_a21oi_1 _2225_ (.A1(_0770_),
    .A2(_0983_),
    .Y(_0469_),
    .B1(net83));
 sg13g2_nand2_1 _2226_ (.Y(_0984_),
    .A(net127),
    .B(\state[86] ));
 sg13g2_a21oi_1 _2227_ (.A1(_0773_),
    .A2(_0984_),
    .Y(_0470_),
    .B1(net83));
 sg13g2_nand2_1 _2228_ (.Y(_0985_),
    .A(net126),
    .B(\state[87] ));
 sg13g2_a21oi_1 _2229_ (.A1(_0776_),
    .A2(_0985_),
    .Y(_0471_),
    .B1(net82));
 sg13g2_nand2_1 _2230_ (.Y(_0986_),
    .A(net125),
    .B(\state[88] ));
 sg13g2_a21oi_1 _2231_ (.A1(_0779_),
    .A2(_0986_),
    .Y(_0472_),
    .B1(net81));
 sg13g2_nand2_1 _2232_ (.Y(_0987_),
    .A(net130),
    .B(\state[89] ));
 sg13g2_a21oi_1 _2233_ (.A1(_0782_),
    .A2(_0987_),
    .Y(_0473_),
    .B1(net86));
 sg13g2_nand2_1 _2234_ (.Y(_0988_),
    .A(net148),
    .B(\state[90] ));
 sg13g2_a21oi_1 _2235_ (.A1(_0785_),
    .A2(_0988_),
    .Y(_0474_),
    .B1(net103));
 sg13g2_nand2_1 _2236_ (.Y(_0989_),
    .A(net149),
    .B(\state[91] ));
 sg13g2_a21oi_1 _2237_ (.A1(_0788_),
    .A2(_0989_),
    .Y(_0475_),
    .B1(net103));
 sg13g2_nand2_1 _2238_ (.Y(_0990_),
    .A(net151),
    .B(\state[92] ));
 sg13g2_a21oi_1 _2239_ (.A1(_0791_),
    .A2(_0990_),
    .Y(_0476_),
    .B1(net105));
 sg13g2_nand2_1 _2240_ (.Y(_0991_),
    .A(net150),
    .B(\state[93] ));
 sg13g2_a21oi_1 _2241_ (.A1(_0794_),
    .A2(_0991_),
    .Y(_0477_),
    .B1(net104));
 sg13g2_nand2_1 _2242_ (.Y(_0992_),
    .A(net134),
    .B(\state[94] ));
 sg13g2_a21oi_1 _2243_ (.A1(_0797_),
    .A2(_0992_),
    .Y(_0478_),
    .B1(net90));
 sg13g2_nand2_1 _2244_ (.Y(_0993_),
    .A(net129),
    .B(\state[95] ));
 sg13g2_a21oi_1 _2245_ (.A1(_0800_),
    .A2(_0993_),
    .Y(_0479_),
    .B1(net85));
 sg13g2_nand2_1 _2246_ (.Y(_0994_),
    .A(net129),
    .B(\state[96] ));
 sg13g2_a21oi_1 _2247_ (.A1(_0803_),
    .A2(_0994_),
    .Y(_0480_),
    .B1(net85));
 sg13g2_nand2_1 _2248_ (.Y(_0995_),
    .A(net128),
    .B(\state[97] ));
 sg13g2_a21oi_1 _2249_ (.A1(_0806_),
    .A2(_0995_),
    .Y(_0481_),
    .B1(net84));
 sg13g2_nand2_1 _2250_ (.Y(_0996_),
    .A(net130),
    .B(\state[98] ));
 sg13g2_a21oi_1 _2251_ (.A1(_0809_),
    .A2(_0996_),
    .Y(_0482_),
    .B1(net86));
 sg13g2_nand2_1 _2252_ (.Y(_0997_),
    .A(net130),
    .B(\state[99] ));
 sg13g2_a21oi_1 _2253_ (.A1(_0812_),
    .A2(_0997_),
    .Y(_0483_),
    .B1(net86));
 sg13g2_nand2_1 _2254_ (.Y(_0998_),
    .A(net133),
    .B(\state[100] ));
 sg13g2_a21oi_1 _2255_ (.A1(_0815_),
    .A2(_0998_),
    .Y(_0484_),
    .B1(net89));
 sg13g2_nand2_1 _2256_ (.Y(_0999_),
    .A(net133),
    .B(\state[101] ));
 sg13g2_a21oi_1 _2257_ (.A1(_0818_),
    .A2(_0999_),
    .Y(_0485_),
    .B1(net89));
 sg13g2_nand2_1 _2258_ (.Y(_1000_),
    .A(net134),
    .B(\state[102] ));
 sg13g2_a21oi_1 _2259_ (.A1(_0821_),
    .A2(_1000_),
    .Y(_0486_),
    .B1(net90));
 sg13g2_nand2_1 _2260_ (.Y(_1001_),
    .A(net132),
    .B(\state[103] ));
 sg13g2_a21oi_1 _2261_ (.A1(_0824_),
    .A2(_1001_),
    .Y(_0487_),
    .B1(net88));
 sg13g2_nand2_1 _2262_ (.Y(_1002_),
    .A(net131),
    .B(\state[104] ));
 sg13g2_a21oi_1 _2263_ (.A1(_0827_),
    .A2(_1002_),
    .Y(_0488_),
    .B1(net87));
 sg13g2_nand2_1 _2264_ (.Y(_1003_),
    .A(net132),
    .B(\state[105] ));
 sg13g2_a21oi_1 _2265_ (.A1(_0830_),
    .A2(_1003_),
    .Y(_0489_),
    .B1(net88));
 sg13g2_nand2_1 _2266_ (.Y(_1004_),
    .A(net132),
    .B(\state[106] ));
 sg13g2_a21oi_1 _2267_ (.A1(_0833_),
    .A2(_1004_),
    .Y(_0490_),
    .B1(net88));
 sg13g2_nand2_1 _2268_ (.Y(_1005_),
    .A(net131),
    .B(\state[107] ));
 sg13g2_a21oi_1 _2269_ (.A1(_0836_),
    .A2(_1005_),
    .Y(_0491_),
    .B1(net88));
 sg13g2_nand2_1 _2270_ (.Y(_1006_),
    .A(net130),
    .B(\state[108] ));
 sg13g2_a21oi_1 _2271_ (.A1(_0839_),
    .A2(_1006_),
    .Y(_0492_),
    .B1(net86));
 sg13g2_nand2_1 _2272_ (.Y(_1007_),
    .A(net130),
    .B(\state[109] ));
 sg13g2_a21oi_1 _2273_ (.A1(_0842_),
    .A2(_1007_),
    .Y(_0493_),
    .B1(net86));
 sg13g2_nand2_1 _2274_ (.Y(_1008_),
    .A(net128),
    .B(\state[110] ));
 sg13g2_a21oi_1 _2275_ (.A1(_0845_),
    .A2(_1008_),
    .Y(_0494_),
    .B1(net84));
 sg13g2_nand2_1 _2276_ (.Y(_1009_),
    .A(net124),
    .B(\state[111] ));
 sg13g2_a21oi_1 _2277_ (.A1(_0848_),
    .A2(_1009_),
    .Y(_0495_),
    .B1(net80));
 sg13g2_nand2_1 _2278_ (.Y(_1010_),
    .A(net124),
    .B(\state[112] ));
 sg13g2_a21oi_1 _2279_ (.A1(_0851_),
    .A2(_1010_),
    .Y(_0496_),
    .B1(net80));
 sg13g2_nand2_1 _2280_ (.Y(_1011_),
    .A(net125),
    .B(\state[113] ));
 sg13g2_a21oi_1 _2281_ (.A1(_0854_),
    .A2(_1011_),
    .Y(_0497_),
    .B1(net81));
 sg13g2_nand2_1 _2282_ (.Y(_1012_),
    .A(net125),
    .B(\state[114] ));
 sg13g2_a21oi_1 _2283_ (.A1(_0857_),
    .A2(_1012_),
    .Y(_0498_),
    .B1(net81));
 sg13g2_nand2_1 _2284_ (.Y(_1013_),
    .A(net131),
    .B(\state[115] ));
 sg13g2_a21oi_1 _2285_ (.A1(_0860_),
    .A2(_1013_),
    .Y(_0499_),
    .B1(net87));
 sg13g2_nand2_1 _2286_ (.Y(_1014_),
    .A(net132),
    .B(\state[116] ));
 sg13g2_a21oi_1 _2287_ (.A1(_0863_),
    .A2(_1014_),
    .Y(_0500_),
    .B1(net88));
 sg13g2_nand2_1 _2288_ (.Y(_1015_),
    .A(net136),
    .B(\state[117] ));
 sg13g2_a21oi_1 _2289_ (.A1(_0866_),
    .A2(_1015_),
    .Y(_0501_),
    .B1(net82));
 sg13g2_nand2_1 _2290_ (.Y(_1016_),
    .A(net127),
    .B(\state[118] ));
 sg13g2_a21oi_1 _2291_ (.A1(_0869_),
    .A2(_1016_),
    .Y(_0502_),
    .B1(net91));
 sg13g2_nand2_1 _2292_ (.Y(_1017_),
    .A(net126),
    .B(\state[119] ));
 sg13g2_a21oi_1 _2293_ (.A1(_0872_),
    .A2(_1017_),
    .Y(_0503_),
    .B1(net82));
 sg13g2_nand2_1 _2294_ (.Y(_1018_),
    .A(net127),
    .B(\state[120] ));
 sg13g2_a21oi_1 _2295_ (.A1(_0875_),
    .A2(_1018_),
    .Y(_0504_),
    .B1(net83));
 sg13g2_nand2_1 _2296_ (.Y(_1019_),
    .A(net113),
    .B(\state[121] ));
 sg13g2_a21oi_1 _2297_ (.A1(_0878_),
    .A2(_1019_),
    .Y(_0505_),
    .B1(net69));
 sg13g2_nand2_1 _2298_ (.Y(_1020_),
    .A(net114),
    .B(\state[122] ));
 sg13g2_a21oi_1 _2299_ (.A1(_0881_),
    .A2(_1020_),
    .Y(_0506_),
    .B1(net70));
 sg13g2_nand2_1 _2300_ (.Y(_1021_),
    .A(net114),
    .B(\state[123] ));
 sg13g2_a21oi_1 _2301_ (.A1(_0884_),
    .A2(_1021_),
    .Y(_0507_),
    .B1(net70));
 sg13g2_nand2_1 _2302_ (.Y(_1022_),
    .A(net115),
    .B(\state[124] ));
 sg13g2_a21oi_1 _2303_ (.A1(_0887_),
    .A2(_1022_),
    .Y(_0508_),
    .B1(net69));
 sg13g2_nand2_1 _2304_ (.Y(_1023_),
    .A(net113),
    .B(\state[125] ));
 sg13g2_a21oi_1 _2305_ (.A1(_0890_),
    .A2(_1023_),
    .Y(_0509_),
    .B1(net69));
 sg13g2_nand2_1 _2306_ (.Y(_1024_),
    .A(net113),
    .B(\state[126] ));
 sg13g2_a21oi_1 _2307_ (.A1(_0893_),
    .A2(_1024_),
    .Y(_0510_),
    .B1(net69));
 sg13g2_nand2_1 _2308_ (.Y(_1025_),
    .A(\state[127] ),
    .B(net115));
 sg13g2_a21oi_1 _2309_ (.A1(_0896_),
    .A2(_1025_),
    .Y(_0511_),
    .B1(net72));
 sg13g2_dfrbpq_1 _2310_ (.RESET_B(net482),
    .D(_0256_),
    .Q(\daisychain[0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2311_ (.RESET_B(net481),
    .D(_0257_),
    .Q(\daisychain[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2312_ (.RESET_B(net479),
    .D(_0258_),
    .Q(\daisychain[2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2313_ (.RESET_B(net477),
    .D(_0259_),
    .Q(\daisychain[3] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2314_ (.RESET_B(net475),
    .D(_0260_),
    .Q(\daisychain[4] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2315_ (.RESET_B(net473),
    .D(_0261_),
    .Q(\daisychain[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2316_ (.RESET_B(net471),
    .D(_0262_),
    .Q(\daisychain[6] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2317_ (.RESET_B(net469),
    .D(_0263_),
    .Q(\daisychain[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2318_ (.RESET_B(net467),
    .D(_0264_),
    .Q(\daisychain[8] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2319_ (.RESET_B(net465),
    .D(_0265_),
    .Q(\daisychain[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2320_ (.RESET_B(net463),
    .D(_0266_),
    .Q(\daisychain[10] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2321_ (.RESET_B(net461),
    .D(_0267_),
    .Q(\daisychain[11] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2322_ (.RESET_B(net459),
    .D(_0268_),
    .Q(\daisychain[12] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2323_ (.RESET_B(net457),
    .D(_0269_),
    .Q(\daisychain[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2324_ (.RESET_B(net455),
    .D(_0270_),
    .Q(\daisychain[14] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2325_ (.RESET_B(net453),
    .D(_0271_),
    .Q(\daisychain[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2326_ (.RESET_B(net451),
    .D(_0272_),
    .Q(\daisychain[16] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2327_ (.RESET_B(net449),
    .D(_0273_),
    .Q(\daisychain[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2328_ (.RESET_B(net447),
    .D(_0274_),
    .Q(\daisychain[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2329_ (.RESET_B(net445),
    .D(_0275_),
    .Q(\daisychain[19] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2330_ (.RESET_B(net443),
    .D(_0276_),
    .Q(\daisychain[20] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2331_ (.RESET_B(net441),
    .D(_0277_),
    .Q(\daisychain[21] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2332_ (.RESET_B(net439),
    .D(_0278_),
    .Q(\daisychain[22] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2333_ (.RESET_B(net437),
    .D(_0279_),
    .Q(\daisychain[23] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2334_ (.RESET_B(net435),
    .D(_0280_),
    .Q(\daisychain[24] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2335_ (.RESET_B(net433),
    .D(_0281_),
    .Q(\daisychain[25] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2336_ (.RESET_B(net431),
    .D(_0282_),
    .Q(\daisychain[26] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2337_ (.RESET_B(net429),
    .D(_0283_),
    .Q(\daisychain[27] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2338_ (.RESET_B(net427),
    .D(_0284_),
    .Q(\daisychain[28] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2339_ (.RESET_B(net425),
    .D(_0285_),
    .Q(\daisychain[29] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2340_ (.RESET_B(net423),
    .D(_0286_),
    .Q(\daisychain[30] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2341_ (.RESET_B(net421),
    .D(_0287_),
    .Q(\daisychain[31] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2342_ (.RESET_B(net419),
    .D(_0288_),
    .Q(\daisychain[32] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2343_ (.RESET_B(net417),
    .D(_0289_),
    .Q(\daisychain[33] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2344_ (.RESET_B(net415),
    .D(_0290_),
    .Q(\daisychain[34] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2345_ (.RESET_B(net413),
    .D(_0291_),
    .Q(\daisychain[35] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2346_ (.RESET_B(net411),
    .D(_0292_),
    .Q(\daisychain[36] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2347_ (.RESET_B(net409),
    .D(_0293_),
    .Q(\daisychain[37] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2348_ (.RESET_B(net407),
    .D(_0294_),
    .Q(\daisychain[38] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2349_ (.RESET_B(net405),
    .D(_0295_),
    .Q(\daisychain[39] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2350_ (.RESET_B(net403),
    .D(_0296_),
    .Q(\daisychain[40] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2351_ (.RESET_B(net401),
    .D(_0297_),
    .Q(\daisychain[41] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2352_ (.RESET_B(net399),
    .D(_0298_),
    .Q(\daisychain[42] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2353_ (.RESET_B(net397),
    .D(_0299_),
    .Q(\daisychain[43] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2354_ (.RESET_B(net395),
    .D(_0300_),
    .Q(\daisychain[44] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2355_ (.RESET_B(net393),
    .D(_0301_),
    .Q(\daisychain[45] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2356_ (.RESET_B(net391),
    .D(_0302_),
    .Q(\daisychain[46] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2357_ (.RESET_B(net389),
    .D(_0303_),
    .Q(\daisychain[47] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2358_ (.RESET_B(net387),
    .D(_0304_),
    .Q(\daisychain[48] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2359_ (.RESET_B(net385),
    .D(_0305_),
    .Q(\daisychain[49] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2360_ (.RESET_B(net383),
    .D(_0306_),
    .Q(\daisychain[50] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2361_ (.RESET_B(net381),
    .D(_0307_),
    .Q(\daisychain[51] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2362_ (.RESET_B(net379),
    .D(_0308_),
    .Q(\daisychain[52] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2363_ (.RESET_B(net377),
    .D(_0309_),
    .Q(\daisychain[53] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2364_ (.RESET_B(net375),
    .D(_0310_),
    .Q(\daisychain[54] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2365_ (.RESET_B(net373),
    .D(_0311_),
    .Q(\daisychain[55] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2366_ (.RESET_B(net371),
    .D(_0312_),
    .Q(\daisychain[56] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2367_ (.RESET_B(net369),
    .D(_0313_),
    .Q(\daisychain[57] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2368_ (.RESET_B(net367),
    .D(_0314_),
    .Q(\daisychain[58] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2369_ (.RESET_B(net365),
    .D(_0315_),
    .Q(\daisychain[59] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2370_ (.RESET_B(net363),
    .D(_0316_),
    .Q(\daisychain[60] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2371_ (.RESET_B(net361),
    .D(_0317_),
    .Q(\daisychain[61] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2372_ (.RESET_B(net359),
    .D(_0318_),
    .Q(\daisychain[62] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2373_ (.RESET_B(net357),
    .D(_0319_),
    .Q(\daisychain[63] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2374_ (.RESET_B(net355),
    .D(_0320_),
    .Q(\daisychain[64] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2375_ (.RESET_B(net353),
    .D(_0321_),
    .Q(\daisychain[65] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2376_ (.RESET_B(net351),
    .D(_0322_),
    .Q(\daisychain[66] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2377_ (.RESET_B(net349),
    .D(_0323_),
    .Q(\daisychain[67] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2378_ (.RESET_B(net347),
    .D(_0324_),
    .Q(\daisychain[68] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2379_ (.RESET_B(net345),
    .D(_0325_),
    .Q(\daisychain[69] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2380_ (.RESET_B(net343),
    .D(_0326_),
    .Q(\daisychain[70] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2381_ (.RESET_B(net341),
    .D(_0327_),
    .Q(\daisychain[71] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2382_ (.RESET_B(net339),
    .D(_0328_),
    .Q(\daisychain[72] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2383_ (.RESET_B(net337),
    .D(_0329_),
    .Q(\daisychain[73] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2384_ (.RESET_B(net335),
    .D(_0330_),
    .Q(\daisychain[74] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2385_ (.RESET_B(net333),
    .D(_0331_),
    .Q(\daisychain[75] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2386_ (.RESET_B(net331),
    .D(_0332_),
    .Q(\daisychain[76] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2387_ (.RESET_B(net329),
    .D(_0333_),
    .Q(\daisychain[77] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2388_ (.RESET_B(net327),
    .D(_0334_),
    .Q(\daisychain[78] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2389_ (.RESET_B(net325),
    .D(_0335_),
    .Q(\daisychain[79] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2390_ (.RESET_B(net323),
    .D(_0336_),
    .Q(\daisychain[80] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2391_ (.RESET_B(net321),
    .D(_0337_),
    .Q(\daisychain[81] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2392_ (.RESET_B(net319),
    .D(_0338_),
    .Q(\daisychain[82] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2393_ (.RESET_B(net317),
    .D(_0339_),
    .Q(\daisychain[83] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2394_ (.RESET_B(net315),
    .D(_0340_),
    .Q(\daisychain[84] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2395_ (.RESET_B(net313),
    .D(_0341_),
    .Q(\daisychain[85] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2396_ (.RESET_B(net311),
    .D(_0342_),
    .Q(\daisychain[86] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2397_ (.RESET_B(net309),
    .D(_0343_),
    .Q(\daisychain[87] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2398_ (.RESET_B(net307),
    .D(_0344_),
    .Q(\daisychain[88] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2399_ (.RESET_B(net305),
    .D(_0345_),
    .Q(\daisychain[89] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2400_ (.RESET_B(net303),
    .D(_0346_),
    .Q(\daisychain[90] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2401_ (.RESET_B(net301),
    .D(_0347_),
    .Q(\daisychain[91] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2402_ (.RESET_B(net299),
    .D(_0348_),
    .Q(\daisychain[92] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2403_ (.RESET_B(net297),
    .D(_0349_),
    .Q(\daisychain[93] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2404_ (.RESET_B(net295),
    .D(_0350_),
    .Q(\daisychain[94] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2405_ (.RESET_B(net293),
    .D(_0351_),
    .Q(\daisychain[95] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2406_ (.RESET_B(net291),
    .D(_0352_),
    .Q(\daisychain[96] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2407_ (.RESET_B(net289),
    .D(_0353_),
    .Q(\daisychain[97] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2408_ (.RESET_B(net287),
    .D(_0354_),
    .Q(\daisychain[98] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2409_ (.RESET_B(net285),
    .D(_0355_),
    .Q(\daisychain[99] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2410_ (.RESET_B(net283),
    .D(_0356_),
    .Q(\daisychain[100] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2411_ (.RESET_B(net281),
    .D(_0357_),
    .Q(\daisychain[101] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2412_ (.RESET_B(net279),
    .D(_0358_),
    .Q(\daisychain[102] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2413_ (.RESET_B(net277),
    .D(_0359_),
    .Q(\daisychain[103] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2414_ (.RESET_B(net275),
    .D(_0360_),
    .Q(\daisychain[104] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2415_ (.RESET_B(net273),
    .D(_0361_),
    .Q(\daisychain[105] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2416_ (.RESET_B(net271),
    .D(_0362_),
    .Q(\daisychain[106] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2417_ (.RESET_B(net269),
    .D(_0363_),
    .Q(\daisychain[107] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2418_ (.RESET_B(net267),
    .D(_0364_),
    .Q(\daisychain[108] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2419_ (.RESET_B(net265),
    .D(_0365_),
    .Q(\daisychain[109] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2420_ (.RESET_B(net263),
    .D(_0366_),
    .Q(\daisychain[110] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2421_ (.RESET_B(net261),
    .D(_0367_),
    .Q(\daisychain[111] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2422_ (.RESET_B(net259),
    .D(_0368_),
    .Q(\daisychain[112] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2423_ (.RESET_B(net257),
    .D(_0369_),
    .Q(\daisychain[113] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2424_ (.RESET_B(net255),
    .D(_0370_),
    .Q(\daisychain[114] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2425_ (.RESET_B(net253),
    .D(_0371_),
    .Q(\daisychain[115] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2426_ (.RESET_B(net251),
    .D(_0372_),
    .Q(\daisychain[116] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2427_ (.RESET_B(net249),
    .D(_0373_),
    .Q(\daisychain[117] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2428_ (.RESET_B(net247),
    .D(_0374_),
    .Q(\daisychain[118] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2429_ (.RESET_B(net245),
    .D(_0375_),
    .Q(\daisychain[119] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2430_ (.RESET_B(net243),
    .D(_0376_),
    .Q(\daisychain[120] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2431_ (.RESET_B(net241),
    .D(_0377_),
    .Q(\daisychain[121] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2432_ (.RESET_B(net239),
    .D(_0378_),
    .Q(\daisychain[122] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2433_ (.RESET_B(net237),
    .D(_0379_),
    .Q(\daisychain[123] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2434_ (.RESET_B(net235),
    .D(_0380_),
    .Q(\daisychain[124] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2435_ (.RESET_B(net233),
    .D(_0381_),
    .Q(\daisychain[125] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2436_ (.RESET_B(net231),
    .D(_0382_),
    .Q(\daisychain[126] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2437_ (.RESET_B(net229),
    .D(_0383_),
    .Q(\daisychain[127] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2438_ (.RESET_B(net483),
    .D(_0384_),
    .Q(\state[0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2439_ (.RESET_B(net480),
    .D(_0385_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2440_ (.RESET_B(net476),
    .D(_0386_),
    .Q(\state[2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2441_ (.RESET_B(net472),
    .D(_0387_),
    .Q(\state[3] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2442_ (.RESET_B(net468),
    .D(_0388_),
    .Q(\state[4] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2443_ (.RESET_B(net464),
    .D(_0389_),
    .Q(\state[5] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2444_ (.RESET_B(net460),
    .D(_0390_),
    .Q(\state[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2445_ (.RESET_B(net456),
    .D(_0391_),
    .Q(\state[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2446_ (.RESET_B(net452),
    .D(_0392_),
    .Q(\state[8] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2447_ (.RESET_B(net448),
    .D(_0393_),
    .Q(\state[9] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2448_ (.RESET_B(net444),
    .D(_0394_),
    .Q(\state[10] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2449_ (.RESET_B(net440),
    .D(_0395_),
    .Q(\state[11] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2450_ (.RESET_B(net436),
    .D(_0396_),
    .Q(\state[12] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2451_ (.RESET_B(net432),
    .D(_0397_),
    .Q(\state[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2452_ (.RESET_B(net428),
    .D(_0398_),
    .Q(\state[14] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2453_ (.RESET_B(net424),
    .D(_0399_),
    .Q(\state[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2454_ (.RESET_B(net420),
    .D(_0400_),
    .Q(\state[16] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2455_ (.RESET_B(net416),
    .D(_0401_),
    .Q(\state[17] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2456_ (.RESET_B(net412),
    .D(_0402_),
    .Q(\state[18] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2457_ (.RESET_B(net408),
    .D(_0403_),
    .Q(\state[19] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2458_ (.RESET_B(net404),
    .D(_0404_),
    .Q(\state[20] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2459_ (.RESET_B(net400),
    .D(_0405_),
    .Q(\state[21] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2460_ (.RESET_B(net396),
    .D(_0406_),
    .Q(\state[22] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2461_ (.RESET_B(net392),
    .D(_0407_),
    .Q(\state[23] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2462_ (.RESET_B(net388),
    .D(_0408_),
    .Q(\state[24] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2463_ (.RESET_B(net384),
    .D(_0409_),
    .Q(\state[25] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2464_ (.RESET_B(net380),
    .D(_0410_),
    .Q(\state[26] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2465_ (.RESET_B(net376),
    .D(_0411_),
    .Q(\state[27] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2466_ (.RESET_B(net372),
    .D(_0412_),
    .Q(\state[28] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2467_ (.RESET_B(net368),
    .D(_0413_),
    .Q(\state[29] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2468_ (.RESET_B(net364),
    .D(_0414_),
    .Q(\state[30] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2469_ (.RESET_B(net360),
    .D(_0415_),
    .Q(\state[31] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2470_ (.RESET_B(net356),
    .D(_0416_),
    .Q(\state[32] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2471_ (.RESET_B(net352),
    .D(_0417_),
    .Q(\state[33] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2472_ (.RESET_B(net348),
    .D(_0418_),
    .Q(\state[34] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2473_ (.RESET_B(net344),
    .D(_0419_),
    .Q(\state[35] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2474_ (.RESET_B(net340),
    .D(_0420_),
    .Q(\state[36] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2475_ (.RESET_B(net336),
    .D(_0421_),
    .Q(\state[37] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2476_ (.RESET_B(net332),
    .D(_0422_),
    .Q(\state[38] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2477_ (.RESET_B(net328),
    .D(_0423_),
    .Q(\state[39] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2478_ (.RESET_B(net324),
    .D(_0424_),
    .Q(\state[40] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2479_ (.RESET_B(net320),
    .D(_0425_),
    .Q(\state[41] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2480_ (.RESET_B(net316),
    .D(_0426_),
    .Q(\state[42] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2481_ (.RESET_B(net312),
    .D(_0427_),
    .Q(\state[43] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2482_ (.RESET_B(net308),
    .D(_0428_),
    .Q(\state[44] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2483_ (.RESET_B(net304),
    .D(_0429_),
    .Q(\state[45] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2484_ (.RESET_B(net300),
    .D(_0430_),
    .Q(\state[46] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2485_ (.RESET_B(net296),
    .D(_0431_),
    .Q(\state[47] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2486_ (.RESET_B(net292),
    .D(_0432_),
    .Q(\state[48] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2487_ (.RESET_B(net288),
    .D(_0433_),
    .Q(\state[49] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2488_ (.RESET_B(net284),
    .D(_0434_),
    .Q(\state[50] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2489_ (.RESET_B(net280),
    .D(_0435_),
    .Q(\state[51] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2490_ (.RESET_B(net276),
    .D(_0436_),
    .Q(\state[52] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2491_ (.RESET_B(net272),
    .D(_0437_),
    .Q(\state[53] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2492_ (.RESET_B(net268),
    .D(_0438_),
    .Q(\state[54] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2493_ (.RESET_B(net264),
    .D(_0439_),
    .Q(\state[55] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2494_ (.RESET_B(net260),
    .D(_0440_),
    .Q(\state[56] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2495_ (.RESET_B(net256),
    .D(_0441_),
    .Q(\state[57] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2496_ (.RESET_B(net252),
    .D(_0442_),
    .Q(\state[58] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2497_ (.RESET_B(net248),
    .D(_0443_),
    .Q(\state[59] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2498_ (.RESET_B(net244),
    .D(_0444_),
    .Q(\state[60] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2499_ (.RESET_B(net240),
    .D(_0445_),
    .Q(\state[61] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2500_ (.RESET_B(net236),
    .D(_0446_),
    .Q(\state[62] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2501_ (.RESET_B(net232),
    .D(_0447_),
    .Q(\state[63] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2502_ (.RESET_B(net),
    .D(_0448_),
    .Q(\state[64] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2503_ (.RESET_B(net478),
    .D(_0449_),
    .Q(\state[65] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2504_ (.RESET_B(net470),
    .D(_0450_),
    .Q(\state[66] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2505_ (.RESET_B(net462),
    .D(_0451_),
    .Q(\state[67] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2506_ (.RESET_B(net454),
    .D(_0452_),
    .Q(\state[68] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2507_ (.RESET_B(net446),
    .D(_0453_),
    .Q(\state[69] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2508_ (.RESET_B(net438),
    .D(_0454_),
    .Q(\state[70] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2509_ (.RESET_B(net430),
    .D(_0455_),
    .Q(\state[71] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2510_ (.RESET_B(net422),
    .D(_0456_),
    .Q(\state[72] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2511_ (.RESET_B(net414),
    .D(_0457_),
    .Q(\state[73] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2512_ (.RESET_B(net406),
    .D(_0458_),
    .Q(\state[74] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2513_ (.RESET_B(net398),
    .D(_0459_),
    .Q(\state[75] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2514_ (.RESET_B(net390),
    .D(_0460_),
    .Q(\state[76] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2515_ (.RESET_B(net382),
    .D(_0461_),
    .Q(\state[77] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2516_ (.RESET_B(net374),
    .D(_0462_),
    .Q(\state[78] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2517_ (.RESET_B(net366),
    .D(_0463_),
    .Q(\state[79] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2518_ (.RESET_B(net358),
    .D(_0464_),
    .Q(\state[80] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2519_ (.RESET_B(net350),
    .D(_0465_),
    .Q(\state[81] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2520_ (.RESET_B(net342),
    .D(_0466_),
    .Q(\state[82] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2521_ (.RESET_B(net334),
    .D(_0467_),
    .Q(\state[83] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2522_ (.RESET_B(net326),
    .D(_0468_),
    .Q(\state[84] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2523_ (.RESET_B(net318),
    .D(_0469_),
    .Q(\state[85] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2524_ (.RESET_B(net310),
    .D(_0470_),
    .Q(\state[86] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2525_ (.RESET_B(net302),
    .D(_0471_),
    .Q(\state[87] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2526_ (.RESET_B(net294),
    .D(_0472_),
    .Q(\state[88] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2527_ (.RESET_B(net286),
    .D(_0473_),
    .Q(\state[89] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2528_ (.RESET_B(net278),
    .D(_0474_),
    .Q(\state[90] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2529_ (.RESET_B(net270),
    .D(_0475_),
    .Q(\state[91] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2530_ (.RESET_B(net262),
    .D(_0476_),
    .Q(\state[92] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2531_ (.RESET_B(net254),
    .D(_0477_),
    .Q(\state[93] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2532_ (.RESET_B(net246),
    .D(_0478_),
    .Q(\state[94] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2533_ (.RESET_B(net238),
    .D(_0479_),
    .Q(\state[95] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2534_ (.RESET_B(net230),
    .D(_0480_),
    .Q(\state[96] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2535_ (.RESET_B(net474),
    .D(_0481_),
    .Q(\state[97] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2536_ (.RESET_B(net458),
    .D(_0482_),
    .Q(\state[98] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2537_ (.RESET_B(net442),
    .D(_0483_),
    .Q(\state[99] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2538_ (.RESET_B(net426),
    .D(_0484_),
    .Q(\state[100] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2539_ (.RESET_B(net410),
    .D(_0485_),
    .Q(\state[101] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2540_ (.RESET_B(net394),
    .D(_0486_),
    .Q(\state[102] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2541_ (.RESET_B(net378),
    .D(_0487_),
    .Q(\state[103] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2542_ (.RESET_B(net362),
    .D(_0488_),
    .Q(\state[104] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2543_ (.RESET_B(net346),
    .D(_0489_),
    .Q(\state[105] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2544_ (.RESET_B(net330),
    .D(_0490_),
    .Q(\state[106] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2545_ (.RESET_B(net314),
    .D(_0491_),
    .Q(\state[107] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2546_ (.RESET_B(net298),
    .D(_0492_),
    .Q(\state[108] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2547_ (.RESET_B(net282),
    .D(_0493_),
    .Q(\state[109] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2548_ (.RESET_B(net266),
    .D(_0494_),
    .Q(\state[110] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2549_ (.RESET_B(net250),
    .D(_0495_),
    .Q(\state[111] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2550_ (.RESET_B(net234),
    .D(_0496_),
    .Q(\state[112] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2551_ (.RESET_B(net466),
    .D(_0497_),
    .Q(\state[113] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2552_ (.RESET_B(net434),
    .D(_0498_),
    .Q(\state[114] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2553_ (.RESET_B(net402),
    .D(_0499_),
    .Q(\state[115] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2554_ (.RESET_B(net370),
    .D(_0500_),
    .Q(\state[116] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2555_ (.RESET_B(net338),
    .D(_0501_),
    .Q(\state[117] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2556_ (.RESET_B(net306),
    .D(_0502_),
    .Q(\state[118] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2557_ (.RESET_B(net274),
    .D(_0503_),
    .Q(\state[119] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2558_ (.RESET_B(net242),
    .D(_0504_),
    .Q(\state[120] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2559_ (.RESET_B(net450),
    .D(_0505_),
    .Q(\state[121] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2560_ (.RESET_B(net386),
    .D(_0506_),
    .Q(\state[122] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2561_ (.RESET_B(net322),
    .D(_0507_),
    .Q(\state[123] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2562_ (.RESET_B(net258),
    .D(_0508_),
    .Q(\state[124] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2563_ (.RESET_B(net418),
    .D(_0509_),
    .Q(\state[125] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2564_ (.RESET_B(net290),
    .D(_0510_),
    .Q(\state[126] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2565_ (.RESET_B(net354),
    .D(_0511_),
    .Q(\state[127] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_tiehi _2437__230 (.L_HI(net229));
 sg13g2_tiehi _2534__231 (.L_HI(net230));
 sg13g2_tiehi _2436__232 (.L_HI(net231));
 sg13g2_tiehi _2501__233 (.L_HI(net232));
 sg13g2_tiehi _2435__234 (.L_HI(net233));
 sg13g2_tiehi _2550__235 (.L_HI(net234));
 sg13g2_tiehi _2434__236 (.L_HI(net235));
 sg13g2_tiehi _2500__237 (.L_HI(net236));
 sg13g2_tiehi _2433__238 (.L_HI(net237));
 sg13g2_tiehi _2533__239 (.L_HI(net238));
 sg13g2_tiehi _2432__240 (.L_HI(net239));
 sg13g2_tiehi _2499__241 (.L_HI(net240));
 sg13g2_tiehi _2431__242 (.L_HI(net241));
 sg13g2_tiehi _2558__243 (.L_HI(net242));
 sg13g2_tiehi _2430__244 (.L_HI(net243));
 sg13g2_tiehi _2498__245 (.L_HI(net244));
 sg13g2_tiehi _2429__246 (.L_HI(net245));
 sg13g2_tiehi _2532__247 (.L_HI(net246));
 sg13g2_tiehi _2428__248 (.L_HI(net247));
 sg13g2_tiehi _2497__249 (.L_HI(net248));
 sg13g2_tiehi _2427__250 (.L_HI(net249));
 sg13g2_tiehi _2549__251 (.L_HI(net250));
 sg13g2_tiehi _2426__252 (.L_HI(net251));
 sg13g2_tiehi _2496__253 (.L_HI(net252));
 sg13g2_tiehi _2425__254 (.L_HI(net253));
 sg13g2_tiehi _2531__255 (.L_HI(net254));
 sg13g2_tiehi _2424__256 (.L_HI(net255));
 sg13g2_tiehi _2495__257 (.L_HI(net256));
 sg13g2_tiehi _2423__258 (.L_HI(net257));
 sg13g2_tiehi _2562__259 (.L_HI(net258));
 sg13g2_tiehi _2422__260 (.L_HI(net259));
 sg13g2_tiehi _2494__261 (.L_HI(net260));
 sg13g2_tiehi _2421__262 (.L_HI(net261));
 sg13g2_tiehi _2530__263 (.L_HI(net262));
 sg13g2_tiehi _2420__264 (.L_HI(net263));
 sg13g2_tiehi _2493__265 (.L_HI(net264));
 sg13g2_tiehi _2419__266 (.L_HI(net265));
 sg13g2_tiehi _2548__267 (.L_HI(net266));
 sg13g2_tiehi _2418__268 (.L_HI(net267));
 sg13g2_tiehi _2492__269 (.L_HI(net268));
 sg13g2_tiehi _2417__270 (.L_HI(net269));
 sg13g2_tiehi _2529__271 (.L_HI(net270));
 sg13g2_tiehi _2416__272 (.L_HI(net271));
 sg13g2_tiehi _2491__273 (.L_HI(net272));
 sg13g2_tiehi _2415__274 (.L_HI(net273));
 sg13g2_tiehi _2557__275 (.L_HI(net274));
 sg13g2_tiehi _2414__276 (.L_HI(net275));
 sg13g2_tiehi _2490__277 (.L_HI(net276));
 sg13g2_tiehi _2413__278 (.L_HI(net277));
 sg13g2_tiehi _2528__279 (.L_HI(net278));
 sg13g2_tiehi _2412__280 (.L_HI(net279));
 sg13g2_tiehi _2489__281 (.L_HI(net280));
 sg13g2_tiehi _2411__282 (.L_HI(net281));
 sg13g2_tiehi _2547__283 (.L_HI(net282));
 sg13g2_tiehi _2410__284 (.L_HI(net283));
 sg13g2_tiehi _2488__285 (.L_HI(net284));
 sg13g2_tiehi _2409__286 (.L_HI(net285));
 sg13g2_tiehi _2527__287 (.L_HI(net286));
 sg13g2_tiehi _2408__288 (.L_HI(net287));
 sg13g2_tiehi _2487__289 (.L_HI(net288));
 sg13g2_tiehi _2407__290 (.L_HI(net289));
 sg13g2_tiehi _2564__291 (.L_HI(net290));
 sg13g2_tiehi _2406__292 (.L_HI(net291));
 sg13g2_tiehi _2486__293 (.L_HI(net292));
 sg13g2_tiehi _2405__294 (.L_HI(net293));
 sg13g2_tiehi _2526__295 (.L_HI(net294));
 sg13g2_tiehi _2404__296 (.L_HI(net295));
 sg13g2_tiehi _2485__297 (.L_HI(net296));
 sg13g2_tiehi _2403__298 (.L_HI(net297));
 sg13g2_tiehi _2546__299 (.L_HI(net298));
 sg13g2_tiehi _2402__300 (.L_HI(net299));
 sg13g2_tiehi _2484__301 (.L_HI(net300));
 sg13g2_tiehi _2401__302 (.L_HI(net301));
 sg13g2_tiehi _2525__303 (.L_HI(net302));
 sg13g2_tiehi _2400__304 (.L_HI(net303));
 sg13g2_tiehi _2483__305 (.L_HI(net304));
 sg13g2_tiehi _2399__306 (.L_HI(net305));
 sg13g2_tiehi _2556__307 (.L_HI(net306));
 sg13g2_tiehi _2398__308 (.L_HI(net307));
 sg13g2_tiehi _2482__309 (.L_HI(net308));
 sg13g2_tiehi _2397__310 (.L_HI(net309));
 sg13g2_tiehi _2524__311 (.L_HI(net310));
 sg13g2_tiehi _2396__312 (.L_HI(net311));
 sg13g2_tiehi _2481__313 (.L_HI(net312));
 sg13g2_tiehi _2395__314 (.L_HI(net313));
 sg13g2_tiehi _2545__315 (.L_HI(net314));
 sg13g2_tiehi _2394__316 (.L_HI(net315));
 sg13g2_tiehi _2480__317 (.L_HI(net316));
 sg13g2_tiehi _2393__318 (.L_HI(net317));
 sg13g2_tiehi _2523__319 (.L_HI(net318));
 sg13g2_tiehi _2392__320 (.L_HI(net319));
 sg13g2_tiehi _2479__321 (.L_HI(net320));
 sg13g2_tiehi _2391__322 (.L_HI(net321));
 sg13g2_tiehi _2561__323 (.L_HI(net322));
 sg13g2_tiehi _2390__324 (.L_HI(net323));
 sg13g2_tiehi _2478__325 (.L_HI(net324));
 sg13g2_tiehi _2389__326 (.L_HI(net325));
 sg13g2_tiehi _2522__327 (.L_HI(net326));
 sg13g2_tiehi _2388__328 (.L_HI(net327));
 sg13g2_tiehi _2477__329 (.L_HI(net328));
 sg13g2_tiehi _2387__330 (.L_HI(net329));
 sg13g2_tiehi _2544__331 (.L_HI(net330));
 sg13g2_tiehi _2386__332 (.L_HI(net331));
 sg13g2_tiehi _2476__333 (.L_HI(net332));
 sg13g2_tiehi _2385__334 (.L_HI(net333));
 sg13g2_tiehi _2521__335 (.L_HI(net334));
 sg13g2_tiehi _2384__336 (.L_HI(net335));
 sg13g2_tiehi _2475__337 (.L_HI(net336));
 sg13g2_tiehi _2383__338 (.L_HI(net337));
 sg13g2_tiehi _2555__339 (.L_HI(net338));
 sg13g2_tiehi _2382__340 (.L_HI(net339));
 sg13g2_tiehi _2474__341 (.L_HI(net340));
 sg13g2_tiehi _2381__342 (.L_HI(net341));
 sg13g2_tiehi _2520__343 (.L_HI(net342));
 sg13g2_tiehi _2380__344 (.L_HI(net343));
 sg13g2_tiehi _2473__345 (.L_HI(net344));
 sg13g2_tiehi _2379__346 (.L_HI(net345));
 sg13g2_tiehi _2543__347 (.L_HI(net346));
 sg13g2_tiehi _2378__348 (.L_HI(net347));
 sg13g2_tiehi _2472__349 (.L_HI(net348));
 sg13g2_tiehi _2377__350 (.L_HI(net349));
 sg13g2_tiehi _2519__351 (.L_HI(net350));
 sg13g2_tiehi _2376__352 (.L_HI(net351));
 sg13g2_tiehi _2471__353 (.L_HI(net352));
 sg13g2_tiehi _2375__354 (.L_HI(net353));
 sg13g2_tiehi _2565__355 (.L_HI(net354));
 sg13g2_tiehi _2374__356 (.L_HI(net355));
 sg13g2_tiehi _2470__357 (.L_HI(net356));
 sg13g2_tiehi _2373__358 (.L_HI(net357));
 sg13g2_tiehi _2518__359 (.L_HI(net358));
 sg13g2_tiehi _2372__360 (.L_HI(net359));
 sg13g2_tiehi _2469__361 (.L_HI(net360));
 sg13g2_tiehi _2371__362 (.L_HI(net361));
 sg13g2_tiehi _2542__363 (.L_HI(net362));
 sg13g2_tiehi _2370__364 (.L_HI(net363));
 sg13g2_tiehi _2468__365 (.L_HI(net364));
 sg13g2_tiehi _2369__366 (.L_HI(net365));
 sg13g2_tiehi _2517__367 (.L_HI(net366));
 sg13g2_tiehi _2368__368 (.L_HI(net367));
 sg13g2_tiehi _2467__369 (.L_HI(net368));
 sg13g2_tiehi _2367__370 (.L_HI(net369));
 sg13g2_tiehi _2554__371 (.L_HI(net370));
 sg13g2_tiehi _2366__372 (.L_HI(net371));
 sg13g2_tiehi _2466__373 (.L_HI(net372));
 sg13g2_tiehi _2365__374 (.L_HI(net373));
 sg13g2_tiehi _2516__375 (.L_HI(net374));
 sg13g2_tiehi _2364__376 (.L_HI(net375));
 sg13g2_tiehi _2465__377 (.L_HI(net376));
 sg13g2_tiehi _2363__378 (.L_HI(net377));
 sg13g2_tiehi _2541__379 (.L_HI(net378));
 sg13g2_tiehi _2362__380 (.L_HI(net379));
 sg13g2_tiehi _2464__381 (.L_HI(net380));
 sg13g2_tiehi _2361__382 (.L_HI(net381));
 sg13g2_tiehi _2515__383 (.L_HI(net382));
 sg13g2_tiehi _2360__384 (.L_HI(net383));
 sg13g2_tiehi _2463__385 (.L_HI(net384));
 sg13g2_tiehi _2359__386 (.L_HI(net385));
 sg13g2_tiehi _2560__387 (.L_HI(net386));
 sg13g2_tiehi _2358__388 (.L_HI(net387));
 sg13g2_tiehi _2462__389 (.L_HI(net388));
 sg13g2_tiehi _2357__390 (.L_HI(net389));
 sg13g2_tiehi _2514__391 (.L_HI(net390));
 sg13g2_tiehi _2356__392 (.L_HI(net391));
 sg13g2_tiehi _2461__393 (.L_HI(net392));
 sg13g2_tiehi _2355__394 (.L_HI(net393));
 sg13g2_tiehi _2540__395 (.L_HI(net394));
 sg13g2_tiehi _2354__396 (.L_HI(net395));
 sg13g2_tiehi _2460__397 (.L_HI(net396));
 sg13g2_tiehi _2353__398 (.L_HI(net397));
 sg13g2_tiehi _2513__399 (.L_HI(net398));
 sg13g2_tiehi _2352__400 (.L_HI(net399));
 sg13g2_tiehi _2459__401 (.L_HI(net400));
 sg13g2_tiehi _2351__402 (.L_HI(net401));
 sg13g2_tiehi _2553__403 (.L_HI(net402));
 sg13g2_tiehi _2350__404 (.L_HI(net403));
 sg13g2_tiehi _2458__405 (.L_HI(net404));
 sg13g2_tiehi _2349__406 (.L_HI(net405));
 sg13g2_tiehi _2512__407 (.L_HI(net406));
 sg13g2_tiehi _2348__408 (.L_HI(net407));
 sg13g2_tiehi _2457__409 (.L_HI(net408));
 sg13g2_tiehi _2347__410 (.L_HI(net409));
 sg13g2_tiehi _2539__411 (.L_HI(net410));
 sg13g2_tiehi _2346__412 (.L_HI(net411));
 sg13g2_tiehi _2456__413 (.L_HI(net412));
 sg13g2_tiehi _2345__414 (.L_HI(net413));
 sg13g2_tiehi _2511__415 (.L_HI(net414));
 sg13g2_tiehi _2344__416 (.L_HI(net415));
 sg13g2_tiehi _2455__417 (.L_HI(net416));
 sg13g2_tiehi _2343__418 (.L_HI(net417));
 sg13g2_tiehi _2563__419 (.L_HI(net418));
 sg13g2_tiehi _2342__420 (.L_HI(net419));
 sg13g2_tiehi _2454__421 (.L_HI(net420));
 sg13g2_tiehi _2341__422 (.L_HI(net421));
 sg13g2_tiehi _2510__423 (.L_HI(net422));
 sg13g2_tiehi _2340__424 (.L_HI(net423));
 sg13g2_tiehi _2453__425 (.L_HI(net424));
 sg13g2_tiehi _2339__426 (.L_HI(net425));
 sg13g2_tiehi _2538__427 (.L_HI(net426));
 sg13g2_tiehi _2338__428 (.L_HI(net427));
 sg13g2_tiehi _2452__429 (.L_HI(net428));
 sg13g2_tiehi _2337__430 (.L_HI(net429));
 sg13g2_tiehi _2509__431 (.L_HI(net430));
 sg13g2_tiehi _2336__432 (.L_HI(net431));
 sg13g2_tiehi _2451__433 (.L_HI(net432));
 sg13g2_tiehi _2335__434 (.L_HI(net433));
 sg13g2_tiehi _2552__435 (.L_HI(net434));
 sg13g2_tiehi _2334__436 (.L_HI(net435));
 sg13g2_tiehi _2450__437 (.L_HI(net436));
 sg13g2_tiehi _2333__438 (.L_HI(net437));
 sg13g2_tiehi _2508__439 (.L_HI(net438));
 sg13g2_tiehi _2332__440 (.L_HI(net439));
 sg13g2_tiehi _2449__441 (.L_HI(net440));
 sg13g2_tiehi _2331__442 (.L_HI(net441));
 sg13g2_tiehi _2537__443 (.L_HI(net442));
 sg13g2_tiehi _2330__444 (.L_HI(net443));
 sg13g2_tiehi _2448__445 (.L_HI(net444));
 sg13g2_tiehi _2329__446 (.L_HI(net445));
 sg13g2_tiehi _2507__447 (.L_HI(net446));
 sg13g2_tiehi _2328__448 (.L_HI(net447));
 sg13g2_tiehi _2447__449 (.L_HI(net448));
 sg13g2_tiehi _2327__450 (.L_HI(net449));
 sg13g2_tiehi _2559__451 (.L_HI(net450));
 sg13g2_tiehi _2326__452 (.L_HI(net451));
 sg13g2_tiehi _2446__453 (.L_HI(net452));
 sg13g2_tiehi _2325__454 (.L_HI(net453));
 sg13g2_tiehi _2506__455 (.L_HI(net454));
 sg13g2_tiehi _2324__456 (.L_HI(net455));
 sg13g2_tiehi _2445__457 (.L_HI(net456));
 sg13g2_tiehi _2323__458 (.L_HI(net457));
 sg13g2_tiehi _2536__459 (.L_HI(net458));
 sg13g2_tiehi _2322__460 (.L_HI(net459));
 sg13g2_tiehi _2444__461 (.L_HI(net460));
 sg13g2_tiehi _2321__462 (.L_HI(net461));
 sg13g2_tiehi _2505__463 (.L_HI(net462));
 sg13g2_tiehi _2320__464 (.L_HI(net463));
 sg13g2_tiehi _2443__465 (.L_HI(net464));
 sg13g2_tiehi _2319__466 (.L_HI(net465));
 sg13g2_tiehi _2551__467 (.L_HI(net466));
 sg13g2_tiehi _2318__468 (.L_HI(net467));
 sg13g2_tiehi _2442__469 (.L_HI(net468));
 sg13g2_tiehi _2317__470 (.L_HI(net469));
 sg13g2_tiehi _2504__471 (.L_HI(net470));
 sg13g2_tiehi _2316__472 (.L_HI(net471));
 sg13g2_tiehi _2441__473 (.L_HI(net472));
 sg13g2_tiehi _2315__474 (.L_HI(net473));
 sg13g2_tiehi _2535__475 (.L_HI(net474));
 sg13g2_tiehi _2314__476 (.L_HI(net475));
 sg13g2_tiehi _2440__477 (.L_HI(net476));
 sg13g2_tiehi _2313__478 (.L_HI(net477));
 sg13g2_tiehi _2503__479 (.L_HI(net478));
 sg13g2_tiehi _2312__480 (.L_HI(net479));
 sg13g2_tiehi _2439__481 (.L_HI(net480));
 sg13g2_tiehi _2311__482 (.L_HI(net481));
 sg13g2_tiehi _2310__483 (.L_HI(net482));
 sg13g2_tiehi _2438__484 (.L_HI(net483));
 sg13g2_tiehi heichips25_pudding (.L_HI(net484));
 sg13g2_tiehi heichips25_pudding_485 (.L_HI(net485));
 sg13g2_tiehi heichips25_pudding_486 (.L_HI(net486));
 sg13g2_tiehi heichips25_pudding_487 (.L_HI(net487));
 sg13g2_tiehi heichips25_pudding_488 (.L_HI(net488));
 sg13g2_tiehi heichips25_pudding_489 (.L_HI(net489));
 sg13g2_tiehi heichips25_pudding_490 (.L_HI(net490));
 sg13g2_tiehi heichips25_pudding_491 (.L_HI(net491));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _2830_ (.A(\state[120] ),
    .X(net8));
 sg13g2_buf_1 _2831_ (.A(\state[121] ),
    .X(net9));
 sg13g2_buf_1 _2832_ (.A(\state[122] ),
    .X(net10));
 sg13g2_buf_1 _2833_ (.A(\state[123] ),
    .X(net11));
 sg13g2_buf_1 _2834_ (.A(\state[124] ),
    .X(net12));
 sg13g2_buf_1 _2835_ (.A(\state[125] ),
    .X(net13));
 sg13g2_buf_1 _2836_ (.A(\state[126] ),
    .X(net14));
 sg13g2_buf_1 _2837_ (.A(\state[127] ),
    .X(net15));
 sg13g2_buf_1 _2838_ (.A(\daisychain[120] ),
    .X(net16));
 sg13g2_buf_1 _2839_ (.A(\daisychain[121] ),
    .X(net17));
 sg13g2_buf_1 _2840_ (.A(\daisychain[122] ),
    .X(net18));
 sg13g2_buf_1 _2841_ (.A(\daisychain[123] ),
    .X(net19));
 sg13g2_buf_1 _2842_ (.A(\daisychain[124] ),
    .X(net20));
 sg13g2_buf_1 _2843_ (.A(\daisychain[125] ),
    .X(net21));
 sg13g2_buf_1 _2844_ (.A(\daisychain[126] ),
    .X(net22));
 sg13g2_buf_1 _2845_ (.A(\daisychain[127] ),
    .X(net23));
 dac128module dacH (.EN({\digitalenH.g[3].u.OUTP ,
    \digitalenH.g[2].u.OUTP ,
    \digitalenH.g[1].u.OUTP ,
    \digitalenH.g[0].u.OUTP }),
    .ENB({\digitalenH.g[3].u.OUTN ,
    \digitalenH.g[2].u.OUTN ,
    \digitalenH.g[1].u.OUTN ,
    \digitalenH.g[0].u.OUTN }),
    .ON({\daisychain[127] ,
    \daisychain[126] ,
    \daisychain[125] ,
    \daisychain[124] ,
    \daisychain[123] ,
    \daisychain[122] ,
    \daisychain[121] ,
    \daisychain[120] ,
    \daisychain[119] ,
    \daisychain[118] ,
    \daisychain[117] ,
    \daisychain[116] ,
    \daisychain[115] ,
    \daisychain[114] ,
    \daisychain[113] ,
    \daisychain[112] ,
    \daisychain[111] ,
    \daisychain[110] ,
    \daisychain[109] ,
    \daisychain[108] ,
    \daisychain[107] ,
    \daisychain[106] ,
    \daisychain[105] ,
    \daisychain[104] ,
    \daisychain[103] ,
    \daisychain[102] ,
    \daisychain[101] ,
    \daisychain[100] ,
    \daisychain[99] ,
    \daisychain[98] ,
    \daisychain[97] ,
    \daisychain[96] ,
    \daisychain[95] ,
    \daisychain[94] ,
    \daisychain[93] ,
    \daisychain[92] ,
    \daisychain[91] ,
    \daisychain[90] ,
    \daisychain[89] ,
    \daisychain[88] ,
    \daisychain[87] ,
    \daisychain[86] ,
    \daisychain[85] ,
    \daisychain[84] ,
    \daisychain[83] ,
    \daisychain[82] ,
    \daisychain[81] ,
    \daisychain[80] ,
    \daisychain[79] ,
    \daisychain[78] ,
    \daisychain[77] ,
    \daisychain[76] ,
    \daisychain[75] ,
    \daisychain[74] ,
    \daisychain[73] ,
    \daisychain[72] ,
    \daisychain[71] ,
    \daisychain[70] ,
    \daisychain[69] ,
    \daisychain[68] ,
    \daisychain[67] ,
    \daisychain[66] ,
    \daisychain[65] ,
    \daisychain[64] ,
    \daisychain[63] ,
    \daisychain[62] ,
    \daisychain[61] ,
    \daisychain[60] ,
    \daisychain[59] ,
    \daisychain[58] ,
    \daisychain[57] ,
    \daisychain[56] ,
    \daisychain[55] ,
    \daisychain[54] ,
    \daisychain[53] ,
    \daisychain[52] ,
    \daisychain[51] ,
    \daisychain[50] ,
    \daisychain[49] ,
    \daisychain[48] ,
    \daisychain[47] ,
    \daisychain[46] ,
    \daisychain[45] ,
    \daisychain[44] ,
    \daisychain[43] ,
    \daisychain[42] ,
    \daisychain[41] ,
    \daisychain[40] ,
    \daisychain[39] ,
    \daisychain[38] ,
    \daisychain[37] ,
    \daisychain[36] ,
    \daisychain[35] ,
    \daisychain[34] ,
    \daisychain[33] ,
    \daisychain[32] ,
    \daisychain[31] ,
    \daisychain[30] ,
    \daisychain[29] ,
    \daisychain[28] ,
    \daisychain[27] ,
    \daisychain[26] ,
    \daisychain[25] ,
    \daisychain[24] ,
    \daisychain[23] ,
    \daisychain[22] ,
    \daisychain[21] ,
    \daisychain[20] ,
    \daisychain[19] ,
    \daisychain[18] ,
    \daisychain[17] ,
    \daisychain[16] ,
    \daisychain[15] ,
    \daisychain[14] ,
    \daisychain[13] ,
    \daisychain[12] ,
    \daisychain[11] ,
    \daisychain[10] ,
    \daisychain[9] ,
    \daisychain[8] ,
    \daisychain[7] ,
    \daisychain[6] ,
    \daisychain[5] ,
    \daisychain[4] ,
    \daisychain[3] ,
    \daisychain[2] ,
    \daisychain[1] ,
    \daisychain[0] }),
    .ONB({_0158_,
    _0157_,
    _0156_,
    _0155_,
    _0154_,
    _0153_,
    _0152_,
    _0151_,
    _0149_,
    _0148_,
    _0147_,
    _0146_,
    _0145_,
    _0144_,
    _0143_,
    _0142_,
    _0141_,
    _0140_,
    _0138_,
    _0137_,
    _0136_,
    _0135_,
    _0134_,
    _0133_,
    _0132_,
    _0131_,
    _0130_,
    _0129_,
    _0254_,
    _0253_,
    _0252_,
    _0251_,
    _0250_,
    _0249_,
    _0248_,
    _0247_,
    _0246_,
    _0245_,
    _0243_,
    _0242_,
    _0241_,
    _0240_,
    _0239_,
    _0238_,
    _0237_,
    _0236_,
    _0235_,
    _0234_,
    _0232_,
    _0231_,
    _0230_,
    _0229_,
    _0228_,
    _0227_,
    _0226_,
    _0225_,
    _0224_,
    _0223_,
    _0221_,
    _0220_,
    _0219_,
    _0218_,
    _0217_,
    _0216_,
    _0215_,
    _0214_,
    _0213_,
    _0212_,
    _0210_,
    _0209_,
    _0208_,
    _0207_,
    _0206_,
    _0205_,
    _0204_,
    _0203_,
    _0202_,
    _0201_,
    _0199_,
    _0198_,
    _0197_,
    _0196_,
    _0195_,
    _0194_,
    _0193_,
    _0192_,
    _0191_,
    _0190_,
    _0188_,
    _0187_,
    _0186_,
    _0185_,
    _0184_,
    _0183_,
    _0182_,
    _0181_,
    _0180_,
    _0179_,
    _0177_,
    _0176_,
    _0175_,
    _0174_,
    _0173_,
    _0172_,
    _0171_,
    _0170_,
    _0169_,
    _0168_,
    _0166_,
    _0165_,
    _0164_,
    _0163_,
    _0162_,
    _0161_,
    _0160_,
    _0159_,
    _0150_,
    _0139_,
    _0255_,
    _0244_,
    _0233_,
    _0222_,
    _0211_,
    _0200_,
    _0189_,
    _0178_,
    _0167_,
    _0128_}));
 dac128module dacL (.EN({\digitalenL.g[3].u.OUTP ,
    \digitalenL.g[2].u.OUTP ,
    \digitalenL.g[1].u.OUTP ,
    \digitalenL.g[0].u.OUTP }),
    .ENB({\digitalenL.g[3].u.OUTN ,
    \digitalenL.g[2].u.OUTN ,
    \digitalenL.g[1].u.OUTN ,
    \digitalenL.g[0].u.OUTN }),
    .ON({\state[127] ,
    \state[126] ,
    \state[125] ,
    \state[124] ,
    \state[123] ,
    \state[122] ,
    \state[121] ,
    \state[120] ,
    \state[119] ,
    \state[118] ,
    \state[117] ,
    \state[116] ,
    \state[115] ,
    \state[114] ,
    \state[113] ,
    \state[112] ,
    \state[111] ,
    \state[110] ,
    \state[109] ,
    \state[108] ,
    \state[107] ,
    \state[106] ,
    \state[105] ,
    \state[104] ,
    \state[103] ,
    \state[102] ,
    \state[101] ,
    \state[100] ,
    \state[99] ,
    \state[98] ,
    \state[97] ,
    \state[96] ,
    \state[95] ,
    \state[94] ,
    \state[93] ,
    \state[92] ,
    \state[91] ,
    \state[90] ,
    \state[89] ,
    \state[88] ,
    \state[87] ,
    \state[86] ,
    \state[85] ,
    \state[84] ,
    \state[83] ,
    \state[82] ,
    \state[81] ,
    \state[80] ,
    \state[79] ,
    \state[78] ,
    \state[77] ,
    \state[76] ,
    \state[75] ,
    \state[74] ,
    \state[73] ,
    \state[72] ,
    \state[71] ,
    \state[70] ,
    \state[69] ,
    \state[68] ,
    \state[67] ,
    \state[66] ,
    \state[65] ,
    \state[64] ,
    \state[63] ,
    \state[62] ,
    \state[61] ,
    \state[60] ,
    \state[59] ,
    \state[58] ,
    \state[57] ,
    \state[56] ,
    \state[55] ,
    \state[54] ,
    \state[53] ,
    \state[52] ,
    \state[51] ,
    \state[50] ,
    \state[49] ,
    \state[48] ,
    \state[47] ,
    \state[46] ,
    \state[45] ,
    \state[44] ,
    \state[43] ,
    \state[42] ,
    \state[41] ,
    \state[40] ,
    \state[39] ,
    \state[38] ,
    \state[37] ,
    \state[36] ,
    \state[35] ,
    \state[34] ,
    \state[33] ,
    \state[32] ,
    \state[31] ,
    \state[30] ,
    \state[29] ,
    \state[28] ,
    \state[27] ,
    \state[26] ,
    \state[25] ,
    \state[24] ,
    \state[23] ,
    \state[22] ,
    \state[21] ,
    \state[20] ,
    \state[19] ,
    \state[18] ,
    \state[17] ,
    \state[16] ,
    \state[15] ,
    \state[14] ,
    \state[13] ,
    \state[12] ,
    \state[11] ,
    \state[10] ,
    \state[9] ,
    \state[8] ,
    \state[7] ,
    \state[6] ,
    \state[5] ,
    \state[4] ,
    \state[3] ,
    \state[2] ,
    \state[1] ,
    \state[0] }),
    .ONB({_0030_,
    _0029_,
    _0028_,
    _0027_,
    _0026_,
    _0025_,
    _0024_,
    _0023_,
    _0021_,
    _0020_,
    _0019_,
    _0018_,
    _0017_,
    _0016_,
    _0015_,
    _0014_,
    _0013_,
    _0012_,
    _0010_,
    _0009_,
    _0008_,
    _0007_,
    _0006_,
    _0005_,
    _0004_,
    _0003_,
    _0002_,
    _0001_,
    _0126_,
    _0125_,
    _0124_,
    _0123_,
    _0122_,
    _0121_,
    _0120_,
    _0119_,
    _0118_,
    _0117_,
    _0115_,
    _0114_,
    _0113_,
    _0112_,
    _0111_,
    _0110_,
    _0109_,
    _0108_,
    _0107_,
    _0106_,
    _0104_,
    _0103_,
    _0102_,
    _0101_,
    _0100_,
    _0099_,
    _0098_,
    _0097_,
    _0096_,
    _0095_,
    _0093_,
    _0092_,
    _0091_,
    _0090_,
    _0089_,
    _0088_,
    _0087_,
    _0086_,
    _0085_,
    _0084_,
    _0082_,
    _0081_,
    _0080_,
    _0079_,
    _0078_,
    _0077_,
    _0076_,
    _0075_,
    _0074_,
    _0073_,
    _0071_,
    _0070_,
    _0069_,
    _0068_,
    _0067_,
    _0066_,
    _0065_,
    _0064_,
    _0063_,
    _0062_,
    _0060_,
    _0059_,
    _0058_,
    _0057_,
    _0056_,
    _0055_,
    _0054_,
    _0053_,
    _0052_,
    _0051_,
    _0049_,
    _0048_,
    _0047_,
    _0046_,
    _0045_,
    _0044_,
    _0043_,
    _0042_,
    _0041_,
    _0040_,
    _0038_,
    _0037_,
    _0036_,
    _0035_,
    _0034_,
    _0033_,
    _0032_,
    _0031_,
    _0022_,
    _0011_,
    _0127_,
    _0116_,
    _0105_,
    _0094_,
    _0083_,
    _0072_,
    _0061_,
    _0050_,
    _0039_,
    _0000_}));
 sg13g2_inv_1 \digitalenH.g[0].u.inv1  (.Y(\digitalenH.g[0].u.OUTN ),
    .A(net7));
 sg13g2_inv_1 \digitalenH.g[0].u.inv2  (.Y(\digitalenH.g[0].u.OUTP ),
    .A(\digitalenH.g[0].u.OUTN ));
 sg13g2_inv_1 \digitalenH.g[1].u.inv1  (.Y(\digitalenH.g[1].u.OUTN ),
    .A(net7));
 sg13g2_inv_1 \digitalenH.g[1].u.inv2  (.Y(\digitalenH.g[1].u.OUTP ),
    .A(\digitalenH.g[1].u.OUTN ));
 sg13g2_inv_1 \digitalenH.g[2].u.inv1  (.Y(\digitalenH.g[2].u.OUTN ),
    .A(net7));
 sg13g2_inv_1 \digitalenH.g[2].u.inv2  (.Y(\digitalenH.g[2].u.OUTP ),
    .A(\digitalenH.g[2].u.OUTN ));
 sg13g2_inv_1 \digitalenH.g[3].u.inv1  (.Y(\digitalenH.g[3].u.OUTN ),
    .A(net7));
 sg13g2_inv_1 \digitalenH.g[3].u.inv2  (.Y(\digitalenH.g[3].u.OUTP ),
    .A(\digitalenH.g[3].u.OUTN ));
 sg13g2_inv_1 \digitalenL.g[0].u.inv1  (.Y(\digitalenL.g[0].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalenL.g[0].u.inv2  (.Y(\digitalenL.g[0].u.OUTP ),
    .A(\digitalenL.g[0].u.OUTN ));
 sg13g2_inv_1 \digitalenL.g[1].u.inv1  (.Y(\digitalenL.g[1].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalenL.g[1].u.inv2  (.Y(\digitalenL.g[1].u.OUTP ),
    .A(\digitalenL.g[1].u.OUTN ));
 sg13g2_inv_1 \digitalenL.g[2].u.inv1  (.Y(\digitalenL.g[2].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalenL.g[2].u.inv2  (.Y(\digitalenL.g[2].u.OUTP ),
    .A(\digitalenL.g[2].u.OUTN ));
 sg13g2_inv_1 \digitalenL.g[3].u.inv1  (.Y(\digitalenL.g[3].u.OUTN ),
    .A(net6));
 sg13g2_inv_1 \digitalenL.g[3].u.inv2  (.Y(\digitalenL.g[3].u.OUTP ),
    .A(\digitalenL.g[3].u.OUTN ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[2]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[3]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[4]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[5]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[6]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[7]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[0]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[1]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[2]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[3]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[4]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[5]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[6]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[7]));
 sg13g2_buf_1 fanout24 (.A(net26),
    .X(net24));
 sg13g2_buf_1 fanout25 (.A(net26),
    .X(net25));
 sg13g2_buf_1 fanout26 (.A(net33),
    .X(net26));
 sg13g2_buf_1 fanout27 (.A(net28),
    .X(net27));
 sg13g2_buf_1 fanout28 (.A(net33),
    .X(net28));
 sg13g2_buf_1 fanout29 (.A(net32),
    .X(net29));
 sg13g2_buf_1 fanout30 (.A(net32),
    .X(net30));
 sg13g2_buf_1 fanout31 (.A(net32),
    .X(net31));
 sg13g2_buf_1 fanout32 (.A(net33),
    .X(net32));
 sg13g2_buf_1 fanout33 (.A(net68),
    .X(net33));
 sg13g2_buf_1 fanout34 (.A(net36),
    .X(net34));
 sg13g2_buf_1 fanout35 (.A(net40),
    .X(net35));
 sg13g2_buf_1 fanout36 (.A(net40),
    .X(net36));
 sg13g2_buf_1 fanout37 (.A(net39),
    .X(net37));
 sg13g2_buf_1 fanout38 (.A(net40),
    .X(net38));
 sg13g2_buf_1 fanout39 (.A(net40),
    .X(net39));
 sg13g2_buf_1 fanout40 (.A(net68),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(net43),
    .X(net41));
 sg13g2_buf_1 fanout42 (.A(net43),
    .X(net42));
 sg13g2_buf_1 fanout43 (.A(net48),
    .X(net43));
 sg13g2_buf_1 fanout44 (.A(net48),
    .X(net44));
 sg13g2_buf_1 fanout45 (.A(net48),
    .X(net45));
 sg13g2_buf_1 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_1 fanout47 (.A(net48),
    .X(net47));
 sg13g2_buf_1 fanout48 (.A(net68),
    .X(net48));
 sg13g2_buf_1 fanout49 (.A(net51),
    .X(net49));
 sg13g2_buf_1 fanout50 (.A(net51),
    .X(net50));
 sg13g2_buf_1 fanout51 (.A(net52),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(net68),
    .X(net52));
 sg13g2_buf_1 fanout53 (.A(net55),
    .X(net53));
 sg13g2_buf_1 fanout54 (.A(net55),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(net56),
    .X(net55));
 sg13g2_buf_1 fanout56 (.A(net68),
    .X(net56));
 sg13g2_buf_1 fanout57 (.A(net67),
    .X(net57));
 sg13g2_buf_1 fanout58 (.A(net67),
    .X(net58));
 sg13g2_buf_1 fanout59 (.A(net61),
    .X(net59));
 sg13g2_buf_1 fanout60 (.A(net61),
    .X(net60));
 sg13g2_buf_1 fanout61 (.A(net67),
    .X(net61));
 sg13g2_buf_1 fanout62 (.A(net64),
    .X(net62));
 sg13g2_buf_1 fanout63 (.A(net64),
    .X(net63));
 sg13g2_buf_1 fanout64 (.A(net67),
    .X(net64));
 sg13g2_buf_1 fanout65 (.A(net67),
    .X(net65));
 sg13g2_buf_1 fanout66 (.A(net67),
    .X(net66));
 sg13g2_buf_1 fanout67 (.A(net68),
    .X(net67));
 sg13g2_buf_1 fanout68 (.A(_0515_),
    .X(net68));
 sg13g2_buf_1 fanout69 (.A(net72),
    .X(net69));
 sg13g2_buf_1 fanout70 (.A(net72),
    .X(net70));
 sg13g2_buf_1 fanout71 (.A(net72),
    .X(net71));
 sg13g2_buf_1 fanout72 (.A(net78),
    .X(net72));
 sg13g2_buf_1 fanout73 (.A(net74),
    .X(net73));
 sg13g2_buf_1 fanout74 (.A(net78),
    .X(net74));
 sg13g2_buf_1 fanout75 (.A(net77),
    .X(net75));
 sg13g2_buf_1 fanout76 (.A(net77),
    .X(net76));
 sg13g2_buf_1 fanout77 (.A(net78),
    .X(net77));
 sg13g2_buf_1 fanout78 (.A(net112),
    .X(net78));
 sg13g2_buf_1 fanout79 (.A(net81),
    .X(net79));
 sg13g2_buf_1 fanout80 (.A(net81),
    .X(net80));
 sg13g2_buf_1 fanout81 (.A(net91),
    .X(net81));
 sg13g2_buf_1 fanout82 (.A(net83),
    .X(net82));
 sg13g2_buf_1 fanout83 (.A(net91),
    .X(net83));
 sg13g2_buf_1 fanout84 (.A(net86),
    .X(net84));
 sg13g2_buf_1 fanout85 (.A(net86),
    .X(net85));
 sg13g2_buf_1 fanout86 (.A(net91),
    .X(net86));
 sg13g2_buf_1 fanout87 (.A(net90),
    .X(net87));
 sg13g2_buf_1 fanout88 (.A(net90),
    .X(net88));
 sg13g2_buf_1 fanout89 (.A(net90),
    .X(net89));
 sg13g2_buf_1 fanout90 (.A(net91),
    .X(net90));
 sg13g2_buf_1 fanout91 (.A(net112),
    .X(net91));
 sg13g2_buf_1 fanout92 (.A(net96),
    .X(net92));
 sg13g2_buf_1 fanout93 (.A(net96),
    .X(net93));
 sg13g2_buf_1 fanout94 (.A(net96),
    .X(net94));
 sg13g2_buf_1 fanout95 (.A(net96),
    .X(net95));
 sg13g2_buf_1 fanout96 (.A(net112),
    .X(net96));
 sg13g2_buf_1 fanout97 (.A(net101),
    .X(net97));
 sg13g2_buf_1 fanout98 (.A(net101),
    .X(net98));
 sg13g2_buf_1 fanout99 (.A(net101),
    .X(net99));
 sg13g2_buf_1 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_1 fanout101 (.A(net112),
    .X(net101));
 sg13g2_buf_1 fanout102 (.A(net103),
    .X(net102));
 sg13g2_buf_1 fanout103 (.A(net111),
    .X(net103));
 sg13g2_buf_1 fanout104 (.A(net111),
    .X(net104));
 sg13g2_buf_1 fanout105 (.A(net111),
    .X(net105));
 sg13g2_buf_1 fanout106 (.A(net110),
    .X(net106));
 sg13g2_buf_1 fanout107 (.A(net110),
    .X(net107));
 sg13g2_buf_1 fanout108 (.A(net110),
    .X(net108));
 sg13g2_buf_1 fanout109 (.A(net110),
    .X(net109));
 sg13g2_buf_1 fanout110 (.A(net111),
    .X(net110));
 sg13g2_buf_1 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_1 fanout112 (.A(_0512_),
    .X(net112));
 sg13g2_buf_1 fanout113 (.A(net115),
    .X(net113));
 sg13g2_buf_1 fanout114 (.A(net115),
    .X(net114));
 sg13g2_buf_1 fanout115 (.A(net137),
    .X(net115));
 sg13g2_buf_1 fanout116 (.A(net117),
    .X(net116));
 sg13g2_buf_1 fanout117 (.A(net122),
    .X(net117));
 sg13g2_buf_1 fanout118 (.A(net121),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(net121),
    .X(net119));
 sg13g2_buf_1 fanout120 (.A(net121),
    .X(net120));
 sg13g2_buf_1 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_1 fanout122 (.A(net137),
    .X(net122));
 sg13g2_buf_1 fanout123 (.A(net125),
    .X(net123));
 sg13g2_buf_1 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_1 fanout125 (.A(net136),
    .X(net125));
 sg13g2_buf_1 fanout126 (.A(net127),
    .X(net126));
 sg13g2_buf_1 fanout127 (.A(net136),
    .X(net127));
 sg13g2_buf_1 fanout128 (.A(net130),
    .X(net128));
 sg13g2_buf_1 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_1 fanout130 (.A(net136),
    .X(net130));
 sg13g2_buf_1 fanout131 (.A(net135),
    .X(net131));
 sg13g2_buf_1 fanout132 (.A(net135),
    .X(net132));
 sg13g2_buf_1 fanout133 (.A(net135),
    .X(net133));
 sg13g2_buf_1 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_1 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_1 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_1 fanout137 (.A(net158),
    .X(net137));
 sg13g2_buf_1 fanout138 (.A(net142),
    .X(net138));
 sg13g2_buf_1 fanout139 (.A(net142),
    .X(net139));
 sg13g2_buf_1 fanout140 (.A(net142),
    .X(net140));
 sg13g2_buf_1 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_1 fanout142 (.A(net147),
    .X(net142));
 sg13g2_buf_1 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_1 fanout144 (.A(net147),
    .X(net144));
 sg13g2_buf_1 fanout145 (.A(net147),
    .X(net145));
 sg13g2_buf_1 fanout146 (.A(net147),
    .X(net146));
 sg13g2_buf_1 fanout147 (.A(net158),
    .X(net147));
 sg13g2_buf_1 fanout148 (.A(net152),
    .X(net148));
 sg13g2_buf_1 fanout149 (.A(net152),
    .X(net149));
 sg13g2_buf_1 fanout150 (.A(net152),
    .X(net150));
 sg13g2_buf_1 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_1 fanout152 (.A(net158),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(net157),
    .X(net153));
 sg13g2_buf_1 fanout154 (.A(net157),
    .X(net154));
 sg13g2_buf_1 fanout155 (.A(net157),
    .X(net155));
 sg13g2_buf_1 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_1 fanout157 (.A(net158),
    .X(net157));
 sg13g2_buf_1 fanout158 (.A(_1026_),
    .X(net158));
 sg13g2_buf_1 fanout159 (.A(net161),
    .X(net159));
 sg13g2_buf_1 fanout160 (.A(net161),
    .X(net160));
 sg13g2_buf_1 fanout161 (.A(net169),
    .X(net161));
 sg13g2_buf_1 fanout162 (.A(net164),
    .X(net162));
 sg13g2_buf_1 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_1 fanout164 (.A(net169),
    .X(net164));
 sg13g2_buf_1 fanout165 (.A(net168),
    .X(net165));
 sg13g2_buf_1 fanout166 (.A(net168),
    .X(net166));
 sg13g2_buf_1 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_1 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_1 fanout169 (.A(net204),
    .X(net169));
 sg13g2_buf_1 fanout170 (.A(net172),
    .X(net170));
 sg13g2_buf_1 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_1 fanout172 (.A(net183),
    .X(net172));
 sg13g2_buf_1 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_1 fanout174 (.A(net183),
    .X(net174));
 sg13g2_buf_1 fanout175 (.A(net178),
    .X(net175));
 sg13g2_buf_1 fanout176 (.A(net178),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_1 fanout178 (.A(net183),
    .X(net178));
 sg13g2_buf_1 fanout179 (.A(net182),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(net182),
    .X(net180));
 sg13g2_buf_1 fanout181 (.A(net182),
    .X(net181));
 sg13g2_buf_1 fanout182 (.A(net183),
    .X(net182));
 sg13g2_buf_1 fanout183 (.A(net204),
    .X(net183));
 sg13g2_buf_1 fanout184 (.A(net186),
    .X(net184));
 sg13g2_buf_1 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_1 fanout186 (.A(net187),
    .X(net186));
 sg13g2_buf_1 fanout187 (.A(net193),
    .X(net187));
 sg13g2_buf_1 fanout188 (.A(net191),
    .X(net188));
 sg13g2_buf_1 fanout189 (.A(net191),
    .X(net189));
 sg13g2_buf_1 fanout190 (.A(net191),
    .X(net190));
 sg13g2_buf_1 fanout191 (.A(net193),
    .X(net191));
 sg13g2_buf_1 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_1 fanout193 (.A(net204),
    .X(net193));
 sg13g2_buf_1 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_1 fanout195 (.A(net198),
    .X(net195));
 sg13g2_buf_1 fanout196 (.A(net198),
    .X(net196));
 sg13g2_buf_1 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_1 fanout198 (.A(net204),
    .X(net198));
 sg13g2_buf_1 fanout199 (.A(net203),
    .X(net199));
 sg13g2_buf_1 fanout200 (.A(net203),
    .X(net200));
 sg13g2_buf_1 fanout201 (.A(net203),
    .X(net201));
 sg13g2_buf_1 fanout202 (.A(net203),
    .X(net202));
 sg13g2_buf_1 fanout203 (.A(net204),
    .X(net203));
 sg13g2_buf_1 fanout204 (.A(net5),
    .X(net204));
 sg13g2_buf_1 fanout205 (.A(net210),
    .X(net205));
 sg13g2_buf_1 fanout206 (.A(net209),
    .X(net206));
 sg13g2_buf_1 fanout207 (.A(net209),
    .X(net207));
 sg13g2_buf_1 fanout208 (.A(net209),
    .X(net208));
 sg13g2_buf_1 fanout209 (.A(net210),
    .X(net209));
 sg13g2_buf_1 fanout210 (.A(net228),
    .X(net210));
 sg13g2_buf_1 fanout211 (.A(net212),
    .X(net211));
 sg13g2_buf_1 fanout212 (.A(net217),
    .X(net212));
 sg13g2_buf_1 fanout213 (.A(net216),
    .X(net213));
 sg13g2_buf_1 fanout214 (.A(net216),
    .X(net214));
 sg13g2_buf_1 fanout215 (.A(net216),
    .X(net215));
 sg13g2_buf_1 fanout216 (.A(net217),
    .X(net216));
 sg13g2_buf_1 fanout217 (.A(net228),
    .X(net217));
 sg13g2_buf_1 fanout218 (.A(net220),
    .X(net218));
 sg13g2_buf_1 fanout219 (.A(net220),
    .X(net219));
 sg13g2_buf_1 fanout220 (.A(net228),
    .X(net220));
 sg13g2_buf_1 fanout221 (.A(net222),
    .X(net221));
 sg13g2_buf_1 fanout222 (.A(net228),
    .X(net222));
 sg13g2_buf_1 fanout223 (.A(net227),
    .X(net223));
 sg13g2_buf_1 fanout224 (.A(net227),
    .X(net224));
 sg13g2_buf_1 fanout225 (.A(net227),
    .X(net225));
 sg13g2_buf_1 fanout226 (.A(net227),
    .X(net226));
 sg13g2_buf_1 fanout227 (.A(net228),
    .X(net227));
 sg13g2_buf_1 fanout228 (.A(net4),
    .X(net228));
 sg13g2_tiehi _2502__229 (.L_HI(net));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_16 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_16 clkbuf_2_0__f_clk (.X(clknet_2_0__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_1__f_clk (.X(clknet_2_1__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_2__f_clk (.X(clknet_2_2__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_16 clkbuf_2_3__f_clk (.X(clknet_2_3__leaf_clk),
    .A(clknet_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_leaf_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_18_clk));
 sg13g2_inv_8 clkload3 (.A(clknet_leaf_19_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_3_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_4_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_7_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_13_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_14_clk));
 sg13g2_inv_8 clkload9 (.A(clknet_leaf_16_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_17_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_8_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_9_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0131_));
 sg13g2_antennanp ANTENNA_2 (.A(_0144_));
 sg13g2_antennanp ANTENNA_3 (.A(_0144_));
 sg13g2_antennanp ANTENNA_4 (.A(_0150_));
 sg13g2_antennanp ANTENNA_5 (.A(_0150_));
 sg13g2_antennanp ANTENNA_6 (.A(_0151_));
 sg13g2_antennanp ANTENNA_7 (.A(_0151_));
 sg13g2_antennanp ANTENNA_8 (.A(_0159_));
 sg13g2_antennanp ANTENNA_9 (.A(_0162_));
 sg13g2_antennanp ANTENNA_10 (.A(_0163_));
 sg13g2_antennanp ANTENNA_11 (.A(_0175_));
 sg13g2_antennanp ANTENNA_12 (.A(_0249_));
 sg13g2_antennanp ANTENNA_13 (.A(_0249_));
 sg13g2_antennanp ANTENNA_14 (.A(\daisychain[110] ));
 sg13g2_antennanp ANTENNA_15 (.A(\daisychain[110] ));
 sg13g2_antennanp ANTENNA_16 (.A(\daisychain[113] ));
 sg13g2_antennanp ANTENNA_17 (.A(\daisychain[27] ));
 sg13g2_antennanp ANTENNA_18 (.A(\daisychain[27] ));
 sg13g2_antennanp ANTENNA_19 (.A(\daisychain[9] ));
 sg13g2_antennanp ANTENNA_20 (.A(_0129_));
 sg13g2_antennanp ANTENNA_21 (.A(_0133_));
 sg13g2_antennanp ANTENNA_22 (.A(_0136_));
 sg13g2_antennanp ANTENNA_23 (.A(_0138_));
 sg13g2_antennanp ANTENNA_24 (.A(_0140_));
 sg13g2_antennanp ANTENNA_25 (.A(_0140_));
 sg13g2_antennanp ANTENNA_26 (.A(_0166_));
 sg13g2_antennanp ANTENNA_27 (.A(_0179_));
 sg13g2_antennanp ANTENNA_28 (.A(_0179_));
 sg13g2_antennanp ANTENNA_29 (.A(_0190_));
 sg13g2_antennanp ANTENNA_30 (.A(_0200_));
 sg13g2_antennanp ANTENNA_31 (.A(_0200_));
 sg13g2_antennanp ANTENNA_32 (.A(_0233_));
 sg13g2_antennanp ANTENNA_33 (.A(_0234_));
 sg13g2_antennanp ANTENNA_34 (.A(_0243_));
 sg13g2_antennanp ANTENNA_35 (.A(_0243_));
 sg13g2_antennanp ANTENNA_36 (.A(_0250_));
 sg13g2_antennanp ANTENNA_37 (.A(_0251_));
 sg13g2_antennanp ANTENNA_38 (.A(_0253_));
 sg13g2_antennanp ANTENNA_39 (.A(_0253_));
 sg13g2_antennanp ANTENNA_40 (.A(\daisychain[104] ));
 sg13g2_antennanp ANTENNA_41 (.A(\daisychain[114] ));
 sg13g2_antennanp ANTENNA_42 (.A(\daisychain[11] ));
 sg13g2_antennanp ANTENNA_43 (.A(\daisychain[11] ));
 sg13g2_antennanp ANTENNA_44 (.A(\daisychain[11] ));
 sg13g2_antennanp ANTENNA_45 (.A(\daisychain[126] ));
 sg13g2_antennanp ANTENNA_46 (.A(\daisychain[127] ));
 sg13g2_antennanp ANTENNA_47 (.A(\daisychain[15] ));
 sg13g2_antennanp ANTENNA_48 (.A(\daisychain[29] ));
 sg13g2_antennanp ANTENNA_49 (.A(\daisychain[29] ));
 sg13g2_antennanp ANTENNA_50 (.A(\daisychain[2] ));
 sg13g2_antennanp ANTENNA_51 (.A(\daisychain[37] ));
 sg13g2_antennanp ANTENNA_52 (.A(\daisychain[41] ));
 sg13g2_antennanp ANTENNA_53 (.A(\daisychain[41] ));
 sg13g2_antennanp ANTENNA_54 (.A(\daisychain[42] ));
 sg13g2_antennanp ANTENNA_55 (.A(\daisychain[79] ));
 sg13g2_antennanp ANTENNA_56 (.A(\daisychain[88] ));
 sg13g2_antennanp ANTENNA_57 (.A(_0187_));
 sg13g2_antennanp ANTENNA_58 (.A(\daisychain[100] ));
 sg13g2_antennanp ANTENNA_59 (.A(\daisychain[126] ));
 sg13g2_antennanp ANTENNA_60 (.A(\daisychain[126] ));
 sg13g2_antennanp ANTENNA_61 (.A(\daisychain[126] ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_4 FILLER_0_709 ();
 sg13g2_fill_2 FILLER_0_713 ();
 sg13g2_decap_4 FILLER_0_720 ();
 sg13g2_fill_1 FILLER_0_724 ();
 sg13g2_decap_4 FILLER_0_729 ();
 sg13g2_fill_2 FILLER_0_733 ();
 sg13g2_fill_2 FILLER_0_762 ();
 sg13g2_decap_8 FILLER_0_768 ();
 sg13g2_fill_2 FILLER_0_775 ();
 sg13g2_decap_8 FILLER_0_786 ();
 sg13g2_decap_8 FILLER_0_793 ();
 sg13g2_decap_8 FILLER_0_800 ();
 sg13g2_decap_8 FILLER_0_807 ();
 sg13g2_fill_2 FILLER_0_814 ();
 sg13g2_fill_1 FILLER_0_816 ();
 sg13g2_decap_8 FILLER_0_830 ();
 sg13g2_decap_8 FILLER_0_837 ();
 sg13g2_fill_2 FILLER_0_844 ();
 sg13g2_fill_1 FILLER_0_846 ();
 sg13g2_fill_2 FILLER_0_851 ();
 sg13g2_fill_1 FILLER_0_853 ();
 sg13g2_decap_8 FILLER_0_863 ();
 sg13g2_decap_4 FILLER_0_870 ();
 sg13g2_fill_2 FILLER_0_874 ();
 sg13g2_fill_1 FILLER_0_880 ();
 sg13g2_decap_4 FILLER_0_890 ();
 sg13g2_decap_8 FILLER_0_901 ();
 sg13g2_decap_8 FILLER_0_912 ();
 sg13g2_decap_8 FILLER_0_919 ();
 sg13g2_decap_4 FILLER_0_926 ();
 sg13g2_fill_1 FILLER_0_930 ();
 sg13g2_decap_8 FILLER_0_944 ();
 sg13g2_decap_8 FILLER_0_951 ();
 sg13g2_decap_8 FILLER_0_958 ();
 sg13g2_decap_4 FILLER_0_965 ();
 sg13g2_fill_1 FILLER_0_969 ();
 sg13g2_fill_2 FILLER_0_974 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_fill_2 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1012 ();
 sg13g2_decap_8 FILLER_0_1019 ();
 sg13g2_fill_2 FILLER_0_1026 ();
 sg13g2_fill_1 FILLER_0_1028 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_fill_2 FILLER_1_693 ();
 sg13g2_fill_1 FILLER_1_695 ();
 sg13g2_fill_1 FILLER_1_750 ();
 sg13g2_fill_2 FILLER_1_810 ();
 sg13g2_fill_1 FILLER_1_812 ();
 sg13g2_fill_2 FILLER_1_840 ();
 sg13g2_fill_2 FILLER_1_869 ();
 sg13g2_decap_4 FILLER_1_898 ();
 sg13g2_fill_1 FILLER_1_902 ();
 sg13g2_decap_4 FILLER_1_957 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_2_410 ();
 sg13g2_decap_8 FILLER_2_417 ();
 sg13g2_decap_8 FILLER_2_424 ();
 sg13g2_decap_8 FILLER_2_431 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_decap_8 FILLER_2_452 ();
 sg13g2_decap_8 FILLER_2_459 ();
 sg13g2_decap_8 FILLER_2_466 ();
 sg13g2_decap_8 FILLER_2_473 ();
 sg13g2_decap_8 FILLER_2_480 ();
 sg13g2_decap_8 FILLER_2_487 ();
 sg13g2_decap_8 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_501 ();
 sg13g2_decap_8 FILLER_2_508 ();
 sg13g2_decap_8 FILLER_2_515 ();
 sg13g2_decap_8 FILLER_2_522 ();
 sg13g2_decap_8 FILLER_2_529 ();
 sg13g2_decap_8 FILLER_2_536 ();
 sg13g2_decap_8 FILLER_2_543 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_599 ();
 sg13g2_decap_8 FILLER_2_606 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_decap_8 FILLER_2_620 ();
 sg13g2_decap_8 FILLER_2_627 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_4 FILLER_2_669 ();
 sg13g2_fill_2 FILLER_2_673 ();
 sg13g2_decap_8 FILLER_2_684 ();
 sg13g2_decap_8 FILLER_2_691 ();
 sg13g2_decap_4 FILLER_2_698 ();
 sg13g2_fill_1 FILLER_2_706 ();
 sg13g2_decap_4 FILLER_2_712 ();
 sg13g2_fill_1 FILLER_2_716 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_fill_1 FILLER_2_735 ();
 sg13g2_fill_1 FILLER_2_745 ();
 sg13g2_decap_8 FILLER_2_750 ();
 sg13g2_fill_2 FILLER_2_757 ();
 sg13g2_fill_1 FILLER_2_759 ();
 sg13g2_decap_4 FILLER_2_774 ();
 sg13g2_fill_2 FILLER_2_778 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_fill_1 FILLER_2_791 ();
 sg13g2_fill_1 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_829 ();
 sg13g2_decap_8 FILLER_2_836 ();
 sg13g2_fill_1 FILLER_2_843 ();
 sg13g2_decap_8 FILLER_2_853 ();
 sg13g2_decap_8 FILLER_2_860 ();
 sg13g2_decap_8 FILLER_2_867 ();
 sg13g2_decap_8 FILLER_2_874 ();
 sg13g2_decap_8 FILLER_2_881 ();
 sg13g2_decap_4 FILLER_2_888 ();
 sg13g2_fill_1 FILLER_2_897 ();
 sg13g2_fill_1 FILLER_2_906 ();
 sg13g2_decap_8 FILLER_2_912 ();
 sg13g2_decap_8 FILLER_2_919 ();
 sg13g2_decap_4 FILLER_2_926 ();
 sg13g2_fill_1 FILLER_2_930 ();
 sg13g2_decap_8 FILLER_2_951 ();
 sg13g2_fill_2 FILLER_2_958 ();
 sg13g2_fill_1 FILLER_2_960 ();
 sg13g2_decap_8 FILLER_2_981 ();
 sg13g2_decap_8 FILLER_2_988 ();
 sg13g2_fill_2 FILLER_2_995 ();
 sg13g2_decap_4 FILLER_2_1002 ();
 sg13g2_fill_1 FILLER_2_1006 ();
 sg13g2_decap_8 FILLER_2_1019 ();
 sg13g2_fill_2 FILLER_2_1026 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_137 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_4 FILLER_3_417 ();
 sg13g2_fill_1 FILLER_3_421 ();
 sg13g2_decap_8 FILLER_3_426 ();
 sg13g2_decap_8 FILLER_3_433 ();
 sg13g2_decap_8 FILLER_3_440 ();
 sg13g2_decap_8 FILLER_3_447 ();
 sg13g2_decap_8 FILLER_3_454 ();
 sg13g2_decap_8 FILLER_3_461 ();
 sg13g2_decap_8 FILLER_3_468 ();
 sg13g2_decap_8 FILLER_3_475 ();
 sg13g2_decap_8 FILLER_3_482 ();
 sg13g2_decap_8 FILLER_3_489 ();
 sg13g2_decap_8 FILLER_3_496 ();
 sg13g2_decap_8 FILLER_3_503 ();
 sg13g2_decap_8 FILLER_3_510 ();
 sg13g2_decap_8 FILLER_3_517 ();
 sg13g2_decap_8 FILLER_3_524 ();
 sg13g2_decap_8 FILLER_3_531 ();
 sg13g2_decap_8 FILLER_3_538 ();
 sg13g2_decap_8 FILLER_3_545 ();
 sg13g2_decap_8 FILLER_3_552 ();
 sg13g2_decap_8 FILLER_3_559 ();
 sg13g2_decap_8 FILLER_3_566 ();
 sg13g2_decap_8 FILLER_3_573 ();
 sg13g2_decap_8 FILLER_3_580 ();
 sg13g2_decap_8 FILLER_3_587 ();
 sg13g2_decap_8 FILLER_3_594 ();
 sg13g2_decap_8 FILLER_3_601 ();
 sg13g2_decap_8 FILLER_3_608 ();
 sg13g2_decap_8 FILLER_3_615 ();
 sg13g2_decap_8 FILLER_3_622 ();
 sg13g2_decap_8 FILLER_3_629 ();
 sg13g2_decap_8 FILLER_3_636 ();
 sg13g2_decap_8 FILLER_3_643 ();
 sg13g2_decap_8 FILLER_3_650 ();
 sg13g2_decap_8 FILLER_3_657 ();
 sg13g2_decap_4 FILLER_3_664 ();
 sg13g2_fill_1 FILLER_3_668 ();
 sg13g2_decap_8 FILLER_3_696 ();
 sg13g2_fill_2 FILLER_3_703 ();
 sg13g2_fill_1 FILLER_3_705 ();
 sg13g2_decap_8 FILLER_3_713 ();
 sg13g2_decap_8 FILLER_3_720 ();
 sg13g2_decap_8 FILLER_3_727 ();
 sg13g2_decap_4 FILLER_3_734 ();
 sg13g2_fill_1 FILLER_3_738 ();
 sg13g2_decap_8 FILLER_3_752 ();
 sg13g2_fill_2 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_fill_1 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_808 ();
 sg13g2_decap_8 FILLER_3_815 ();
 sg13g2_decap_4 FILLER_3_829 ();
 sg13g2_fill_1 FILLER_3_833 ();
 sg13g2_fill_2 FILLER_3_865 ();
 sg13g2_fill_1 FILLER_3_867 ();
 sg13g2_fill_1 FILLER_3_900 ();
 sg13g2_decap_8 FILLER_3_914 ();
 sg13g2_fill_2 FILLER_3_921 ();
 sg13g2_fill_1 FILLER_3_923 ();
 sg13g2_decap_8 FILLER_3_955 ();
 sg13g2_decap_8 FILLER_3_962 ();
 sg13g2_decap_4 FILLER_3_969 ();
 sg13g2_fill_1 FILLER_3_1008 ();
 sg13g2_decap_8 FILLER_3_1013 ();
 sg13g2_decap_8 FILLER_3_1020 ();
 sg13g2_fill_2 FILLER_3_1027 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_decap_8 FILLER_4_39 ();
 sg13g2_decap_8 FILLER_4_46 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_decap_8 FILLER_4_67 ();
 sg13g2_decap_8 FILLER_4_74 ();
 sg13g2_decap_8 FILLER_4_81 ();
 sg13g2_decap_8 FILLER_4_88 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_179 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_decap_8 FILLER_4_214 ();
 sg13g2_decap_8 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_228 ();
 sg13g2_decap_8 FILLER_4_235 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_decap_8 FILLER_4_249 ();
 sg13g2_decap_8 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_263 ();
 sg13g2_decap_8 FILLER_4_270 ();
 sg13g2_decap_8 FILLER_4_277 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_8 FILLER_4_424 ();
 sg13g2_decap_8 FILLER_4_431 ();
 sg13g2_decap_8 FILLER_4_438 ();
 sg13g2_decap_8 FILLER_4_445 ();
 sg13g2_decap_8 FILLER_4_452 ();
 sg13g2_decap_8 FILLER_4_459 ();
 sg13g2_decap_4 FILLER_4_466 ();
 sg13g2_fill_2 FILLER_4_470 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_4 FILLER_4_637 ();
 sg13g2_fill_2 FILLER_4_650 ();
 sg13g2_fill_1 FILLER_4_652 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_fill_2 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_690 ();
 sg13g2_decap_4 FILLER_4_697 ();
 sg13g2_fill_2 FILLER_4_701 ();
 sg13g2_fill_2 FILLER_4_738 ();
 sg13g2_fill_1 FILLER_4_740 ();
 sg13g2_decap_8 FILLER_4_775 ();
 sg13g2_decap_8 FILLER_4_782 ();
 sg13g2_decap_8 FILLER_4_789 ();
 sg13g2_fill_2 FILLER_4_796 ();
 sg13g2_decap_8 FILLER_4_823 ();
 sg13g2_decap_8 FILLER_4_830 ();
 sg13g2_decap_4 FILLER_4_846 ();
 sg13g2_decap_8 FILLER_4_857 ();
 sg13g2_decap_4 FILLER_4_864 ();
 sg13g2_fill_2 FILLER_4_868 ();
 sg13g2_decap_8 FILLER_4_883 ();
 sg13g2_fill_2 FILLER_4_890 ();
 sg13g2_decap_8 FILLER_4_896 ();
 sg13g2_decap_4 FILLER_4_903 ();
 sg13g2_fill_2 FILLER_4_907 ();
 sg13g2_decap_8 FILLER_4_918 ();
 sg13g2_decap_8 FILLER_4_925 ();
 sg13g2_fill_2 FILLER_4_932 ();
 sg13g2_fill_1 FILLER_4_934 ();
 sg13g2_decap_8 FILLER_4_952 ();
 sg13g2_decap_4 FILLER_4_959 ();
 sg13g2_fill_1 FILLER_4_963 ();
 sg13g2_decap_4 FILLER_4_973 ();
 sg13g2_fill_1 FILLER_4_977 ();
 sg13g2_decap_8 FILLER_4_982 ();
 sg13g2_decap_8 FILLER_4_989 ();
 sg13g2_fill_1 FILLER_4_996 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_165 ();
 sg13g2_decap_8 FILLER_5_172 ();
 sg13g2_decap_8 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_200 ();
 sg13g2_decap_8 FILLER_5_207 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_decap_8 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_8 FILLER_5_298 ();
 sg13g2_decap_8 FILLER_5_305 ();
 sg13g2_decap_8 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_361 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_8 FILLER_5_403 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_8 FILLER_5_424 ();
 sg13g2_decap_8 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_438 ();
 sg13g2_decap_8 FILLER_5_445 ();
 sg13g2_decap_8 FILLER_5_452 ();
 sg13g2_decap_8 FILLER_5_459 ();
 sg13g2_decap_8 FILLER_5_466 ();
 sg13g2_decap_8 FILLER_5_473 ();
 sg13g2_decap_8 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_494 ();
 sg13g2_decap_8 FILLER_5_501 ();
 sg13g2_fill_1 FILLER_5_508 ();
 sg13g2_decap_8 FILLER_5_513 ();
 sg13g2_decap_8 FILLER_5_520 ();
 sg13g2_decap_8 FILLER_5_527 ();
 sg13g2_decap_8 FILLER_5_534 ();
 sg13g2_decap_8 FILLER_5_541 ();
 sg13g2_decap_8 FILLER_5_548 ();
 sg13g2_decap_8 FILLER_5_555 ();
 sg13g2_decap_8 FILLER_5_562 ();
 sg13g2_decap_8 FILLER_5_569 ();
 sg13g2_decap_8 FILLER_5_576 ();
 sg13g2_decap_8 FILLER_5_583 ();
 sg13g2_decap_8 FILLER_5_590 ();
 sg13g2_decap_8 FILLER_5_597 ();
 sg13g2_decap_8 FILLER_5_604 ();
 sg13g2_decap_8 FILLER_5_611 ();
 sg13g2_decap_8 FILLER_5_618 ();
 sg13g2_decap_8 FILLER_5_625 ();
 sg13g2_decap_4 FILLER_5_632 ();
 sg13g2_fill_1 FILLER_5_636 ();
 sg13g2_decap_8 FILLER_5_668 ();
 sg13g2_decap_8 FILLER_5_675 ();
 sg13g2_fill_1 FILLER_5_682 ();
 sg13g2_decap_8 FILLER_5_696 ();
 sg13g2_fill_2 FILLER_5_703 ();
 sg13g2_fill_1 FILLER_5_705 ();
 sg13g2_fill_2 FILLER_5_711 ();
 sg13g2_fill_1 FILLER_5_713 ();
 sg13g2_decap_8 FILLER_5_722 ();
 sg13g2_decap_8 FILLER_5_729 ();
 sg13g2_fill_2 FILLER_5_736 ();
 sg13g2_decap_8 FILLER_5_754 ();
 sg13g2_decap_8 FILLER_5_761 ();
 sg13g2_decap_4 FILLER_5_768 ();
 sg13g2_fill_2 FILLER_5_772 ();
 sg13g2_decap_4 FILLER_5_828 ();
 sg13g2_decap_4 FILLER_5_900 ();
 sg13g2_fill_2 FILLER_5_931 ();
 sg13g2_decap_8 FILLER_5_1018 ();
 sg13g2_decap_4 FILLER_5_1025 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_25 ();
 sg13g2_decap_8 FILLER_6_32 ();
 sg13g2_decap_8 FILLER_6_39 ();
 sg13g2_decap_8 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_decap_8 FILLER_6_60 ();
 sg13g2_decap_8 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_74 ();
 sg13g2_decap_8 FILLER_6_81 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_decap_8 FILLER_6_95 ();
 sg13g2_decap_8 FILLER_6_102 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_decap_8 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_137 ();
 sg13g2_decap_8 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_158 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_decap_8 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_207 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_403 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_decap_8 FILLER_6_424 ();
 sg13g2_decap_8 FILLER_6_431 ();
 sg13g2_decap_8 FILLER_6_438 ();
 sg13g2_decap_8 FILLER_6_445 ();
 sg13g2_decap_8 FILLER_6_452 ();
 sg13g2_decap_8 FILLER_6_459 ();
 sg13g2_decap_8 FILLER_6_466 ();
 sg13g2_decap_8 FILLER_6_473 ();
 sg13g2_decap_8 FILLER_6_480 ();
 sg13g2_decap_8 FILLER_6_487 ();
 sg13g2_decap_8 FILLER_6_494 ();
 sg13g2_decap_8 FILLER_6_501 ();
 sg13g2_decap_8 FILLER_6_508 ();
 sg13g2_decap_8 FILLER_6_515 ();
 sg13g2_decap_8 FILLER_6_522 ();
 sg13g2_decap_8 FILLER_6_529 ();
 sg13g2_decap_8 FILLER_6_536 ();
 sg13g2_decap_8 FILLER_6_543 ();
 sg13g2_decap_8 FILLER_6_550 ();
 sg13g2_decap_8 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_564 ();
 sg13g2_decap_8 FILLER_6_571 ();
 sg13g2_decap_8 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_592 ();
 sg13g2_fill_2 FILLER_6_599 ();
 sg13g2_fill_1 FILLER_6_601 ();
 sg13g2_decap_8 FILLER_6_622 ();
 sg13g2_decap_8 FILLER_6_633 ();
 sg13g2_decap_4 FILLER_6_640 ();
 sg13g2_fill_1 FILLER_6_659 ();
 sg13g2_decap_8 FILLER_6_726 ();
 sg13g2_decap_4 FILLER_6_733 ();
 sg13g2_fill_2 FILLER_6_737 ();
 sg13g2_decap_8 FILLER_6_748 ();
 sg13g2_decap_8 FILLER_6_755 ();
 sg13g2_decap_8 FILLER_6_762 ();
 sg13g2_fill_2 FILLER_6_769 ();
 sg13g2_fill_1 FILLER_6_771 ();
 sg13g2_decap_8 FILLER_6_790 ();
 sg13g2_decap_8 FILLER_6_797 ();
 sg13g2_fill_1 FILLER_6_804 ();
 sg13g2_decap_4 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_829 ();
 sg13g2_decap_8 FILLER_6_836 ();
 sg13g2_fill_1 FILLER_6_843 ();
 sg13g2_decap_8 FILLER_6_853 ();
 sg13g2_fill_2 FILLER_6_860 ();
 sg13g2_fill_2 FILLER_6_867 ();
 sg13g2_fill_2 FILLER_6_892 ();
 sg13g2_fill_1 FILLER_6_894 ();
 sg13g2_decap_8 FILLER_6_900 ();
 sg13g2_fill_2 FILLER_6_907 ();
 sg13g2_decap_8 FILLER_6_925 ();
 sg13g2_decap_4 FILLER_6_932 ();
 sg13g2_decap_8 FILLER_6_952 ();
 sg13g2_decap_4 FILLER_6_959 ();
 sg13g2_fill_1 FILLER_6_963 ();
 sg13g2_decap_8 FILLER_6_980 ();
 sg13g2_fill_2 FILLER_6_987 ();
 sg13g2_fill_1 FILLER_6_998 ();
 sg13g2_fill_1 FILLER_6_1003 ();
 sg13g2_fill_2 FILLER_6_1009 ();
 sg13g2_decap_4 FILLER_6_1023 ();
 sg13g2_fill_2 FILLER_6_1027 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_fill_2 FILLER_7_595 ();
 sg13g2_fill_1 FILLER_7_660 ();
 sg13g2_decap_8 FILLER_7_682 ();
 sg13g2_fill_1 FILLER_7_693 ();
 sg13g2_decap_4 FILLER_7_698 ();
 sg13g2_decap_8 FILLER_7_711 ();
 sg13g2_fill_2 FILLER_7_718 ();
 sg13g2_fill_1 FILLER_7_720 ();
 sg13g2_decap_4 FILLER_7_725 ();
 sg13g2_fill_1 FILLER_7_729 ();
 sg13g2_decap_8 FILLER_7_762 ();
 sg13g2_decap_8 FILLER_7_769 ();
 sg13g2_decap_8 FILLER_7_776 ();
 sg13g2_decap_4 FILLER_7_783 ();
 sg13g2_fill_2 FILLER_7_787 ();
 sg13g2_decap_8 FILLER_7_792 ();
 sg13g2_decap_8 FILLER_7_799 ();
 sg13g2_decap_8 FILLER_7_806 ();
 sg13g2_decap_8 FILLER_7_813 ();
 sg13g2_fill_1 FILLER_7_820 ();
 sg13g2_decap_8 FILLER_7_825 ();
 sg13g2_decap_8 FILLER_7_832 ();
 sg13g2_decap_8 FILLER_7_839 ();
 sg13g2_decap_4 FILLER_7_846 ();
 sg13g2_fill_1 FILLER_7_850 ();
 sg13g2_decap_8 FILLER_7_855 ();
 sg13g2_decap_8 FILLER_7_862 ();
 sg13g2_decap_8 FILLER_7_869 ();
 sg13g2_decap_4 FILLER_7_876 ();
 sg13g2_decap_8 FILLER_7_884 ();
 sg13g2_decap_8 FILLER_7_891 ();
 sg13g2_decap_8 FILLER_7_898 ();
 sg13g2_decap_8 FILLER_7_905 ();
 sg13g2_decap_8 FILLER_7_912 ();
 sg13g2_decap_8 FILLER_7_919 ();
 sg13g2_decap_8 FILLER_7_926 ();
 sg13g2_decap_8 FILLER_7_933 ();
 sg13g2_decap_4 FILLER_7_940 ();
 sg13g2_decap_8 FILLER_7_948 ();
 sg13g2_decap_8 FILLER_7_955 ();
 sg13g2_decap_8 FILLER_7_962 ();
 sg13g2_decap_8 FILLER_7_969 ();
 sg13g2_decap_8 FILLER_7_976 ();
 sg13g2_decap_8 FILLER_7_983 ();
 sg13g2_decap_8 FILLER_7_990 ();
 sg13g2_fill_2 FILLER_7_997 ();
 sg13g2_fill_1 FILLER_7_999 ();
 sg13g2_decap_8 FILLER_7_1011 ();
 sg13g2_decap_8 FILLER_7_1018 ();
 sg13g2_decap_4 FILLER_7_1025 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_8 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_decap_8 FILLER_8_46 ();
 sg13g2_decap_8 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_8 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_decap_8 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_109 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_8 FILLER_8_137 ();
 sg13g2_decap_8 FILLER_8_144 ();
 sg13g2_decap_8 FILLER_8_151 ();
 sg13g2_decap_8 FILLER_8_158 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_decap_8 FILLER_8_193 ();
 sg13g2_decap_8 FILLER_8_200 ();
 sg13g2_decap_8 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_221 ();
 sg13g2_decap_8 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_235 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_270 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_8 FILLER_8_291 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_8 FILLER_8_424 ();
 sg13g2_decap_8 FILLER_8_431 ();
 sg13g2_decap_4 FILLER_8_438 ();
 sg13g2_decap_8 FILLER_8_446 ();
 sg13g2_decap_8 FILLER_8_453 ();
 sg13g2_decap_8 FILLER_8_460 ();
 sg13g2_decap_8 FILLER_8_467 ();
 sg13g2_decap_8 FILLER_8_474 ();
 sg13g2_decap_8 FILLER_8_481 ();
 sg13g2_decap_8 FILLER_8_488 ();
 sg13g2_decap_8 FILLER_8_495 ();
 sg13g2_decap_8 FILLER_8_502 ();
 sg13g2_decap_8 FILLER_8_509 ();
 sg13g2_decap_8 FILLER_8_516 ();
 sg13g2_decap_8 FILLER_8_523 ();
 sg13g2_decap_8 FILLER_8_530 ();
 sg13g2_decap_8 FILLER_8_537 ();
 sg13g2_decap_8 FILLER_8_544 ();
 sg13g2_decap_8 FILLER_8_551 ();
 sg13g2_decap_8 FILLER_8_558 ();
 sg13g2_decap_8 FILLER_8_565 ();
 sg13g2_decap_8 FILLER_8_572 ();
 sg13g2_decap_8 FILLER_8_579 ();
 sg13g2_decap_8 FILLER_8_586 ();
 sg13g2_fill_1 FILLER_8_593 ();
 sg13g2_decap_8 FILLER_8_598 ();
 sg13g2_decap_4 FILLER_8_605 ();
 sg13g2_fill_2 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_624 ();
 sg13g2_decap_8 FILLER_8_631 ();
 sg13g2_decap_8 FILLER_8_638 ();
 sg13g2_decap_8 FILLER_8_645 ();
 sg13g2_decap_4 FILLER_8_652 ();
 sg13g2_fill_1 FILLER_8_688 ();
 sg13g2_decap_8 FILLER_8_716 ();
 sg13g2_decap_8 FILLER_8_723 ();
 sg13g2_decap_4 FILLER_8_730 ();
 sg13g2_fill_2 FILLER_8_734 ();
 sg13g2_decap_8 FILLER_8_744 ();
 sg13g2_fill_2 FILLER_8_754 ();
 sg13g2_fill_1 FILLER_8_756 ();
 sg13g2_fill_2 FILLER_8_760 ();
 sg13g2_fill_1 FILLER_8_762 ();
 sg13g2_fill_2 FILLER_8_766 ();
 sg13g2_fill_1 FILLER_8_771 ();
 sg13g2_fill_1 FILLER_8_775 ();
 sg13g2_fill_1 FILLER_8_779 ();
 sg13g2_fill_1 FILLER_8_783 ();
 sg13g2_decap_8 FILLER_8_787 ();
 sg13g2_fill_1 FILLER_8_797 ();
 sg13g2_fill_1 FILLER_8_801 ();
 sg13g2_fill_1 FILLER_8_805 ();
 sg13g2_fill_1 FILLER_8_812 ();
 sg13g2_fill_2 FILLER_8_816 ();
 sg13g2_fill_1 FILLER_8_821 ();
 sg13g2_fill_1 FILLER_8_825 ();
 sg13g2_fill_2 FILLER_8_829 ();
 sg13g2_fill_1 FILLER_8_834 ();
 sg13g2_fill_1 FILLER_8_838 ();
 sg13g2_fill_1 FILLER_8_842 ();
 sg13g2_fill_2 FILLER_8_846 ();
 sg13g2_fill_1 FILLER_8_851 ();
 sg13g2_fill_1 FILLER_8_855 ();
 sg13g2_fill_2 FILLER_8_859 ();
 sg13g2_fill_1 FILLER_8_864 ();
 sg13g2_fill_1 FILLER_8_868 ();
 sg13g2_fill_2 FILLER_8_872 ();
 sg13g2_fill_1 FILLER_8_877 ();
 sg13g2_fill_1 FILLER_8_881 ();
 sg13g2_fill_1 FILLER_8_885 ();
 sg13g2_fill_2 FILLER_8_889 ();
 sg13g2_fill_1 FILLER_8_894 ();
 sg13g2_fill_1 FILLER_8_898 ();
 sg13g2_fill_1 FILLER_8_902 ();
 sg13g2_fill_1 FILLER_8_906 ();
 sg13g2_fill_1 FILLER_8_910 ();
 sg13g2_fill_2 FILLER_8_914 ();
 sg13g2_fill_1 FILLER_8_919 ();
 sg13g2_fill_1 FILLER_8_923 ();
 sg13g2_fill_1 FILLER_8_927 ();
 sg13g2_fill_1 FILLER_8_931 ();
 sg13g2_fill_1 FILLER_8_935 ();
 sg13g2_fill_1 FILLER_8_939 ();
 sg13g2_fill_1 FILLER_8_943 ();
 sg13g2_fill_2 FILLER_8_947 ();
 sg13g2_fill_1 FILLER_8_952 ();
 sg13g2_fill_1 FILLER_8_956 ();
 sg13g2_fill_1 FILLER_8_960 ();
 sg13g2_fill_1 FILLER_8_964 ();
 sg13g2_fill_1 FILLER_8_968 ();
 sg13g2_fill_2 FILLER_8_972 ();
 sg13g2_fill_2 FILLER_8_977 ();
 sg13g2_fill_1 FILLER_8_985 ();
 sg13g2_fill_1 FILLER_8_989 ();
 sg13g2_fill_2 FILLER_8_993 ();
 sg13g2_decap_4 FILLER_8_998 ();
 sg13g2_fill_1 FILLER_8_1002 ();
 sg13g2_fill_2 FILLER_8_1006 ();
 sg13g2_fill_1 FILLER_8_1014 ();
 sg13g2_decap_4 FILLER_8_1024 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_18 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_39 ();
 sg13g2_decap_8 FILLER_9_46 ();
 sg13g2_decap_8 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_67 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_109 ();
 sg13g2_decap_8 FILLER_9_116 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_decap_8 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_172 ();
 sg13g2_decap_8 FILLER_9_179 ();
 sg13g2_decap_8 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_221 ();
 sg13g2_decap_8 FILLER_9_228 ();
 sg13g2_decap_8 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_8 FILLER_9_424 ();
 sg13g2_decap_8 FILLER_9_431 ();
 sg13g2_decap_8 FILLER_9_438 ();
 sg13g2_decap_8 FILLER_9_445 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_8 FILLER_9_466 ();
 sg13g2_decap_8 FILLER_9_473 ();
 sg13g2_decap_8 FILLER_9_480 ();
 sg13g2_decap_8 FILLER_9_487 ();
 sg13g2_decap_8 FILLER_9_494 ();
 sg13g2_decap_8 FILLER_9_501 ();
 sg13g2_decap_8 FILLER_9_508 ();
 sg13g2_decap_8 FILLER_9_515 ();
 sg13g2_decap_8 FILLER_9_522 ();
 sg13g2_decap_8 FILLER_9_529 ();
 sg13g2_decap_8 FILLER_9_536 ();
 sg13g2_decap_8 FILLER_9_543 ();
 sg13g2_decap_8 FILLER_9_550 ();
 sg13g2_decap_8 FILLER_9_557 ();
 sg13g2_decap_8 FILLER_9_568 ();
 sg13g2_fill_2 FILLER_9_575 ();
 sg13g2_fill_1 FILLER_9_577 ();
 sg13g2_decap_8 FILLER_9_605 ();
 sg13g2_decap_4 FILLER_9_612 ();
 sg13g2_fill_2 FILLER_9_616 ();
 sg13g2_decap_4 FILLER_9_623 ();
 sg13g2_fill_1 FILLER_9_627 ();
 sg13g2_fill_2 FILLER_9_659 ();
 sg13g2_decap_8 FILLER_9_677 ();
 sg13g2_decap_8 FILLER_9_684 ();
 sg13g2_decap_8 FILLER_9_691 ();
 sg13g2_decap_4 FILLER_9_698 ();
 sg13g2_fill_1 FILLER_9_702 ();
 sg13g2_fill_2 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_725 ();
 sg13g2_fill_1 FILLER_9_732 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_32 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_decap_8 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_8 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_decap_8 FILLER_10_424 ();
 sg13g2_decap_8 FILLER_10_431 ();
 sg13g2_decap_8 FILLER_10_438 ();
 sg13g2_decap_8 FILLER_10_445 ();
 sg13g2_decap_8 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_459 ();
 sg13g2_decap_8 FILLER_10_466 ();
 sg13g2_decap_8 FILLER_10_473 ();
 sg13g2_decap_8 FILLER_10_480 ();
 sg13g2_decap_8 FILLER_10_487 ();
 sg13g2_decap_8 FILLER_10_494 ();
 sg13g2_decap_8 FILLER_10_501 ();
 sg13g2_decap_8 FILLER_10_508 ();
 sg13g2_decap_8 FILLER_10_515 ();
 sg13g2_decap_8 FILLER_10_522 ();
 sg13g2_decap_8 FILLER_10_529 ();
 sg13g2_decap_8 FILLER_10_536 ();
 sg13g2_decap_8 FILLER_10_543 ();
 sg13g2_decap_8 FILLER_10_550 ();
 sg13g2_fill_2 FILLER_10_593 ();
 sg13g2_fill_1 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_612 ();
 sg13g2_decap_8 FILLER_10_619 ();
 sg13g2_fill_1 FILLER_10_626 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_8 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_decap_4 FILLER_10_662 ();
 sg13g2_decap_8 FILLER_10_678 ();
 sg13g2_decap_8 FILLER_10_685 ();
 sg13g2_fill_2 FILLER_10_692 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_4 FILLER_10_728 ();
 sg13g2_fill_1 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_18 ();
 sg13g2_decap_8 FILLER_11_25 ();
 sg13g2_decap_8 FILLER_11_32 ();
 sg13g2_decap_8 FILLER_11_39 ();
 sg13g2_decap_8 FILLER_11_46 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_decap_8 FILLER_11_60 ();
 sg13g2_decap_8 FILLER_11_67 ();
 sg13g2_decap_8 FILLER_11_74 ();
 sg13g2_decap_8 FILLER_11_81 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_decap_8 FILLER_11_95 ();
 sg13g2_decap_8 FILLER_11_102 ();
 sg13g2_decap_8 FILLER_11_109 ();
 sg13g2_decap_8 FILLER_11_116 ();
 sg13g2_decap_8 FILLER_11_123 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_137 ();
 sg13g2_decap_8 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_186 ();
 sg13g2_decap_8 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_decap_8 FILLER_11_249 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_decap_8 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_decap_8 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_decap_8 FILLER_11_431 ();
 sg13g2_decap_8 FILLER_11_438 ();
 sg13g2_decap_8 FILLER_11_445 ();
 sg13g2_decap_8 FILLER_11_452 ();
 sg13g2_decap_8 FILLER_11_459 ();
 sg13g2_decap_8 FILLER_11_466 ();
 sg13g2_decap_8 FILLER_11_473 ();
 sg13g2_decap_8 FILLER_11_480 ();
 sg13g2_decap_8 FILLER_11_487 ();
 sg13g2_decap_8 FILLER_11_494 ();
 sg13g2_decap_8 FILLER_11_501 ();
 sg13g2_decap_8 FILLER_11_508 ();
 sg13g2_decap_8 FILLER_11_515 ();
 sg13g2_decap_8 FILLER_11_522 ();
 sg13g2_decap_8 FILLER_11_529 ();
 sg13g2_decap_8 FILLER_11_536 ();
 sg13g2_decap_8 FILLER_11_543 ();
 sg13g2_decap_4 FILLER_11_550 ();
 sg13g2_fill_1 FILLER_11_554 ();
 sg13g2_fill_1 FILLER_11_564 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_4 FILLER_11_581 ();
 sg13g2_fill_2 FILLER_11_585 ();
 sg13g2_fill_1 FILLER_11_626 ();
 sg13g2_decap_8 FILLER_11_647 ();
 sg13g2_decap_4 FILLER_11_654 ();
 sg13g2_fill_1 FILLER_11_658 ();
 sg13g2_decap_4 FILLER_11_694 ();
 sg13g2_decap_8 FILLER_11_724 ();
 sg13g2_decap_8 FILLER_11_731 ();
 sg13g2_fill_1 FILLER_11_738 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_32 ();
 sg13g2_decap_8 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_53 ();
 sg13g2_decap_8 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_67 ();
 sg13g2_decap_8 FILLER_12_74 ();
 sg13g2_decap_8 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_95 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_decap_8 FILLER_12_109 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_decap_8 FILLER_12_130 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_decap_8 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_8 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_410 ();
 sg13g2_decap_8 FILLER_12_416 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_8 FILLER_12_430 ();
 sg13g2_decap_8 FILLER_12_437 ();
 sg13g2_decap_8 FILLER_12_444 ();
 sg13g2_decap_8 FILLER_12_451 ();
 sg13g2_decap_8 FILLER_12_458 ();
 sg13g2_decap_8 FILLER_12_465 ();
 sg13g2_decap_8 FILLER_12_472 ();
 sg13g2_decap_8 FILLER_12_479 ();
 sg13g2_decap_8 FILLER_12_486 ();
 sg13g2_decap_8 FILLER_12_493 ();
 sg13g2_decap_8 FILLER_12_500 ();
 sg13g2_decap_8 FILLER_12_507 ();
 sg13g2_decap_8 FILLER_12_514 ();
 sg13g2_decap_8 FILLER_12_521 ();
 sg13g2_decap_8 FILLER_12_528 ();
 sg13g2_decap_8 FILLER_12_535 ();
 sg13g2_decap_8 FILLER_12_542 ();
 sg13g2_decap_8 FILLER_12_549 ();
 sg13g2_decap_4 FILLER_12_556 ();
 sg13g2_decap_8 FILLER_12_575 ();
 sg13g2_decap_8 FILLER_12_582 ();
 sg13g2_decap_4 FILLER_12_589 ();
 sg13g2_fill_1 FILLER_12_593 ();
 sg13g2_decap_4 FILLER_12_611 ();
 sg13g2_fill_2 FILLER_12_615 ();
 sg13g2_decap_8 FILLER_12_626 ();
 sg13g2_decap_8 FILLER_12_633 ();
 sg13g2_fill_1 FILLER_12_671 ();
 sg13g2_fill_2 FILLER_12_676 ();
 sg13g2_decap_8 FILLER_12_690 ();
 sg13g2_decap_4 FILLER_12_697 ();
 sg13g2_fill_1 FILLER_12_701 ();
 sg13g2_fill_1 FILLER_12_706 ();
 sg13g2_decap_8 FILLER_12_723 ();
 sg13g2_decap_8 FILLER_12_730 ();
 sg13g2_fill_2 FILLER_12_737 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_25 ();
 sg13g2_decap_8 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_39 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_decap_8 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_decap_8 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_109 ();
 sg13g2_decap_8 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_144 ();
 sg13g2_decap_8 FILLER_13_151 ();
 sg13g2_decap_8 FILLER_13_158 ();
 sg13g2_decap_8 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_decap_8 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_13_424 ();
 sg13g2_decap_8 FILLER_13_431 ();
 sg13g2_decap_8 FILLER_13_438 ();
 sg13g2_decap_8 FILLER_13_445 ();
 sg13g2_decap_4 FILLER_13_452 ();
 sg13g2_fill_1 FILLER_13_456 ();
 sg13g2_fill_2 FILLER_13_461 ();
 sg13g2_fill_1 FILLER_13_467 ();
 sg13g2_decap_8 FILLER_13_472 ();
 sg13g2_decap_8 FILLER_13_479 ();
 sg13g2_decap_8 FILLER_13_486 ();
 sg13g2_decap_8 FILLER_13_493 ();
 sg13g2_decap_8 FILLER_13_500 ();
 sg13g2_decap_4 FILLER_13_511 ();
 sg13g2_fill_2 FILLER_13_528 ();
 sg13g2_fill_1 FILLER_13_530 ();
 sg13g2_decap_8 FILLER_13_558 ();
 sg13g2_fill_2 FILLER_13_592 ();
 sg13g2_fill_1 FILLER_13_594 ();
 sg13g2_decap_8 FILLER_13_600 ();
 sg13g2_decap_8 FILLER_13_638 ();
 sg13g2_decap_4 FILLER_13_649 ();
 sg13g2_fill_1 FILLER_13_653 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_fill_2 FILLER_13_665 ();
 sg13g2_fill_2 FILLER_13_694 ();
 sg13g2_fill_1 FILLER_13_696 ();
 sg13g2_decap_8 FILLER_13_729 ();
 sg13g2_fill_2 FILLER_13_736 ();
 sg13g2_fill_1 FILLER_13_738 ();
 sg13g2_decap_8 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_46 ();
 sg13g2_decap_8 FILLER_14_53 ();
 sg13g2_decap_8 FILLER_14_60 ();
 sg13g2_decap_8 FILLER_14_67 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_decap_8 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_88 ();
 sg13g2_decap_8 FILLER_14_95 ();
 sg13g2_decap_8 FILLER_14_102 ();
 sg13g2_decap_8 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_decap_8 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_8 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_235 ();
 sg13g2_decap_8 FILLER_14_242 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_decap_8 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_8 FILLER_14_403 ();
 sg13g2_decap_8 FILLER_14_410 ();
 sg13g2_decap_8 FILLER_14_417 ();
 sg13g2_decap_8 FILLER_14_424 ();
 sg13g2_decap_8 FILLER_14_431 ();
 sg13g2_decap_8 FILLER_14_438 ();
 sg13g2_decap_8 FILLER_14_445 ();
 sg13g2_decap_4 FILLER_14_452 ();
 sg13g2_fill_2 FILLER_14_456 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_4 FILLER_14_504 ();
 sg13g2_fill_1 FILLER_14_508 ();
 sg13g2_decap_4 FILLER_14_557 ();
 sg13g2_decap_4 FILLER_14_566 ();
 sg13g2_decap_4 FILLER_14_574 ();
 sg13g2_fill_2 FILLER_14_578 ();
 sg13g2_decap_8 FILLER_14_611 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_fill_1 FILLER_14_637 ();
 sg13g2_fill_2 FILLER_14_665 ();
 sg13g2_fill_1 FILLER_14_667 ();
 sg13g2_fill_2 FILLER_14_677 ();
 sg13g2_fill_1 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_685 ();
 sg13g2_decap_8 FILLER_14_692 ();
 sg13g2_decap_4 FILLER_14_699 ();
 sg13g2_fill_2 FILLER_14_703 ();
 sg13g2_fill_2 FILLER_14_710 ();
 sg13g2_decap_8 FILLER_14_725 ();
 sg13g2_decap_8 FILLER_14_732 ();
 sg13g2_decap_8 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_88 ();
 sg13g2_decap_8 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_130 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_decap_8 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_decap_8 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_249 ();
 sg13g2_decap_8 FILLER_15_256 ();
 sg13g2_decap_8 FILLER_15_263 ();
 sg13g2_decap_8 FILLER_15_270 ();
 sg13g2_decap_8 FILLER_15_277 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_8 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_305 ();
 sg13g2_decap_8 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_319 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_8 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_4 FILLER_15_452 ();
 sg13g2_fill_1 FILLER_15_456 ();
 sg13g2_decap_4 FILLER_15_477 ();
 sg13g2_decap_8 FILLER_15_489 ();
 sg13g2_decap_4 FILLER_15_496 ();
 sg13g2_fill_2 FILLER_15_504 ();
 sg13g2_fill_1 FILLER_15_506 ();
 sg13g2_decap_4 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_550 ();
 sg13g2_decap_8 FILLER_15_557 ();
 sg13g2_fill_2 FILLER_15_564 ();
 sg13g2_fill_1 FILLER_15_566 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_decap_4 FILLER_15_578 ();
 sg13g2_fill_2 FILLER_15_582 ();
 sg13g2_decap_4 FILLER_15_600 ();
 sg13g2_fill_1 FILLER_15_604 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_fill_2 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_4 FILLER_15_637 ();
 sg13g2_fill_2 FILLER_15_641 ();
 sg13g2_fill_2 FILLER_15_647 ();
 sg13g2_fill_2 FILLER_15_654 ();
 sg13g2_decap_8 FILLER_15_661 ();
 sg13g2_decap_8 FILLER_15_668 ();
 sg13g2_fill_2 FILLER_15_675 ();
 sg13g2_fill_1 FILLER_15_677 ();
 sg13g2_decap_8 FILLER_15_685 ();
 sg13g2_decap_8 FILLER_15_692 ();
 sg13g2_decap_8 FILLER_15_726 ();
 sg13g2_fill_2 FILLER_15_733 ();
 sg13g2_fill_1 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_11 ();
 sg13g2_decap_8 FILLER_16_18 ();
 sg13g2_decap_8 FILLER_16_25 ();
 sg13g2_decap_8 FILLER_16_32 ();
 sg13g2_decap_8 FILLER_16_39 ();
 sg13g2_decap_8 FILLER_16_46 ();
 sg13g2_decap_8 FILLER_16_53 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_67 ();
 sg13g2_decap_8 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_88 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_109 ();
 sg13g2_decap_8 FILLER_16_116 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_decap_8 FILLER_16_130 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_144 ();
 sg13g2_decap_8 FILLER_16_151 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_179 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_decap_8 FILLER_16_221 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_decap_8 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_277 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_312 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_8 FILLER_16_403 ();
 sg13g2_decap_8 FILLER_16_410 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_8 FILLER_16_424 ();
 sg13g2_fill_2 FILLER_16_435 ();
 sg13g2_decap_8 FILLER_16_450 ();
 sg13g2_decap_8 FILLER_16_457 ();
 sg13g2_decap_4 FILLER_16_464 ();
 sg13g2_fill_1 FILLER_16_468 ();
 sg13g2_decap_4 FILLER_16_474 ();
 sg13g2_fill_2 FILLER_16_478 ();
 sg13g2_decap_8 FILLER_16_516 ();
 sg13g2_decap_8 FILLER_16_523 ();
 sg13g2_decap_4 FILLER_16_530 ();
 sg13g2_fill_1 FILLER_16_534 ();
 sg13g2_fill_2 FILLER_16_589 ();
 sg13g2_fill_1 FILLER_16_591 ();
 sg13g2_decap_8 FILLER_16_639 ();
 sg13g2_fill_1 FILLER_16_646 ();
 sg13g2_decap_8 FILLER_16_662 ();
 sg13g2_decap_8 FILLER_16_669 ();
 sg13g2_decap_8 FILLER_16_684 ();
 sg13g2_decap_8 FILLER_16_691 ();
 sg13g2_decap_4 FILLER_16_698 ();
 sg13g2_fill_2 FILLER_16_702 ();
 sg13g2_fill_2 FILLER_16_708 ();
 sg13g2_decap_8 FILLER_16_717 ();
 sg13g2_decap_4 FILLER_16_724 ();
 sg13g2_fill_2 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_4 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_431 ();
 sg13g2_fill_2 FILLER_17_468 ();
 sg13g2_fill_1 FILLER_17_470 ();
 sg13g2_fill_2 FILLER_17_498 ();
 sg13g2_fill_1 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_550 ();
 sg13g2_fill_2 FILLER_17_557 ();
 sg13g2_fill_1 FILLER_17_559 ();
 sg13g2_fill_1 FILLER_17_565 ();
 sg13g2_decap_8 FILLER_17_570 ();
 sg13g2_fill_2 FILLER_17_577 ();
 sg13g2_fill_1 FILLER_17_579 ();
 sg13g2_fill_2 FILLER_17_589 ();
 sg13g2_decap_4 FILLER_17_596 ();
 sg13g2_fill_1 FILLER_17_600 ();
 sg13g2_decap_8 FILLER_17_606 ();
 sg13g2_decap_8 FILLER_17_613 ();
 sg13g2_decap_4 FILLER_17_620 ();
 sg13g2_fill_1 FILLER_17_624 ();
 sg13g2_decap_8 FILLER_17_718 ();
 sg13g2_decap_8 FILLER_17_725 ();
 sg13g2_decap_4 FILLER_17_732 ();
 sg13g2_decap_8 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_25 ();
 sg13g2_decap_8 FILLER_18_32 ();
 sg13g2_decap_8 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_decap_8 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_decap_8 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_186 ();
 sg13g2_decap_8 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_4 FILLER_18_375 ();
 sg13g2_fill_2 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_4 FILLER_18_434 ();
 sg13g2_fill_2 FILLER_18_438 ();
 sg13g2_decap_8 FILLER_18_447 ();
 sg13g2_fill_1 FILLER_18_454 ();
 sg13g2_decap_4 FILLER_18_459 ();
 sg13g2_fill_2 FILLER_18_463 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_4 FILLER_18_497 ();
 sg13g2_fill_2 FILLER_18_501 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_fill_1 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_544 ();
 sg13g2_fill_2 FILLER_18_551 ();
 sg13g2_decap_4 FILLER_18_580 ();
 sg13g2_fill_2 FILLER_18_604 ();
 sg13g2_decap_8 FILLER_18_611 ();
 sg13g2_fill_2 FILLER_18_618 ();
 sg13g2_decap_8 FILLER_18_647 ();
 sg13g2_decap_4 FILLER_18_654 ();
 sg13g2_fill_1 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_668 ();
 sg13g2_fill_2 FILLER_18_684 ();
 sg13g2_fill_1 FILLER_18_686 ();
 sg13g2_fill_1 FILLER_18_691 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_fill_2 FILLER_18_756 ();
 sg13g2_fill_1 FILLER_18_761 ();
 sg13g2_fill_1 FILLER_18_765 ();
 sg13g2_fill_1 FILLER_18_769 ();
 sg13g2_fill_2 FILLER_18_773 ();
 sg13g2_fill_1 FILLER_18_775 ();
 sg13g2_fill_2 FILLER_18_779 ();
 sg13g2_fill_1 FILLER_18_784 ();
 sg13g2_fill_1 FILLER_18_788 ();
 sg13g2_fill_1 FILLER_18_792 ();
 sg13g2_fill_2 FILLER_18_796 ();
 sg13g2_fill_1 FILLER_18_801 ();
 sg13g2_fill_1 FILLER_18_805 ();
 sg13g2_fill_1 FILLER_18_809 ();
 sg13g2_fill_1 FILLER_18_813 ();
 sg13g2_fill_1 FILLER_18_817 ();
 sg13g2_fill_2 FILLER_18_821 ();
 sg13g2_fill_1 FILLER_18_826 ();
 sg13g2_fill_1 FILLER_18_830 ();
 sg13g2_fill_1 FILLER_18_834 ();
 sg13g2_fill_1 FILLER_18_838 ();
 sg13g2_fill_2 FILLER_18_842 ();
 sg13g2_fill_1 FILLER_18_847 ();
 sg13g2_fill_1 FILLER_18_851 ();
 sg13g2_fill_1 FILLER_18_855 ();
 sg13g2_fill_1 FILLER_18_859 ();
 sg13g2_fill_2 FILLER_18_909 ();
 sg13g2_fill_1 FILLER_18_914 ();
 sg13g2_fill_1 FILLER_18_918 ();
 sg13g2_fill_1 FILLER_18_922 ();
 sg13g2_fill_1 FILLER_18_926 ();
 sg13g2_fill_1 FILLER_18_930 ();
 sg13g2_fill_2 FILLER_18_934 ();
 sg13g2_fill_1 FILLER_18_939 ();
 sg13g2_fill_1 FILLER_18_943 ();
 sg13g2_fill_1 FILLER_18_947 ();
 sg13g2_fill_1 FILLER_18_951 ();
 sg13g2_fill_2 FILLER_18_955 ();
 sg13g2_fill_1 FILLER_18_960 ();
 sg13g2_fill_1 FILLER_18_964 ();
 sg13g2_fill_1 FILLER_18_985 ();
 sg13g2_fill_1 FILLER_18_1028 ();
 sg13g2_decap_8 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_46 ();
 sg13g2_decap_8 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_60 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_decap_8 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_88 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_130 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_decap_8 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_decap_8 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_8 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_decap_4 FILLER_19_410 ();
 sg13g2_fill_2 FILLER_19_414 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_4 FILLER_19_427 ();
 sg13g2_fill_2 FILLER_19_431 ();
 sg13g2_fill_2 FILLER_19_446 ();
 sg13g2_decap_8 FILLER_19_452 ();
 sg13g2_decap_8 FILLER_19_459 ();
 sg13g2_fill_2 FILLER_19_466 ();
 sg13g2_decap_8 FILLER_19_492 ();
 sg13g2_decap_4 FILLER_19_499 ();
 sg13g2_fill_2 FILLER_19_503 ();
 sg13g2_fill_2 FILLER_19_522 ();
 sg13g2_decap_8 FILLER_19_545 ();
 sg13g2_decap_4 FILLER_19_552 ();
 sg13g2_fill_2 FILLER_19_556 ();
 sg13g2_decap_4 FILLER_19_562 ();
 sg13g2_decap_8 FILLER_19_578 ();
 sg13g2_decap_4 FILLER_19_585 ();
 sg13g2_fill_2 FILLER_19_589 ();
 sg13g2_fill_2 FILLER_19_622 ();
 sg13g2_decap_4 FILLER_19_647 ();
 sg13g2_fill_2 FILLER_19_651 ();
 sg13g2_fill_1 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_668 ();
 sg13g2_decap_4 FILLER_19_675 ();
 sg13g2_fill_1 FILLER_19_710 ();
 sg13g2_fill_1 FILLER_19_747 ();
 sg13g2_decap_8 FILLER_19_761 ();
 sg13g2_fill_2 FILLER_19_768 ();
 sg13g2_decap_8 FILLER_19_785 ();
 sg13g2_decap_8 FILLER_19_792 ();
 sg13g2_fill_2 FILLER_19_799 ();
 sg13g2_fill_1 FILLER_19_801 ();
 sg13g2_decap_8 FILLER_19_810 ();
 sg13g2_decap_8 FILLER_19_817 ();
 sg13g2_fill_2 FILLER_19_824 ();
 sg13g2_fill_1 FILLER_19_826 ();
 sg13g2_decap_4 FILLER_19_854 ();
 sg13g2_fill_2 FILLER_19_858 ();
 sg13g2_fill_1 FILLER_19_863 ();
 sg13g2_fill_2 FILLER_19_867 ();
 sg13g2_fill_1 FILLER_19_883 ();
 sg13g2_decap_4 FILLER_19_888 ();
 sg13g2_fill_1 FILLER_19_892 ();
 sg13g2_decap_8 FILLER_19_900 ();
 sg13g2_fill_2 FILLER_19_907 ();
 sg13g2_fill_1 FILLER_19_909 ();
 sg13g2_decap_8 FILLER_19_922 ();
 sg13g2_decap_8 FILLER_19_929 ();
 sg13g2_fill_1 FILLER_19_936 ();
 sg13g2_decap_8 FILLER_19_947 ();
 sg13g2_decap_8 FILLER_19_954 ();
 sg13g2_fill_1 FILLER_19_994 ();
 sg13g2_fill_1 FILLER_19_1028 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_39 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_102 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_decap_8 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_8 FILLER_20_403 ();
 sg13g2_decap_8 FILLER_20_410 ();
 sg13g2_decap_8 FILLER_20_417 ();
 sg13g2_decap_8 FILLER_20_424 ();
 sg13g2_decap_8 FILLER_20_431 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_4 FILLER_20_476 ();
 sg13g2_fill_2 FILLER_20_480 ();
 sg13g2_fill_2 FILLER_20_509 ();
 sg13g2_fill_1 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_578 ();
 sg13g2_fill_2 FILLER_20_615 ();
 sg13g2_decap_4 FILLER_20_641 ();
 sg13g2_fill_2 FILLER_20_676 ();
 sg13g2_fill_1 FILLER_20_687 ();
 sg13g2_fill_2 FILLER_20_697 ();
 sg13g2_fill_1 FILLER_20_699 ();
 sg13g2_decap_4 FILLER_20_735 ();
 sg13g2_fill_1 FILLER_20_739 ();
 sg13g2_decap_4 FILLER_20_747 ();
 sg13g2_fill_1 FILLER_20_751 ();
 sg13g2_fill_2 FILLER_20_779 ();
 sg13g2_fill_1 FILLER_20_781 ();
 sg13g2_decap_4 FILLER_20_841 ();
 sg13g2_fill_1 FILLER_20_907 ();
 sg13g2_decap_8 FILLER_20_948 ();
 sg13g2_decap_8 FILLER_20_955 ();
 sg13g2_decap_8 FILLER_20_975 ();
 sg13g2_decap_8 FILLER_20_982 ();
 sg13g2_fill_2 FILLER_20_989 ();
 sg13g2_decap_8 FILLER_20_1012 ();
 sg13g2_decap_8 FILLER_20_1019 ();
 sg13g2_fill_2 FILLER_20_1026 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_32 ();
 sg13g2_decap_8 FILLER_21_39 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_decap_8 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_decap_8 FILLER_21_81 ();
 sg13g2_decap_8 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_decap_8 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_179 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_decap_8 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_221 ();
 sg13g2_decap_8 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_decap_8 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_8 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_417 ();
 sg13g2_decap_8 FILLER_21_424 ();
 sg13g2_decap_8 FILLER_21_431 ();
 sg13g2_decap_8 FILLER_21_438 ();
 sg13g2_fill_2 FILLER_21_445 ();
 sg13g2_decap_8 FILLER_21_451 ();
 sg13g2_fill_2 FILLER_21_458 ();
 sg13g2_decap_8 FILLER_21_468 ();
 sg13g2_decap_8 FILLER_21_475 ();
 sg13g2_fill_2 FILLER_21_482 ();
 sg13g2_fill_1 FILLER_21_484 ();
 sg13g2_fill_2 FILLER_21_521 ();
 sg13g2_fill_1 FILLER_21_523 ();
 sg13g2_fill_1 FILLER_21_541 ();
 sg13g2_decap_8 FILLER_21_551 ();
 sg13g2_fill_1 FILLER_21_558 ();
 sg13g2_fill_2 FILLER_21_617 ();
 sg13g2_decap_8 FILLER_21_636 ();
 sg13g2_decap_8 FILLER_21_643 ();
 sg13g2_fill_2 FILLER_21_650 ();
 sg13g2_fill_1 FILLER_21_652 ();
 sg13g2_fill_1 FILLER_21_664 ();
 sg13g2_decap_8 FILLER_21_673 ();
 sg13g2_decap_4 FILLER_21_680 ();
 sg13g2_fill_2 FILLER_21_684 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_fill_1 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_717 ();
 sg13g2_decap_8 FILLER_21_724 ();
 sg13g2_decap_8 FILLER_21_731 ();
 sg13g2_decap_4 FILLER_21_738 ();
 sg13g2_decap_8 FILLER_21_762 ();
 sg13g2_fill_2 FILLER_21_769 ();
 sg13g2_fill_1 FILLER_21_771 ();
 sg13g2_fill_2 FILLER_21_785 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_4 FILLER_21_798 ();
 sg13g2_fill_2 FILLER_21_802 ();
 sg13g2_decap_4 FILLER_21_817 ();
 sg13g2_fill_2 FILLER_21_821 ();
 sg13g2_fill_1 FILLER_21_831 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_fill_1 FILLER_21_847 ();
 sg13g2_fill_2 FILLER_21_855 ();
 sg13g2_decap_4 FILLER_21_866 ();
 sg13g2_fill_2 FILLER_21_870 ();
 sg13g2_decap_8 FILLER_21_885 ();
 sg13g2_fill_1 FILLER_21_892 ();
 sg13g2_fill_2 FILLER_21_897 ();
 sg13g2_decap_8 FILLER_21_903 ();
 sg13g2_decap_8 FILLER_21_910 ();
 sg13g2_decap_8 FILLER_21_917 ();
 sg13g2_decap_4 FILLER_21_924 ();
 sg13g2_fill_1 FILLER_21_928 ();
 sg13g2_decap_8 FILLER_21_983 ();
 sg13g2_decap_8 FILLER_22_4 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_18 ();
 sg13g2_decap_8 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_32 ();
 sg13g2_decap_8 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_46 ();
 sg13g2_decap_8 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_60 ();
 sg13g2_decap_8 FILLER_22_67 ();
 sg13g2_decap_8 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_123 ();
 sg13g2_decap_8 FILLER_22_130 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_200 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_decap_8 FILLER_22_424 ();
 sg13g2_decap_8 FILLER_22_431 ();
 sg13g2_decap_8 FILLER_22_438 ();
 sg13g2_decap_8 FILLER_22_445 ();
 sg13g2_fill_2 FILLER_22_452 ();
 sg13g2_fill_1 FILLER_22_486 ();
 sg13g2_decap_8 FILLER_22_503 ();
 sg13g2_decap_8 FILLER_22_510 ();
 sg13g2_fill_2 FILLER_22_517 ();
 sg13g2_fill_2 FILLER_22_550 ();
 sg13g2_fill_1 FILLER_22_552 ();
 sg13g2_fill_2 FILLER_22_558 ();
 sg13g2_fill_2 FILLER_22_565 ();
 sg13g2_fill_1 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_573 ();
 sg13g2_decap_8 FILLER_22_580 ();
 sg13g2_decap_4 FILLER_22_587 ();
 sg13g2_fill_1 FILLER_22_591 ();
 sg13g2_fill_1 FILLER_22_600 ();
 sg13g2_decap_8 FILLER_22_612 ();
 sg13g2_decap_8 FILLER_22_619 ();
 sg13g2_fill_1 FILLER_22_626 ();
 sg13g2_fill_2 FILLER_22_654 ();
 sg13g2_fill_2 FILLER_22_673 ();
 sg13g2_fill_1 FILLER_22_675 ();
 sg13g2_decap_4 FILLER_22_715 ();
 sg13g2_fill_2 FILLER_22_773 ();
 sg13g2_fill_1 FILLER_22_775 ();
 sg13g2_fill_2 FILLER_22_781 ();
 sg13g2_decap_8 FILLER_22_810 ();
 sg13g2_fill_2 FILLER_22_817 ();
 sg13g2_fill_1 FILLER_22_819 ();
 sg13g2_fill_2 FILLER_22_833 ();
 sg13g2_fill_1 FILLER_22_835 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_decap_8 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_22_868 ();
 sg13g2_decap_8 FILLER_22_875 ();
 sg13g2_decap_4 FILLER_22_882 ();
 sg13g2_decap_4 FILLER_22_921 ();
 sg13g2_fill_1 FILLER_22_925 ();
 sg13g2_decap_8 FILLER_22_944 ();
 sg13g2_decap_8 FILLER_22_951 ();
 sg13g2_fill_1 FILLER_22_958 ();
 sg13g2_decap_8 FILLER_22_981 ();
 sg13g2_fill_2 FILLER_22_988 ();
 sg13g2_fill_1 FILLER_22_990 ();
 sg13g2_decap_8 FILLER_22_1018 ();
 sg13g2_decap_4 FILLER_22_1025 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_25 ();
 sg13g2_decap_8 FILLER_23_32 ();
 sg13g2_decap_8 FILLER_23_39 ();
 sg13g2_decap_8 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_60 ();
 sg13g2_decap_8 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_decap_8 FILLER_23_81 ();
 sg13g2_decap_8 FILLER_23_88 ();
 sg13g2_decap_8 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_decap_8 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_172 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_decap_8 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_8 FILLER_23_403 ();
 sg13g2_decap_8 FILLER_23_410 ();
 sg13g2_decap_8 FILLER_23_417 ();
 sg13g2_decap_8 FILLER_23_424 ();
 sg13g2_decap_8 FILLER_23_431 ();
 sg13g2_decap_8 FILLER_23_438 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_4 FILLER_23_483 ();
 sg13g2_fill_2 FILLER_23_500 ();
 sg13g2_fill_1 FILLER_23_502 ();
 sg13g2_decap_8 FILLER_23_507 ();
 sg13g2_decap_8 FILLER_23_514 ();
 sg13g2_fill_2 FILLER_23_521 ();
 sg13g2_fill_1 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_538 ();
 sg13g2_fill_1 FILLER_23_603 ();
 sg13g2_decap_8 FILLER_23_620 ();
 sg13g2_decap_4 FILLER_23_627 ();
 sg13g2_fill_2 FILLER_23_631 ();
 sg13g2_decap_8 FILLER_23_646 ();
 sg13g2_fill_2 FILLER_23_653 ();
 sg13g2_fill_1 FILLER_23_655 ();
 sg13g2_fill_2 FILLER_23_683 ();
 sg13g2_fill_2 FILLER_23_690 ();
 sg13g2_fill_1 FILLER_23_692 ();
 sg13g2_decap_8 FILLER_23_697 ();
 sg13g2_decap_8 FILLER_23_704 ();
 sg13g2_fill_2 FILLER_23_711 ();
 sg13g2_fill_2 FILLER_23_726 ();
 sg13g2_fill_1 FILLER_23_728 ();
 sg13g2_fill_2 FILLER_23_746 ();
 sg13g2_decap_8 FILLER_23_761 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_4 FILLER_23_784 ();
 sg13g2_decap_4 FILLER_23_792 ();
 sg13g2_fill_2 FILLER_23_801 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_fill_2 FILLER_23_819 ();
 sg13g2_fill_1 FILLER_23_821 ();
 sg13g2_decap_4 FILLER_23_857 ();
 sg13g2_decap_4 FILLER_23_868 ();
 sg13g2_fill_2 FILLER_23_903 ();
 sg13g2_fill_1 FILLER_23_905 ();
 sg13g2_decap_8 FILLER_23_911 ();
 sg13g2_decap_4 FILLER_23_918 ();
 sg13g2_decap_8 FILLER_23_925 ();
 sg13g2_fill_1 FILLER_23_932 ();
 sg13g2_decap_8 FILLER_23_940 ();
 sg13g2_decap_8 FILLER_23_947 ();
 sg13g2_decap_8 FILLER_23_954 ();
 sg13g2_fill_2 FILLER_23_961 ();
 sg13g2_decap_8 FILLER_23_978 ();
 sg13g2_decap_8 FILLER_23_985 ();
 sg13g2_fill_2 FILLER_23_1000 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_32 ();
 sg13g2_decap_8 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_53 ();
 sg13g2_decap_8 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_decap_8 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_172 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_417 ();
 sg13g2_decap_8 FILLER_24_424 ();
 sg13g2_fill_2 FILLER_24_431 ();
 sg13g2_decap_8 FILLER_24_437 ();
 sg13g2_decap_8 FILLER_24_444 ();
 sg13g2_fill_2 FILLER_24_451 ();
 sg13g2_fill_1 FILLER_24_453 ();
 sg13g2_decap_8 FILLER_24_479 ();
 sg13g2_decap_8 FILLER_24_486 ();
 sg13g2_fill_1 FILLER_24_497 ();
 sg13g2_decap_4 FILLER_24_525 ();
 sg13g2_fill_2 FILLER_24_529 ();
 sg13g2_decap_8 FILLER_24_542 ();
 sg13g2_decap_4 FILLER_24_549 ();
 sg13g2_fill_1 FILLER_24_553 ();
 sg13g2_fill_1 FILLER_24_558 ();
 sg13g2_decap_8 FILLER_24_566 ();
 sg13g2_fill_1 FILLER_24_573 ();
 sg13g2_fill_1 FILLER_24_582 ();
 sg13g2_fill_1 FILLER_24_605 ();
 sg13g2_fill_2 FILLER_24_660 ();
 sg13g2_fill_1 FILLER_24_666 ();
 sg13g2_decap_8 FILLER_24_698 ();
 sg13g2_fill_1 FILLER_24_710 ();
 sg13g2_fill_2 FILLER_24_716 ();
 sg13g2_fill_1 FILLER_24_737 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_839 ();
 sg13g2_decap_4 FILLER_24_846 ();
 sg13g2_fill_2 FILLER_24_881 ();
 sg13g2_fill_1 FILLER_24_883 ();
 sg13g2_fill_2 FILLER_24_893 ();
 sg13g2_fill_1 FILLER_24_895 ();
 sg13g2_decap_8 FILLER_24_912 ();
 sg13g2_fill_2 FILLER_24_919 ();
 sg13g2_fill_1 FILLER_24_921 ();
 sg13g2_decap_8 FILLER_24_926 ();
 sg13g2_fill_1 FILLER_24_933 ();
 sg13g2_decap_4 FILLER_24_950 ();
 sg13g2_fill_2 FILLER_24_954 ();
 sg13g2_decap_8 FILLER_24_987 ();
 sg13g2_decap_4 FILLER_24_994 ();
 sg13g2_fill_1 FILLER_24_998 ();
 sg13g2_decap_8 FILLER_24_1021 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_decap_8 FILLER_25_32 ();
 sg13g2_decap_8 FILLER_25_39 ();
 sg13g2_decap_8 FILLER_25_46 ();
 sg13g2_decap_8 FILLER_25_53 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_decap_8 FILLER_25_67 ();
 sg13g2_decap_8 FILLER_25_74 ();
 sg13g2_decap_8 FILLER_25_81 ();
 sg13g2_decap_8 FILLER_25_88 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_decap_8 FILLER_25_102 ();
 sg13g2_decap_8 FILLER_25_109 ();
 sg13g2_decap_8 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_179 ();
 sg13g2_decap_8 FILLER_25_186 ();
 sg13g2_decap_8 FILLER_25_193 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_decap_8 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_221 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_decap_8 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_242 ();
 sg13g2_decap_8 FILLER_25_249 ();
 sg13g2_decap_8 FILLER_25_256 ();
 sg13g2_decap_8 FILLER_25_263 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_284 ();
 sg13g2_decap_8 FILLER_25_291 ();
 sg13g2_decap_8 FILLER_25_298 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_8 FILLER_25_424 ();
 sg13g2_decap_8 FILLER_25_431 ();
 sg13g2_decap_4 FILLER_25_438 ();
 sg13g2_fill_1 FILLER_25_442 ();
 sg13g2_decap_8 FILLER_25_516 ();
 sg13g2_decap_8 FILLER_25_523 ();
 sg13g2_decap_8 FILLER_25_543 ();
 sg13g2_decap_8 FILLER_25_550 ();
 sg13g2_decap_8 FILLER_25_565 ();
 sg13g2_decap_4 FILLER_25_572 ();
 sg13g2_fill_2 FILLER_25_607 ();
 sg13g2_decap_8 FILLER_25_622 ();
 sg13g2_decap_4 FILLER_25_629 ();
 sg13g2_decap_8 FILLER_25_645 ();
 sg13g2_decap_8 FILLER_25_652 ();
 sg13g2_decap_8 FILLER_25_659 ();
 sg13g2_decap_4 FILLER_25_691 ();
 sg13g2_fill_2 FILLER_25_695 ();
 sg13g2_fill_1 FILLER_25_728 ();
 sg13g2_fill_1 FILLER_25_737 ();
 sg13g2_decap_4 FILLER_25_771 ();
 sg13g2_decap_8 FILLER_25_780 ();
 sg13g2_decap_4 FILLER_25_787 ();
 sg13g2_fill_2 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_fill_1 FILLER_25_826 ();
 sg13g2_fill_1 FILLER_25_854 ();
 sg13g2_fill_2 FILLER_25_859 ();
 sg13g2_decap_8 FILLER_25_874 ();
 sg13g2_decap_8 FILLER_25_881 ();
 sg13g2_decap_8 FILLER_25_908 ();
 sg13g2_fill_2 FILLER_25_915 ();
 sg13g2_fill_2 FILLER_25_976 ();
 sg13g2_fill_1 FILLER_25_978 ();
 sg13g2_decap_8 FILLER_25_988 ();
 sg13g2_fill_2 FILLER_25_995 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_decap_8 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_39 ();
 sg13g2_decap_8 FILLER_26_46 ();
 sg13g2_decap_8 FILLER_26_53 ();
 sg13g2_decap_8 FILLER_26_60 ();
 sg13g2_decap_8 FILLER_26_67 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_decap_8 FILLER_26_81 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_109 ();
 sg13g2_decap_8 FILLER_26_116 ();
 sg13g2_decap_8 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_284 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_326 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_8 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_410 ();
 sg13g2_decap_8 FILLER_26_417 ();
 sg13g2_decap_8 FILLER_26_424 ();
 sg13g2_decap_8 FILLER_26_431 ();
 sg13g2_decap_8 FILLER_26_438 ();
 sg13g2_decap_8 FILLER_26_445 ();
 sg13g2_decap_8 FILLER_26_472 ();
 sg13g2_decap_8 FILLER_26_479 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_fill_2 FILLER_26_511 ();
 sg13g2_decap_4 FILLER_26_625 ();
 sg13g2_fill_1 FILLER_26_629 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_fill_2 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_687 ();
 sg13g2_decap_8 FILLER_26_694 ();
 sg13g2_decap_4 FILLER_26_701 ();
 sg13g2_decap_8 FILLER_26_716 ();
 sg13g2_fill_1 FILLER_26_723 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_fill_2 FILLER_26_735 ();
 sg13g2_fill_1 FILLER_26_737 ();
 sg13g2_decap_8 FILLER_26_759 ();
 sg13g2_decap_4 FILLER_26_766 ();
 sg13g2_fill_2 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_787 ();
 sg13g2_decap_4 FILLER_26_794 ();
 sg13g2_fill_1 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_815 ();
 sg13g2_decap_8 FILLER_26_822 ();
 sg13g2_fill_2 FILLER_26_829 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_4 FILLER_26_854 ();
 sg13g2_fill_1 FILLER_26_858 ();
 sg13g2_decap_4 FILLER_26_890 ();
 sg13g2_decap_8 FILLER_26_921 ();
 sg13g2_decap_4 FILLER_26_928 ();
 sg13g2_fill_2 FILLER_26_932 ();
 sg13g2_fill_2 FILLER_26_942 ();
 sg13g2_fill_1 FILLER_26_944 ();
 sg13g2_decap_8 FILLER_26_949 ();
 sg13g2_decap_8 FILLER_26_956 ();
 sg13g2_decap_8 FILLER_26_963 ();
 sg13g2_fill_1 FILLER_26_970 ();
 sg13g2_decap_4 FILLER_26_1003 ();
 sg13g2_fill_1 FILLER_26_1007 ();
 sg13g2_decap_8 FILLER_26_1015 ();
 sg13g2_decap_8 FILLER_26_1022 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_fill_2 FILLER_27_448 ();
 sg13g2_fill_1 FILLER_27_450 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_fill_2 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_499 ();
 sg13g2_decap_4 FILLER_27_506 ();
 sg13g2_fill_1 FILLER_27_510 ();
 sg13g2_fill_2 FILLER_27_520 ();
 sg13g2_decap_4 FILLER_27_535 ();
 sg13g2_fill_2 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_545 ();
 sg13g2_decap_8 FILLER_27_552 ();
 sg13g2_fill_2 FILLER_27_564 ();
 sg13g2_fill_1 FILLER_27_566 ();
 sg13g2_decap_8 FILLER_27_571 ();
 sg13g2_decap_8 FILLER_27_578 ();
 sg13g2_decap_4 FILLER_27_585 ();
 sg13g2_fill_2 FILLER_27_606 ();
 sg13g2_decap_4 FILLER_27_635 ();
 sg13g2_fill_1 FILLER_27_639 ();
 sg13g2_decap_8 FILLER_27_657 ();
 sg13g2_decap_8 FILLER_27_664 ();
 sg13g2_fill_2 FILLER_27_714 ();
 sg13g2_decap_4 FILLER_27_733 ();
 sg13g2_fill_2 FILLER_27_839 ();
 sg13g2_fill_2 FILLER_27_859 ();
 sg13g2_decap_8 FILLER_27_878 ();
 sg13g2_fill_2 FILLER_27_885 ();
 sg13g2_fill_1 FILLER_27_887 ();
 sg13g2_fill_1 FILLER_27_897 ();
 sg13g2_decap_8 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_910 ();
 sg13g2_decap_4 FILLER_27_917 ();
 sg13g2_fill_2 FILLER_27_921 ();
 sg13g2_fill_1 FILLER_27_928 ();
 sg13g2_decap_8 FILLER_27_938 ();
 sg13g2_decap_8 FILLER_27_945 ();
 sg13g2_fill_1 FILLER_27_957 ();
 sg13g2_fill_1 FILLER_27_976 ();
 sg13g2_decap_8 FILLER_27_988 ();
 sg13g2_fill_2 FILLER_27_995 ();
 sg13g2_decap_4 FILLER_27_1002 ();
 sg13g2_fill_2 FILLER_27_1006 ();
 sg13g2_decap_8 FILLER_27_1012 ();
 sg13g2_decap_8 FILLER_27_1019 ();
 sg13g2_fill_2 FILLER_27_1026 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_decap_8 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_39 ();
 sg13g2_decap_8 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_53 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_decap_8 FILLER_28_74 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_95 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_109 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_decap_8 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_144 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_172 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_decap_8 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_decap_8 FILLER_28_270 ();
 sg13g2_decap_8 FILLER_28_277 ();
 sg13g2_decap_8 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_decap_8 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_319 ();
 sg13g2_decap_8 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_28_333 ();
 sg13g2_decap_8 FILLER_28_340 ();
 sg13g2_decap_8 FILLER_28_347 ();
 sg13g2_decap_8 FILLER_28_354 ();
 sg13g2_decap_8 FILLER_28_361 ();
 sg13g2_decap_8 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_396 ();
 sg13g2_decap_8 FILLER_28_403 ();
 sg13g2_decap_8 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_417 ();
 sg13g2_decap_8 FILLER_28_424 ();
 sg13g2_decap_8 FILLER_28_435 ();
 sg13g2_decap_8 FILLER_28_442 ();
 sg13g2_decap_4 FILLER_28_449 ();
 sg13g2_fill_2 FILLER_28_453 ();
 sg13g2_decap_8 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_496 ();
 sg13g2_decap_8 FILLER_28_503 ();
 sg13g2_decap_8 FILLER_28_529 ();
 sg13g2_decap_4 FILLER_28_536 ();
 sg13g2_decap_8 FILLER_28_549 ();
 sg13g2_decap_8 FILLER_28_556 ();
 sg13g2_fill_2 FILLER_28_590 ();
 sg13g2_fill_2 FILLER_28_609 ();
 sg13g2_fill_1 FILLER_28_611 ();
 sg13g2_fill_2 FILLER_28_617 ();
 sg13g2_decap_8 FILLER_28_624 ();
 sg13g2_decap_8 FILLER_28_631 ();
 sg13g2_decap_4 FILLER_28_638 ();
 sg13g2_fill_1 FILLER_28_642 ();
 sg13g2_fill_2 FILLER_28_648 ();
 sg13g2_decap_8 FILLER_28_659 ();
 sg13g2_fill_1 FILLER_28_666 ();
 sg13g2_decap_8 FILLER_28_694 ();
 sg13g2_fill_2 FILLER_28_701 ();
 sg13g2_fill_1 FILLER_28_703 ();
 sg13g2_decap_8 FILLER_28_762 ();
 sg13g2_decap_4 FILLER_28_769 ();
 sg13g2_fill_1 FILLER_28_773 ();
 sg13g2_decap_8 FILLER_28_783 ();
 sg13g2_decap_8 FILLER_28_790 ();
 sg13g2_decap_4 FILLER_28_797 ();
 sg13g2_decap_8 FILLER_28_811 ();
 sg13g2_decap_8 FILLER_28_818 ();
 sg13g2_fill_2 FILLER_28_825 ();
 sg13g2_fill_1 FILLER_28_827 ();
 sg13g2_fill_2 FILLER_28_916 ();
 sg13g2_fill_1 FILLER_28_918 ();
 sg13g2_decap_8 FILLER_28_973 ();
 sg13g2_decap_8 FILLER_28_988 ();
 sg13g2_decap_8 FILLER_28_995 ();
 sg13g2_decap_8 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_11 ();
 sg13g2_decap_8 FILLER_29_18 ();
 sg13g2_decap_8 FILLER_29_25 ();
 sg13g2_decap_8 FILLER_29_32 ();
 sg13g2_decap_8 FILLER_29_39 ();
 sg13g2_decap_8 FILLER_29_46 ();
 sg13g2_decap_8 FILLER_29_53 ();
 sg13g2_decap_8 FILLER_29_60 ();
 sg13g2_decap_8 FILLER_29_67 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_decap_8 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_95 ();
 sg13g2_decap_8 FILLER_29_102 ();
 sg13g2_decap_8 FILLER_29_109 ();
 sg13g2_decap_8 FILLER_29_116 ();
 sg13g2_decap_8 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_137 ();
 sg13g2_decap_8 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_151 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_165 ();
 sg13g2_decap_8 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_decap_8 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_200 ();
 sg13g2_decap_8 FILLER_29_207 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_decap_8 FILLER_29_249 ();
 sg13g2_decap_8 FILLER_29_256 ();
 sg13g2_decap_8 FILLER_29_263 ();
 sg13g2_decap_8 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_277 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_decap_8 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_305 ();
 sg13g2_decap_8 FILLER_29_312 ();
 sg13g2_decap_8 FILLER_29_319 ();
 sg13g2_decap_8 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_354 ();
 sg13g2_decap_8 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_368 ();
 sg13g2_decap_8 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_403 ();
 sg13g2_decap_4 FILLER_29_410 ();
 sg13g2_fill_1 FILLER_29_414 ();
 sg13g2_decap_8 FILLER_29_451 ();
 sg13g2_decap_4 FILLER_29_458 ();
 sg13g2_decap_8 FILLER_29_473 ();
 sg13g2_decap_8 FILLER_29_480 ();
 sg13g2_fill_1 FILLER_29_487 ();
 sg13g2_fill_2 FILLER_29_579 ();
 sg13g2_fill_2 FILLER_29_612 ();
 sg13g2_fill_1 FILLER_29_614 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_4 FILLER_29_664 ();
 sg13g2_fill_2 FILLER_29_677 ();
 sg13g2_decap_8 FILLER_29_684 ();
 sg13g2_decap_8 FILLER_29_691 ();
 sg13g2_decap_8 FILLER_29_698 ();
 sg13g2_decap_4 FILLER_29_705 ();
 sg13g2_fill_1 FILLER_29_718 ();
 sg13g2_decap_8 FILLER_29_744 ();
 sg13g2_decap_4 FILLER_29_751 ();
 sg13g2_fill_1 FILLER_29_755 ();
 sg13g2_decap_4 FILLER_29_761 ();
 sg13g2_fill_1 FILLER_29_765 ();
 sg13g2_decap_8 FILLER_29_771 ();
 sg13g2_decap_8 FILLER_29_778 ();
 sg13g2_decap_4 FILLER_29_785 ();
 sg13g2_fill_1 FILLER_29_789 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_fill_2 FILLER_29_833 ();
 sg13g2_fill_1 FILLER_29_835 ();
 sg13g2_decap_8 FILLER_29_844 ();
 sg13g2_decap_8 FILLER_29_851 ();
 sg13g2_fill_2 FILLER_29_858 ();
 sg13g2_fill_1 FILLER_29_860 ();
 sg13g2_decap_4 FILLER_29_885 ();
 sg13g2_fill_2 FILLER_29_889 ();
 sg13g2_decap_8 FILLER_29_903 ();
 sg13g2_decap_8 FILLER_29_910 ();
 sg13g2_decap_4 FILLER_29_917 ();
 sg13g2_fill_2 FILLER_29_921 ();
 sg13g2_decap_8 FILLER_29_934 ();
 sg13g2_decap_8 FILLER_29_941 ();
 sg13g2_fill_2 FILLER_29_948 ();
 sg13g2_decap_8 FILLER_29_969 ();
 sg13g2_fill_2 FILLER_29_976 ();
 sg13g2_fill_1 FILLER_29_978 ();
 sg13g2_decap_4 FILLER_29_1024 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_decap_8 FILLER_30_4 ();
 sg13g2_decap_8 FILLER_30_11 ();
 sg13g2_decap_8 FILLER_30_18 ();
 sg13g2_decap_8 FILLER_30_25 ();
 sg13g2_decap_8 FILLER_30_32 ();
 sg13g2_decap_8 FILLER_30_39 ();
 sg13g2_decap_8 FILLER_30_46 ();
 sg13g2_decap_8 FILLER_30_53 ();
 sg13g2_decap_8 FILLER_30_60 ();
 sg13g2_decap_8 FILLER_30_67 ();
 sg13g2_decap_8 FILLER_30_74 ();
 sg13g2_decap_8 FILLER_30_81 ();
 sg13g2_decap_8 FILLER_30_88 ();
 sg13g2_decap_8 FILLER_30_95 ();
 sg13g2_decap_8 FILLER_30_102 ();
 sg13g2_decap_8 FILLER_30_109 ();
 sg13g2_decap_8 FILLER_30_116 ();
 sg13g2_decap_8 FILLER_30_123 ();
 sg13g2_decap_8 FILLER_30_130 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_decap_8 FILLER_30_151 ();
 sg13g2_decap_8 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_186 ();
 sg13g2_decap_8 FILLER_30_193 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_decap_8 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_228 ();
 sg13g2_decap_8 FILLER_30_235 ();
 sg13g2_decap_8 FILLER_30_242 ();
 sg13g2_decap_8 FILLER_30_249 ();
 sg13g2_decap_8 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_263 ();
 sg13g2_decap_8 FILLER_30_270 ();
 sg13g2_decap_8 FILLER_30_277 ();
 sg13g2_decap_8 FILLER_30_284 ();
 sg13g2_decap_8 FILLER_30_291 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_8 FILLER_30_403 ();
 sg13g2_decap_8 FILLER_30_410 ();
 sg13g2_fill_2 FILLER_30_425 ();
 sg13g2_fill_1 FILLER_30_427 ();
 sg13g2_decap_8 FILLER_30_437 ();
 sg13g2_decap_8 FILLER_30_444 ();
 sg13g2_decap_8 FILLER_30_451 ();
 sg13g2_decap_4 FILLER_30_458 ();
 sg13g2_fill_1 FILLER_30_462 ();
 sg13g2_decap_4 FILLER_30_471 ();
 sg13g2_fill_2 FILLER_30_475 ();
 sg13g2_decap_8 FILLER_30_501 ();
 sg13g2_fill_2 FILLER_30_508 ();
 sg13g2_fill_2 FILLER_30_519 ();
 sg13g2_decap_8 FILLER_30_529 ();
 sg13g2_fill_2 FILLER_30_536 ();
 sg13g2_fill_1 FILLER_30_538 ();
 sg13g2_decap_4 FILLER_30_555 ();
 sg13g2_fill_2 FILLER_30_559 ();
 sg13g2_fill_2 FILLER_30_584 ();
 sg13g2_fill_1 FILLER_30_591 ();
 sg13g2_decap_8 FILLER_30_601 ();
 sg13g2_decap_4 FILLER_30_608 ();
 sg13g2_fill_2 FILLER_30_639 ();
 sg13g2_fill_1 FILLER_30_641 ();
 sg13g2_fill_2 FILLER_30_646 ();
 sg13g2_fill_1 FILLER_30_648 ();
 sg13g2_decap_8 FILLER_30_664 ();
 sg13g2_decap_4 FILLER_30_671 ();
 sg13g2_fill_1 FILLER_30_675 ();
 sg13g2_decap_8 FILLER_30_691 ();
 sg13g2_decap_4 FILLER_30_698 ();
 sg13g2_fill_2 FILLER_30_702 ();
 sg13g2_fill_1 FILLER_30_741 ();
 sg13g2_decap_4 FILLER_30_776 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_817 ();
 sg13g2_decap_4 FILLER_30_824 ();
 sg13g2_fill_1 FILLER_30_860 ();
 sg13g2_decap_8 FILLER_30_907 ();
 sg13g2_decap_8 FILLER_30_914 ();
 sg13g2_decap_4 FILLER_30_921 ();
 sg13g2_fill_2 FILLER_30_933 ();
 sg13g2_decap_8 FILLER_30_938 ();
 sg13g2_decap_8 FILLER_30_945 ();
 sg13g2_decap_8 FILLER_30_952 ();
 sg13g2_decap_8 FILLER_30_972 ();
 sg13g2_decap_4 FILLER_30_979 ();
 sg13g2_fill_1 FILLER_30_983 ();
 sg13g2_decap_8 FILLER_30_988 ();
 sg13g2_decap_8 FILLER_30_1015 ();
 sg13g2_decap_8 FILLER_30_1022 ();
 sg13g2_decap_8 FILLER_31_4 ();
 sg13g2_decap_8 FILLER_31_11 ();
 sg13g2_decap_8 FILLER_31_18 ();
 sg13g2_decap_8 FILLER_31_25 ();
 sg13g2_decap_8 FILLER_31_32 ();
 sg13g2_decap_8 FILLER_31_39 ();
 sg13g2_decap_8 FILLER_31_46 ();
 sg13g2_decap_8 FILLER_31_53 ();
 sg13g2_decap_8 FILLER_31_60 ();
 sg13g2_decap_8 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_74 ();
 sg13g2_decap_8 FILLER_31_81 ();
 sg13g2_decap_8 FILLER_31_88 ();
 sg13g2_decap_8 FILLER_31_95 ();
 sg13g2_decap_8 FILLER_31_102 ();
 sg13g2_decap_8 FILLER_31_109 ();
 sg13g2_decap_8 FILLER_31_116 ();
 sg13g2_decap_8 FILLER_31_123 ();
 sg13g2_decap_8 FILLER_31_130 ();
 sg13g2_decap_8 FILLER_31_137 ();
 sg13g2_decap_8 FILLER_31_144 ();
 sg13g2_decap_8 FILLER_31_151 ();
 sg13g2_decap_8 FILLER_31_158 ();
 sg13g2_decap_8 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_172 ();
 sg13g2_decap_8 FILLER_31_179 ();
 sg13g2_decap_8 FILLER_31_186 ();
 sg13g2_decap_8 FILLER_31_193 ();
 sg13g2_decap_8 FILLER_31_200 ();
 sg13g2_decap_8 FILLER_31_207 ();
 sg13g2_decap_8 FILLER_31_214 ();
 sg13g2_decap_8 FILLER_31_221 ();
 sg13g2_decap_8 FILLER_31_228 ();
 sg13g2_decap_8 FILLER_31_235 ();
 sg13g2_decap_8 FILLER_31_242 ();
 sg13g2_decap_8 FILLER_31_249 ();
 sg13g2_decap_8 FILLER_31_256 ();
 sg13g2_decap_8 FILLER_31_263 ();
 sg13g2_decap_8 FILLER_31_270 ();
 sg13g2_decap_8 FILLER_31_277 ();
 sg13g2_decap_8 FILLER_31_284 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_decap_8 FILLER_31_298 ();
 sg13g2_decap_8 FILLER_31_305 ();
 sg13g2_decap_8 FILLER_31_312 ();
 sg13g2_decap_8 FILLER_31_319 ();
 sg13g2_decap_8 FILLER_31_326 ();
 sg13g2_decap_8 FILLER_31_333 ();
 sg13g2_decap_8 FILLER_31_340 ();
 sg13g2_decap_8 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_354 ();
 sg13g2_decap_8 FILLER_31_361 ();
 sg13g2_decap_8 FILLER_31_368 ();
 sg13g2_decap_8 FILLER_31_375 ();
 sg13g2_decap_8 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_31_389 ();
 sg13g2_decap_8 FILLER_31_396 ();
 sg13g2_decap_8 FILLER_31_403 ();
 sg13g2_decap_8 FILLER_31_410 ();
 sg13g2_fill_2 FILLER_31_417 ();
 sg13g2_fill_2 FILLER_31_427 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_31_445 ();
 sg13g2_decap_8 FILLER_31_452 ();
 sg13g2_decap_4 FILLER_31_459 ();
 sg13g2_decap_8 FILLER_31_468 ();
 sg13g2_fill_1 FILLER_31_475 ();
 sg13g2_fill_2 FILLER_31_503 ();
 sg13g2_decap_8 FILLER_31_518 ();
 sg13g2_decap_8 FILLER_31_525 ();
 sg13g2_decap_4 FILLER_31_532 ();
 sg13g2_fill_2 FILLER_31_536 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_fill_2 FILLER_31_560 ();
 sg13g2_fill_1 FILLER_31_562 ();
 sg13g2_decap_8 FILLER_31_603 ();
 sg13g2_decap_8 FILLER_31_610 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_4 FILLER_31_644 ();
 sg13g2_fill_1 FILLER_31_648 ();
 sg13g2_decap_8 FILLER_31_661 ();
 sg13g2_decap_8 FILLER_31_668 ();
 sg13g2_fill_1 FILLER_31_675 ();
 sg13g2_fill_2 FILLER_31_681 ();
 sg13g2_fill_2 FILLER_31_714 ();
 sg13g2_fill_1 FILLER_31_716 ();
 sg13g2_fill_2 FILLER_31_726 ();
 sg13g2_fill_2 FILLER_31_744 ();
 sg13g2_fill_1 FILLER_31_746 ();
 sg13g2_decap_8 FILLER_31_751 ();
 sg13g2_fill_2 FILLER_31_758 ();
 sg13g2_fill_2 FILLER_31_764 ();
 sg13g2_fill_1 FILLER_31_766 ();
 sg13g2_fill_1 FILLER_31_807 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_fill_1 FILLER_31_857 ();
 sg13g2_fill_1 FILLER_31_893 ();
 sg13g2_fill_2 FILLER_31_921 ();
 sg13g2_fill_1 FILLER_31_953 ();
 sg13g2_fill_2 FILLER_31_957 ();
 sg13g2_fill_1 FILLER_31_959 ();
 sg13g2_decap_8 FILLER_31_991 ();
 sg13g2_fill_2 FILLER_31_998 ();
 sg13g2_fill_2 FILLER_31_1027 ();
 sg13g2_decap_8 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_18 ();
 sg13g2_decap_8 FILLER_32_25 ();
 sg13g2_decap_8 FILLER_32_32 ();
 sg13g2_decap_8 FILLER_32_39 ();
 sg13g2_decap_8 FILLER_32_46 ();
 sg13g2_decap_8 FILLER_32_53 ();
 sg13g2_decap_8 FILLER_32_60 ();
 sg13g2_decap_8 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_74 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_decap_8 FILLER_32_88 ();
 sg13g2_decap_8 FILLER_32_95 ();
 sg13g2_decap_8 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_109 ();
 sg13g2_decap_8 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_123 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_144 ();
 sg13g2_decap_8 FILLER_32_151 ();
 sg13g2_decap_8 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_172 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_186 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_decap_8 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_decap_8 FILLER_32_312 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_8 FILLER_32_403 ();
 sg13g2_decap_8 FILLER_32_410 ();
 sg13g2_decap_8 FILLER_32_417 ();
 sg13g2_decap_4 FILLER_32_424 ();
 sg13g2_fill_2 FILLER_32_436 ();
 sg13g2_decap_8 FILLER_32_442 ();
 sg13g2_decap_8 FILLER_32_449 ();
 sg13g2_decap_8 FILLER_32_456 ();
 sg13g2_decap_8 FILLER_32_463 ();
 sg13g2_fill_2 FILLER_32_470 ();
 sg13g2_fill_1 FILLER_32_472 ();
 sg13g2_fill_1 FILLER_32_477 ();
 sg13g2_decap_8 FILLER_32_482 ();
 sg13g2_decap_8 FILLER_32_489 ();
 sg13g2_fill_1 FILLER_32_496 ();
 sg13g2_decap_4 FILLER_32_524 ();
 sg13g2_fill_2 FILLER_32_555 ();
 sg13g2_fill_1 FILLER_32_557 ();
 sg13g2_fill_2 FILLER_32_585 ();
 sg13g2_fill_1 FILLER_32_587 ();
 sg13g2_decap_4 FILLER_32_615 ();
 sg13g2_fill_2 FILLER_32_619 ();
 sg13g2_fill_2 FILLER_32_648 ();
 sg13g2_fill_1 FILLER_32_650 ();
 sg13g2_fill_2 FILLER_32_678 ();
 sg13g2_fill_1 FILLER_32_680 ();
 sg13g2_decap_8 FILLER_32_698 ();
 sg13g2_decap_8 FILLER_32_705 ();
 sg13g2_decap_4 FILLER_32_712 ();
 sg13g2_fill_1 FILLER_32_716 ();
 sg13g2_decap_8 FILLER_32_720 ();
 sg13g2_fill_2 FILLER_32_727 ();
 sg13g2_fill_1 FILLER_32_729 ();
 sg13g2_decap_8 FILLER_32_742 ();
 sg13g2_fill_1 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_753 ();
 sg13g2_decap_8 FILLER_32_760 ();
 sg13g2_decap_4 FILLER_32_767 ();
 sg13g2_fill_1 FILLER_32_776 ();
 sg13g2_decap_4 FILLER_32_789 ();
 sg13g2_fill_1 FILLER_32_793 ();
 sg13g2_fill_1 FILLER_32_797 ();
 sg13g2_fill_2 FILLER_32_801 ();
 sg13g2_fill_1 FILLER_32_842 ();
 sg13g2_decap_4 FILLER_32_852 ();
 sg13g2_fill_2 FILLER_32_874 ();
 sg13g2_decap_4 FILLER_32_915 ();
 sg13g2_fill_1 FILLER_32_919 ();
 sg13g2_fill_1 FILLER_32_923 ();
 sg13g2_fill_1 FILLER_32_945 ();
 sg13g2_fill_1 FILLER_32_949 ();
 sg13g2_fill_1 FILLER_32_982 ();
 sg13g2_decap_8 FILLER_32_986 ();
 sg13g2_fill_1 FILLER_32_993 ();
 sg13g2_decap_4 FILLER_32_997 ();
 sg13g2_fill_1 FILLER_32_1001 ();
 sg13g2_decap_4 FILLER_32_1024 ();
 sg13g2_fill_1 FILLER_32_1028 ();
 sg13g2_decap_8 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_11 ();
 sg13g2_decap_8 FILLER_33_18 ();
 sg13g2_decap_8 FILLER_33_25 ();
 sg13g2_decap_8 FILLER_33_32 ();
 sg13g2_decap_8 FILLER_33_39 ();
 sg13g2_decap_8 FILLER_33_46 ();
 sg13g2_decap_8 FILLER_33_53 ();
 sg13g2_decap_8 FILLER_33_60 ();
 sg13g2_decap_8 FILLER_33_67 ();
 sg13g2_decap_8 FILLER_33_74 ();
 sg13g2_decap_8 FILLER_33_81 ();
 sg13g2_decap_8 FILLER_33_88 ();
 sg13g2_decap_8 FILLER_33_95 ();
 sg13g2_decap_8 FILLER_33_102 ();
 sg13g2_decap_8 FILLER_33_109 ();
 sg13g2_decap_8 FILLER_33_116 ();
 sg13g2_decap_8 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_130 ();
 sg13g2_decap_8 FILLER_33_137 ();
 sg13g2_decap_8 FILLER_33_144 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_decap_8 FILLER_33_158 ();
 sg13g2_decap_8 FILLER_33_165 ();
 sg13g2_decap_8 FILLER_33_172 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_decap_8 FILLER_33_200 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_8 FILLER_33_214 ();
 sg13g2_decap_8 FILLER_33_221 ();
 sg13g2_decap_8 FILLER_33_228 ();
 sg13g2_decap_8 FILLER_33_235 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_decap_8 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_284 ();
 sg13g2_decap_8 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_decap_8 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_8 FILLER_33_403 ();
 sg13g2_decap_8 FILLER_33_410 ();
 sg13g2_decap_4 FILLER_33_417 ();
 sg13g2_decap_8 FILLER_33_460 ();
 sg13g2_fill_1 FILLER_33_467 ();
 sg13g2_fill_2 FILLER_33_500 ();
 sg13g2_fill_1 FILLER_33_506 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_fill_1 FILLER_33_532 ();
 sg13g2_fill_2 FILLER_33_537 ();
 sg13g2_fill_1 FILLER_33_539 ();
 sg13g2_fill_1 FILLER_33_543 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_fill_2 FILLER_33_570 ();
 sg13g2_decap_8 FILLER_33_580 ();
 sg13g2_decap_4 FILLER_33_606 ();
 sg13g2_fill_2 FILLER_33_613 ();
 sg13g2_fill_1 FILLER_33_618 ();
 sg13g2_decap_8 FILLER_33_642 ();
 sg13g2_fill_1 FILLER_33_655 ();
 sg13g2_fill_2 FILLER_33_667 ();
 sg13g2_fill_1 FILLER_33_669 ();
 sg13g2_fill_2 FILLER_33_673 ();
 sg13g2_decap_4 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_34_4 ();
 sg13g2_decap_8 FILLER_34_11 ();
 sg13g2_decap_8 FILLER_34_18 ();
 sg13g2_decap_8 FILLER_34_25 ();
 sg13g2_decap_8 FILLER_34_32 ();
 sg13g2_decap_8 FILLER_34_39 ();
 sg13g2_decap_8 FILLER_34_46 ();
 sg13g2_decap_8 FILLER_34_53 ();
 sg13g2_decap_8 FILLER_34_60 ();
 sg13g2_decap_8 FILLER_34_67 ();
 sg13g2_decap_8 FILLER_34_74 ();
 sg13g2_decap_8 FILLER_34_81 ();
 sg13g2_decap_8 FILLER_34_88 ();
 sg13g2_decap_8 FILLER_34_95 ();
 sg13g2_decap_8 FILLER_34_102 ();
 sg13g2_decap_8 FILLER_34_109 ();
 sg13g2_decap_8 FILLER_34_116 ();
 sg13g2_decap_8 FILLER_34_123 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_decap_8 FILLER_34_137 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_decap_8 FILLER_34_158 ();
 sg13g2_decap_8 FILLER_34_165 ();
 sg13g2_decap_8 FILLER_34_172 ();
 sg13g2_decap_8 FILLER_34_179 ();
 sg13g2_decap_8 FILLER_34_186 ();
 sg13g2_decap_8 FILLER_34_193 ();
 sg13g2_decap_8 FILLER_34_200 ();
 sg13g2_decap_8 FILLER_34_207 ();
 sg13g2_decap_8 FILLER_34_214 ();
 sg13g2_decap_8 FILLER_34_221 ();
 sg13g2_decap_8 FILLER_34_228 ();
 sg13g2_decap_8 FILLER_34_235 ();
 sg13g2_decap_8 FILLER_34_242 ();
 sg13g2_decap_8 FILLER_34_249 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_270 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_decap_8 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_298 ();
 sg13g2_decap_8 FILLER_34_305 ();
 sg13g2_decap_8 FILLER_34_312 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_decap_8 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_decap_8 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_347 ();
 sg13g2_decap_8 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_8 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_34_410 ();
 sg13g2_decap_8 FILLER_34_417 ();
 sg13g2_decap_4 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_34_442 ();
 sg13g2_decap_8 FILLER_34_449 ();
 sg13g2_decap_8 FILLER_34_456 ();
 sg13g2_decap_8 FILLER_34_463 ();
 sg13g2_fill_1 FILLER_34_470 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_decap_8 FILLER_34_483 ();
 sg13g2_fill_2 FILLER_34_490 ();
 sg13g2_fill_1 FILLER_34_492 ();
 sg13g2_decap_8 FILLER_34_497 ();
 sg13g2_decap_8 FILLER_34_504 ();
 sg13g2_decap_8 FILLER_34_524 ();
 sg13g2_decap_4 FILLER_34_531 ();
 sg13g2_decap_8 FILLER_34_562 ();
 sg13g2_fill_1 FILLER_34_569 ();
 sg13g2_fill_1 FILLER_34_573 ();
 sg13g2_decap_8 FILLER_34_587 ();
 sg13g2_decap_4 FILLER_34_594 ();
 sg13g2_decap_4 FILLER_34_602 ();
 sg13g2_fill_1 FILLER_34_606 ();
 sg13g2_decap_8 FILLER_34_611 ();
 sg13g2_decap_8 FILLER_34_618 ();
 sg13g2_fill_1 FILLER_34_625 ();
 sg13g2_decap_8 FILLER_34_633 ();
 sg13g2_decap_8 FILLER_34_640 ();
 sg13g2_decap_4 FILLER_34_647 ();
 sg13g2_fill_2 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_662 ();
 sg13g2_decap_8 FILLER_34_669 ();
 sg13g2_decap_4 FILLER_34_676 ();
 sg13g2_decap_8 FILLER_34_695 ();
 sg13g2_decap_4 FILLER_34_702 ();
 sg13g2_fill_2 FILLER_34_706 ();
 sg13g2_fill_1 FILLER_34_735 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_fill_2 FILLER_35_420 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_fill_2 FILLER_35_430 ();
 sg13g2_decap_8 FILLER_35_437 ();
 sg13g2_decap_8 FILLER_35_444 ();
 sg13g2_decap_8 FILLER_35_451 ();
 sg13g2_decap_8 FILLER_35_458 ();
 sg13g2_fill_1 FILLER_35_465 ();
 sg13g2_decap_8 FILLER_35_473 ();
 sg13g2_fill_1 FILLER_35_480 ();
 sg13g2_decap_4 FILLER_35_513 ();
 sg13g2_fill_2 FILLER_35_517 ();
 sg13g2_decap_8 FILLER_35_523 ();
 sg13g2_decap_4 FILLER_35_530 ();
 sg13g2_fill_2 FILLER_35_534 ();
 sg13g2_fill_2 FILLER_35_545 ();
 sg13g2_fill_1 FILLER_35_547 ();
 sg13g2_decap_8 FILLER_35_553 ();
 sg13g2_fill_2 FILLER_35_560 ();
 sg13g2_fill_1 FILLER_35_562 ();
 sg13g2_decap_4 FILLER_35_639 ();
 sg13g2_fill_2 FILLER_35_643 ();
 sg13g2_decap_8 FILLER_35_676 ();
 sg13g2_fill_1 FILLER_35_683 ();
 sg13g2_decap_8 FILLER_35_695 ();
 sg13g2_decap_4 FILLER_35_702 ();
 sg13g2_fill_2 FILLER_35_706 ();
 sg13g2_decap_8 FILLER_35_726 ();
 sg13g2_fill_2 FILLER_35_733 ();
 sg13g2_fill_1 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_36_406 ();
 sg13g2_decap_4 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_444 ();
 sg13g2_decap_8 FILLER_36_451 ();
 sg13g2_fill_1 FILLER_36_458 ();
 sg13g2_decap_8 FILLER_36_472 ();
 sg13g2_decap_8 FILLER_36_479 ();
 sg13g2_fill_1 FILLER_36_486 ();
 sg13g2_decap_8 FILLER_36_507 ();
 sg13g2_decap_4 FILLER_36_541 ();
 sg13g2_fill_1 FILLER_36_545 ();
 sg13g2_decap_8 FILLER_36_553 ();
 sg13g2_decap_8 FILLER_36_560 ();
 sg13g2_fill_2 FILLER_36_582 ();
 sg13g2_decap_4 FILLER_36_618 ();
 sg13g2_fill_2 FILLER_36_622 ();
 sg13g2_fill_1 FILLER_36_655 ();
 sg13g2_fill_2 FILLER_36_676 ();
 sg13g2_decap_4 FILLER_36_713 ();
 sg13g2_decap_8 FILLER_36_732 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_fill_2 FILLER_37_420 ();
 sg13g2_fill_1 FILLER_37_422 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_501 ();
 sg13g2_decap_8 FILLER_37_508 ();
 sg13g2_decap_4 FILLER_37_515 ();
 sg13g2_fill_2 FILLER_37_519 ();
 sg13g2_decap_4 FILLER_37_534 ();
 sg13g2_fill_2 FILLER_37_551 ();
 sg13g2_decap_8 FILLER_37_557 ();
 sg13g2_decap_8 FILLER_37_564 ();
 sg13g2_fill_2 FILLER_37_571 ();
 sg13g2_fill_1 FILLER_37_600 ();
 sg13g2_decap_8 FILLER_37_613 ();
 sg13g2_decap_8 FILLER_37_620 ();
 sg13g2_decap_8 FILLER_37_627 ();
 sg13g2_decap_8 FILLER_37_643 ();
 sg13g2_fill_2 FILLER_37_663 ();
 sg13g2_fill_1 FILLER_37_673 ();
 sg13g2_fill_2 FILLER_37_678 ();
 sg13g2_decap_4 FILLER_37_685 ();
 sg13g2_fill_1 FILLER_37_689 ();
 sg13g2_fill_1 FILLER_37_699 ();
 sg13g2_decap_4 FILLER_37_704 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_4 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_410 ();
 sg13g2_decap_4 FILLER_38_443 ();
 sg13g2_fill_2 FILLER_38_447 ();
 sg13g2_decap_4 FILLER_38_476 ();
 sg13g2_fill_1 FILLER_38_480 ();
 sg13g2_fill_2 FILLER_38_575 ();
 sg13g2_decap_8 FILLER_38_594 ();
 sg13g2_fill_2 FILLER_38_601 ();
 sg13g2_decap_4 FILLER_38_619 ();
 sg13g2_fill_2 FILLER_38_623 ();
 sg13g2_fill_2 FILLER_38_652 ();
 sg13g2_fill_1 FILLER_38_654 ();
 sg13g2_fill_2 FILLER_38_686 ();
 sg13g2_fill_1 FILLER_38_688 ();
 sg13g2_decap_4 FILLER_38_733 ();
 sg13g2_fill_2 FILLER_38_737 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_4 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_433 ();
 sg13g2_decap_4 FILLER_39_440 ();
 sg13g2_fill_1 FILLER_39_456 ();
 sg13g2_decap_8 FILLER_39_466 ();
 sg13g2_decap_8 FILLER_39_479 ();
 sg13g2_decap_4 FILLER_39_491 ();
 sg13g2_fill_1 FILLER_39_495 ();
 sg13g2_decap_8 FILLER_39_503 ();
 sg13g2_decap_4 FILLER_39_510 ();
 sg13g2_decap_4 FILLER_39_520 ();
 sg13g2_fill_1 FILLER_39_524 ();
 sg13g2_decap_4 FILLER_39_528 ();
 sg13g2_fill_1 FILLER_39_532 ();
 sg13g2_decap_8 FILLER_39_540 ();
 sg13g2_fill_1 FILLER_39_547 ();
 sg13g2_decap_8 FILLER_39_551 ();
 sg13g2_decap_8 FILLER_39_558 ();
 sg13g2_fill_1 FILLER_39_584 ();
 sg13g2_decap_4 FILLER_39_592 ();
 sg13g2_fill_2 FILLER_39_596 ();
 sg13g2_fill_2 FILLER_39_628 ();
 sg13g2_fill_2 FILLER_39_634 ();
 sg13g2_fill_1 FILLER_39_663 ();
 sg13g2_decap_8 FILLER_39_668 ();
 sg13g2_decap_4 FILLER_39_675 ();
 sg13g2_fill_2 FILLER_39_679 ();
 sg13g2_decap_8 FILLER_39_704 ();
 sg13g2_decap_8 FILLER_39_711 ();
 sg13g2_fill_2 FILLER_39_718 ();
 sg13g2_decap_8 FILLER_39_723 ();
 sg13g2_decap_8 FILLER_39_730 ();
 sg13g2_fill_2 FILLER_39_737 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_fill_2 FILLER_40_413 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_438 ();
 sg13g2_decap_8 FILLER_40_445 ();
 sg13g2_decap_4 FILLER_40_452 ();
 sg13g2_fill_2 FILLER_40_456 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_485 ();
 sg13g2_fill_1 FILLER_40_492 ();
 sg13g2_fill_2 FILLER_40_501 ();
 sg13g2_decap_8 FILLER_40_512 ();
 sg13g2_decap_8 FILLER_40_519 ();
 sg13g2_decap_4 FILLER_40_526 ();
 sg13g2_fill_2 FILLER_40_530 ();
 sg13g2_fill_1 FILLER_40_547 ();
 sg13g2_decap_8 FILLER_40_551 ();
 sg13g2_fill_2 FILLER_40_594 ();
 sg13g2_decap_4 FILLER_40_599 ();
 sg13g2_fill_2 FILLER_40_603 ();
 sg13g2_fill_2 FILLER_40_616 ();
 sg13g2_fill_1 FILLER_40_618 ();
 sg13g2_decap_8 FILLER_40_622 ();
 sg13g2_decap_4 FILLER_40_629 ();
 sg13g2_fill_1 FILLER_40_633 ();
 sg13g2_fill_2 FILLER_40_637 ();
 sg13g2_fill_1 FILLER_40_639 ();
 sg13g2_decap_8 FILLER_40_652 ();
 sg13g2_decap_8 FILLER_40_659 ();
 sg13g2_decap_8 FILLER_40_666 ();
 sg13g2_decap_4 FILLER_40_673 ();
 sg13g2_fill_1 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_684 ();
 sg13g2_decap_4 FILLER_40_691 ();
 sg13g2_decap_8 FILLER_40_725 ();
 sg13g2_fill_2 FILLER_40_732 ();
 sg13g2_fill_2 FILLER_40_737 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_fill_2 FILLER_41_413 ();
 sg13g2_fill_1 FILLER_41_415 ();
 sg13g2_fill_2 FILLER_41_447 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_4 FILLER_41_476 ();
 sg13g2_fill_1 FILLER_41_480 ();
 sg13g2_decap_8 FILLER_41_527 ();
 sg13g2_decap_8 FILLER_41_561 ();
 sg13g2_fill_2 FILLER_41_589 ();
 sg13g2_fill_1 FILLER_41_591 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_fill_2 FILLER_41_602 ();
 sg13g2_decap_4 FILLER_41_639 ();
 sg13g2_decap_8 FILLER_41_673 ();
 sg13g2_fill_1 FILLER_41_680 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_709 ();
 sg13g2_decap_4 FILLER_41_716 ();
 sg13g2_fill_2 FILLER_41_733 ();
 sg13g2_fill_1 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_413 ();
 sg13g2_fill_1 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_429 ();
 sg13g2_decap_8 FILLER_42_436 ();
 sg13g2_decap_8 FILLER_42_443 ();
 sg13g2_decap_4 FILLER_42_450 ();
 sg13g2_fill_2 FILLER_42_535 ();
 sg13g2_fill_2 FILLER_42_542 ();
 sg13g2_fill_1 FILLER_42_544 ();
 sg13g2_decap_8 FILLER_42_557 ();
 sg13g2_decap_4 FILLER_42_564 ();
 sg13g2_fill_1 FILLER_42_568 ();
 sg13g2_decap_4 FILLER_42_573 ();
 sg13g2_decap_4 FILLER_42_581 ();
 sg13g2_decap_8 FILLER_42_626 ();
 sg13g2_decap_8 FILLER_42_633 ();
 sg13g2_decap_8 FILLER_42_640 ();
 sg13g2_fill_1 FILLER_42_652 ();
 sg13g2_decap_4 FILLER_42_661 ();
 sg13g2_fill_1 FILLER_42_665 ();
 sg13g2_fill_2 FILLER_42_693 ();
 sg13g2_fill_1 FILLER_42_695 ();
 sg13g2_fill_1 FILLER_42_704 ();
 sg13g2_decap_8 FILLER_42_709 ();
 sg13g2_decap_8 FILLER_42_716 ();
 sg13g2_decap_4 FILLER_42_723 ();
 sg13g2_fill_2 FILLER_42_727 ();
 sg13g2_decap_4 FILLER_42_732 ();
 sg13g2_fill_2 FILLER_42_736 ();
 sg13g2_decap_8 FILLER_42_742 ();
 sg13g2_decap_8 FILLER_42_749 ();
 sg13g2_fill_1 FILLER_42_756 ();
 sg13g2_decap_8 FILLER_42_760 ();
 sg13g2_fill_2 FILLER_42_775 ();
 sg13g2_decap_4 FILLER_42_789 ();
 sg13g2_fill_1 FILLER_42_793 ();
 sg13g2_fill_2 FILLER_42_799 ();
 sg13g2_fill_1 FILLER_42_801 ();
 sg13g2_decap_8 FILLER_42_815 ();
 sg13g2_decap_4 FILLER_42_851 ();
 sg13g2_fill_1 FILLER_42_858 ();
 sg13g2_decap_8 FILLER_42_862 ();
 sg13g2_fill_1 FILLER_42_878 ();
 sg13g2_fill_1 FILLER_42_888 ();
 sg13g2_fill_2 FILLER_42_908 ();
 sg13g2_fill_1 FILLER_42_916 ();
 sg13g2_decap_4 FILLER_42_923 ();
 sg13g2_fill_2 FILLER_42_927 ();
 sg13g2_fill_2 FILLER_42_932 ();
 sg13g2_fill_2 FILLER_42_937 ();
 sg13g2_fill_1 FILLER_42_939 ();
 sg13g2_fill_2 FILLER_42_943 ();
 sg13g2_fill_1 FILLER_42_945 ();
 sg13g2_fill_1 FILLER_42_967 ();
 sg13g2_fill_1 FILLER_42_971 ();
 sg13g2_decap_8 FILLER_42_975 ();
 sg13g2_decap_4 FILLER_42_982 ();
 sg13g2_fill_1 FILLER_42_986 ();
 sg13g2_fill_1 FILLER_42_992 ();
 sg13g2_decap_4 FILLER_42_999 ();
 sg13g2_decap_8 FILLER_42_1020 ();
 sg13g2_fill_2 FILLER_42_1027 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_fill_2 FILLER_43_462 ();
 sg13g2_fill_1 FILLER_43_464 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_decap_8 FILLER_43_476 ();
 sg13g2_decap_4 FILLER_43_483 ();
 sg13g2_decap_8 FILLER_43_491 ();
 sg13g2_decap_8 FILLER_43_498 ();
 sg13g2_decap_8 FILLER_43_505 ();
 sg13g2_fill_1 FILLER_43_512 ();
 sg13g2_decap_4 FILLER_43_517 ();
 sg13g2_fill_1 FILLER_43_521 ();
 sg13g2_decap_8 FILLER_43_526 ();
 sg13g2_decap_8 FILLER_43_533 ();
 sg13g2_fill_2 FILLER_43_540 ();
 sg13g2_decap_8 FILLER_43_562 ();
 sg13g2_fill_1 FILLER_43_600 ();
 sg13g2_decap_8 FILLER_43_610 ();
 sg13g2_decap_8 FILLER_43_617 ();
 sg13g2_decap_8 FILLER_43_624 ();
 sg13g2_decap_8 FILLER_43_631 ();
 sg13g2_fill_2 FILLER_43_638 ();
 sg13g2_fill_1 FILLER_43_640 ();
 sg13g2_decap_8 FILLER_43_661 ();
 sg13g2_decap_4 FILLER_43_668 ();
 sg13g2_decap_4 FILLER_43_676 ();
 sg13g2_fill_1 FILLER_43_680 ();
 sg13g2_fill_2 FILLER_43_690 ();
 sg13g2_fill_1 FILLER_43_692 ();
 sg13g2_fill_2 FILLER_43_698 ();
 sg13g2_decap_4 FILLER_43_727 ();
 sg13g2_fill_2 FILLER_43_731 ();
 sg13g2_fill_1 FILLER_43_760 ();
 sg13g2_fill_1 FILLER_43_780 ();
 sg13g2_decap_4 FILLER_43_784 ();
 sg13g2_decap_4 FILLER_43_827 ();
 sg13g2_fill_2 FILLER_43_834 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_decap_8 FILLER_43_875 ();
 sg13g2_fill_2 FILLER_43_914 ();
 sg13g2_fill_2 FILLER_43_971 ();
 sg13g2_fill_1 FILLER_43_973 ();
 sg13g2_fill_1 FILLER_43_978 ();
 sg13g2_fill_1 FILLER_43_984 ();
 sg13g2_fill_2 FILLER_43_1000 ();
 sg13g2_fill_1 FILLER_43_1002 ();
 sg13g2_decap_8 FILLER_43_1018 ();
 sg13g2_decap_4 FILLER_43_1025 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_8 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_301 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_44_406 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_decap_8 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_4 FILLER_44_462 ();
 sg13g2_fill_1 FILLER_44_466 ();
 sg13g2_decap_8 FILLER_44_471 ();
 sg13g2_decap_8 FILLER_44_478 ();
 sg13g2_fill_1 FILLER_44_485 ();
 sg13g2_decap_8 FILLER_44_491 ();
 sg13g2_decap_8 FILLER_44_498 ();
 sg13g2_decap_8 FILLER_44_508 ();
 sg13g2_fill_2 FILLER_44_515 ();
 sg13g2_decap_8 FILLER_44_593 ();
 sg13g2_decap_8 FILLER_44_600 ();
 sg13g2_fill_2 FILLER_44_620 ();
 sg13g2_fill_1 FILLER_44_622 ();
 sg13g2_fill_1 FILLER_44_653 ();
 sg13g2_decap_8 FILLER_44_697 ();
 sg13g2_decap_8 FILLER_44_704 ();
 sg13g2_fill_1 FILLER_44_711 ();
 sg13g2_decap_4 FILLER_44_717 ();
 sg13g2_decap_8 FILLER_44_741 ();
 sg13g2_decap_4 FILLER_44_748 ();
 sg13g2_decap_8 FILLER_44_783 ();
 sg13g2_decap_4 FILLER_44_790 ();
 sg13g2_fill_2 FILLER_44_794 ();
 sg13g2_decap_4 FILLER_44_816 ();
 sg13g2_fill_1 FILLER_44_820 ();
 sg13g2_fill_2 FILLER_44_848 ();
 sg13g2_fill_1 FILLER_44_850 ();
 sg13g2_fill_2 FILLER_44_886 ();
 sg13g2_fill_1 FILLER_44_888 ();
 sg13g2_decap_8 FILLER_44_929 ();
 sg13g2_decap_4 FILLER_44_936 ();
 sg13g2_fill_2 FILLER_44_940 ();
 sg13g2_fill_1 FILLER_44_996 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_fill_1 FILLER_45_489 ();
 sg13g2_decap_8 FILLER_45_498 ();
 sg13g2_decap_8 FILLER_45_517 ();
 sg13g2_decap_8 FILLER_45_524 ();
 sg13g2_decap_8 FILLER_45_531 ();
 sg13g2_decap_8 FILLER_45_538 ();
 sg13g2_decap_8 FILLER_45_554 ();
 sg13g2_decap_8 FILLER_45_561 ();
 sg13g2_decap_8 FILLER_45_568 ();
 sg13g2_fill_1 FILLER_45_575 ();
 sg13g2_decap_8 FILLER_45_594 ();
 sg13g2_decap_4 FILLER_45_601 ();
 sg13g2_fill_2 FILLER_45_636 ();
 sg13g2_fill_1 FILLER_45_647 ();
 sg13g2_fill_2 FILLER_45_656 ();
 sg13g2_fill_1 FILLER_45_658 ();
 sg13g2_decap_8 FILLER_45_663 ();
 sg13g2_decap_4 FILLER_45_670 ();
 sg13g2_fill_1 FILLER_45_674 ();
 sg13g2_fill_1 FILLER_45_729 ();
 sg13g2_decap_4 FILLER_45_757 ();
 sg13g2_fill_1 FILLER_45_761 ();
 sg13g2_decap_8 FILLER_45_767 ();
 sg13g2_decap_8 FILLER_45_779 ();
 sg13g2_decap_4 FILLER_45_786 ();
 sg13g2_fill_1 FILLER_45_790 ();
 sg13g2_fill_2 FILLER_45_823 ();
 sg13g2_fill_1 FILLER_45_825 ();
 sg13g2_decap_8 FILLER_45_830 ();
 sg13g2_decap_4 FILLER_45_846 ();
 sg13g2_fill_2 FILLER_45_850 ();
 sg13g2_decap_8 FILLER_45_868 ();
 sg13g2_decap_4 FILLER_45_875 ();
 sg13g2_fill_1 FILLER_45_879 ();
 sg13g2_decap_8 FILLER_45_915 ();
 sg13g2_fill_2 FILLER_45_922 ();
 sg13g2_fill_1 FILLER_45_924 ();
 sg13g2_decap_8 FILLER_45_930 ();
 sg13g2_decap_4 FILLER_45_937 ();
 sg13g2_fill_1 FILLER_45_941 ();
 sg13g2_decap_8 FILLER_45_955 ();
 sg13g2_decap_8 FILLER_45_962 ();
 sg13g2_decap_8 FILLER_45_969 ();
 sg13g2_decap_8 FILLER_45_976 ();
 sg13g2_fill_1 FILLER_45_983 ();
 sg13g2_decap_8 FILLER_45_988 ();
 sg13g2_decap_8 FILLER_45_995 ();
 sg13g2_decap_4 FILLER_45_1002 ();
 sg13g2_fill_2 FILLER_45_1006 ();
 sg13g2_decap_8 FILLER_45_1015 ();
 sg13g2_decap_8 FILLER_45_1022 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_533 ();
 sg13g2_decap_8 FILLER_46_540 ();
 sg13g2_fill_2 FILLER_46_547 ();
 sg13g2_fill_1 FILLER_46_549 ();
 sg13g2_decap_4 FILLER_46_566 ();
 sg13g2_fill_1 FILLER_46_570 ();
 sg13g2_decap_8 FILLER_46_622 ();
 sg13g2_decap_8 FILLER_46_629 ();
 sg13g2_fill_2 FILLER_46_636 ();
 sg13g2_fill_2 FILLER_46_654 ();
 sg13g2_fill_1 FILLER_46_656 ();
 sg13g2_decap_8 FILLER_46_660 ();
 sg13g2_decap_8 FILLER_46_667 ();
 sg13g2_decap_8 FILLER_46_693 ();
 sg13g2_fill_2 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_706 ();
 sg13g2_fill_2 FILLER_46_713 ();
 sg13g2_fill_1 FILLER_46_715 ();
 sg13g2_fill_2 FILLER_46_720 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_749 ();
 sg13g2_fill_1 FILLER_46_756 ();
 sg13g2_decap_8 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_fill_1 FILLER_46_806 ();
 sg13g2_decap_8 FILLER_46_820 ();
 sg13g2_decap_8 FILLER_46_827 ();
 sg13g2_decap_8 FILLER_46_834 ();
 sg13g2_decap_8 FILLER_46_841 ();
 sg13g2_fill_2 FILLER_46_853 ();
 sg13g2_decap_8 FILLER_46_859 ();
 sg13g2_decap_4 FILLER_46_866 ();
 sg13g2_fill_2 FILLER_46_870 ();
 sg13g2_fill_2 FILLER_46_875 ();
 sg13g2_decap_4 FILLER_46_880 ();
 sg13g2_fill_2 FILLER_46_884 ();
 sg13g2_fill_2 FILLER_46_891 ();
 sg13g2_fill_1 FILLER_46_893 ();
 sg13g2_fill_2 FILLER_46_898 ();
 sg13g2_decap_8 FILLER_46_904 ();
 sg13g2_decap_4 FILLER_46_911 ();
 sg13g2_fill_2 FILLER_46_915 ();
 sg13g2_fill_2 FILLER_46_937 ();
 sg13g2_decap_8 FILLER_46_943 ();
 sg13g2_fill_2 FILLER_46_950 ();
 sg13g2_fill_1 FILLER_46_965 ();
 sg13g2_decap_8 FILLER_46_969 ();
 sg13g2_fill_1 FILLER_46_976 ();
 sg13g2_fill_1 FILLER_46_980 ();
 sg13g2_decap_4 FILLER_46_994 ();
 sg13g2_fill_2 FILLER_46_998 ();
 sg13g2_fill_2 FILLER_46_1027 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_4 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_516 ();
 sg13g2_fill_2 FILLER_47_523 ();
 sg13g2_fill_1 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_565 ();
 sg13g2_decap_4 FILLER_47_572 ();
 sg13g2_decap_8 FILLER_47_590 ();
 sg13g2_decap_8 FILLER_47_597 ();
 sg13g2_fill_1 FILLER_47_604 ();
 sg13g2_decap_8 FILLER_47_614 ();
 sg13g2_decap_4 FILLER_47_621 ();
 sg13g2_fill_2 FILLER_47_625 ();
 sg13g2_fill_2 FILLER_47_667 ();
 sg13g2_fill_1 FILLER_47_669 ();
 sg13g2_fill_2 FILLER_47_675 ();
 sg13g2_fill_1 FILLER_47_677 ();
 sg13g2_decap_8 FILLER_47_683 ();
 sg13g2_decap_8 FILLER_47_690 ();
 sg13g2_fill_2 FILLER_47_701 ();
 sg13g2_fill_1 FILLER_47_703 ();
 sg13g2_fill_2 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_752 ();
 sg13g2_fill_2 FILLER_47_759 ();
 sg13g2_fill_1 FILLER_47_761 ();
 sg13g2_decap_4 FILLER_47_766 ();
 sg13g2_fill_1 FILLER_47_770 ();
 sg13g2_fill_2 FILLER_47_776 ();
 sg13g2_fill_1 FILLER_47_806 ();
 sg13g2_decap_8 FILLER_47_810 ();
 sg13g2_decap_4 FILLER_47_817 ();
 sg13g2_fill_1 FILLER_47_821 ();
 sg13g2_fill_2 FILLER_47_825 ();
 sg13g2_fill_2 FILLER_47_847 ();
 sg13g2_fill_1 FILLER_47_849 ();
 sg13g2_decap_4 FILLER_47_877 ();
 sg13g2_decap_8 FILLER_47_901 ();
 sg13g2_fill_2 FILLER_47_908 ();
 sg13g2_decap_8 FILLER_47_913 ();
 sg13g2_decap_8 FILLER_47_925 ();
 sg13g2_fill_2 FILLER_47_932 ();
 sg13g2_decap_8 FILLER_47_961 ();
 sg13g2_decap_4 FILLER_47_968 ();
 sg13g2_decap_8 FILLER_47_991 ();
 sg13g2_fill_2 FILLER_47_998 ();
 sg13g2_fill_1 FILLER_47_1000 ();
 sg13g2_fill_2 FILLER_47_1010 ();
 sg13g2_decap_8 FILLER_47_1017 ();
 sg13g2_decap_4 FILLER_47_1024 ();
 sg13g2_fill_1 FILLER_47_1028 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_4 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_4 FILLER_48_525 ();
 sg13g2_fill_2 FILLER_48_529 ();
 sg13g2_decap_8 FILLER_48_535 ();
 sg13g2_fill_2 FILLER_48_542 ();
 sg13g2_fill_1 FILLER_48_544 ();
 sg13g2_fill_2 FILLER_48_572 ();
 sg13g2_fill_1 FILLER_48_628 ();
 sg13g2_decap_8 FILLER_48_656 ();
 sg13g2_fill_2 FILLER_48_690 ();
 sg13g2_decap_4 FILLER_48_719 ();
 sg13g2_fill_2 FILLER_48_723 ();
 sg13g2_fill_2 FILLER_48_745 ();
 sg13g2_decap_8 FILLER_48_752 ();
 sg13g2_decap_4 FILLER_48_786 ();
 sg13g2_decap_4 FILLER_48_848 ();
 sg13g2_fill_2 FILLER_48_852 ();
 sg13g2_decap_4 FILLER_48_885 ();
 sg13g2_fill_2 FILLER_48_889 ();
 sg13g2_fill_2 FILLER_48_918 ();
 sg13g2_fill_1 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_18 ();
 sg13g2_decap_8 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_8 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_74 ();
 sg13g2_decap_8 FILLER_49_81 ();
 sg13g2_decap_8 FILLER_49_88 ();
 sg13g2_decap_8 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_102 ();
 sg13g2_decap_8 FILLER_49_109 ();
 sg13g2_decap_8 FILLER_49_116 ();
 sg13g2_decap_8 FILLER_49_123 ();
 sg13g2_decap_8 FILLER_49_130 ();
 sg13g2_decap_8 FILLER_49_137 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_decap_8 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_decap_8 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_8 FILLER_49_179 ();
 sg13g2_decap_8 FILLER_49_186 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_8 FILLER_49_214 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_228 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_256 ();
 sg13g2_decap_8 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_270 ();
 sg13g2_decap_8 FILLER_49_277 ();
 sg13g2_decap_8 FILLER_49_284 ();
 sg13g2_decap_8 FILLER_49_291 ();
 sg13g2_decap_8 FILLER_49_298 ();
 sg13g2_decap_8 FILLER_49_305 ();
 sg13g2_decap_8 FILLER_49_312 ();
 sg13g2_decap_8 FILLER_49_319 ();
 sg13g2_decap_8 FILLER_49_326 ();
 sg13g2_decap_8 FILLER_49_333 ();
 sg13g2_decap_8 FILLER_49_340 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_decap_8 FILLER_49_354 ();
 sg13g2_decap_8 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_8 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_410 ();
 sg13g2_decap_8 FILLER_49_417 ();
 sg13g2_decap_8 FILLER_49_424 ();
 sg13g2_decap_8 FILLER_49_431 ();
 sg13g2_decap_8 FILLER_49_438 ();
 sg13g2_decap_8 FILLER_49_445 ();
 sg13g2_decap_8 FILLER_49_452 ();
 sg13g2_decap_8 FILLER_49_459 ();
 sg13g2_decap_8 FILLER_49_466 ();
 sg13g2_decap_8 FILLER_49_473 ();
 sg13g2_decap_8 FILLER_49_480 ();
 sg13g2_decap_8 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_494 ();
 sg13g2_decap_8 FILLER_49_501 ();
 sg13g2_decap_8 FILLER_49_508 ();
 sg13g2_decap_8 FILLER_49_515 ();
 sg13g2_decap_8 FILLER_49_522 ();
 sg13g2_decap_8 FILLER_49_529 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_fill_1 FILLER_49_543 ();
 sg13g2_decap_8 FILLER_49_557 ();
 sg13g2_decap_8 FILLER_49_564 ();
 sg13g2_fill_2 FILLER_49_571 ();
 sg13g2_decap_8 FILLER_49_589 ();
 sg13g2_decap_8 FILLER_49_596 ();
 sg13g2_fill_2 FILLER_49_603 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_4 FILLER_49_623 ();
 sg13g2_fill_2 FILLER_49_627 ();
 sg13g2_fill_2 FILLER_49_642 ();
 sg13g2_fill_1 FILLER_49_644 ();
 sg13g2_decap_8 FILLER_49_649 ();
 sg13g2_decap_8 FILLER_49_656 ();
 sg13g2_decap_4 FILLER_49_663 ();
 sg13g2_fill_1 FILLER_49_667 ();
 sg13g2_fill_2 FILLER_49_672 ();
 sg13g2_fill_1 FILLER_49_674 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_fill_2 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_713 ();
 sg13g2_decap_8 FILLER_49_720 ();
 sg13g2_fill_2 FILLER_49_727 ();
 sg13g2_fill_1 FILLER_49_729 ();
 sg13g2_decap_8 FILLER_49_738 ();
 sg13g2_decap_8 FILLER_49_745 ();
 sg13g2_decap_8 FILLER_49_752 ();
 sg13g2_decap_4 FILLER_49_759 ();
 sg13g2_fill_1 FILLER_49_763 ();
 sg13g2_fill_1 FILLER_49_768 ();
 sg13g2_decap_4 FILLER_49_772 ();
 sg13g2_fill_2 FILLER_49_780 ();
 sg13g2_decap_8 FILLER_49_785 ();
 sg13g2_fill_1 FILLER_49_792 ();
 sg13g2_decap_8 FILLER_49_803 ();
 sg13g2_decap_8 FILLER_49_810 ();
 sg13g2_fill_2 FILLER_49_817 ();
 sg13g2_fill_1 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_836 ();
 sg13g2_decap_8 FILLER_49_843 ();
 sg13g2_decap_8 FILLER_49_850 ();
 sg13g2_fill_2 FILLER_49_857 ();
 sg13g2_fill_2 FILLER_49_863 ();
 sg13g2_decap_8 FILLER_49_881 ();
 sg13g2_decap_8 FILLER_49_888 ();
 sg13g2_fill_1 FILLER_49_895 ();
 sg13g2_decap_8 FILLER_49_900 ();
 sg13g2_decap_8 FILLER_49_907 ();
 sg13g2_decap_8 FILLER_49_914 ();
 sg13g2_fill_2 FILLER_49_921 ();
 sg13g2_fill_1 FILLER_49_923 ();
 sg13g2_decap_8 FILLER_49_932 ();
 sg13g2_decap_8 FILLER_49_939 ();
 sg13g2_decap_4 FILLER_49_946 ();
 sg13g2_decap_8 FILLER_49_957 ();
 sg13g2_decap_4 FILLER_49_964 ();
 sg13g2_fill_2 FILLER_49_968 ();
 sg13g2_fill_1 FILLER_49_979 ();
 sg13g2_decap_8 FILLER_49_984 ();
 sg13g2_decap_8 FILLER_49_991 ();
 sg13g2_decap_8 FILLER_49_998 ();
 sg13g2_decap_8 FILLER_49_1013 ();
 sg13g2_decap_8 FILLER_49_1020 ();
 sg13g2_fill_2 FILLER_49_1027 ();
 assign uio_oe[0] = net484;
 assign uio_oe[1] = net485;
 assign uio_oe[2] = net486;
 assign uio_oe[3] = net487;
 assign uio_oe[4] = net488;
 assign uio_oe[5] = net489;
 assign uio_oe[6] = net490;
 assign uio_oe[7] = net491;
endmodule
