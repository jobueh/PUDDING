* NGSPICE file created from heichips25_pudding.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for dac128module abstract view
.subckt dac128module ON[64] ONB[64] ON[65] ONB[65] ON[66] ONB[66] ON[67] ONB[67] ON[68]
+ ONB[68] ON[69] ONB[69] ON[70] ONB[70] ON[71] ONB[71] ON[72] ONB[72] EN[2] ENB[2]
+ ON[73] ONB[73] ON[74] ONB[74] ON[75] ONB[75] ON[76] ONB[76] ON[77] ONB[77] ON[78]
+ ONB[78] ON[79] ONB[79] ON[80] ONB[80] ON[81] ONB[81] ON[82] ONB[82] ON[83] ONB[83]
+ ON[84] ONB[84] ON[85] ONB[85] ON[86] ONB[86] ON[87] ONB[87] ON[88] ONB[88] ON[89]
+ ONB[89] ON[90] ONB[90] ON[91] ONB[91] ON[92] ONB[92] ON[93] ONB[93] ON[94] ONB[94]
+ ON[95] ONB[95] ON[96] ONB[96] ON[97] ONB[97] ON[98] ONB[98] ON[99] ONB[99] ON[100]
+ ONB[100] ON[101] ONB[101] ON[102] ONB[102] ON[103] ONB[103] ON[104] ONB[104] ON[105]
+ ONB[105] ON[106] ONB[106] ON[107] ONB[107] ON[108] ONB[108] ON[109] ONB[109] ON[110]
+ ONB[110] ON[111] ONB[111] ON[112] ONB[112] ON[113] ONB[113] ON[114] ONB[114] ON[115]
+ ONB[115] ON[116] ONB[116] ON[117] ONB[117] ON[118] ONB[118] ON[119] ONB[119] ON[120]
+ ONB[120] ON[121] ONB[121] ON[122] ONB[122] EN[3] ENB[3] ON[123] ONB[123] ON[124]
+ ONB[124] ON[125] ONB[125] ON[126] ONB[126] ON[127] ONB[127] ON[0] ONB[0] ON[1] ONB[1]
+ ON[2] ONB[2] ON[3] ONB[3] ON[4] ONB[4] ON[5] ONB[5] ON[6] EN[0] ENB[0] ONB[6] ON[7]
+ ONB[7] ON[8] ONB[8] ON[9] ONB[9] ON[10] ONB[10] ON[11] ONB[11] ON[12] ONB[12] ON[13]
+ ONB[13] ON[14] ONB[14] ON[15] ONB[15] ON[16] ONB[16] ON[17] ONB[17] ON[18] ONB[18]
+ ON[19] ONB[19] ON[20] ONB[20] ON[21] ONB[21] ON[22] ONB[22] ON[23] ONB[23] ON[24]
+ ONB[24] ON[25] ONB[25] ON[26] ONB[26] ON[27] ONB[27] ON[28] ONB[28] ON[29] ONB[29]
+ ON[30] ONB[30] ON[31] ONB[31] ON[33] ONB[33] ON[32] ONB[32] ON[34] ONB[34] ON[35]
+ ONB[35] ON[36] ONB[36] ON[37] ONB[37] ON[38] ONB[38] ON[39] ONB[39] ON[40] ONB[40]
+ ON[41] ONB[41] ON[42] ONB[42] ON[43] ONB[43] ON[44] ONB[44] ON[45] ONB[45] ON[46]
+ ONB[46] ON[47] ONB[47] ON[48] ONB[48] ON[49] ONB[49] ON[50] ONB[50] ON[51] ONB[51]
+ ON[52] ONB[52] ON[53] ONB[53] ON[54] ONB[54] ON[55] ONB[55] ON[56] ONB[56] ON[57]
+ ONB[57] ON[58] ONB[58] ON[59] ONB[59] ON[60] ONB[60] ON[61] ONB[61] ON[62] ONB[62]
+ ON[63] ONB[63] EN[1] ENB[1] VSS VDD
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

.subckt heichips25_pudding VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_266 VPWR VGND sg13g2_decap_8
XFILLER_28_918 VPWR VGND sg13g2_fill_1
XFILLER_27_406 VPWR VGND sg13g2_decap_8
X_2106_ _0924_ net119 state\[26\] VPWR VGND sg13g2_nand2_1
X_2037_ VPWR VGND _0885_ net71 _0884_ _0154_ _0379_ net25 sg13g2_a221oi_1
XFILLER_22_144 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_19_907 VPWR VGND sg13g2_fill_2
XFILLER_18_406 VPWR VGND sg13g2_decap_8
XFILLER_46_715 VPWR VGND sg13g2_fill_1
XFILLER_19_929 VPWR VGND sg13g2_decap_8
XFILLER_45_203 VPWR VGND sg13g2_decap_8
XFILLER_42_932 VPWR VGND sg13g2_fill_2
XFILLER_27_995 VPWR VGND sg13g2_fill_2
XFILLER_26_74 VPWR VGND sg13g2_decap_8
XFILLER_26_472 VPWR VGND sg13g2_decap_8
XFILLER_42_943 VPWR VGND sg13g2_fill_2
XFILLER_13_144 VPWR VGND sg13g2_decap_8
XFILLER_14_667 VPWR VGND sg13g2_fill_1
XFILLER_9_137 VPWR VGND sg13g2_decap_8
XFILLER_42_84 VPWR VGND sg13g2_decap_8
XFILLER_5_354 VPWR VGND sg13g2_decap_8
XFILLER_1_560 VPWR VGND sg13g2_decap_8
XFILLER_3_67 VPWR VGND sg13g2_decap_8
XFILLER_49_564 VPWR VGND sg13g2_decap_8
XFILLER_37_704 VPWR VGND sg13g2_decap_4
XFILLER_36_203 VPWR VGND sg13g2_decap_8
XFILLER_18_951 VPWR VGND sg13g2_fill_1
XFILLER_44_280 VPWR VGND sg13g2_decap_8
XFILLER_32_442 VPWR VGND sg13g2_decap_8
XFILLER_20_615 VPWR VGND sg13g2_fill_2
X_1606_ net213 VPWR _0562_ VGND state\[16\] net177 sg13g2_o21ai_1
Xfanout138 net142 net138 VPWR VGND sg13g2_buf_1
Xfanout127 net136 net127 VPWR VGND sg13g2_buf_1
Xfanout116 net117 net116 VPWR VGND sg13g2_buf_1
Xfanout105 net111 net105 VPWR VGND sg13g2_buf_1
X_1537_ VPWR _0178_ daisychain\[2\] VGND sg13g2_inv_1
Xfanout149 net152 net149 VPWR VGND sg13g2_buf_1
X_1468_ VPWR _0224_ daisychain\[71\] VGND sg13g2_inv_1
X_1399_ VPWR _0031_ state\[12\] VGND sg13g2_inv_1
XFILLER_27_203 VPWR VGND sg13g2_decap_8
XFILLER_42_217 VPWR VGND sg13g2_decap_8
XFILLER_24_921 VPWR VGND sg13g2_fill_1
XFILLER_35_280 VPWR VGND sg13g2_decap_8
XFILLER_24_954 VPWR VGND sg13g2_fill_2
XFILLER_23_431 VPWR VGND sg13g2_decap_8
XFILLER_24_998 VPWR VGND sg13g2_fill_1
XFILLER_24_987 VPWR VGND sg13g2_decap_8
XFILLER_11_626 VPWR VGND sg13g2_fill_1
XFILLER_10_158 VPWR VGND sg13g2_decap_8
XFILLER_12_32 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_2_368 VPWR VGND sg13g2_decap_8
X_2400__304 VPWR VGND net303 sg13g2_tiehi
XFILLER_18_214 VPWR VGND sg13g2_decap_8
XFILLER_37_84 VPWR VGND sg13g2_decap_8
XFILLER_14_431 VPWR VGND sg13g2_decap_8
XFILLER_33_228 VPWR VGND sg13g2_decap_8
XFILLER_26_291 VPWR VGND sg13g2_decap_8
XFILLER_14_497 VPWR VGND sg13g2_decap_8
XFILLER_41_294 VPWR VGND sg13g2_decap_8
XFILLER_30_979 VPWR VGND sg13g2_decap_4
XFILLER_10_692 VPWR VGND sg13g2_fill_2
X_2440_ net476 VGND VPWR _0386_ state\[2\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_5_151 VPWR VGND sg13g2_decap_8
X_2371_ net361 VGND VPWR _0317_ daisychain\[61\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1322_ VPWR _0115_ state\[89\] VGND sg13g2_inv_1
XFILLER_49_361 VPWR VGND sg13g2_decap_8
XFILLER_37_534 VPWR VGND sg13g2_decap_4
XFILLER_37_501 VPWR VGND sg13g2_decap_8
XFILLER_17_280 VPWR VGND sg13g2_decap_8
XFILLER_18_792 VPWR VGND sg13g2_fill_1
XFILLER_24_228 VPWR VGND sg13g2_decap_8
XFILLER_21_924 VPWR VGND sg13g2_decap_4
XFILLER_28_556 VPWR VGND sg13g2_decap_8
XFILLER_43_526 VPWR VGND sg13g2_decap_8
XFILLER_15_228 VPWR VGND sg13g2_decap_8
XFILLER_11_445 VPWR VGND sg13g2_decap_8
XFILLER_8_939 VPWR VGND sg13g2_fill_1
XFILLER_8_906 VPWR VGND sg13g2_fill_1
XFILLER_23_53 VPWR VGND sg13g2_decap_8
XFILLER_7_427 VPWR VGND sg13g2_decap_8
X_2428__248 VPWR VGND net247 sg13g2_tiehi
XFILLER_3_622 VPWR VGND sg13g2_decap_8
XFILLER_2_165 VPWR VGND sg13g2_decap_8
XFILLER_47_821 VPWR VGND sg13g2_fill_1
XFILLER_47_810 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_19_556 VPWR VGND sg13g2_fill_2
XFILLER_19_545 VPWR VGND sg13g2_decap_8
XFILLER_46_364 VPWR VGND sg13g2_decap_8
XFILLER_34_504 VPWR VGND sg13g2_decap_8
XFILLER_19_589 VPWR VGND sg13g2_fill_2
XFILLER_19_578 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_8
X_1940_ VGND VPWR net133 daisychain\[98\] _0813_ net46 sg13g2_a21oi_1
XFILLER_42_581 VPWR VGND sg13g2_decap_4
X_1871_ net172 _0236_ _0760_ _0761_ VPWR VGND sg13g2_a21o_1
XFILLER_9_88 VPWR VGND sg13g2_decap_8
XFILLER_30_776 VPWR VGND sg13g2_decap_4
XFILLER_7_983 VPWR VGND sg13g2_decap_8
X_2423_ net257 VGND VPWR _0369_ daisychain\[113\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2354_ net395 VGND VPWR _0300_ daisychain\[44\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1305_ VPWR _0007_ state\[106\] VGND sg13g2_inv_1
X_2285_ VGND VPWR _0860_ _1013_ _0499_ net87 sg13g2_a21oi_1
XFILLER_37_364 VPWR VGND sg13g2_decap_8
XFILLER_33_570 VPWR VGND sg13g2_fill_2
XFILLER_20_242 VPWR VGND sg13g2_decap_8
XFILLER_21_798 VPWR VGND sg13g2_decap_4
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_18_53 VPWR VGND sg13g2_decap_8
XFILLER_43_301 VPWR VGND sg13g2_decap_8
XFILLER_28_375 VPWR VGND sg13g2_decap_8
XFILLER_31_518 VPWR VGND sg13g2_decap_8
XFILLER_43_378 VPWR VGND sg13g2_decap_8
XFILLER_34_74 VPWR VGND sg13g2_decap_8
XFILLER_11_242 VPWR VGND sg13g2_decap_8
XFILLER_7_224 VPWR VGND sg13g2_decap_8
XFILLER_3_496 VPWR VGND sg13g2_decap_8
X_2070_ _0906_ net137 state\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_19_375 VPWR VGND sg13g2_decap_8
XFILLER_46_161 VPWR VGND sg13g2_decap_8
XFILLER_34_312 VPWR VGND sg13g2_decap_8
XFILLER_34_389 VPWR VGND sg13g2_decap_8
X_1923_ net177 _0250_ _0799_ _0800_ VPWR VGND sg13g2_a21o_1
X_1854_ net224 VPWR _0748_ VGND state\[78\] net196 sg13g2_o21ai_1
XFILLER_30_584 VPWR VGND sg13g2_fill_2
X_1785_ VPWR VGND _0696_ net98 _0695_ _0212_ _0316_ net56 sg13g2_a221oi_1
X_2406_ net291 VGND VPWR _0352_ daisychain\[96\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2337_ net429 VGND VPWR _0283_ daisychain\[27\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2268_ _1005_ net131 state\[107\] VPWR VGND sg13g2_nand2_1
X_2199_ VGND VPWR _0731_ _0970_ _0456_ net108 sg13g2_a21oi_1
XFILLER_37_161 VPWR VGND sg13g2_decap_8
XFILLER_25_312 VPWR VGND sg13g2_decap_8
XFILLER_40_315 VPWR VGND sg13g2_decap_8
XFILLER_25_389 VPWR VGND sg13g2_decap_8
XFILLER_21_551 VPWR VGND sg13g2_decap_8
XFILLER_4_249 VPWR VGND sg13g2_decap_8
XFILLER_20_32 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_48_448 VPWR VGND sg13g2_decap_8
XFILLER_29_74 VPWR VGND sg13g2_decap_8
XFILLER_16_312 VPWR VGND sg13g2_decap_8
XFILLER_29_684 VPWR VGND sg13g2_decap_8
XFILLER_28_172 VPWR VGND sg13g2_decap_8
XFILLER_16_389 VPWR VGND sg13g2_decap_8
XFILLER_45_84 VPWR VGND sg13g2_decap_8
XFILLER_43_175 VPWR VGND sg13g2_decap_8
XFILLER_31_326 VPWR VGND sg13g2_decap_8
XFILLER_8_544 VPWR VGND sg13g2_decap_8
XANTENNA_5 VPWR VGND _0150_ sg13g2_antennanp
X_1570_ net205 VPWR _0535_ VGND state\[7\] net160 sg13g2_o21ai_1
XFILLER_6_67 VPWR VGND sg13g2_decap_8
XFILLER_6_1027 VPWR VGND sg13g2_fill_2
XFILLER_20_4 VPWR VGND sg13g2_decap_8
X_2122_ _0932_ net117 state\[34\] VPWR VGND sg13g2_nand2_1
XFILLER_26_109 VPWR VGND sg13g2_decap_8
XFILLER_19_172 VPWR VGND sg13g2_decap_8
X_2053_ VPWR VGND _0897_ net69 _0896_ _0158_ _0383_ net26 sg13g2_a221oi_1
XFILLER_35_643 VPWR VGND sg13g2_fill_2
XFILLER_35_676 VPWR VGND sg13g2_decap_8
XFILLER_34_186 VPWR VGND sg13g2_decap_8
XFILLER_22_326 VPWR VGND sg13g2_decap_8
X_1906_ net223 VPWR _0787_ VGND state\[91\] net198 sg13g2_o21ai_1
X_2487__289 VPWR VGND net288 sg13g2_tiehi
XFILLER_31_893 VPWR VGND sg13g2_fill_1
X_1837_ VPWR VGND _0735_ net109 _0734_ _0226_ _0329_ net66 sg13g2_a221oi_1
X_1768_ VGND VPWR net145 daisychain\[55\] _0684_ net53 sg13g2_a21oi_1
X_1699_ net195 _0188_ _0631_ _0632_ VPWR VGND sg13g2_a21o_1
XFILLER_26_665 VPWR VGND sg13g2_decap_8
XFILLER_15_32 VPWR VGND sg13g2_decap_8
XFILLER_41_602 VPWR VGND sg13g2_fill_2
XFILLER_26_687 VPWR VGND sg13g2_decap_8
XFILLER_13_326 VPWR VGND sg13g2_decap_8
XFILLER_40_112 VPWR VGND sg13g2_decap_8
XFILLER_25_186 VPWR VGND sg13g2_decap_8
XFILLER_9_319 VPWR VGND sg13g2_decap_8
XFILLER_40_189 VPWR VGND sg13g2_decap_8
XFILLER_22_882 VPWR VGND sg13g2_decap_4
XFILLER_31_53 VPWR VGND sg13g2_decap_8
XFILLER_5_569 VPWR VGND sg13g2_decap_8
Xoutput20 net20 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_49_713 VPWR VGND sg13g2_decap_8
XFILLER_49_768 VPWR VGND sg13g2_fill_1
XdigitalenH.g\[1\].u.inv1 VPWR digitalenH.g\[1\].u.OUTN net7 VGND sg13g2_inv_1
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_45_941 VPWR VGND sg13g2_fill_1
XFILLER_45_930 VPWR VGND sg13g2_decap_8
XFILLER_44_462 VPWR VGND sg13g2_decap_4
XFILLER_16_186 VPWR VGND sg13g2_decap_8
XFILLER_31_123 VPWR VGND sg13g2_decap_8
X_1622_ net207 VPWR _0574_ VGND state\[20\] net165 sg13g2_o21ai_1
XFILLER_8_396 VPWR VGND sg13g2_decap_8
X_1553_ VPWR VGND _0522_ net80 _0521_ _0178_ _0258_ net34 sg13g2_a221oi_1
X_1484_ VPWR _0206_ daisychain\[55\] VGND sg13g2_inv_1
XFILLER_39_245 VPWR VGND sg13g2_decap_8
X_2105_ VGND VPWR _0590_ _0923_ _0409_ net102 sg13g2_a21oi_1
X_2036_ VGND VPWR net115 daisychain\[122\] _0885_ net25 sg13g2_a21oi_1
XFILLER_35_473 VPWR VGND sg13g2_decap_8
XFILLER_35_451 VPWR VGND sg13g2_decap_8
XFILLER_23_646 VPWR VGND sg13g2_decap_8
XFILLER_22_123 VPWR VGND sg13g2_decap_8
X_2361__382 VPWR VGND net381 sg13g2_tiehi
XFILLER_46_749 VPWR VGND sg13g2_decap_8
XFILLER_45_259 VPWR VGND sg13g2_decap_8
XFILLER_26_53 VPWR VGND sg13g2_decap_8
XFILLER_13_123 VPWR VGND sg13g2_decap_8
XFILLER_14_679 VPWR VGND sg13g2_fill_1
XFILLER_9_116 VPWR VGND sg13g2_decap_8
XFILLER_42_999 VPWR VGND sg13g2_decap_4
XFILLER_41_476 VPWR VGND sg13g2_decap_4
XFILLER_42_63 VPWR VGND sg13g2_decap_8
XFILLER_6_867 VPWR VGND sg13g2_fill_2
XFILLER_5_333 VPWR VGND sg13g2_decap_8
X_2407__290 VPWR VGND net289 sg13g2_tiehi
XFILLER_3_46 VPWR VGND sg13g2_decap_8
XFILLER_49_543 VPWR VGND sg13g2_fill_1
XFILLER_3_1008 VPWR VGND sg13g2_fill_1
XFILLER_18_930 VPWR VGND sg13g2_fill_1
XFILLER_36_259 VPWR VGND sg13g2_decap_8
XFILLER_18_985 VPWR VGND sg13g2_fill_1
XFILLER_32_410 VPWR VGND sg13g2_decap_8
XFILLER_8_193 VPWR VGND sg13g2_decap_8
X_1605_ VPWR VGND _0561_ net76 _0560_ _0162_ _0271_ net30 sg13g2_a221oi_1
X_1536_ VPWR _0189_ daisychain\[3\] VGND sg13g2_inv_1
Xfanout128 net130 net128 VPWR VGND sg13g2_buf_1
Xfanout117 net122 net117 VPWR VGND sg13g2_buf_1
Xfanout106 net110 net106 VPWR VGND sg13g2_buf_1
Xfanout139 net142 net139 VPWR VGND sg13g2_buf_1
X_1467_ VPWR _0225_ daisychain\[72\] VGND sg13g2_inv_1
X_1398_ VPWR _0032_ state\[13\] VGND sg13g2_inv_1
XFILLER_27_259 VPWR VGND sg13g2_decap_8
X_2019_ net173 _0149_ _0871_ _0872_ VPWR VGND sg13g2_a21o_1
XFILLER_24_933 VPWR VGND sg13g2_fill_1
XFILLER_23_410 VPWR VGND sg13g2_decap_8
XFILLER_23_476 VPWR VGND sg13g2_decap_8
XFILLER_10_137 VPWR VGND sg13g2_decap_8
XFILLER_12_11 VPWR VGND sg13g2_decap_8
XFILLER_12_88 VPWR VGND sg13g2_decap_8
XFILLER_3_815 VPWR VGND sg13g2_decap_8
XFILLER_2_347 VPWR VGND sg13g2_decap_8
XFILLER_37_63 VPWR VGND sg13g2_decap_8
XFILLER_33_207 VPWR VGND sg13g2_decap_8
XFILLER_14_410 VPWR VGND sg13g2_decap_8
XFILLER_26_270 VPWR VGND sg13g2_decap_8
XFILLER_30_914 VPWR VGND sg13g2_decap_8
XFILLER_41_273 VPWR VGND sg13g2_decap_8
X_2548__267 VPWR VGND net266 sg13g2_tiehi
XFILLER_5_130 VPWR VGND sg13g2_decap_8
X_2370_ net363 VGND VPWR _0316_ daisychain\[60\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1321_ VPWR _0117_ state\[90\] VGND sg13g2_inv_1
XFILLER_2_881 VPWR VGND sg13g2_decap_8
XFILLER_49_340 VPWR VGND sg13g2_decap_8
XFILLER_37_557 VPWR VGND sg13g2_decap_8
XFILLER_24_207 VPWR VGND sg13g2_decap_8
XFILLER_21_903 VPWR VGND sg13g2_decap_8
XFILLER_32_284 VPWR VGND sg13g2_decap_8
XFILLER_20_424 VPWR VGND sg13g2_decap_8
XFILLER_9_480 VPWR VGND sg13g2_decap_8
XFILLER_0_807 VPWR VGND sg13g2_decap_8
X_2499_ net240 VGND VPWR _0445_ state\[61\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1519_ VPWR _0168_ daisychain\[20\] VGND sg13g2_inv_1
XFILLER_15_207 VPWR VGND sg13g2_decap_8
XFILLER_16_708 VPWR VGND sg13g2_fill_2
XFILLER_43_505 VPWR VGND sg13g2_decap_8
XFILLER_11_424 VPWR VGND sg13g2_decap_8
XFILLER_7_406 VPWR VGND sg13g2_decap_8
XFILLER_23_32 VPWR VGND sg13g2_decap_8
XFILLER_23_284 VPWR VGND sg13g2_decap_8
XFILLER_3_601 VPWR VGND sg13g2_decap_8
XFILLER_2_144 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_46_343 VPWR VGND sg13g2_decap_8
XFILLER_47_877 VPWR VGND sg13g2_decap_4
XFILLER_14_284 VPWR VGND sg13g2_decap_8
X_1870_ net211 VPWR _0760_ VGND state\[82\] net172 sg13g2_o21ai_1
XFILLER_9_67 VPWR VGND sg13g2_decap_8
XFILLER_7_962 VPWR VGND sg13g2_decap_8
XFILLER_7_940 VPWR VGND sg13g2_decap_4
XFILLER_6_494 VPWR VGND sg13g2_decap_8
X_2422_ net259 VGND VPWR _0368_ daisychain\[112\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2353_ net397 VGND VPWR _0299_ daisychain\[43\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1304_ VPWR _0008_ state\[107\] VGND sg13g2_inv_1
X_2284_ _1013_ net131 state\[115\] VPWR VGND sg13g2_nand2_1
XFILLER_37_343 VPWR VGND sg13g2_decap_8
XFILLER_25_516 VPWR VGND sg13g2_decap_8
XFILLER_40_519 VPWR VGND sg13g2_decap_8
XFILLER_21_700 VPWR VGND sg13g2_decap_8
XFILLER_20_221 VPWR VGND sg13g2_decap_8
X_1999_ net171 _0144_ _0856_ _0857_ VPWR VGND sg13g2_a21o_1
XFILLER_20_298 VPWR VGND sg13g2_decap_8
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_18_32 VPWR VGND sg13g2_decap_8
XFILLER_29_844 VPWR VGND sg13g2_decap_8
XFILLER_29_833 VPWR VGND sg13g2_fill_2
XFILLER_16_516 VPWR VGND sg13g2_decap_8
XFILLER_28_354 VPWR VGND sg13g2_decap_8
XFILLER_43_357 VPWR VGND sg13g2_decap_8
XFILLER_34_53 VPWR VGND sg13g2_decap_8
XFILLER_24_582 VPWR VGND sg13g2_fill_1
XFILLER_11_221 VPWR VGND sg13g2_decap_8
XFILLER_7_203 VPWR VGND sg13g2_decap_8
XFILLER_11_298 VPWR VGND sg13g2_decap_8
XFILLER_4_932 VPWR VGND sg13g2_fill_2
XFILLER_3_475 VPWR VGND sg13g2_decap_8
XFILLER_19_354 VPWR VGND sg13g2_decap_8
XFILLER_46_140 VPWR VGND sg13g2_decap_8
XFILLER_34_368 VPWR VGND sg13g2_decap_8
XFILLER_15_571 VPWR VGND sg13g2_decap_8
XFILLER_15_582 VPWR VGND sg13g2_fill_2
X_1922_ net214 VPWR _0799_ VGND state\[95\] net177 sg13g2_o21ai_1
X_1853_ VPWR VGND _0747_ net108 _0746_ _0230_ _0333_ net65 sg13g2_a221oi_1
X_1784_ VGND VPWR net143 daisychain\[59\] _0696_ net56 sg13g2_a21oi_1
XFILLER_7_792 VPWR VGND sg13g2_decap_8
XFILLER_6_291 VPWR VGND sg13g2_decap_8
X_2405_ net293 VGND VPWR _0351_ daisychain\[95\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_41_0 VPWR VGND sg13g2_decap_8
X_2336_ net431 VGND VPWR _0282_ daisychain\[26\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2267_ VGND VPWR _0833_ _1004_ _0490_ net88 sg13g2_a21oi_1
X_2320__464 VPWR VGND net463 sg13g2_tiehi
XFILLER_38_652 VPWR VGND sg13g2_fill_2
XFILLER_37_140 VPWR VGND sg13g2_decap_8
X_2198_ _0970_ net155 state\[72\] VPWR VGND sg13g2_nand2_1
XFILLER_26_847 VPWR VGND sg13g2_decap_8
XFILLER_26_858 VPWR VGND sg13g2_fill_1
XFILLER_25_368 VPWR VGND sg13g2_decap_8
XFILLER_21_541 VPWR VGND sg13g2_fill_1
XFILLER_5_729 VPWR VGND sg13g2_decap_8
XFILLER_4_228 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_1_902 VPWR VGND sg13g2_fill_1
XFILLER_20_88 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_1_957 VPWR VGND sg13g2_decap_4
XFILLER_49_939 VPWR VGND sg13g2_decap_8
XFILLER_48_427 VPWR VGND sg13g2_decap_8
XFILLER_29_53 VPWR VGND sg13g2_decap_8
XFILLER_29_630 VPWR VGND sg13g2_decap_8
XFILLER_44_622 VPWR VGND sg13g2_fill_1
XFILLER_44_600 VPWR VGND sg13g2_decap_8
XFILLER_28_151 VPWR VGND sg13g2_decap_8
XFILLER_45_63 VPWR VGND sg13g2_decap_8
XFILLER_16_368 VPWR VGND sg13g2_decap_8
X_2371__362 VPWR VGND net361 sg13g2_tiehi
XFILLER_43_154 VPWR VGND sg13g2_decap_8
XFILLER_31_305 VPWR VGND sg13g2_decap_8
XFILLER_8_523 VPWR VGND sg13g2_decap_8
XANTENNA_6 VPWR VGND _0151_ sg13g2_antennanp
XFILLER_6_46 VPWR VGND sg13g2_decap_8
XFILLER_4_740 VPWR VGND sg13g2_fill_1
XFILLER_13_4 VPWR VGND sg13g2_decap_8
X_2121_ VGND VPWR _0614_ _0931_ _0417_ net78 sg13g2_a21oi_1
X_2052_ VGND VPWR net113 daisychain\[126\] _0897_ net26 sg13g2_a21oi_1
XFILLER_19_151 VPWR VGND sg13g2_decap_8
X_2417__270 VPWR VGND net269 sg13g2_tiehi
XFILLER_34_165 VPWR VGND sg13g2_decap_8
XFILLER_22_305 VPWR VGND sg13g2_decap_8
XFILLER_31_850 VPWR VGND sg13g2_decap_8
X_1905_ VPWR VGND _0786_ net104 _0785_ _0245_ _0346_ net59 sg13g2_a221oi_1
XFILLER_30_382 VPWR VGND sg13g2_decap_8
X_1836_ VGND VPWR net156 daisychain\[72\] _0735_ net66 sg13g2_a21oi_1
X_1767_ net189 _0207_ _0682_ _0683_ VPWR VGND sg13g2_a21o_1
X_1698_ net223 VPWR _0631_ VGND state\[39\] net195 sg13g2_o21ai_1
X_2319_ net465 VGND VPWR _0265_ daisychain\[9\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_13_305 VPWR VGND sg13g2_decap_8
XFILLER_15_11 VPWR VGND sg13g2_decap_8
XFILLER_25_165 VPWR VGND sg13g2_decap_8
XFILLER_15_88 VPWR VGND sg13g2_decap_8
XFILLER_40_168 VPWR VGND sg13g2_decap_8
XFILLER_22_861 VPWR VGND sg13g2_decap_8
XFILLER_21_382 VPWR VGND sg13g2_decap_8
XFILLER_31_32 VPWR VGND sg13g2_decap_8
XFILLER_5_548 VPWR VGND sg13g2_decap_8
Xoutput10 net10 uio_out[2] VPWR VGND sg13g2_buf_1
Xoutput21 net21 uo_out[5] VPWR VGND sg13g2_buf_1
Xoutput8 net8 uio_out[0] VPWR VGND sg13g2_buf_1
XFILLER_0_231 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XdigitalenH.g\[1\].u.inv2 VPWR digitalenH.g\[1\].u.OUTP digitalenH.g\[1\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_17_600 VPWR VGND sg13g2_fill_1
XFILLER_44_441 VPWR VGND sg13g2_decap_8
XFILLER_16_165 VPWR VGND sg13g2_decap_8
XFILLER_44_485 VPWR VGND sg13g2_fill_1
XFILLER_31_102 VPWR VGND sg13g2_decap_8
XFILLER_12_382 VPWR VGND sg13g2_decap_8
XFILLER_31_179 VPWR VGND sg13g2_decap_8
XFILLER_40_691 VPWR VGND sg13g2_decap_4
X_1621_ VPWR VGND _0573_ net84 _0572_ _0166_ _0275_ net41 sg13g2_a221oi_1
XFILLER_8_375 VPWR VGND sg13g2_decap_8
X_1552_ VGND VPWR net124 daisychain\[1\] _0522_ net34 sg13g2_a21oi_1
X_1483_ VPWR _0207_ daisychain\[56\] VGND sg13g2_inv_1
XFILLER_4_581 VPWR VGND sg13g2_decap_8
XFILLER_39_224 VPWR VGND sg13g2_decap_8
X_2104_ _0923_ net140 state\[25\] VPWR VGND sg13g2_nand2_1
X_2035_ net160 _0154_ _0883_ _0884_ VPWR VGND sg13g2_a21o_1
XFILLER_35_430 VPWR VGND sg13g2_fill_2
XFILLER_23_603 VPWR VGND sg13g2_fill_1
XFILLER_22_102 VPWR VGND sg13g2_decap_8
XFILLER_10_319 VPWR VGND sg13g2_decap_8
XFILLER_22_179 VPWR VGND sg13g2_decap_8
X_1819_ net202 _0221_ _0721_ _0722_ VPWR VGND sg13g2_a21o_1
XFILLER_2_529 VPWR VGND sg13g2_decap_8
XFILLER_46_706 VPWR VGND sg13g2_decap_8
XFILLER_19_909 VPWR VGND sg13g2_fill_1
XFILLER_45_238 VPWR VGND sg13g2_decap_8
XFILLER_26_32 VPWR VGND sg13g2_decap_8
XFILLER_42_923 VPWR VGND sg13g2_decap_4
XFILLER_13_102 VPWR VGND sg13g2_decap_8
XFILLER_42_945 VPWR VGND sg13g2_fill_1
XFILLER_42_967 VPWR VGND sg13g2_fill_1
XFILLER_13_179 VPWR VGND sg13g2_decap_8
XFILLER_42_42 VPWR VGND sg13g2_decap_8
XFILLER_5_312 VPWR VGND sg13g2_decap_8
XFILLER_5_389 VPWR VGND sg13g2_decap_8
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_49_522 VPWR VGND sg13g2_decap_8
XFILLER_1_595 VPWR VGND sg13g2_decap_8
XFILLER_18_964 VPWR VGND sg13g2_fill_1
XFILLER_36_238 VPWR VGND sg13g2_decap_8
XFILLER_45_761 VPWR VGND sg13g2_fill_1
XFILLER_32_477 VPWR VGND sg13g2_fill_1
XFILLER_9_684 VPWR VGND sg13g2_decap_8
XFILLER_8_172 VPWR VGND sg13g2_decap_8
X_1604_ VGND VPWR net119 daisychain\[14\] _0561_ net30 sg13g2_a21oi_1
X_1535_ VPWR _0200_ daisychain\[4\] VGND sg13g2_inv_1
Xfanout129 net130 net129 VPWR VGND sg13g2_buf_1
Xfanout118 net121 net118 VPWR VGND sg13g2_buf_1
Xfanout107 net110 net107 VPWR VGND sg13g2_buf_1
X_1466_ VPWR _0226_ daisychain\[73\] VGND sg13g2_inv_1
X_1397_ VPWR _0033_ state\[14\] VGND sg13g2_inv_1
XFILLER_27_238 VPWR VGND sg13g2_decap_8
X_2018_ net217 VPWR _0871_ VGND state\[119\] net173 sg13g2_o21ai_1
XFILLER_24_912 VPWR VGND sg13g2_decap_8
XFILLER_10_116 VPWR VGND sg13g2_decap_8
XFILLER_6_109 VPWR VGND sg13g2_decap_8
XFILLER_12_67 VPWR VGND sg13g2_decap_8
XFILLER_2_326 VPWR VGND sg13g2_decap_8
XFILLER_37_42 VPWR VGND sg13g2_decap_8
XFILLER_18_249 VPWR VGND sg13g2_decap_8
XFILLER_46_547 VPWR VGND sg13g2_fill_2
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_42_742 VPWR VGND sg13g2_decap_8
XFILLER_42_775 VPWR VGND sg13g2_fill_2
XFILLER_41_252 VPWR VGND sg13g2_decap_8
XFILLER_5_186 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
X_1320_ VPWR _0118_ state\[91\] VGND sg13g2_inv_1
XFILLER_2_860 VPWR VGND sg13g2_decap_8
XFILLER_1_392 VPWR VGND sg13g2_decap_8
XFILLER_49_396 VPWR VGND sg13g2_decap_8
XFILLER_18_761 VPWR VGND sg13g2_fill_1
XFILLER_32_263 VPWR VGND sg13g2_decap_8
XFILLER_20_403 VPWR VGND sg13g2_decap_8
XFILLER_20_469 VPWR VGND sg13g2_decap_8
X_2498_ net244 VGND VPWR _0444_ state\[60\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1518_ VPWR _0169_ daisychain\[21\] VGND sg13g2_inv_1
X_1449_ VPWR _0245_ daisychain\[90\] VGND sg13g2_inv_1
XFILLER_28_503 VPWR VGND sg13g2_decap_8
XFILLER_28_536 VPWR VGND sg13g2_decap_4
XFILLER_43_517 VPWR VGND sg13g2_decap_4
XFILLER_11_403 VPWR VGND sg13g2_decap_8
XFILLER_23_263 VPWR VGND sg13g2_decap_8
XFILLER_23_11 VPWR VGND sg13g2_decap_8
X_2330__444 VPWR VGND net443 sg13g2_tiehi
XFILLER_8_919 VPWR VGND sg13g2_fill_1
XFILLER_23_88 VPWR VGND sg13g2_decap_8
XFILLER_3_668 VPWR VGND sg13g2_fill_1
XFILLER_3_657 VPWR VGND sg13g2_decap_8
XFILLER_2_123 VPWR VGND sg13g2_decap_8
XFILLER_24_1021 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_19_503 VPWR VGND sg13g2_fill_2
XFILLER_46_322 VPWR VGND sg13g2_decap_8
XFILLER_46_399 VPWR VGND sg13g2_decap_8
XFILLER_14_263 VPWR VGND sg13g2_decap_8
XFILLER_9_46 VPWR VGND sg13g2_decap_8
XFILLER_10_480 VPWR VGND sg13g2_decap_8
X_2381__342 VPWR VGND net341 sg13g2_tiehi
XFILLER_6_473 VPWR VGND sg13g2_decap_8
X_2421_ net261 VGND VPWR _0367_ daisychain\[111\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2352_ net399 VGND VPWR _0298_ daisychain\[42\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2283_ VGND VPWR _0857_ _1012_ _0498_ net81 sg13g2_a21oi_1
X_1303_ VPWR _0009_ state\[108\] VGND sg13g2_inv_1
XFILLER_49_193 VPWR VGND sg13g2_decap_8
XFILLER_37_322 VPWR VGND sg13g2_decap_8
XFILLER_18_580 VPWR VGND sg13g2_decap_4
XFILLER_37_399 VPWR VGND sg13g2_decap_8
XFILLER_20_200 VPWR VGND sg13g2_decap_8
X_1998_ net212 VPWR _0856_ VGND state\[114\] net171 sg13g2_o21ai_1
XFILLER_20_277 VPWR VGND sg13g2_decap_8
X_2427__250 VPWR VGND net249 sg13g2_tiehi
XFILLER_47_1010 VPWR VGND sg13g2_fill_2
XFILLER_0_616 VPWR VGND sg13g2_decap_8
XFILLER_47_119 VPWR VGND sg13g2_decap_8
XFILLER_18_11 VPWR VGND sg13g2_decap_8
XFILLER_28_333 VPWR VGND sg13g2_decap_8
X_2358__388 VPWR VGND net387 sg13g2_tiehi
XFILLER_29_889 VPWR VGND sg13g2_fill_2
XFILLER_18_88 VPWR VGND sg13g2_decap_8
X_2512__407 VPWR VGND net406 sg13g2_tiehi
XFILLER_44_848 VPWR VGND sg13g2_fill_2
X_2551__467 VPWR VGND net466 sg13g2_tiehi
XFILLER_43_336 VPWR VGND sg13g2_decap_8
XFILLER_12_701 VPWR VGND sg13g2_fill_1
XFILLER_34_32 VPWR VGND sg13g2_decap_8
XFILLER_11_200 VPWR VGND sg13g2_decap_8
XFILLER_12_723 VPWR VGND sg13g2_decap_8
XFILLER_8_716 VPWR VGND sg13g2_decap_8
XFILLER_11_277 VPWR VGND sg13g2_decap_8
XFILLER_7_259 VPWR VGND sg13g2_decap_8
XFILLER_3_421 VPWR VGND sg13g2_fill_1
XFILLER_3_410 VPWR VGND sg13g2_decap_8
XFILLER_4_977 VPWR VGND sg13g2_fill_1
XFILLER_3_454 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_38_119 VPWR VGND sg13g2_decap_8
XFILLER_19_333 VPWR VGND sg13g2_decap_8
XFILLER_47_675 VPWR VGND sg13g2_fill_2
XFILLER_46_196 VPWR VGND sg13g2_decap_8
XFILLER_34_347 VPWR VGND sg13g2_decap_8
XFILLER_15_550 VPWR VGND sg13g2_decap_8
X_1921_ VPWR VGND _0798_ net89 _0797_ _0249_ _0350_ net47 sg13g2_a221oi_1
X_1852_ VGND VPWR net155 daisychain\[76\] _0747_ net65 sg13g2_a21oi_1
X_1783_ net189 _0212_ _0694_ _0695_ VPWR VGND sg13g2_a21o_1
XFILLER_6_270 VPWR VGND sg13g2_decap_8
X_2404_ net295 VGND VPWR _0350_ daisychain\[94\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2335_ net433 VGND VPWR _0281_ daisychain\[25\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2266_ _1004_ net132 state\[106\] VPWR VGND sg13g2_nand2_1
X_2197_ VGND VPWR _0728_ _0969_ _0455_ net105 sg13g2_a21oi_1
XFILLER_26_815 VPWR VGND sg13g2_decap_8
XFILLER_38_686 VPWR VGND sg13g2_fill_2
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_37_196 VPWR VGND sg13g2_decap_8
XFILLER_25_347 VPWR VGND sg13g2_decap_8
XFILLER_4_207 VPWR VGND sg13g2_decap_8
XFILLER_20_67 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_49_907 VPWR VGND sg13g2_decap_8
XFILLER_48_406 VPWR VGND sg13g2_decap_4
XFILLER_29_32 VPWR VGND sg13g2_decap_8
XFILLER_29_664 VPWR VGND sg13g2_decap_4
XFILLER_28_130 VPWR VGND sg13g2_decap_8
XFILLER_16_347 VPWR VGND sg13g2_decap_8
XFILLER_45_42 VPWR VGND sg13g2_decap_8
XFILLER_43_133 VPWR VGND sg13g2_decap_8
XFILLER_25_881 VPWR VGND sg13g2_decap_8
XFILLER_12_542 VPWR VGND sg13g2_decap_8
XFILLER_8_502 VPWR VGND sg13g2_decap_8
XFILLER_12_575 VPWR VGND sg13g2_decap_8
XFILLER_8_579 VPWR VGND sg13g2_decap_8
XFILLER_6_25 VPWR VGND sg13g2_decap_8
XANTENNA_7 VPWR VGND _0151_ sg13g2_antennanp
XFILLER_4_796 VPWR VGND sg13g2_fill_2
XFILLER_3_284 VPWR VGND sg13g2_decap_8
XFILLER_39_406 VPWR VGND sg13g2_decap_4
XFILLER_0_980 VPWR VGND sg13g2_decap_8
X_2120_ _0931_ net122 state\[33\] VPWR VGND sg13g2_nand2_1
XFILLER_19_130 VPWR VGND sg13g2_decap_8
X_2051_ net161 _0158_ _0895_ _0896_ VPWR VGND sg13g2_a21o_1
XFILLER_47_483 VPWR VGND sg13g2_decap_8
XFILLER_34_144 VPWR VGND sg13g2_decap_8
X_1904_ VGND VPWR net150 daisychain\[89\] _0786_ net59 sg13g2_a21oi_1
XFILLER_30_361 VPWR VGND sg13g2_decap_8
X_1835_ net202 _0226_ _0733_ _0734_ VPWR VGND sg13g2_a21o_1
X_1766_ net221 VPWR _0682_ VGND state\[56\] net189 sg13g2_o21ai_1
X_1697_ VPWR VGND _0630_ net94 _0629_ _0187_ _0294_ net49 sg13g2_a221oi_1
X_2318_ net467 VGND VPWR _0264_ daisychain\[8\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2249_ VGND VPWR _0806_ _0995_ _0481_ net84 sg13g2_a21oi_1
XFILLER_25_144 VPWR VGND sg13g2_decap_8
XFILLER_15_67 VPWR VGND sg13g2_decap_8
XFILLER_40_147 VPWR VGND sg13g2_decap_8
XFILLER_21_361 VPWR VGND sg13g2_decap_8
XFILLER_31_11 VPWR VGND sg13g2_decap_8
XFILLER_5_527 VPWR VGND sg13g2_decap_8
XFILLER_31_88 VPWR VGND sg13g2_decap_8
Xoutput11 net11 uio_out[3] VPWR VGND sg13g2_buf_1
Xoutput22 net22 uo_out[6] VPWR VGND sg13g2_buf_1
Xoutput9 net9 uio_out[1] VPWR VGND sg13g2_buf_1
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_49_759 VPWR VGND sg13g2_decap_4
XFILLER_48_203 VPWR VGND sg13g2_decap_8
XFILLER_44_420 VPWR VGND sg13g2_decap_8
XFILLER_16_144 VPWR VGND sg13g2_decap_8
XFILLER_45_976 VPWR VGND sg13g2_decap_8
XFILLER_32_615 VPWR VGND sg13g2_decap_4
XFILLER_32_648 VPWR VGND sg13g2_fill_2
XFILLER_31_158 VPWR VGND sg13g2_decap_8
XFILLER_12_361 VPWR VGND sg13g2_decap_8
XFILLER_8_354 VPWR VGND sg13g2_decap_8
X_1620_ VGND VPWR net129 daisychain\[18\] _0573_ net42 sg13g2_a21oi_1
X_1551_ net160 _0178_ _0520_ _0521_ VPWR VGND sg13g2_a21o_1
XFILLER_4_560 VPWR VGND sg13g2_decap_8
X_1482_ VPWR _0208_ daisychain\[57\] VGND sg13g2_inv_1
XFILLER_39_203 VPWR VGND sg13g2_decap_8
X_2103_ VGND VPWR _0587_ _0922_ _0408_ net103 sg13g2_a21oi_1
X_2034_ net210 VPWR _0883_ VGND state\[123\] net160 sg13g2_o21ai_1
XFILLER_47_280 VPWR VGND sg13g2_decap_8
XFILLER_35_420 VPWR VGND sg13g2_fill_2
XFILLER_22_158 VPWR VGND sg13g2_decap_8
XFILLER_31_681 VPWR VGND sg13g2_fill_2
X_1818_ net226 VPWR _0721_ VGND state\[69\] net202 sg13g2_o21ai_1
X_1749_ VPWR VGND _0669_ net99 _0668_ _0202_ _0307_ net55 sg13g2_a221oi_1
XFILLER_2_508 VPWR VGND sg13g2_decap_8
XFILLER_45_217 VPWR VGND sg13g2_decap_8
XFILLER_27_921 VPWR VGND sg13g2_fill_2
XFILLER_27_910 VPWR VGND sg13g2_decap_8
XFILLER_38_280 VPWR VGND sg13g2_decap_8
XFILLER_26_431 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_27_976 VPWR VGND sg13g2_fill_1
XFILLER_14_637 VPWR VGND sg13g2_fill_1
XFILLER_26_88 VPWR VGND sg13g2_decap_8
XFILLER_13_158 VPWR VGND sg13g2_decap_8
XFILLER_42_21 VPWR VGND sg13g2_decap_8
XFILLER_6_836 VPWR VGND sg13g2_decap_8
XFILLER_42_98 VPWR VGND sg13g2_decap_8
XFILLER_5_368 VPWR VGND sg13g2_decap_8
X_2340__424 VPWR VGND net423 sg13g2_tiehi
XFILLER_49_501 VPWR VGND sg13g2_decap_8
XFILLER_1_574 VPWR VGND sg13g2_decap_8
XFILLER_49_589 VPWR VGND sg13g2_decap_8
XFILLER_36_217 VPWR VGND sg13g2_decap_8
XFILLER_17_420 VPWR VGND sg13g2_decap_8
XFILLER_17_431 VPWR VGND sg13g2_fill_1
XFILLER_18_943 VPWR VGND sg13g2_fill_1
XFILLER_29_291 VPWR VGND sg13g2_decap_8
XFILLER_44_294 VPWR VGND sg13g2_decap_8
XFILLER_32_456 VPWR VGND sg13g2_decap_8
XFILLER_32_489 VPWR VGND sg13g2_decap_8
XFILLER_8_151 VPWR VGND sg13g2_decap_8
X_1603_ net167 _0162_ _0559_ _0560_ VPWR VGND sg13g2_a21o_1
X_1534_ VPWR _0211_ daisychain\[5\] VGND sg13g2_inv_1
Xfanout119 net121 net119 VPWR VGND sg13g2_buf_1
Xfanout108 net110 net108 VPWR VGND sg13g2_buf_1
X_1465_ VPWR _0227_ daisychain\[74\] VGND sg13g2_inv_1
X_1396_ VPWR _0034_ state\[15\] VGND sg13g2_inv_1
XFILLER_27_217 VPWR VGND sg13g2_decap_8
X_2391__322 VPWR VGND net321 sg13g2_tiehi
X_2017_ VPWR VGND _0870_ net82 _0869_ _0148_ _0374_ net39 sg13g2_a221oi_1
XFILLER_35_294 VPWR VGND sg13g2_decap_8
XFILLER_23_445 VPWR VGND sg13g2_decap_8
XFILLER_12_46 VPWR VGND sg13g2_decap_8
X_2543__347 VPWR VGND net346 sg13g2_tiehi
XFILLER_2_305 VPWR VGND sg13g2_decap_8
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_18_228 VPWR VGND sg13g2_decap_8
X_2437__230 VPWR VGND net229 sg13g2_tiehi
XFILLER_37_98 VPWR VGND sg13g2_decap_8
XFILLER_42_732 VPWR VGND sg13g2_decap_4
XFILLER_14_445 VPWR VGND sg13g2_decap_8
XFILLER_14_456 VPWR VGND sg13g2_fill_2
XFILLER_41_231 VPWR VGND sg13g2_decap_8
XFILLER_30_938 VPWR VGND sg13g2_decap_8
XFILLER_10_662 VPWR VGND sg13g2_decap_4
X_2368__368 VPWR VGND net367 sg13g2_tiehi
XFILLER_6_633 VPWR VGND sg13g2_decap_8
XFILLER_6_622 VPWR VGND sg13g2_decap_8
XFILLER_5_165 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_8
XFILLER_1_371 VPWR VGND sg13g2_decap_8
XFILLER_49_375 VPWR VGND sg13g2_decap_8
XFILLER_37_515 VPWR VGND sg13g2_decap_4
XFILLER_18_773 VPWR VGND sg13g2_fill_2
XFILLER_18_784 VPWR VGND sg13g2_fill_1
XFILLER_17_294 VPWR VGND sg13g2_decap_8
XFILLER_32_242 VPWR VGND sg13g2_decap_8
X_2462__389 VPWR VGND net388 sg13g2_tiehi
X_2497_ net248 VGND VPWR _0443_ state\[59\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1517_ VPWR _0170_ daisychain\[22\] VGND sg13g2_inv_1
X_2538__427 VPWR VGND net426 sg13g2_tiehi
X_1448_ VPWR _0246_ daisychain\[91\] VGND sg13g2_inv_1
X_1379_ VPWR _0053_ state\[32\] VGND sg13g2_inv_1
XFILLER_24_710 VPWR VGND sg13g2_fill_1
XFILLER_23_242 VPWR VGND sg13g2_decap_8
XFILLER_11_459 VPWR VGND sg13g2_decap_8
XFILLER_23_67 VPWR VGND sg13g2_decap_8
XFILLER_20_982 VPWR VGND sg13g2_decap_8
XFILLER_3_636 VPWR VGND sg13g2_decap_8
XFILLER_2_102 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_179 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_46_301 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_46_378 VPWR VGND sg13g2_decap_8
XFILLER_14_242 VPWR VGND sg13g2_decap_8
XFILLER_9_25 VPWR VGND sg13g2_decap_8
XFILLER_42_573 VPWR VGND sg13g2_decap_4
XFILLER_30_702 VPWR VGND sg13g2_fill_2
Xfanout90 net91 net90 VPWR VGND sg13g2_buf_1
XFILLER_6_452 VPWR VGND sg13g2_decap_8
X_2420_ net263 VGND VPWR _0366_ daisychain\[110\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_7_997 VPWR VGND sg13g2_fill_2
X_2351_ net401 VGND VPWR _0297_ daisychain\[41\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2282_ _1012_ net125 state\[114\] VPWR VGND sg13g2_nand2_1
X_1302_ VPWR _0010_ state\[109\] VGND sg13g2_inv_1
XFILLER_2_691 VPWR VGND sg13g2_decap_8
XFILLER_49_172 VPWR VGND sg13g2_decap_8
XFILLER_37_301 VPWR VGND sg13g2_decap_8
XFILLER_37_378 VPWR VGND sg13g2_decap_8
XFILLER_21_724 VPWR VGND sg13g2_decap_8
X_1997_ VPWR VGND _0855_ net81 _0854_ _0143_ _0369_ net36 sg13g2_a221oi_1
XFILLER_20_256 VPWR VGND sg13g2_decap_8
XFILLER_47_1000 VPWR VGND sg13g2_fill_1
X_2549_ net250 VGND VPWR _0495_ state\[111\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2497__249 VPWR VGND net248 sg13g2_tiehi
XFILLER_29_835 VPWR VGND sg13g2_fill_1
XFILLER_28_312 VPWR VGND sg13g2_decap_8
XFILLER_18_67 VPWR VGND sg13g2_decap_8
XFILLER_44_816 VPWR VGND sg13g2_decap_4
XFILLER_43_315 VPWR VGND sg13g2_decap_8
XFILLER_28_389 VPWR VGND sg13g2_decap_8
XFILLER_34_11 VPWR VGND sg13g2_decap_8
XFILLER_24_573 VPWR VGND sg13g2_fill_1
XFILLER_34_88 VPWR VGND sg13g2_decap_8
XFILLER_11_256 VPWR VGND sg13g2_decap_8
XFILLER_7_238 VPWR VGND sg13g2_decap_8
XFILLER_4_934 VPWR VGND sg13g2_fill_1
XFILLER_3_433 VPWR VGND sg13g2_decap_8
XFILLER_4_989 VPWR VGND sg13g2_decap_8
XFILLER_19_312 VPWR VGND sg13g2_decap_8
XFILLER_47_621 VPWR VGND sg13g2_decap_4
XFILLER_19_389 VPWR VGND sg13g2_decap_8
XFILLER_46_175 VPWR VGND sg13g2_decap_8
XFILLER_34_326 VPWR VGND sg13g2_decap_8
X_1920_ VGND VPWR net134 daisychain\[93\] _0798_ net47 sg13g2_a21oi_1
X_1851_ net201 _0230_ _0745_ _0746_ VPWR VGND sg13g2_a21o_1
XFILLER_42_392 VPWR VGND sg13g2_decap_8
X_1782_ net222 VPWR _0694_ VGND state\[60\] net189 sg13g2_o21ai_1
XFILLER_7_783 VPWR VGND sg13g2_decap_4
X_2403_ net297 VGND VPWR _0349_ daisychain\[93\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2334_ net435 VGND VPWR _0280_ daisychain\[24\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_29_109 VPWR VGND sg13g2_decap_8
XFILLER_27_0 VPWR VGND sg13g2_decap_8
X_2265_ VGND VPWR _0830_ _1003_ _0489_ net88 sg13g2_a21oi_1
X_2196_ _0969_ net151 state\[71\] VPWR VGND sg13g2_nand2_1
XFILLER_38_654 VPWR VGND sg13g2_fill_1
XFILLER_37_175 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_25_326 VPWR VGND sg13g2_decap_8
XFILLER_40_329 VPWR VGND sg13g2_decap_8
XFILLER_21_521 VPWR VGND sg13g2_fill_2
XFILLER_20_46 VPWR VGND sg13g2_decap_8
XFILLER_29_11 VPWR VGND sg13g2_decap_8
XFILLER_0_469 VPWR VGND sg13g2_decap_8
XFILLER_29_88 VPWR VGND sg13g2_decap_8
XFILLER_45_21 VPWR VGND sg13g2_decap_8
XFILLER_29_698 VPWR VGND sg13g2_decap_8
XFILLER_16_326 VPWR VGND sg13g2_decap_8
XFILLER_43_112 VPWR VGND sg13g2_decap_8
XFILLER_28_186 VPWR VGND sg13g2_decap_8
XFILLER_45_98 VPWR VGND sg13g2_decap_8
XFILLER_12_521 VPWR VGND sg13g2_decap_8
XFILLER_43_189 VPWR VGND sg13g2_decap_8
XFILLER_8_558 VPWR VGND sg13g2_decap_8
XANTENNA_8 VPWR VGND _0159_ sg13g2_antennanp
XFILLER_4_775 VPWR VGND sg13g2_decap_8
XFILLER_3_263 VPWR VGND sg13g2_decap_8
X_2050_ net205 VPWR _0895_ VGND state\[127\] net159 sg13g2_o21ai_1
XFILLER_47_462 VPWR VGND sg13g2_decap_8
XFILLER_19_186 VPWR VGND sg13g2_decap_8
XFILLER_34_123 VPWR VGND sg13g2_decap_8
X_2350__404 VPWR VGND net403 sg13g2_tiehi
XFILLER_23_819 VPWR VGND sg13g2_fill_2
XFILLER_43_690 VPWR VGND sg13g2_fill_2
X_1903_ net195 _0245_ _0784_ _0785_ VPWR VGND sg13g2_a21o_1
XFILLER_30_340 VPWR VGND sg13g2_decap_8
X_1834_ net226 VPWR _0733_ VGND state\[73\] net202 sg13g2_o21ai_1
X_1765_ VPWR VGND _0681_ net99 _0680_ _0206_ _0311_ net53 sg13g2_a221oi_1
X_1696_ VGND VPWR net140 daisychain\[37\] _0630_ net49 sg13g2_a21oi_1
X_2317_ net469 VGND VPWR _0263_ daisychain\[7\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2248_ _0995_ net128 state\[97\] VPWR VGND sg13g2_nand2_1
X_2179_ VGND VPWR _0701_ _0960_ _0446_ net98 sg13g2_a21oi_1
XFILLER_25_123 VPWR VGND sg13g2_decap_8
XFILLER_15_46 VPWR VGND sg13g2_decap_8
XFILLER_40_126 VPWR VGND sg13g2_decap_8
XFILLER_21_340 VPWR VGND sg13g2_decap_8
XFILLER_31_67 VPWR VGND sg13g2_decap_8
Xoutput12 net12 uio_out[4] VPWR VGND sg13g2_buf_1
Xoutput23 net23 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_49_738 VPWR VGND sg13g2_decap_8
XFILLER_49_727 VPWR VGND sg13g2_fill_2
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_17_613 VPWR VGND sg13g2_decap_8
XFILLER_45_922 VPWR VGND sg13g2_fill_2
XFILLER_29_473 VPWR VGND sg13g2_decap_8
XFILLER_29_451 VPWR VGND sg13g2_decap_8
XFILLER_16_123 VPWR VGND sg13g2_decap_8
XFILLER_17_624 VPWR VGND sg13g2_fill_1
XFILLER_45_955 VPWR VGND sg13g2_decap_8
XFILLER_45_988 VPWR VGND sg13g2_decap_8
XFILLER_44_498 VPWR VGND sg13g2_decap_8
XFILLER_31_137 VPWR VGND sg13g2_decap_8
XFILLER_12_340 VPWR VGND sg13g2_decap_8
XFILLER_8_333 VPWR VGND sg13g2_decap_8
X_1550_ net205 VPWR _0520_ VGND state\[2\] net160 sg13g2_o21ai_1
X_1481_ VPWR _0209_ daisychain\[58\] VGND sg13g2_inv_1
X_2102_ _0922_ net149 state\[24\] VPWR VGND sg13g2_nand2_1
X_2378__348 VPWR VGND net347 sg13g2_tiehi
XFILLER_39_259 VPWR VGND sg13g2_decap_8
X_2033_ VPWR VGND _0882_ net70 _0881_ _0153_ _0378_ net25 sg13g2_a221oi_1
XFILLER_35_465 VPWR VGND sg13g2_fill_1
XFILLER_23_627 VPWR VGND sg13g2_decap_4
XFILLER_22_137 VPWR VGND sg13g2_decap_8
X_1817_ VPWR VGND _0720_ net108 _0719_ _0220_ _0324_ net66 sg13g2_a221oi_1
XFILLER_7_91 VPWR VGND sg13g2_decap_8
X_1748_ VGND VPWR net145 daisychain\[50\] _0669_ net55 sg13g2_a21oi_1
X_1679_ net164 _0183_ _0616_ _0617_ VPWR VGND sg13g2_a21o_1
XFILLER_26_410 VPWR VGND sg13g2_decap_8
XFILLER_27_988 VPWR VGND sg13g2_decap_8
XFILLER_41_413 VPWR VGND sg13g2_fill_2
XFILLER_26_67 VPWR VGND sg13g2_decap_8
XFILLER_13_137 VPWR VGND sg13g2_decap_8
X_2513__399 VPWR VGND net398 sg13g2_tiehi
XFILLER_42_77 VPWR VGND sg13g2_decap_8
XFILLER_6_804 VPWR VGND sg13g2_fill_1
XFILLER_5_347 VPWR VGND sg13g2_decap_8
XFILLER_1_553 VPWR VGND sg13g2_decap_8
XFILLER_49_557 VPWR VGND sg13g2_decap_8
XFILLER_18_922 VPWR VGND sg13g2_fill_1
XFILLER_18_955 VPWR VGND sg13g2_fill_2
XFILLER_29_270 VPWR VGND sg13g2_decap_8
XFILLER_17_498 VPWR VGND sg13g2_fill_2
XFILLER_44_273 VPWR VGND sg13g2_decap_8
XFILLER_32_424 VPWR VGND sg13g2_decap_4
XFILLER_8_130 VPWR VGND sg13g2_decap_8
X_1602_ net207 VPWR _0559_ VGND state\[15\] net167 sg13g2_o21ai_1
X_1533_ VPWR _0222_ daisychain\[6\] VGND sg13g2_inv_1
Xfanout109 net110 net109 VPWR VGND sg13g2_buf_1
X_1464_ VPWR _0228_ daisychain\[75\] VGND sg13g2_inv_1
X_1395_ VPWR _0035_ state\[16\] VGND sg13g2_inv_1
X_2016_ VGND VPWR net126 daisychain\[117\] _0870_ net39 sg13g2_a21oi_1
XFILLER_35_273 VPWR VGND sg13g2_decap_8
XFILLER_23_424 VPWR VGND sg13g2_decap_8
XFILLER_12_25 VPWR VGND sg13g2_decap_8
XFILLER_3_829 VPWR VGND sg13g2_decap_4
XFILLER_18_207 VPWR VGND sg13g2_decap_8
XFILLER_46_549 VPWR VGND sg13g2_fill_1
XFILLER_37_77 VPWR VGND sg13g2_decap_8
XFILLER_14_424 VPWR VGND sg13g2_decap_8
XFILLER_41_210 VPWR VGND sg13g2_decap_8
XFILLER_26_284 VPWR VGND sg13g2_decap_8
XFILLER_42_799 VPWR VGND sg13g2_fill_2
XFILLER_41_287 VPWR VGND sg13g2_decap_8
XFILLER_10_641 VPWR VGND sg13g2_decap_8
XFILLER_6_601 VPWR VGND sg13g2_fill_1
XFILLER_10_685 VPWR VGND sg13g2_decap_8
XFILLER_5_144 VPWR VGND sg13g2_decap_8
XFILLER_1_350 VPWR VGND sg13g2_decap_8
XFILLER_49_354 VPWR VGND sg13g2_decap_8
XFILLER_17_273 VPWR VGND sg13g2_decap_8
XFILLER_18_796 VPWR VGND sg13g2_fill_2
X_2490__277 VPWR VGND net276 sg13g2_tiehi
XFILLER_32_221 VPWR VGND sg13g2_decap_8
XFILLER_21_928 VPWR VGND sg13g2_fill_1
XFILLER_21_917 VPWR VGND sg13g2_decap_8
XFILLER_32_298 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_12_clk clknet_2_3__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
XFILLER_9_494 VPWR VGND sg13g2_decap_8
X_2565_ net354 VGND VPWR _0511_ state\[127\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1516_ VPWR _0171_ daisychain\[23\] VGND sg13g2_inv_1
X_2496_ net252 VGND VPWR _0442_ state\[58\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1447_ VPWR _0247_ daisychain\[92\] VGND sg13g2_inv_1
XFILLER_4_81 VPWR VGND sg13g2_decap_8
X_1378_ VPWR _0054_ state\[33\] VGND sg13g2_inv_1
XFILLER_28_549 VPWR VGND sg13g2_decap_8
XFILLER_36_560 VPWR VGND sg13g2_decap_8
XFILLER_36_582 VPWR VGND sg13g2_fill_2
XFILLER_23_221 VPWR VGND sg13g2_decap_8
XFILLER_11_438 VPWR VGND sg13g2_decap_8
XFILLER_23_46 VPWR VGND sg13g2_decap_8
XFILLER_23_298 VPWR VGND sg13g2_decap_8
XFILLER_3_615 VPWR VGND sg13g2_decap_8
XFILLER_2_158 VPWR VGND sg13g2_decap_8
X_2404__296 VPWR VGND net295 sg13g2_tiehi
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_47_847 VPWR VGND sg13g2_fill_2
XFILLER_47_825 VPWR VGND sg13g2_fill_2
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_46_357 VPWR VGND sg13g2_decap_8
XFILLER_27_571 VPWR VGND sg13g2_decap_8
XFILLER_14_221 VPWR VGND sg13g2_decap_8
XFILLER_15_733 VPWR VGND sg13g2_fill_2
XFILLER_14_298 VPWR VGND sg13g2_decap_8
Xfanout80 net81 net80 VPWR VGND sg13g2_buf_1
Xfanout91 net112 net91 VPWR VGND sg13g2_buf_1
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_7_976 VPWR VGND sg13g2_decap_8
XFILLER_6_431 VPWR VGND sg13g2_decap_8
X_2350_ net403 VGND VPWR _0296_ daisychain\[40\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2281_ VGND VPWR _0854_ _1011_ _0497_ net81 sg13g2_a21oi_1
X_1301_ VPWR _0012_ state\[110\] VGND sg13g2_inv_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
XFILLER_29_4 VPWR VGND sg13g2_decap_8
XFILLER_49_151 VPWR VGND sg13g2_decap_8
XFILLER_37_357 VPWR VGND sg13g2_decap_8
XFILLER_46_880 VPWR VGND sg13g2_decap_4
XFILLER_46_891 VPWR VGND sg13g2_fill_2
X_1996_ VGND VPWR net124 daisychain\[112\] _0855_ net36 sg13g2_a21oi_1
XFILLER_21_769 VPWR VGND sg13g2_fill_2
XFILLER_20_235 VPWR VGND sg13g2_decap_8
XFILLER_9_291 VPWR VGND sg13g2_decap_8
X_2548_ net266 VGND VPWR _0494_ state\[110\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2479_ net320 VGND VPWR _0425_ state\[41\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_18_46 VPWR VGND sg13g2_decap_8
XFILLER_29_858 VPWR VGND sg13g2_fill_2
XFILLER_28_368 VPWR VGND sg13g2_decap_8
XFILLER_34_67 VPWR VGND sg13g2_decap_8
XFILLER_11_235 VPWR VGND sg13g2_decap_8
Xclkload0 clknet_leaf_0_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_7_217 VPWR VGND sg13g2_decap_8
XFILLER_3_489 VPWR VGND sg13g2_decap_8
XFILLER_19_368 VPWR VGND sg13g2_decap_8
XFILLER_47_677 VPWR VGND sg13g2_fill_1
XFILLER_46_154 VPWR VGND sg13g2_decap_8
XFILLER_34_305 VPWR VGND sg13g2_decap_8
XFILLER_42_371 VPWR VGND sg13g2_decap_8
X_1850_ net226 VPWR _0745_ VGND state\[77\] net201 sg13g2_o21ai_1
XFILLER_30_555 VPWR VGND sg13g2_decap_4
X_1781_ VPWR VGND _0693_ net97 _0692_ _0210_ _0315_ net56 sg13g2_a221oi_1
XFILLER_7_762 VPWR VGND sg13g2_decap_8
X_2402_ net299 VGND VPWR _0348_ daisychain\[92\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2333_ net437 VGND VPWR _0279_ daisychain\[23\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2504__471 VPWR VGND net470 sg13g2_tiehi
X_2264_ _1003_ net132 state\[105\] VPWR VGND sg13g2_nand2_1
X_2195_ VGND VPWR _0725_ _0968_ _0454_ net108 sg13g2_a21oi_1
XFILLER_38_688 VPWR VGND sg13g2_fill_1
XFILLER_37_154 VPWR VGND sg13g2_decap_8
XFILLER_25_305 VPWR VGND sg13g2_decap_8
X_2357__390 VPWR VGND net389 sg13g2_tiehi
XFILLER_40_308 VPWR VGND sg13g2_decap_8
XFILLER_33_382 VPWR VGND sg13g2_decap_8
X_2388__328 VPWR VGND net327 sg13g2_tiehi
X_1979_ net176 _0138_ _0841_ _0842_ VPWR VGND sg13g2_a21o_1
XFILLER_20_25 VPWR VGND sg13g2_decap_8
XFILLER_0_448 VPWR VGND sg13g2_decap_8
XFILLER_29_67 VPWR VGND sg13g2_decap_8
XFILLER_16_305 VPWR VGND sg13g2_decap_8
XFILLER_29_677 VPWR VGND sg13g2_fill_2
XFILLER_28_165 VPWR VGND sg13g2_decap_8
X_2516__375 VPWR VGND net374 sg13g2_tiehi
XFILLER_45_77 VPWR VGND sg13g2_decap_8
XFILLER_43_168 VPWR VGND sg13g2_decap_8
XFILLER_12_500 VPWR VGND sg13g2_decap_8
XFILLER_31_319 VPWR VGND sg13g2_decap_8
XFILLER_24_382 VPWR VGND sg13g2_decap_8
XFILLER_8_537 VPWR VGND sg13g2_decap_8
XANTENNA_9 VPWR VGND _0162_ sg13g2_antennanp
XFILLER_3_242 VPWR VGND sg13g2_decap_8
XFILLER_6_1009 VPWR VGND sg13g2_fill_2
XFILLER_47_441 VPWR VGND sg13g2_decap_8
XFILLER_19_165 VPWR VGND sg13g2_decap_8
XFILLER_34_102 VPWR VGND sg13g2_decap_8
XFILLER_43_680 VPWR VGND sg13g2_fill_1
XFILLER_34_179 VPWR VGND sg13g2_decap_8
XFILLER_22_319 VPWR VGND sg13g2_decap_8
XFILLER_15_382 VPWR VGND sg13g2_decap_8
X_1902_ net223 VPWR _0784_ VGND state\[90\] net195 sg13g2_o21ai_1
X_1833_ VPWR VGND _0732_ net108 _0731_ _0225_ _0328_ net65 sg13g2_a221oi_1
XFILLER_30_396 VPWR VGND sg13g2_decap_8
X_1764_ VGND VPWR net153 daisychain\[54\] _0681_ net53 sg13g2_a21oi_1
X_2528__279 VPWR VGND net278 sg13g2_tiehi
XFILLER_7_581 VPWR VGND sg13g2_decap_8
X_1695_ net187 _0187_ _0628_ _0629_ VPWR VGND sg13g2_a21o_1
X_2316_ net471 VGND VPWR _0262_ daisychain\[6\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2247_ VGND VPWR _0803_ _0994_ _0480_ net85 sg13g2_a21oi_1
X_2178_ _0960_ net144 state\[62\] VPWR VGND sg13g2_nand2_1
XFILLER_26_625 VPWR VGND sg13g2_decap_4
XFILLER_25_102 VPWR VGND sg13g2_decap_8
XFILLER_13_319 VPWR VGND sg13g2_decap_8
XFILLER_15_25 VPWR VGND sg13g2_decap_8
XFILLER_41_639 VPWR VGND sg13g2_decap_4
XFILLER_40_105 VPWR VGND sg13g2_decap_8
XFILLER_25_179 VPWR VGND sg13g2_decap_8
XFILLER_22_875 VPWR VGND sg13g2_decap_8
XFILLER_21_396 VPWR VGND sg13g2_decap_8
XFILLER_31_46 VPWR VGND sg13g2_decap_8
Xoutput13 net13 uio_out[5] VPWR VGND sg13g2_buf_1
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_16_102 VPWR VGND sg13g2_decap_8
XFILLER_44_466 VPWR VGND sg13g2_fill_1
XFILLER_44_455 VPWR VGND sg13g2_decap_8
XFILLER_16_179 VPWR VGND sg13g2_decap_8
XFILLER_31_116 VPWR VGND sg13g2_decap_8
XFILLER_25_691 VPWR VGND sg13g2_decap_4
XFILLER_8_312 VPWR VGND sg13g2_decap_8
XFILLER_12_396 VPWR VGND sg13g2_decap_8
X_2486__293 VPWR VGND net292 sg13g2_tiehi
XFILLER_8_389 VPWR VGND sg13g2_decap_8
X_1480_ VPWR _0210_ daisychain\[59\] VGND sg13g2_inv_1
XFILLER_4_595 VPWR VGND sg13g2_decap_8
X_2101_ VGND VPWR _0584_ _0921_ _0407_ net102 sg13g2_a21oi_1
XFILLER_39_238 VPWR VGND sg13g2_decap_8
XFILLER_11_4 VPWR VGND sg13g2_decap_8
X_2032_ VGND VPWR net114 daisychain\[121\] _0882_ net25 sg13g2_a21oi_1
XFILLER_35_444 VPWR VGND sg13g2_decap_8
XFILLER_22_116 VPWR VGND sg13g2_decap_8
XFILLER_16_691 VPWR VGND sg13g2_decap_8
XFILLER_31_661 VPWR VGND sg13g2_decap_8
X_1816_ VGND VPWR net155 daisychain\[67\] _0720_ net66 sg13g2_a21oi_1
XFILLER_30_193 VPWR VGND sg13g2_decap_8
X_2465__377 VPWR VGND net376 sg13g2_tiehi
XFILLER_7_70 VPWR VGND sg13g2_decap_8
X_1747_ net188 _0202_ _0667_ _0668_ VPWR VGND sg13g2_a21o_1
X_1678_ net206 VPWR _0616_ VGND state\[34\] net164 sg13g2_o21ai_1
XFILLER_27_945 VPWR VGND sg13g2_decap_8
XFILLER_26_46 VPWR VGND sg13g2_decap_8
XFILLER_42_937 VPWR VGND sg13g2_fill_2
XFILLER_13_116 VPWR VGND sg13g2_decap_8
XFILLER_41_447 VPWR VGND sg13g2_fill_2
XFILLER_9_109 VPWR VGND sg13g2_decap_8
XFILLER_41_469 VPWR VGND sg13g2_decap_8
XFILLER_42_56 VPWR VGND sg13g2_decap_8
XFILLER_21_193 VPWR VGND sg13g2_decap_8
XFILLER_5_326 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_49_536 VPWR VGND sg13g2_decap_8
XFILLER_18_934 VPWR VGND sg13g2_fill_2
XFILLER_45_786 VPWR VGND sg13g2_decap_4
XFILLER_44_252 VPWR VGND sg13g2_decap_8
XFILLER_32_403 VPWR VGND sg13g2_decap_8
XFILLER_32_436 VPWR VGND sg13g2_fill_2
X_2414__276 VPWR VGND net275 sg13g2_tiehi
XFILLER_13_694 VPWR VGND sg13g2_fill_2
XFILLER_12_193 VPWR VGND sg13g2_decap_8
X_1601_ VPWR VGND _0558_ net73 _0557_ _0161_ _0270_ net27 sg13g2_a221oi_1
XFILLER_9_698 VPWR VGND sg13g2_decap_4
XFILLER_8_186 VPWR VGND sg13g2_decap_8
X_1532_ VPWR _0233_ daisychain\[7\] VGND sg13g2_inv_1
X_1463_ VPWR _0229_ daisychain\[76\] VGND sg13g2_inv_1
X_1394_ VPWR _0036_ state\[17\] VGND sg13g2_inv_1
X_2015_ net174 _0148_ _0868_ _0869_ VPWR VGND sg13g2_a21o_1
XFILLER_35_252 VPWR VGND sg13g2_decap_8
XFILLER_24_926 VPWR VGND sg13g2_decap_8
XFILLER_23_403 VPWR VGND sg13g2_decap_8
XFILLER_3_808 VPWR VGND sg13g2_decap_8
XFILLER_37_56 VPWR VGND sg13g2_decap_8
XFILLER_14_403 VPWR VGND sg13g2_decap_8
XFILLER_42_723 VPWR VGND sg13g2_decap_4
XFILLER_26_263 VPWR VGND sg13g2_decap_8
XFILLER_42_756 VPWR VGND sg13g2_fill_1
XFILLER_42_789 VPWR VGND sg13g2_decap_4
XFILLER_41_266 VPWR VGND sg13g2_decap_8
XFILLER_30_907 VPWR VGND sg13g2_decap_8
XFILLER_5_123 VPWR VGND sg13g2_decap_8
XFILLER_2_874 VPWR VGND sg13g2_decap_8
XFILLER_49_333 VPWR VGND sg13g2_decap_8
XFILLER_18_742 VPWR VGND sg13g2_decap_8
XFILLER_17_252 VPWR VGND sg13g2_decap_8
XFILLER_18_775 VPWR VGND sg13g2_fill_1
XFILLER_45_561 VPWR VGND sg13g2_decap_8
XFILLER_45_594 VPWR VGND sg13g2_decap_8
XFILLER_32_200 VPWR VGND sg13g2_decap_8
X_2316__472 VPWR VGND net471 sg13g2_tiehi
XFILLER_32_277 VPWR VGND sg13g2_decap_8
XFILLER_20_417 VPWR VGND sg13g2_decap_8
XFILLER_9_473 VPWR VGND sg13g2_decap_8
X_2564_ net290 VGND VPWR _0510_ state\[126\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1515_ VPWR _0172_ daisychain\[24\] VGND sg13g2_inv_1
X_2495_ net256 VGND VPWR _0441_ state\[57\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_4_60 VPWR VGND sg13g2_decap_8
X_1446_ VPWR _0248_ daisychain\[93\] VGND sg13g2_inv_1
X_1377_ VPWR _0055_ state\[34\] VGND sg13g2_inv_1
XFILLER_23_200 VPWR VGND sg13g2_decap_8
XFILLER_11_417 VPWR VGND sg13g2_decap_8
XFILLER_23_277 VPWR VGND sg13g2_decap_8
XFILLER_23_25 VPWR VGND sg13g2_decap_8
X_2367__370 VPWR VGND net369 sg13g2_tiehi
XFILLER_2_137 VPWR VGND sg13g2_decap_8
X_2398__308 VPWR VGND net307 sg13g2_tiehi
X_2519__351 VPWR VGND net350 sg13g2_tiehi
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_46_336 VPWR VGND sg13g2_decap_8
XFILLER_14_200 VPWR VGND sg13g2_decap_8
XFILLER_42_564 VPWR VGND sg13g2_decap_4
XFILLER_42_542 VPWR VGND sg13g2_fill_2
XFILLER_14_277 VPWR VGND sg13g2_decap_8
Xfanout70 net72 net70 VPWR VGND sg13g2_buf_1
Xfanout81 net91 net81 VPWR VGND sg13g2_buf_1
Xfanout92 net96 net92 VPWR VGND sg13g2_buf_1
XFILLER_7_933 VPWR VGND sg13g2_decap_8
XFILLER_6_410 VPWR VGND sg13g2_decap_8
XFILLER_10_494 VPWR VGND sg13g2_decap_8
XFILLER_7_955 VPWR VGND sg13g2_decap_8
XFILLER_7_999 VPWR VGND sg13g2_fill_1
XFILLER_6_487 VPWR VGND sg13g2_decap_8
XFILLER_43_7 VPWR VGND sg13g2_decap_8
X_2280_ _1011_ net125 state\[113\] VPWR VGND sg13g2_nand2_1
X_1300_ VPWR _0013_ state\[111\] VGND sg13g2_inv_1
XFILLER_49_130 VPWR VGND sg13g2_decap_8
XFILLER_37_336 VPWR VGND sg13g2_decap_8
XFILLER_46_870 VPWR VGND sg13g2_fill_2
XFILLER_33_553 VPWR VGND sg13g2_decap_8
XFILLER_20_214 VPWR VGND sg13g2_decap_8
X_1995_ net171 _0143_ _0853_ _0854_ VPWR VGND sg13g2_a21o_1
XFILLER_9_270 VPWR VGND sg13g2_decap_8
X_2547_ net282 VGND VPWR _0493_ state\[109\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_47_1024 VPWR VGND sg13g2_decap_4
X_2478_ net324 VGND VPWR _0424_ state\[40\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1429_ VPWR _0140_ daisychain\[110\] VGND sg13g2_inv_1
XFILLER_18_25 VPWR VGND sg13g2_decap_8
XFILLER_29_826 VPWR VGND sg13g2_decap_8
XFILLER_28_347 VPWR VGND sg13g2_decap_8
XFILLER_34_46 VPWR VGND sg13g2_decap_8
XFILLER_24_553 VPWR VGND sg13g2_fill_1
XFILLER_24_542 VPWR VGND sg13g2_decap_8
XFILLER_11_214 VPWR VGND sg13g2_decap_8
XFILLER_12_737 VPWR VGND sg13g2_fill_2
Xclkload1 clknet_leaf_1_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_20_781 VPWR VGND sg13g2_fill_1
XFILLER_4_925 VPWR VGND sg13g2_decap_8
XFILLER_4_903 VPWR VGND sg13g2_decap_4
XFILLER_3_468 VPWR VGND sg13g2_decap_8
XFILLER_19_347 VPWR VGND sg13g2_decap_8
XFILLER_46_133 VPWR VGND sg13g2_decap_8
XFILLER_47_667 VPWR VGND sg13g2_fill_2
XFILLER_15_564 VPWR VGND sg13g2_fill_2
XFILLER_42_350 VPWR VGND sg13g2_decap_8
XFILLER_30_501 VPWR VGND sg13g2_decap_8
X_1780_ VGND VPWR net143 daisychain\[58\] _0693_ net56 sg13g2_a21oi_1
XFILLER_10_291 VPWR VGND sg13g2_decap_8
XFILLER_6_284 VPWR VGND sg13g2_decap_8
X_2401_ net301 VGND VPWR _0347_ daisychain\[91\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2332_ net439 VGND VPWR _0278_ daisychain\[22\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2263_ VGND VPWR _0827_ _1002_ _0488_ net87 sg13g2_a21oi_1
XFILLER_38_623 VPWR VGND sg13g2_fill_2
XFILLER_38_601 VPWR VGND sg13g2_fill_2
X_2194_ _0968_ net155 state\[70\] VPWR VGND sg13g2_nand2_1
XFILLER_37_133 VPWR VGND sg13g2_decap_8
XFILLER_26_829 VPWR VGND sg13g2_fill_2
XFILLER_19_892 VPWR VGND sg13g2_fill_1
XFILLER_33_361 VPWR VGND sg13g2_decap_8
XFILLER_21_523 VPWR VGND sg13g2_fill_1
X_1978_ net213 VPWR _0841_ VGND state\[109\] net176 sg13g2_o21ai_1
XFILLER_0_427 VPWR VGND sg13g2_decap_8
XFILLER_29_612 VPWR VGND sg13g2_fill_2
XFILLER_29_46 VPWR VGND sg13g2_decap_8
XFILLER_28_144 VPWR VGND sg13g2_decap_8
XFILLER_45_56 VPWR VGND sg13g2_decap_8
XFILLER_43_147 VPWR VGND sg13g2_decap_8
XFILLER_24_361 VPWR VGND sg13g2_decap_8
XFILLER_12_556 VPWR VGND sg13g2_decap_4
XFILLER_12_589 VPWR VGND sg13g2_decap_4
XFILLER_8_516 VPWR VGND sg13g2_decap_8
XFILLER_6_39 VPWR VGND sg13g2_decap_8
XFILLER_3_221 VPWR VGND sg13g2_decap_8
XFILLER_10_81 VPWR VGND sg13g2_decap_8
XFILLER_3_298 VPWR VGND sg13g2_decap_8
XFILLER_0_994 VPWR VGND sg13g2_decap_8
XFILLER_47_420 VPWR VGND sg13g2_decap_8
XFILLER_19_144 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_34_158 VPWR VGND sg13g2_decap_8
XFILLER_15_361 VPWR VGND sg13g2_decap_8
X_1901_ VPWR VGND _0783_ net85 _0782_ _0243_ _0345_ net42 sg13g2_a221oi_1
XFILLER_43_692 VPWR VGND sg13g2_fill_1
X_1832_ VGND VPWR net155 daisychain\[71\] _0732_ net65 sg13g2_a21oi_1
XFILLER_30_375 VPWR VGND sg13g2_decap_8
X_1763_ net192 _0206_ _0679_ _0680_ VPWR VGND sg13g2_a21o_1
XFILLER_7_560 VPWR VGND sg13g2_decap_8
X_1694_ net218 VPWR _0628_ VGND state\[38\] net184 sg13g2_o21ai_1
X_2424__256 VPWR VGND net255 sg13g2_tiehi
X_2315_ net473 VGND VPWR _0261_ daisychain\[5\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2246_ _0994_ net129 state\[96\] VPWR VGND sg13g2_nand2_1
X_2177_ VGND VPWR _0698_ _0959_ _0445_ net98 sg13g2_a21oi_1
XFILLER_25_158 VPWR VGND sg13g2_decap_8
XFILLER_22_810 VPWR VGND sg13g2_decap_8
XFILLER_22_854 VPWR VGND sg13g2_decap_8
XFILLER_31_25 VPWR VGND sg13g2_decap_8
XFILLER_21_375 VPWR VGND sg13g2_decap_8
XFILLER_5_508 VPWR VGND sg13g2_fill_1
Xoutput14 net14 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_49_707 VPWR VGND sg13g2_fill_2
XFILLER_49_729 VPWR VGND sg13g2_fill_1
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_45_924 VPWR VGND sg13g2_fill_1
XFILLER_44_434 VPWR VGND sg13g2_decap_8
XFILLER_16_158 VPWR VGND sg13g2_decap_8
XFILLER_44_478 VPWR VGND sg13g2_decap_8
XFILLER_12_375 VPWR VGND sg13g2_decap_8
XFILLER_40_684 VPWR VGND sg13g2_decap_8
XFILLER_40_673 VPWR VGND sg13g2_decap_4
XFILLER_8_368 VPWR VGND sg13g2_decap_8
XFILLER_4_574 VPWR VGND sg13g2_decap_8
X_2100_ _0921_ net148 state\[23\] VPWR VGND sg13g2_nand2_1
XFILLER_39_217 VPWR VGND sg13g2_decap_8
X_2031_ net160 _0153_ _0880_ _0881_ VPWR VGND sg13g2_a21o_1
X_2493__265 VPWR VGND net264 sg13g2_tiehi
XFILLER_47_294 VPWR VGND sg13g2_decap_8
XFILLER_30_172 VPWR VGND sg13g2_decap_8
X_1815_ net202 _0220_ _0718_ _0719_ VPWR VGND sg13g2_a21o_1
X_1746_ net221 VPWR _0667_ VGND state\[51\] net188 sg13g2_o21ai_1
X_1677_ VPWR VGND _0615_ net73 _0614_ _0182_ _0289_ net27 sg13g2_a221oi_1
X_2326__452 VPWR VGND net451 sg13g2_tiehi
X_2229_ VGND VPWR _0776_ _0985_ _0471_ net82 sg13g2_a21oi_1
X_2472__349 VPWR VGND net348 sg13g2_tiehi
XFILLER_38_294 VPWR VGND sg13g2_decap_8
XFILLER_27_957 VPWR VGND sg13g2_fill_1
XFILLER_26_445 VPWR VGND sg13g2_decap_8
XFILLER_26_25 VPWR VGND sg13g2_decap_8
XFILLER_42_927 VPWR VGND sg13g2_fill_2
XFILLER_42_916 VPWR VGND sg13g2_fill_1
XFILLER_41_415 VPWR VGND sg13g2_fill_1
XFILLER_42_35 VPWR VGND sg13g2_decap_8
XFILLER_22_673 VPWR VGND sg13g2_fill_2
XFILLER_21_172 VPWR VGND sg13g2_decap_8
XFILLER_5_305 VPWR VGND sg13g2_decap_8
XFILLER_1_511 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_49_515 VPWR VGND sg13g2_decap_8
XFILLER_1_588 VPWR VGND sg13g2_decap_8
X_2377__350 VPWR VGND net349 sg13g2_tiehi
XFILLER_44_231 VPWR VGND sg13g2_decap_8
XFILLER_12_172 VPWR VGND sg13g2_decap_8
XFILLER_9_677 VPWR VGND sg13g2_decap_8
XFILLER_40_492 VPWR VGND sg13g2_fill_1
X_1600_ VGND VPWR net116 daisychain\[13\] _0558_ net27 sg13g2_a21oi_1
XFILLER_8_165 VPWR VGND sg13g2_decap_8
X_1531_ VPWR _0244_ daisychain\[8\] VGND sg13g2_inv_1
X_1462_ VPWR _0230_ daisychain\[77\] VGND sg13g2_inv_1
XFILLER_4_382 VPWR VGND sg13g2_decap_8
X_1393_ VPWR _0037_ state\[18\] VGND sg13g2_inv_1
X_2014_ net217 VPWR _0868_ VGND state\[118\] net174 sg13g2_o21ai_1
XFILLER_36_732 VPWR VGND sg13g2_decap_8
XFILLER_35_231 VPWR VGND sg13g2_decap_8
XFILLER_10_109 VPWR VGND sg13g2_decap_8
XFILLER_32_993 VPWR VGND sg13g2_fill_1
XFILLER_32_982 VPWR VGND sg13g2_fill_1
X_1729_ VPWR VGND _0654_ net95 _0653_ _0196_ _0302_ net50 sg13g2_a221oi_1
XFILLER_2_319 VPWR VGND sg13g2_decap_8
XFILLER_37_35 VPWR VGND sg13g2_decap_8
XFILLER_2_1002 VPWR VGND sg13g2_decap_4
XFILLER_39_592 VPWR VGND sg13g2_decap_4
XFILLER_26_242 VPWR VGND sg13g2_decap_8
XFILLER_41_245 VPWR VGND sg13g2_decap_8
XFILLER_5_102 VPWR VGND sg13g2_decap_8
XFILLER_5_179 VPWR VGND sg13g2_decap_8
XFILLER_2_853 VPWR VGND sg13g2_decap_8
XFILLER_49_312 VPWR VGND sg13g2_decap_8
XFILLER_2_897 VPWR VGND sg13g2_fill_1
XFILLER_1_385 VPWR VGND sg13g2_decap_8
XFILLER_49_389 VPWR VGND sg13g2_decap_8
XFILLER_17_231 VPWR VGND sg13g2_decap_8
XFILLER_18_765 VPWR VGND sg13g2_fill_1
XFILLER_32_256 VPWR VGND sg13g2_decap_8
XFILLER_9_452 VPWR VGND sg13g2_decap_8
X_2563_ net418 VGND VPWR _0509_ state\[125\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_1514_ VPWR _0173_ daisychain\[25\] VGND sg13g2_inv_1
X_2494_ net260 VGND VPWR _0440_ state\[56\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1445_ VPWR _0249_ daisychain\[94\] VGND sg13g2_inv_1
X_1376_ VPWR _0056_ state\[35\] VGND sg13g2_inv_1
XFILLER_28_529 VPWR VGND sg13g2_decap_8
XFILLER_23_256 VPWR VGND sg13g2_decap_8
X_2547__283 VPWR VGND net282 sg13g2_tiehi
XFILLER_2_116 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_46_315 VPWR VGND sg13g2_decap_8
XFILLER_47_849 VPWR VGND sg13g2_fill_1
XFILLER_15_735 VPWR VGND sg13g2_fill_1
XFILLER_14_256 VPWR VGND sg13g2_decap_8
XFILLER_9_39 VPWR VGND sg13g2_decap_8
Xfanout60 net61 net60 VPWR VGND sg13g2_buf_1
Xfanout71 net72 net71 VPWR VGND sg13g2_buf_1
Xfanout82 net83 net82 VPWR VGND sg13g2_buf_1
Xfanout93 net96 net93 VPWR VGND sg13g2_buf_1
XFILLER_7_912 VPWR VGND sg13g2_decap_8
XFILLER_10_473 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_decap_8
XFILLER_6_466 VPWR VGND sg13g2_decap_8
XFILLER_36_7 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_37_315 VPWR VGND sg13g2_decap_8
XFILLER_49_186 VPWR VGND sg13g2_decap_8
XFILLER_18_551 VPWR VGND sg13g2_fill_2
XFILLER_46_893 VPWR VGND sg13g2_fill_1
XFILLER_45_392 VPWR VGND sg13g2_decap_8
XFILLER_33_543 VPWR VGND sg13g2_fill_1
XFILLER_33_532 VPWR VGND sg13g2_fill_1
XFILLER_21_738 VPWR VGND sg13g2_decap_4
X_1994_ net212 VPWR _0853_ VGND state\[113\] net171 sg13g2_o21ai_1
XFILLER_0_609 VPWR VGND sg13g2_decap_8
X_2546_ net298 VGND VPWR _0492_ state\[108\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2477_ net328 VGND VPWR _0423_ state\[39\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1428_ VPWR _0141_ daisychain\[111\] VGND sg13g2_inv_1
X_1359_ VPWR _0075_ state\[52\] VGND sg13g2_inv_1
XFILLER_28_326 VPWR VGND sg13g2_decap_8
X_2434__236 VPWR VGND net235 sg13g2_tiehi
XFILLER_43_329 VPWR VGND sg13g2_decap_8
XFILLER_36_392 VPWR VGND sg13g2_decap_8
XFILLER_34_25 VPWR VGND sg13g2_decap_8
Xclkload2 VPWR clkload2/Y clknet_leaf_18_clk VGND sg13g2_inv_1
XFILLER_3_403 VPWR VGND sg13g2_decap_8
XFILLER_4_959 VPWR VGND sg13g2_decap_4
XFILLER_3_447 VPWR VGND sg13g2_decap_8
XFILLER_19_326 VPWR VGND sg13g2_decap_8
XFILLER_46_112 VPWR VGND sg13g2_decap_8
XFILLER_46_189 VPWR VGND sg13g2_decap_8
XFILLER_27_392 VPWR VGND sg13g2_decap_8
X_2489__281 VPWR VGND net280 sg13g2_tiehi
XFILLER_10_270 VPWR VGND sg13g2_decap_8
XFILLER_7_720 VPWR VGND sg13g2_fill_1
X_2400_ net303 VGND VPWR _0346_ daisychain\[90\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_6_263 VPWR VGND sg13g2_decap_8
X_2331_ net441 VGND VPWR _0277_ daisychain\[21\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_34_4 VPWR VGND sg13g2_decap_8
X_2262_ _1002_ net131 state\[104\] VPWR VGND sg13g2_nand2_1
XFILLER_2_480 VPWR VGND sg13g2_decap_8
X_2193_ VGND VPWR _0722_ _0967_ _0453_ net109 sg13g2_a21oi_1
XFILLER_37_112 VPWR VGND sg13g2_decap_8
XFILLER_37_189 VPWR VGND sg13g2_decap_8
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_18_392 VPWR VGND sg13g2_decap_8
XFILLER_33_340 VPWR VGND sg13g2_decap_8
X_1977_ VPWR VGND _0840_ net87 _0839_ _0137_ _0364_ net44 sg13g2_a221oi_1
X_2468__365 VPWR VGND net364 sg13g2_tiehi
XFILLER_0_406 VPWR VGND sg13g2_decap_8
X_2529_ net270 VGND VPWR _0475_ state\[91\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_29_25 VPWR VGND sg13g2_decap_8
XFILLER_28_123 VPWR VGND sg13g2_decap_8
X_2336__432 VPWR VGND net431 sg13g2_tiehi
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_43_126 VPWR VGND sg13g2_decap_8
XFILLER_25_874 VPWR VGND sg13g2_decap_8
XFILLER_24_340 VPWR VGND sg13g2_decap_8
XFILLER_12_535 VPWR VGND sg13g2_decap_8
X_2447__449 VPWR VGND net448 sg13g2_tiehi
XFILLER_6_18 VPWR VGND sg13g2_decap_8
XFILLER_4_701 VPWR VGND sg13g2_fill_2
XFILLER_3_200 VPWR VGND sg13g2_decap_8
XFILLER_10_60 VPWR VGND sg13g2_decap_8
XFILLER_4_789 VPWR VGND sg13g2_decap_8
XFILLER_3_277 VPWR VGND sg13g2_decap_8
XFILLER_0_951 VPWR VGND sg13g2_decap_8
XFILLER_19_123 VPWR VGND sg13g2_decap_8
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_34_137 VPWR VGND sg13g2_decap_8
XFILLER_15_340 VPWR VGND sg13g2_decap_8
X_1900_ VGND VPWR net133 daisychain\[88\] _0783_ net46 sg13g2_a21oi_1
X_1831_ net201 _0225_ _0730_ _0731_ VPWR VGND sg13g2_a21o_1
X_2387__330 VPWR VGND net329 sg13g2_tiehi
XFILLER_30_354 VPWR VGND sg13g2_decap_8
X_1762_ net222 VPWR _0679_ VGND state\[55\] net192 sg13g2_o21ai_1
X_1693_ VPWR VGND _0627_ net94 _0626_ _0186_ _0293_ net49 sg13g2_a221oi_1
X_2314_ net475 VGND VPWR _0260_ daisychain\[4\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2245_ VGND VPWR _0800_ _0993_ _0479_ net85 sg13g2_a21oi_1
XFILLER_38_410 VPWR VGND sg13g2_fill_1
X_2176_ _0959_ net143 state\[61\] VPWR VGND sg13g2_nand2_1
XFILLER_38_443 VPWR VGND sg13g2_decap_4
XFILLER_38_476 VPWR VGND sg13g2_decap_4
XFILLER_25_137 VPWR VGND sg13g2_decap_8
XFILLER_22_833 VPWR VGND sg13g2_fill_2
XFILLER_21_354 VPWR VGND sg13g2_decap_8
Xoutput15 net15 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_0_203 VPWR VGND sg13g2_decap_8
XFILLER_29_410 VPWR VGND sg13g2_decap_4
XFILLER_44_413 VPWR VGND sg13g2_decap_8
XFILLER_29_487 VPWR VGND sg13g2_fill_1
XFILLER_16_137 VPWR VGND sg13g2_decap_8
XFILLER_45_969 VPWR VGND sg13g2_decap_8
XFILLER_32_619 VPWR VGND sg13g2_fill_2
XFILLER_12_354 VPWR VGND sg13g2_decap_8
XFILLER_40_652 VPWR VGND sg13g2_decap_8
XFILLER_8_347 VPWR VGND sg13g2_decap_8
XFILLER_21_81 VPWR VGND sg13g2_decap_8
XFILLER_4_553 VPWR VGND sg13g2_decap_8
X_2030_ net205 VPWR _0880_ VGND state\[122\] net160 sg13g2_o21ai_1
XFILLER_48_752 VPWR VGND sg13g2_decap_8
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_35_413 VPWR VGND sg13g2_decap_8
XFILLER_31_630 VPWR VGND sg13g2_decap_8
XFILLER_30_151 VPWR VGND sg13g2_decap_8
X_1814_ net225 VPWR _0718_ VGND state\[68\] net202 sg13g2_o21ai_1
X_1745_ VPWR VGND _0666_ net95 _0665_ _0201_ _0306_ net51 sg13g2_a221oi_1
XFILLER_8_881 VPWR VGND sg13g2_fill_1
X_1676_ VGND VPWR net116 daisychain\[32\] _0615_ net27 sg13g2_a21oi_1
X_2502__229 VPWR VGND net sg13g2_tiehi
XFILLER_39_730 VPWR VGND sg13g2_decap_8
XFILLER_27_903 VPWR VGND sg13g2_decap_8
X_2228_ _0985_ net126 state\[87\] VPWR VGND sg13g2_nand2_1
XFILLER_38_273 VPWR VGND sg13g2_decap_8
X_2159_ VGND VPWR _0671_ _0950_ _0436_ net97 sg13g2_a21oi_1
XFILLER_26_424 VPWR VGND sg13g2_decap_8
XFILLER_42_939 VPWR VGND sg13g2_fill_1
XFILLER_26_479 VPWR VGND sg13g2_decap_8
XFILLER_42_14 VPWR VGND sg13g2_decap_8
XFILLER_34_490 VPWR VGND sg13g2_fill_2
XFILLER_21_151 VPWR VGND sg13g2_decap_8
XFILLER_6_829 VPWR VGND sg13g2_decap_8
XFILLER_27_1012 VPWR VGND sg13g2_decap_8
XFILLER_1_567 VPWR VGND sg13g2_decap_8
XFILLER_17_413 VPWR VGND sg13g2_decap_8
XFILLER_18_914 VPWR VGND sg13g2_fill_1
XFILLER_18_947 VPWR VGND sg13g2_fill_1
XFILLER_44_210 VPWR VGND sg13g2_decap_8
XFILLER_29_284 VPWR VGND sg13g2_decap_8
XFILLER_17_468 VPWR VGND sg13g2_fill_2
XFILLER_44_287 VPWR VGND sg13g2_decap_8
XFILLER_16_81 VPWR VGND sg13g2_decap_8
XFILLER_32_449 VPWR VGND sg13g2_decap_8
XFILLER_12_151 VPWR VGND sg13g2_decap_8
XFILLER_13_696 VPWR VGND sg13g2_fill_1
XFILLER_9_623 VPWR VGND sg13g2_decap_4
XFILLER_9_612 VPWR VGND sg13g2_decap_4
XFILLER_8_144 VPWR VGND sg13g2_decap_8
X_1530_ VPWR _0255_ daisychain\[9\] VGND sg13g2_inv_1
XFILLER_4_361 VPWR VGND sg13g2_decap_8
X_1461_ VPWR _0231_ daisychain\[78\] VGND sg13g2_inv_1
X_1392_ VPWR _0038_ state\[19\] VGND sg13g2_inv_1
X_2013_ VPWR VGND _0867_ net82 _0866_ _0147_ _0373_ net39 sg13g2_a221oi_1
XFILLER_35_210 VPWR VGND sg13g2_decap_8
XFILLER_35_287 VPWR VGND sg13g2_decap_8
XFILLER_23_438 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk clknet_2_2__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
XFILLER_12_39 VPWR VGND sg13g2_decap_8
X_1728_ VGND VPWR net141 daisychain\[45\] _0654_ net50 sg13g2_a21oi_1
X_1659_ net166 _0177_ _0601_ _0602_ VPWR VGND sg13g2_a21o_1
XFILLER_37_14 VPWR VGND sg13g2_decap_8
XFILLER_27_733 VPWR VGND sg13g2_decap_4
XFILLER_26_221 VPWR VGND sg13g2_decap_8
XFILLER_14_438 VPWR VGND sg13g2_decap_8
XFILLER_42_736 VPWR VGND sg13g2_fill_2
XFILLER_41_224 VPWR VGND sg13g2_decap_8
XFILLER_26_298 VPWR VGND sg13g2_decap_8
XFILLER_23_961 VPWR VGND sg13g2_fill_2
XFILLER_10_655 VPWR VGND sg13g2_decap_8
XFILLER_6_659 VPWR VGND sg13g2_fill_1
XFILLER_5_158 VPWR VGND sg13g2_decap_8
XFILLER_2_843 VPWR VGND sg13g2_fill_1
XFILLER_1_364 VPWR VGND sg13g2_decap_8
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_37_519 VPWR VGND sg13g2_fill_2
XFILLER_37_508 VPWR VGND sg13g2_decap_8
XFILLER_17_210 VPWR VGND sg13g2_decap_8
XFILLER_18_788 VPWR VGND sg13g2_fill_1
XFILLER_17_287 VPWR VGND sg13g2_decap_8
X_2531__255 VPWR VGND net254 sg13g2_tiehi
XFILLER_27_91 VPWR VGND sg13g2_decap_8
XFILLER_32_235 VPWR VGND sg13g2_decap_8
XFILLER_13_493 VPWR VGND sg13g2_decap_8
XFILLER_9_431 VPWR VGND sg13g2_decap_8
X_2562_ net258 VGND VPWR _0508_ state\[124\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1513_ VPWR _0174_ daisychain\[26\] VGND sg13g2_inv_1
X_2493_ net264 VGND VPWR _0439_ state\[55\] clknet_leaf_14_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_4_clk clknet_2_1__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_1444_ VPWR _0250_ daisychain\[95\] VGND sg13g2_inv_1
XFILLER_4_95 VPWR VGND sg13g2_decap_8
X_1375_ VPWR _0057_ state\[36\] VGND sg13g2_inv_1
XFILLER_36_541 VPWR VGND sg13g2_decap_4
XFILLER_23_235 VPWR VGND sg13g2_decap_8
XFILLER_20_975 VPWR VGND sg13g2_decap_8
XFILLER_3_629 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_47_806 VPWR VGND sg13g2_fill_1
XFILLER_47_817 VPWR VGND sg13g2_decap_4
XFILLER_27_552 VPWR VGND sg13g2_decap_8
XFILLER_27_585 VPWR VGND sg13g2_decap_4
XFILLER_14_235 VPWR VGND sg13g2_decap_8
XFILLER_9_18 VPWR VGND sg13g2_decap_8
XFILLER_42_544 VPWR VGND sg13g2_fill_1
Xfanout50 net51 net50 VPWR VGND sg13g2_buf_1
Xfanout61 net67 net61 VPWR VGND sg13g2_buf_1
Xfanout72 net78 net72 VPWR VGND sg13g2_buf_1
Xfanout83 net91 net83 VPWR VGND sg13g2_buf_1
XFILLER_10_452 VPWR VGND sg13g2_decap_8
XFILLER_13_60 VPWR VGND sg13g2_decap_8
Xfanout94 net96 net94 VPWR VGND sg13g2_buf_1
X_2346__412 VPWR VGND net411 sg13g2_tiehi
XFILLER_6_445 VPWR VGND sg13g2_decap_8
X_2461__393 VPWR VGND net392 sg13g2_tiehi
XFILLER_2_684 VPWR VGND sg13g2_decap_8
XFILLER_2_673 VPWR VGND sg13g2_fill_2
XFILLER_2_662 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_49_165 VPWR VGND sg13g2_decap_8
XFILLER_45_371 VPWR VGND sg13g2_decap_8
XFILLER_33_500 VPWR VGND sg13g2_fill_2
XFILLER_21_717 VPWR VGND sg13g2_decap_8
X_1993_ VPWR VGND _0852_ net80 _0851_ _0142_ _0368_ net36 sg13g2_a221oi_1
XFILLER_20_249 VPWR VGND sg13g2_decap_8
X_2545_ net314 VGND VPWR _0491_ state\[107\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2476_ net332 VGND VPWR _0422_ state\[38\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2397__310 VPWR VGND net309 sg13g2_tiehi
X_2440__477 VPWR VGND net476 sg13g2_tiehi
X_1427_ VPWR _0142_ daisychain\[112\] VGND sg13g2_inv_1
XFILLER_28_305 VPWR VGND sg13g2_decap_8
X_1358_ VPWR _0076_ state\[53\] VGND sg13g2_inv_1
X_1289_ VPWR _0025_ state\[122\] VGND sg13g2_inv_1
XFILLER_43_308 VPWR VGND sg13g2_decap_8
XFILLER_36_371 VPWR VGND sg13g2_decap_8
XFILLER_12_706 VPWR VGND sg13g2_fill_1
XFILLER_24_566 VPWR VGND sg13g2_decap_8
XFILLER_11_249 VPWR VGND sg13g2_decap_8
Xclkload3 clkload3/Y clknet_leaf_19_clk VPWR VGND sg13g2_inv_8
XFILLER_3_426 VPWR VGND sg13g2_decap_8
XFILLER_19_305 VPWR VGND sg13g2_decap_8
XFILLER_47_614 VPWR VGND sg13g2_decap_8
XFILLER_47_625 VPWR VGND sg13g2_fill_2
XFILLER_47_669 VPWR VGND sg13g2_fill_1
XFILLER_15_511 VPWR VGND sg13g2_decap_4
XFILLER_46_168 VPWR VGND sg13g2_decap_8
XFILLER_34_319 VPWR VGND sg13g2_decap_8
XFILLER_27_371 VPWR VGND sg13g2_decap_8
XFILLER_15_566 VPWR VGND sg13g2_fill_1
XFILLER_43_875 VPWR VGND sg13g2_decap_8
XFILLER_42_385 VPWR VGND sg13g2_decap_8
XFILLER_30_536 VPWR VGND sg13g2_fill_2
XFILLER_24_81 VPWR VGND sg13g2_decap_8
XFILLER_7_776 VPWR VGND sg13g2_decap_8
XFILLER_6_242 VPWR VGND sg13g2_decap_8
XFILLER_7_787 VPWR VGND sg13g2_fill_2
XFILLER_40_91 VPWR VGND sg13g2_decap_8
X_2330_ net443 VGND VPWR _0276_ daisychain\[20\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2261_ VGND VPWR _0824_ _1001_ _0487_ net88 sg13g2_a21oi_1
X_2496__253 VPWR VGND net252 sg13g2_tiehi
X_2192_ _0967_ net156 state\[69\] VPWR VGND sg13g2_nand2_1
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_37_168 VPWR VGND sg13g2_decap_8
XFILLER_25_319 VPWR VGND sg13g2_decap_8
XFILLER_19_883 VPWR VGND sg13g2_fill_1
XFILLER_33_396 VPWR VGND sg13g2_decap_8
X_1976_ VGND VPWR net131 daisychain\[107\] _0840_ net44 sg13g2_a21oi_1
XFILLER_21_558 VPWR VGND sg13g2_fill_1
XFILLER_20_39 VPWR VGND sg13g2_decap_8
X_2528_ net278 VGND VPWR _0474_ state\[90\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2459_ net400 VGND VPWR _0405_ state\[21\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2475__337 VPWR VGND net336 sg13g2_tiehi
XFILLER_29_614 VPWR VGND sg13g2_fill_1
XFILLER_28_102 VPWR VGND sg13g2_decap_8
XFILLER_16_319 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_43_105 VPWR VGND sg13g2_decap_8
XFILLER_28_179 VPWR VGND sg13g2_decap_8
XFILLER_12_514 VPWR VGND sg13g2_decap_8
XFILLER_24_396 VPWR VGND sg13g2_decap_8
XFILLER_3_256 VPWR VGND sg13g2_decap_8
XFILLER_0_930 VPWR VGND sg13g2_fill_1
XFILLER_0_974 VPWR VGND sg13g2_fill_2
XFILLER_19_102 VPWR VGND sg13g2_decap_8
XFILLER_47_455 VPWR VGND sg13g2_decap_8
XFILLER_19_81 VPWR VGND sg13g2_decap_8
XFILLER_19_179 VPWR VGND sg13g2_decap_8
XFILLER_35_639 VPWR VGND sg13g2_decap_4
XFILLER_34_116 VPWR VGND sg13g2_decap_8
XFILLER_43_661 VPWR VGND sg13g2_decap_8
XFILLER_15_396 VPWR VGND sg13g2_decap_8
XFILLER_42_182 VPWR VGND sg13g2_decap_8
XFILLER_35_91 VPWR VGND sg13g2_decap_8
X_1830_ net226 VPWR _0730_ VGND state\[72\] net201 sg13g2_o21ai_1
XFILLER_30_333 VPWR VGND sg13g2_decap_8
X_1761_ VPWR VGND _0678_ net107 _0677_ _0205_ _0310_ net53 sg13g2_a221oi_1
X_1692_ VGND VPWR net140 daisychain\[36\] _0627_ net49 sg13g2_a21oi_1
XFILLER_7_595 VPWR VGND sg13g2_fill_2
X_2313_ net477 VGND VPWR _0259_ daisychain\[3\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2244_ _0993_ net129 state\[95\] VPWR VGND sg13g2_nand2_1
X_2175_ VGND VPWR _0695_ _0958_ _0444_ net98 sg13g2_a21oi_1
XFILLER_25_116 VPWR VGND sg13g2_decap_8
XFILLER_15_39 VPWR VGND sg13g2_decap_8
XFILLER_40_119 VPWR VGND sg13g2_decap_8
XFILLER_33_193 VPWR VGND sg13g2_decap_8
XFILLER_21_333 VPWR VGND sg13g2_decap_8
X_1959_ net180 _0133_ _0826_ _0827_ VPWR VGND sg13g2_a21o_1
Xoutput16 net16 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_0_259 VPWR VGND sg13g2_decap_8
XFILLER_17_606 VPWR VGND sg13g2_decap_8
XFILLER_45_937 VPWR VGND sg13g2_decap_4
XFILLER_45_915 VPWR VGND sg13g2_decap_8
XFILLER_16_116 VPWR VGND sg13g2_decap_8
XFILLER_12_333 VPWR VGND sg13g2_decap_8
XFILLER_24_193 VPWR VGND sg13g2_decap_8
XFILLER_8_326 VPWR VGND sg13g2_decap_8
XFILLER_4_532 VPWR VGND sg13g2_decap_8
XFILLER_21_60 VPWR VGND sg13g2_decap_8
XFILLER_0_793 VPWR VGND sg13g2_decap_8
X_2534__231 VPWR VGND net230 sg13g2_tiehi
XFILLER_48_786 VPWR VGND sg13g2_decap_4
XFILLER_47_252 VPWR VGND sg13g2_decap_8
XFILLER_35_458 VPWR VGND sg13g2_decap_8
X_2354__396 VPWR VGND net395 sg13g2_tiehi
XFILLER_15_193 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clknet_0_clk clk VPWR VGND sg13g2_buf_16
XFILLER_43_491 VPWR VGND sg13g2_decap_8
XFILLER_30_130 VPWR VGND sg13g2_decap_8
XFILLER_31_675 VPWR VGND sg13g2_fill_1
X_1813_ VPWR VGND _0717_ net108 _0716_ _0219_ _0323_ net65 sg13g2_a221oi_1
X_1744_ VGND VPWR net141 daisychain\[49\] _0666_ net51 sg13g2_a21oi_1
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_7_392 VPWR VGND sg13g2_decap_8
X_1675_ net163 _0182_ _0613_ _0614_ VPWR VGND sg13g2_a21o_1
X_2227_ VGND VPWR _0773_ _0984_ _0470_ net83 sg13g2_a21oi_1
XFILLER_38_252 VPWR VGND sg13g2_decap_8
XFILLER_26_403 VPWR VGND sg13g2_decap_8
X_2158_ _0950_ net144 state\[52\] VPWR VGND sg13g2_nand2_1
X_2089_ VGND VPWR _0566_ _0915_ _0401_ net94 sg13g2_a21oi_1
XFILLER_41_406 VPWR VGND sg13g2_decap_8
XFILLER_21_130 VPWR VGND sg13g2_decap_8
XFILLER_22_675 VPWR VGND sg13g2_fill_1
XFILLER_27_1002 VPWR VGND sg13g2_decap_4
XFILLER_1_546 VPWR VGND sg13g2_decap_8
X_2557__275 VPWR VGND net274 sg13g2_tiehi
XFILLER_18_926 VPWR VGND sg13g2_fill_1
XFILLER_29_263 VPWR VGND sg13g2_decap_8
XFILLER_45_767 VPWR VGND sg13g2_decap_8
XFILLER_16_60 VPWR VGND sg13g2_decap_8
XFILLER_44_266 VPWR VGND sg13g2_decap_8
XFILLER_32_417 VPWR VGND sg13g2_decap_8
XFILLER_26_970 VPWR VGND sg13g2_fill_1
XFILLER_13_653 VPWR VGND sg13g2_fill_1
XFILLER_12_130 VPWR VGND sg13g2_decap_8
XFILLER_8_123 VPWR VGND sg13g2_decap_8
XFILLER_32_81 VPWR VGND sg13g2_decap_8
XFILLER_4_340 VPWR VGND sg13g2_decap_8
X_1460_ VPWR _0232_ daisychain\[79\] VGND sg13g2_inv_1
X_1391_ VPWR _0040_ state\[20\] VGND sg13g2_inv_1
XFILLER_48_572 VPWR VGND sg13g2_fill_2
X_2012_ VGND VPWR net126 daisychain\[116\] _0867_ net37 sg13g2_a21oi_1
XFILLER_35_266 VPWR VGND sg13g2_decap_8
XFILLER_23_417 VPWR VGND sg13g2_decap_8
XFILLER_12_18 VPWR VGND sg13g2_decap_8
X_2845_ daisychain\[127\] net23 VPWR VGND sg13g2_buf_1
X_2508__439 VPWR VGND net438 sg13g2_tiehi
X_1727_ net187 _0196_ _0652_ _0653_ VPWR VGND sg13g2_a21o_1
X_1658_ net207 VPWR _0601_ VGND state\[29\] net166 sg13g2_o21ai_1
X_1589_ VPWR VGND _0549_ net73 _0548_ _0150_ _0267_ net27 sg13g2_a221oi_1
XFILLER_2_1026 VPWR VGND sg13g2_fill_2
XFILLER_26_200 VPWR VGND sg13g2_decap_8
XFILLER_42_704 VPWR VGND sg13g2_fill_1
XFILLER_14_417 VPWR VGND sg13g2_decap_8
XFILLER_41_203 VPWR VGND sg13g2_decap_8
XFILLER_26_277 VPWR VGND sg13g2_decap_8
XFILLER_23_940 VPWR VGND sg13g2_decap_8
XFILLER_10_612 VPWR VGND sg13g2_decap_8
XFILLER_10_678 VPWR VGND sg13g2_decap_8
XFILLER_5_137 VPWR VGND sg13g2_decap_8
XFILLER_1_343 VPWR VGND sg13g2_decap_8
XFILLER_2_888 VPWR VGND sg13g2_decap_4
XFILLER_49_347 VPWR VGND sg13g2_decap_8
XFILLER_18_756 VPWR VGND sg13g2_fill_2
XFILLER_45_531 VPWR VGND sg13g2_decap_8
XFILLER_27_70 VPWR VGND sg13g2_decap_8
XFILLER_17_266 VPWR VGND sg13g2_decap_8
XFILLER_45_575 VPWR VGND sg13g2_fill_1
XFILLER_32_214 VPWR VGND sg13g2_decap_8
XFILLER_13_461 VPWR VGND sg13g2_fill_2
XFILLER_9_410 VPWR VGND sg13g2_decap_8
XFILLER_13_472 VPWR VGND sg13g2_decap_8
XFILLER_43_91 VPWR VGND sg13g2_decap_8
XFILLER_40_280 VPWR VGND sg13g2_decap_8
XFILLER_9_487 VPWR VGND sg13g2_decap_8
X_2561_ net322 VGND VPWR _0507_ state\[123\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2492_ net268 VGND VPWR _0438_ state\[54\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2542__363 VPWR VGND net362 sg13g2_tiehi
X_1512_ VPWR _0175_ daisychain\[27\] VGND sg13g2_inv_1
XFILLER_5_682 VPWR VGND sg13g2_fill_1
X_1443_ VPWR _0251_ daisychain\[96\] VGND sg13g2_inv_1
XFILLER_4_74 VPWR VGND sg13g2_decap_8
X_1374_ VPWR _0058_ state\[37\] VGND sg13g2_inv_1
XFILLER_49_881 VPWR VGND sg13g2_decap_8
XFILLER_36_553 VPWR VGND sg13g2_decap_8
XFILLER_24_737 VPWR VGND sg13g2_fill_1
XFILLER_23_214 VPWR VGND sg13g2_decap_8
XFILLER_23_39 VPWR VGND sg13g2_decap_8
XFILLER_31_291 VPWR VGND sg13g2_decap_8
XFILLER_3_608 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_27_520 VPWR VGND sg13g2_fill_2
XFILLER_15_726 VPWR VGND sg13g2_decap_8
XFILLER_27_564 VPWR VGND sg13g2_fill_2
XFILLER_14_214 VPWR VGND sg13g2_decap_8
Xfanout40 net68 net40 VPWR VGND sg13g2_buf_1
Xfanout51 net52 net51 VPWR VGND sg13g2_buf_1
Xfanout62 net64 net62 VPWR VGND sg13g2_buf_1
Xfanout73 net74 net73 VPWR VGND sg13g2_buf_1
XFILLER_23_792 VPWR VGND sg13g2_decap_4
XFILLER_10_431 VPWR VGND sg13g2_decap_8
Xfanout84 net86 net84 VPWR VGND sg13g2_buf_1
Xfanout95 net96 net95 VPWR VGND sg13g2_buf_1
XFILLER_22_291 VPWR VGND sg13g2_decap_8
XFILLER_6_424 VPWR VGND sg13g2_decap_8
XFILLER_7_969 VPWR VGND sg13g2_decap_8
XFILLER_2_641 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_49_144 VPWR VGND sg13g2_decap_8
X_2537__443 VPWR VGND net442 sg13g2_tiehi
XFILLER_38_91 VPWR VGND sg13g2_decap_8
XFILLER_46_884 VPWR VGND sg13g2_fill_2
XFILLER_45_350 VPWR VGND sg13g2_decap_8
XFILLER_21_707 VPWR VGND sg13g2_fill_1
X_1992_ VGND VPWR net124 daisychain\[111\] _0852_ net34 sg13g2_a21oi_1
XFILLER_20_228 VPWR VGND sg13g2_decap_8
XFILLER_13_291 VPWR VGND sg13g2_decap_8
Xclkload10 VPWR clkload10/Y clknet_leaf_17_clk VGND sg13g2_inv_1
XFILLER_9_284 VPWR VGND sg13g2_decap_8
X_2544_ net330 VGND VPWR _0490_ state\[106\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_6_980 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_2475_ net336 VGND VPWR _0421_ state\[37\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1426_ VPWR _0143_ daisychain\[113\] VGND sg13g2_inv_1
X_1357_ VPWR _0077_ state\[54\] VGND sg13g2_inv_1
XFILLER_18_39 VPWR VGND sg13g2_decap_8
X_1288_ VPWR _0026_ state\[123\] VGND sg13g2_inv_1
XFILLER_36_350 VPWR VGND sg13g2_decap_8
XFILLER_11_228 VPWR VGND sg13g2_decap_8
Xclkload4 VPWR clkload4/Y clknet_leaf_3_clk VGND sg13g2_inv_1
XFILLER_20_751 VPWR VGND sg13g2_fill_1
X_2556__307 VPWR VGND net306 sg13g2_tiehi
XFILLER_47_604 VPWR VGND sg13g2_fill_1
XFILLER_46_147 VPWR VGND sg13g2_decap_8
XFILLER_27_350 VPWR VGND sg13g2_decap_8
XFILLER_15_578 VPWR VGND sg13g2_decap_4
XFILLER_42_364 VPWR VGND sg13g2_decap_8
XFILLER_24_60 VPWR VGND sg13g2_decap_8
X_2313__478 VPWR VGND net477 sg13g2_tiehi
XFILLER_30_559 VPWR VGND sg13g2_fill_2
XFILLER_7_711 VPWR VGND sg13g2_decap_8
XFILLER_6_221 VPWR VGND sg13g2_decap_8
XFILLER_7_799 VPWR VGND sg13g2_decap_8
XFILLER_40_70 VPWR VGND sg13g2_decap_8
XFILLER_6_298 VPWR VGND sg13g2_decap_8
XFILLER_41_7 VPWR VGND sg13g2_decap_8
X_2260_ _1001_ net132 state\[103\] VPWR VGND sg13g2_nand2_1
X_2191_ VGND VPWR _0719_ _0966_ _0452_ net109 sg13g2_a21oi_1
XFILLER_37_147 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_18_361 VPWR VGND sg13g2_decap_8
XFILLER_33_375 VPWR VGND sg13g2_decap_8
X_1975_ net179 _0137_ _0838_ _0839_ VPWR VGND sg13g2_a21o_1
XFILLER_20_18 VPWR VGND sg13g2_decap_8
X_2364__376 VPWR VGND net375 sg13g2_tiehi
X_2527_ net286 VGND VPWR _0473_ state\[89\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2458_ net404 VGND VPWR _0404_ state\[20\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1409_ VPWR _0050_ state\[2\] VGND sg13g2_inv_1
X_2389_ net325 VGND VPWR _0335_ daisychain\[79\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_28_158 VPWR VGND sg13g2_decap_8
XFILLER_25_854 VPWR VGND sg13g2_fill_1
XFILLER_24_375 VPWR VGND sg13g2_decap_8
X_2482__309 VPWR VGND net308 sg13g2_tiehi
XFILLER_3_235 VPWR VGND sg13g2_decap_8
XFILLER_10_95 VPWR VGND sg13g2_decap_8
XFILLER_47_434 VPWR VGND sg13g2_decap_8
XFILLER_19_60 VPWR VGND sg13g2_decap_8
XFILLER_19_158 VPWR VGND sg13g2_decap_8
XFILLER_43_640 VPWR VGND sg13g2_fill_1
XFILLER_35_70 VPWR VGND sg13g2_decap_8
XFILLER_15_375 VPWR VGND sg13g2_decap_8
XFILLER_42_161 VPWR VGND sg13g2_decap_8
XFILLER_30_312 VPWR VGND sg13g2_decap_8
XFILLER_31_857 VPWR VGND sg13g2_fill_1
X_1760_ VGND VPWR net153 daisychain\[53\] _0678_ net63 sg13g2_a21oi_1
XFILLER_30_389 VPWR VGND sg13g2_decap_8
XFILLER_11_581 VPWR VGND sg13g2_decap_4
X_1691_ net184 _0186_ _0625_ _0626_ VPWR VGND sg13g2_a21o_1
XFILLER_7_574 VPWR VGND sg13g2_decap_8
X_2312_ net479 VGND VPWR _0258_ daisychain\[2\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_3_791 VPWR VGND sg13g2_decap_8
X_2243_ VGND VPWR _0797_ _0992_ _0478_ net90 sg13g2_a21oi_1
X_2174_ _0958_ net143 state\[60\] VPWR VGND sg13g2_nand2_1
XFILLER_26_629 VPWR VGND sg13g2_fill_1
XFILLER_15_18 VPWR VGND sg13g2_decap_8
XFILLER_34_662 VPWR VGND sg13g2_decap_8
XFILLER_34_651 VPWR VGND sg13g2_fill_2
XFILLER_34_640 VPWR VGND sg13g2_decap_8
XFILLER_34_695 VPWR VGND sg13g2_decap_8
XFILLER_33_172 VPWR VGND sg13g2_decap_8
XFILLER_22_835 VPWR VGND sg13g2_fill_1
XFILLER_21_312 VPWR VGND sg13g2_decap_8
XFILLER_22_868 VPWR VGND sg13g2_decap_8
XFILLER_21_389 VPWR VGND sg13g2_decap_8
X_1958_ net216 VPWR _0826_ VGND state\[104\] net180 sg13g2_o21ai_1
XFILLER_31_39 VPWR VGND sg13g2_decap_8
X_1889_ VPWR VGND _0774_ net83 _0773_ _0240_ _0342_ net38 sg13g2_a221oi_1
Xoutput17 net17 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_44_448 VPWR VGND sg13g2_decap_8
XFILLER_12_312 VPWR VGND sg13g2_decap_8
XFILLER_31_109 VPWR VGND sg13g2_decap_8
XFILLER_25_695 VPWR VGND sg13g2_fill_2
XFILLER_24_172 VPWR VGND sg13g2_decap_8
XFILLER_8_305 VPWR VGND sg13g2_decap_8
XFILLER_12_389 VPWR VGND sg13g2_decap_8
XdigitalenL.g\[2\].u.inv1 VPWR digitalenL.g\[2\].u.OUTN net6 VGND sg13g2_inv_1
XFILLER_4_511 VPWR VGND sg13g2_decap_8
XFILLER_4_588 VPWR VGND sg13g2_decap_8
XFILLER_47_231 VPWR VGND sg13g2_decap_8
XFILLER_35_437 VPWR VGND sg13g2_decap_8
XFILLER_35_426 VPWR VGND sg13g2_decap_4
XFILLER_46_91 VPWR VGND sg13g2_decap_8
XFILLER_16_662 VPWR VGND sg13g2_decap_8
XFILLER_16_684 VPWR VGND sg13g2_decap_8
XFILLER_31_610 VPWR VGND sg13g2_decap_8
XFILLER_22_109 VPWR VGND sg13g2_decap_8
XFILLER_15_172 VPWR VGND sg13g2_decap_8
X_1812_ VGND VPWR net155 daisychain\[66\] _0717_ net65 sg13g2_a21oi_1
XFILLER_30_186 VPWR VGND sg13g2_decap_8
X_1743_ net186 _0201_ _0664_ _0665_ VPWR VGND sg13g2_a21o_1
XFILLER_8_872 VPWR VGND sg13g2_fill_2
XFILLER_7_63 VPWR VGND sg13g2_decap_8
X_1674_ net209 VPWR _0613_ VGND state\[33\] net163 sg13g2_o21ai_1
XFILLER_8_894 VPWR VGND sg13g2_fill_1
XFILLER_7_371 VPWR VGND sg13g2_decap_8
X_2226_ _0984_ net127 state\[86\] VPWR VGND sg13g2_nand2_1
XFILLER_38_231 VPWR VGND sg13g2_decap_8
X_2157_ VGND VPWR _0668_ _0949_ _0435_ net97 sg13g2_a21oi_1
XFILLER_27_938 VPWR VGND sg13g2_decap_8
XFILLER_26_39 VPWR VGND sg13g2_decap_8
X_2088_ _0915_ net140 state\[17\] VPWR VGND sg13g2_nand2_1
XFILLER_42_908 VPWR VGND sg13g2_fill_2
XFILLER_13_109 VPWR VGND sg13g2_decap_8
XFILLER_34_470 VPWR VGND sg13g2_fill_1
XFILLER_34_492 VPWR VGND sg13g2_fill_1
XFILLER_42_49 VPWR VGND sg13g2_decap_8
XFILLER_22_654 VPWR VGND sg13g2_fill_2
XFILLER_6_809 VPWR VGND sg13g2_decap_4
XFILLER_21_186 VPWR VGND sg13g2_decap_8
XFILLER_5_319 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_49_529 VPWR VGND sg13g2_decap_8
XFILLER_29_242 VPWR VGND sg13g2_decap_8
XFILLER_45_779 VPWR VGND sg13g2_decap_8
XFILLER_45_757 VPWR VGND sg13g2_decap_4
XFILLER_44_245 VPWR VGND sg13g2_decap_8
XFILLER_13_665 VPWR VGND sg13g2_fill_2
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_40_462 VPWR VGND sg13g2_decap_8
XFILLER_12_186 VPWR VGND sg13g2_decap_8
XFILLER_8_179 VPWR VGND sg13g2_decap_8
XFILLER_32_60 VPWR VGND sg13g2_decap_8
X_2464__381 VPWR VGND net380 sg13g2_tiehi
X_1390_ VPWR _0041_ state\[21\] VGND sg13g2_inv_1
XFILLER_4_396 VPWR VGND sg13g2_decap_8
X_2011_ net174 _0147_ _0865_ _0866_ VPWR VGND sg13g2_a21o_1
XFILLER_36_713 VPWR VGND sg13g2_decap_4
XFILLER_35_245 VPWR VGND sg13g2_decap_8
XFILLER_24_919 VPWR VGND sg13g2_fill_2
XFILLER_44_790 VPWR VGND sg13g2_decap_4
X_2844_ daisychain\[126\] net22 VPWR VGND sg13g2_buf_1
X_1726_ net219 VPWR _0652_ VGND state\[46\] net185 sg13g2_o21ai_1
X_1657_ VPWR VGND _0600_ net75 _0599_ _0176_ _0284_ net29 sg13g2_a221oi_1
X_2443__465 VPWR VGND net464 sg13g2_tiehi
X_1588_ VGND VPWR net116 daisychain\[10\] _0549_ net27 sg13g2_a21oi_1
XFILLER_39_551 VPWR VGND sg13g2_decap_8
XFILLER_39_540 VPWR VGND sg13g2_decap_8
XFILLER_37_49 VPWR VGND sg13g2_decap_8
X_2209_ VGND VPWR _0746_ _0975_ _0461_ net108 sg13g2_a21oi_1
XFILLER_39_584 VPWR VGND sg13g2_fill_1
XFILLER_42_727 VPWR VGND sg13g2_fill_2
XFILLER_42_716 VPWR VGND sg13g2_decap_8
XFILLER_26_256 VPWR VGND sg13g2_decap_8
XFILLER_42_749 VPWR VGND sg13g2_decap_8
XFILLER_41_259 VPWR VGND sg13g2_decap_8
XFILLER_23_985 VPWR VGND sg13g2_decap_8
XFILLER_5_116 VPWR VGND sg13g2_decap_8
XFILLER_2_823 VPWR VGND sg13g2_fill_1
XFILLER_2_867 VPWR VGND sg13g2_decap_8
XFILLER_1_322 VPWR VGND sg13g2_decap_8
XFILLER_49_326 VPWR VGND sg13g2_decap_8
XFILLER_1_399 VPWR VGND sg13g2_decap_8
XFILLER_18_735 VPWR VGND sg13g2_decap_8
XFILLER_17_245 VPWR VGND sg13g2_decap_8
XFILLER_45_554 VPWR VGND sg13g2_decap_8
XFILLER_18_779 VPWR VGND sg13g2_fill_2
Xclkbuf_2_0__f_clk clknet_2_0__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_43_70 VPWR VGND sg13g2_decap_8
XFILLER_9_466 VPWR VGND sg13g2_decap_8
X_2560_ net386 VGND VPWR _0506_ state\[122\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_2491_ net272 VGND VPWR _0437_ state\[53\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1511_ VPWR _0176_ daisychain\[28\] VGND sg13g2_inv_1
X_2499__241 VPWR VGND net240 sg13g2_tiehi
X_1442_ VPWR _0252_ daisychain\[97\] VGND sg13g2_inv_1
XFILLER_4_193 VPWR VGND sg13g2_decap_8
X_2323__458 VPWR VGND net457 sg13g2_tiehi
XFILLER_4_53 VPWR VGND sg13g2_decap_8
X_1373_ VPWR _0059_ state\[38\] VGND sg13g2_inv_1
XFILLER_48_392 VPWR VGND sg13g2_decap_8
XFILLER_24_716 VPWR VGND sg13g2_fill_2
XFILLER_32_760 VPWR VGND sg13g2_decap_8
XFILLER_23_18 VPWR VGND sg13g2_decap_8
XFILLER_32_793 VPWR VGND sg13g2_fill_1
XFILLER_31_270 VPWR VGND sg13g2_decap_8
XFILLER_20_955 VPWR VGND sg13g2_decap_8
X_1709_ VPWR VGND _0639_ net94 _0638_ _0191_ _0297_ net49 sg13g2_a221oi_1
X_2478__325 VPWR VGND net324 sg13g2_tiehi
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_329 VPWR VGND sg13g2_decap_8
XFILLER_27_510 VPWR VGND sg13g2_fill_1
X_2374__356 VPWR VGND net355 sg13g2_tiehi
XFILLER_39_392 VPWR VGND sg13g2_decap_8
XFILLER_42_535 VPWR VGND sg13g2_fill_2
Xfanout30 net32 net30 VPWR VGND sg13g2_buf_1
XFILLER_42_568 VPWR VGND sg13g2_fill_1
XFILLER_42_557 VPWR VGND sg13g2_decap_8
XFILLER_10_410 VPWR VGND sg13g2_decap_8
Xfanout41 net43 net41 VPWR VGND sg13g2_buf_1
Xfanout52 net68 net52 VPWR VGND sg13g2_buf_1
Xfanout63 net64 net63 VPWR VGND sg13g2_buf_1
Xfanout74 net78 net74 VPWR VGND sg13g2_buf_1
XFILLER_22_270 VPWR VGND sg13g2_decap_8
Xfanout85 net86 net85 VPWR VGND sg13g2_buf_1
Xfanout96 net112 net96 VPWR VGND sg13g2_buf_1
XFILLER_7_926 VPWR VGND sg13g2_decap_8
XFILLER_10_487 VPWR VGND sg13g2_decap_8
XFILLER_7_948 VPWR VGND sg13g2_decap_8
XFILLER_6_403 VPWR VGND sg13g2_decap_8
XFILLER_13_95 VPWR VGND sg13g2_decap_8
XFILLER_2_620 VPWR VGND sg13g2_decap_8
X_2457__409 VPWR VGND net408 sg13g2_tiehi
XFILLER_49_123 VPWR VGND sg13g2_decap_8
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_38_70 VPWR VGND sg13g2_decap_8
XFILLER_37_329 VPWR VGND sg13g2_decap_8
XFILLER_18_532 VPWR VGND sg13g2_decap_8
XFILLER_46_841 VPWR VGND sg13g2_decap_8
XFILLER_13_270 VPWR VGND sg13g2_decap_8
X_1991_ net170 _0142_ _0850_ _0851_ VPWR VGND sg13g2_a21o_1
XFILLER_20_207 VPWR VGND sg13g2_decap_8
XFILLER_9_263 VPWR VGND sg13g2_decap_8
Xclkload11 clknet_leaf_8_clk clkload11/Y VPWR VGND sg13g2_inv_4
X_2543_ net346 VGND VPWR _0489_ state\[105\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_5_480 VPWR VGND sg13g2_decap_8
XFILLER_47_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_1017 VPWR VGND sg13g2_decap_8
X_2474_ net340 VGND VPWR _0420_ state\[36\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_1425_ VPWR _0144_ daisychain\[114\] VGND sg13g2_inv_1
X_1356_ VPWR _0078_ state\[55\] VGND sg13g2_inv_1
XFILLER_18_18 VPWR VGND sg13g2_decap_8
X_1287_ VPWR _0027_ state\[124\] VGND sg13g2_inv_1
XFILLER_34_39 VPWR VGND sg13g2_decap_8
XFILLER_11_207 VPWR VGND sg13g2_decap_8
Xclkload5 clkload5/Y clknet_leaf_4_clk VPWR VGND sg13g2_inv_2
XFILLER_4_907 VPWR VGND sg13g2_fill_2
XFILLER_4_918 VPWR VGND sg13g2_decap_8
XFILLER_3_417 VPWR VGND sg13g2_decap_4
XFILLER_1_7 VPWR VGND sg13g2_decap_8
Xfanout220 net228 net220 VPWR VGND sg13g2_buf_1
XFILLER_46_126 VPWR VGND sg13g2_decap_8
XFILLER_15_557 VPWR VGND sg13g2_decap_8
XFILLER_42_343 VPWR VGND sg13g2_decap_8
XFILLER_30_538 VPWR VGND sg13g2_fill_1
XFILLER_6_200 VPWR VGND sg13g2_decap_8
XFILLER_10_284 VPWR VGND sg13g2_decap_8
XFILLER_6_277 VPWR VGND sg13g2_decap_8
XFILLER_3_962 VPWR VGND sg13g2_decap_8
X_2190_ _0966_ net156 state\[68\] VPWR VGND sg13g2_nand2_1
XFILLER_2_494 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_decap_8
XFILLER_18_340 VPWR VGND sg13g2_decap_8
XFILLER_46_660 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_19_863 VPWR VGND sg13g2_fill_1
XFILLER_46_693 VPWR VGND sg13g2_decap_8
XFILLER_33_354 VPWR VGND sg13g2_decap_8
X_1974_ net215 VPWR _0838_ VGND state\[108\] net179 sg13g2_o21ai_1
X_2526_ net294 VGND VPWR _0472_ state\[88\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2457_ net408 VGND VPWR _0403_ state\[19\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_1408_ VPWR _0061_ state\[3\] VGND sg13g2_inv_1
XFILLER_29_39 VPWR VGND sg13g2_decap_8
X_2388_ net327 VGND VPWR _0334_ daisychain\[78\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1339_ VPWR _0097_ state\[72\] VGND sg13g2_inv_1
XFILLER_28_137 VPWR VGND sg13g2_decap_8
XFILLER_45_49 VPWR VGND sg13g2_decap_8
XFILLER_24_354 VPWR VGND sg13g2_decap_8
XFILLER_12_549 VPWR VGND sg13g2_decap_8
XFILLER_8_509 VPWR VGND sg13g2_decap_8
XFILLER_3_214 VPWR VGND sg13g2_decap_8
XFILLER_10_74 VPWR VGND sg13g2_decap_8
XFILLER_0_965 VPWR VGND sg13g2_decap_4
XFILLER_0_987 VPWR VGND sg13g2_decap_8
XFILLER_47_413 VPWR VGND sg13g2_decap_8
XFILLER_19_137 VPWR VGND sg13g2_decap_8
XFILLER_15_354 VPWR VGND sg13g2_decap_8
XFILLER_42_140 VPWR VGND sg13g2_decap_8
XFILLER_30_368 VPWR VGND sg13g2_decap_8
X_1690_ net218 VPWR _0625_ VGND state\[37\] net184 sg13g2_o21ai_1
XFILLER_7_553 VPWR VGND sg13g2_decap_8
X_2311_ net481 VGND VPWR _0257_ daisychain\[1\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_32_4 VPWR VGND sg13g2_decap_8
XFILLER_2_291 VPWR VGND sg13g2_decap_8
X_2242_ _0992_ net134 state\[94\] VPWR VGND sg13g2_nand2_1
X_2173_ VGND VPWR _0692_ _0957_ _0443_ net98 sg13g2_a21oi_1
X_2439__481 VPWR VGND net480 sg13g2_tiehi
XFILLER_47_991 VPWR VGND sg13g2_decap_8
XFILLER_46_490 VPWR VGND sg13g2_decap_8
XFILLER_33_151 VPWR VGND sg13g2_decap_8
XFILLER_21_368 VPWR VGND sg13g2_decap_8
X_1957_ VPWR VGND _0825_ net87 _0824_ _0132_ _0359_ net44 sg13g2_a221oi_1
XFILLER_31_18 VPWR VGND sg13g2_decap_8
X_1888_ VGND VPWR net127 daisychain\[85\] _0774_ net38 sg13g2_a21oi_1
Xoutput18 net18 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_0_217 VPWR VGND sg13g2_decap_8
X_2509_ net430 VGND VPWR _0455_ state\[71\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_5_1025 VPWR VGND sg13g2_decap_4
XFILLER_44_427 VPWR VGND sg13g2_decap_8
XFILLER_37_490 VPWR VGND sg13g2_decap_8
XFILLER_25_652 VPWR VGND sg13g2_decap_8
XFILLER_24_151 VPWR VGND sg13g2_decap_8
XFILLER_40_633 VPWR VGND sg13g2_fill_1
XFILLER_40_622 VPWR VGND sg13g2_decap_8
XFILLER_12_368 VPWR VGND sg13g2_decap_8
XFILLER_40_677 VPWR VGND sg13g2_fill_1
XFILLER_40_666 VPWR VGND sg13g2_decap_8
XdigitalenL.g\[2\].u.inv2 VPWR digitalenL.g\[2\].u.OUTP digitalenL.g\[2\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_4_567 VPWR VGND sg13g2_decap_8
XFILLER_21_95 VPWR VGND sg13g2_decap_8
XFILLER_0_762 VPWR VGND sg13g2_fill_2
XFILLER_47_210 VPWR VGND sg13g2_decap_8
XFILLER_47_287 VPWR VGND sg13g2_decap_8
XFILLER_46_70 VPWR VGND sg13g2_decap_8
XFILLER_15_151 VPWR VGND sg13g2_decap_8
XFILLER_31_644 VPWR VGND sg13g2_decap_4
X_1811_ net201 _0219_ _0715_ _0716_ VPWR VGND sg13g2_a21o_1
XFILLER_30_165 VPWR VGND sg13g2_decap_8
X_1742_ net219 VPWR _0664_ VGND state\[50\] net186 sg13g2_o21ai_1
XFILLER_8_851 VPWR VGND sg13g2_fill_1
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_7_350 VPWR VGND sg13g2_decap_8
X_1673_ VPWR VGND _0612_ net76 _0611_ _0181_ _0288_ net30 sg13g2_a221oi_1
X_2402__300 VPWR VGND net299 sg13g2_tiehi
XFILLER_39_711 VPWR VGND sg13g2_decap_8
X_2225_ VGND VPWR _0770_ _0983_ _0469_ net83 sg13g2_a21oi_1
XFILLER_38_210 VPWR VGND sg13g2_decap_8
XFILLER_27_928 VPWR VGND sg13g2_fill_1
XFILLER_27_917 VPWR VGND sg13g2_decap_4
X_2156_ _0949_ net144 state\[51\] VPWR VGND sg13g2_nand2_1
XFILLER_38_287 VPWR VGND sg13g2_decap_8
XFILLER_26_438 VPWR VGND sg13g2_decap_8
XFILLER_26_18 VPWR VGND sg13g2_decap_8
X_2087_ VGND VPWR _0563_ _0914_ _0400_ net85 sg13g2_a21oi_1
Xclkbuf_leaf_18_clk clknet_2_0__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
X_2333__438 VPWR VGND net437 sg13g2_tiehi
XFILLER_22_600 VPWR VGND sg13g2_fill_1
XFILLER_42_28 VPWR VGND sg13g2_decap_8
XFILLER_21_165 VPWR VGND sg13g2_decap_8
XFILLER_1_504 VPWR VGND sg13g2_decap_8
XFILLER_27_1026 VPWR VGND sg13g2_fill_2
XFILLER_49_508 VPWR VGND sg13g2_decap_8
XFILLER_29_221 VPWR VGND sg13g2_decap_8
XFILLER_17_427 VPWR VGND sg13g2_decap_4
XFILLER_18_939 VPWR VGND sg13g2_fill_1
XFILLER_44_224 VPWR VGND sg13g2_decap_8
XFILLER_29_298 VPWR VGND sg13g2_decap_8
XFILLER_13_600 VPWR VGND sg13g2_decap_8
XFILLER_16_95 VPWR VGND sg13g2_decap_8
XFILLER_40_452 VPWR VGND sg13g2_decap_4
XFILLER_12_165 VPWR VGND sg13g2_decap_8
XFILLER_9_659 VPWR VGND sg13g2_fill_2
XFILLER_40_485 VPWR VGND sg13g2_decap_8
X_2384__336 VPWR VGND net335 sg13g2_tiehi
XFILLER_8_158 VPWR VGND sg13g2_decap_8
XFILLER_4_375 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
X_2010_ net212 VPWR _0865_ VGND state\[117\] net173 sg13g2_o21ai_1
X_2471__353 VPWR VGND net352 sg13g2_tiehi
XFILLER_35_224 VPWR VGND sg13g2_decap_8
XFILLER_32_986 VPWR VGND sg13g2_decap_8
XFILLER_31_452 VPWR VGND sg13g2_decap_8
X_2843_ daisychain\[125\] net21 VPWR VGND sg13g2_buf_1
XFILLER_32_997 VPWR VGND sg13g2_decap_4
X_1725_ VPWR VGND _0651_ net95 _0650_ _0195_ _0301_ net50 sg13g2_a221oi_1
X_1656_ VGND VPWR net118 daisychain\[27\] _0600_ net29 sg13g2_a21oi_1
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
X_1587_ net162 _0150_ _0547_ _0548_ VPWR VGND sg13g2_a21o_1
XFILLER_37_28 VPWR VGND sg13g2_decap_8
X_2208_ _0975_ net155 state\[77\] VPWR VGND sg13g2_nand2_1
XFILLER_39_596 VPWR VGND sg13g2_fill_2
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_1006 VPWR VGND sg13g2_fill_1
XFILLER_27_714 VPWR VGND sg13g2_fill_2
X_2139_ VGND VPWR _0641_ _0940_ _0426_ net92 sg13g2_a21oi_1
XFILLER_26_235 VPWR VGND sg13g2_decap_8
X_2450__437 VPWR VGND net436 sg13g2_tiehi
XFILLER_41_238 VPWR VGND sg13g2_decap_8
XFILLER_22_452 VPWR VGND sg13g2_fill_2
XFILLER_1_301 VPWR VGND sg13g2_decap_8
XFILLER_49_305 VPWR VGND sg13g2_decap_8
XFILLER_1_378 VPWR VGND sg13g2_decap_8
XFILLER_17_224 VPWR VGND sg13g2_decap_8
XFILLER_18_769 VPWR VGND sg13g2_fill_1
XFILLER_13_452 VPWR VGND sg13g2_decap_4
XFILLER_32_249 VPWR VGND sg13g2_decap_8
XFILLER_9_445 VPWR VGND sg13g2_decap_8
X_2490_ net276 VGND VPWR _0436_ state\[52\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1510_ VPWR _0177_ daisychain\[29\] VGND sg13g2_inv_1
X_1441_ VPWR _0253_ daisychain\[98\] VGND sg13g2_inv_1
XFILLER_4_32 VPWR VGND sg13g2_decap_8
XFILLER_4_172 VPWR VGND sg13g2_decap_8
X_1372_ VPWR _0060_ state\[39\] VGND sg13g2_inv_1
XFILLER_49_850 VPWR VGND sg13g2_decap_8
XFILLER_48_371 VPWR VGND sg13g2_decap_8
XFILLER_23_249 VPWR VGND sg13g2_decap_8
XFILLER_20_989 VPWR VGND sg13g2_fill_2
X_1708_ VGND VPWR net140 daisychain\[40\] _0639_ net49 sg13g2_a21oi_1
XFILLER_2_109 VPWR VGND sg13g2_decap_8
X_1639_ net195 _0172_ _0586_ _0587_ VPWR VGND sg13g2_a21o_1
XFILLER_48_49 VPWR VGND sg13g2_decap_8
XFILLER_46_308 VPWR VGND sg13g2_decap_8
XFILLER_39_371 VPWR VGND sg13g2_decap_8
XFILLER_27_566 VPWR VGND sg13g2_fill_1
XFILLER_14_249 VPWR VGND sg13g2_decap_8
Xfanout31 net32 net31 VPWR VGND sg13g2_buf_1
Xfanout42 net43 net42 VPWR VGND sg13g2_buf_1
Xfanout53 net55 net53 VPWR VGND sg13g2_buf_1
Xfanout64 net67 net64 VPWR VGND sg13g2_buf_1
XFILLER_23_761 VPWR VGND sg13g2_decap_8
Xfanout75 net77 net75 VPWR VGND sg13g2_buf_1
Xfanout86 net91 net86 VPWR VGND sg13g2_buf_1
Xfanout97 net101 net97 VPWR VGND sg13g2_buf_1
XFILLER_7_905 VPWR VGND sg13g2_decap_8
XFILLER_10_466 VPWR VGND sg13g2_decap_8
XFILLER_13_74 VPWR VGND sg13g2_decap_8
XFILLER_6_459 VPWR VGND sg13g2_decap_8
XFILLER_49_102 VPWR VGND sg13g2_decap_8
XFILLER_2_698 VPWR VGND sg13g2_decap_4
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_49_179 VPWR VGND sg13g2_decap_8
XFILLER_46_820 VPWR VGND sg13g2_decap_8
XFILLER_37_308 VPWR VGND sg13g2_decap_8
XFILLER_18_544 VPWR VGND sg13g2_decap_8
XFILLER_46_853 VPWR VGND sg13g2_fill_2
XFILLER_46_875 VPWR VGND sg13g2_fill_2
XFILLER_45_385 VPWR VGND sg13g2_decap_8
XFILLER_33_525 VPWR VGND sg13g2_decap_8
X_1990_ net212 VPWR _0850_ VGND state\[112\] net170 sg13g2_o21ai_1
XFILLER_9_242 VPWR VGND sg13g2_decap_8
XFILLER_41_591 VPWR VGND sg13g2_fill_1
Xclkload12 VPWR clkload12/Y clknet_leaf_9_clk VGND sg13g2_inv_1
X_2542_ net362 VGND VPWR _0488_ state\[104\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2473_ net344 VGND VPWR _0419_ state\[35\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1424_ VPWR _0145_ daisychain\[115\] VGND sg13g2_inv_1
X_1355_ VPWR _0079_ state\[56\] VGND sg13g2_inv_1
XFILLER_28_319 VPWR VGND sg13g2_decap_8
X_1286_ VPWR _0028_ state\[125\] VGND sg13g2_inv_1
XFILLER_36_385 VPWR VGND sg13g2_decap_8
XFILLER_34_18 VPWR VGND sg13g2_decap_8
XFILLER_24_525 VPWR VGND sg13g2_decap_4
XFILLER_24_558 VPWR VGND sg13g2_fill_1
X_2410__284 VPWR VGND net283 sg13g2_tiehi
Xclkload6 VPWR clkload6/Y clknet_leaf_7_clk VGND sg13g2_inv_1
XFILLER_30_1022 VPWR VGND sg13g2_decap_8
Xfanout221 net222 net221 VPWR VGND sg13g2_buf_1
Xfanout210 net228 net210 VPWR VGND sg13g2_buf_1
XFILLER_19_319 VPWR VGND sg13g2_decap_8
XFILLER_46_105 VPWR VGND sg13g2_decap_8
XFILLER_43_834 VPWR VGND sg13g2_fill_2
XFILLER_27_385 VPWR VGND sg13g2_decap_8
XFILLER_42_322 VPWR VGND sg13g2_decap_8
XFILLER_11_731 VPWR VGND sg13g2_decap_8
XFILLER_42_399 VPWR VGND sg13g2_decap_8
XFILLER_24_95 VPWR VGND sg13g2_decap_8
XFILLER_10_263 VPWR VGND sg13g2_decap_8
XFILLER_6_256 VPWR VGND sg13g2_decap_8
XFILLER_2_473 VPWR VGND sg13g2_decap_8
XFILLER_49_81 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_18_385 VPWR VGND sg13g2_decap_8
X_2511__415 VPWR VGND net414 sg13g2_tiehi
XFILLER_45_182 VPWR VGND sg13g2_decap_8
XFILLER_33_333 VPWR VGND sg13g2_decap_8
X_1973_ VPWR VGND _0837_ net87 _0836_ _0136_ _0363_ net44 sg13g2_a221oi_1
XFILLER_6_790 VPWR VGND sg13g2_decap_8
X_2525_ net302 VGND VPWR _0471_ state\[87\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2456_ net412 VGND VPWR _0402_ state\[18\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_1407_ VPWR _0072_ state\[4\] VGND sg13g2_inv_1
XFILLER_29_18 VPWR VGND sg13g2_decap_8
X_2387_ net329 VGND VPWR _0333_ daisychain\[77\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1338_ VPWR _0098_ state\[73\] VGND sg13g2_inv_1
XFILLER_28_116 VPWR VGND sg13g2_decap_8
XFILLER_45_28 VPWR VGND sg13g2_decap_8
XFILLER_43_119 VPWR VGND sg13g2_decap_8
XFILLER_25_812 VPWR VGND sg13g2_decap_8
XFILLER_36_182 VPWR VGND sg13g2_decap_8
XFILLER_24_333 VPWR VGND sg13g2_decap_8
XFILLER_12_528 VPWR VGND sg13g2_decap_8
X_2312__480 VPWR VGND net479 sg13g2_tiehi
X_2343__418 VPWR VGND net417 sg13g2_tiehi
X_2523__319 VPWR VGND net318 sg13g2_tiehi
XFILLER_4_738 VPWR VGND sg13g2_fill_2
XFILLER_10_53 VPWR VGND sg13g2_decap_8
XFILLER_0_944 VPWR VGND sg13g2_decap_8
XFILLER_19_116 VPWR VGND sg13g2_decap_8
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_19_95 VPWR VGND sg13g2_decap_8
XFILLER_28_694 VPWR VGND sg13g2_decap_8
XFILLER_15_333 VPWR VGND sg13g2_decap_8
XFILLER_43_631 VPWR VGND sg13g2_decap_8
XFILLER_27_182 VPWR VGND sg13g2_decap_8
XFILLER_42_196 VPWR VGND sg13g2_decap_8
XFILLER_11_550 VPWR VGND sg13g2_decap_4
XFILLER_30_347 VPWR VGND sg13g2_decap_8
XFILLER_7_532 VPWR VGND sg13g2_decap_8
X_2310_ net482 VGND VPWR _0256_ daisychain\[0\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2241_ VGND VPWR _0794_ _0991_ _0477_ net104 sg13g2_a21oi_1
XFILLER_2_270 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
X_2172_ _0957_ net143 state\[59\] VPWR VGND sg13g2_nand2_1
X_2394__316 VPWR VGND net315 sg13g2_tiehi
XFILLER_38_447 VPWR VGND sg13g2_fill_2
XFILLER_18_193 VPWR VGND sg13g2_decap_8
XFILLER_33_130 VPWR VGND sg13g2_decap_8
X_1956_ VGND VPWR net134 daisychain\[102\] _0825_ net47 sg13g2_a21oi_1
XFILLER_21_347 VPWR VGND sg13g2_decap_8
X_1887_ net174 _0240_ _0772_ _0773_ VPWR VGND sg13g2_a21o_1
X_2446__453 VPWR VGND net452 sg13g2_tiehi
Xoutput19 net19 uo_out[3] VPWR VGND sg13g2_buf_1
X_2508_ net438 VGND VPWR _0454_ state\[70\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2439_ net480 VGND VPWR _0385_ state\[1\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_29_403 VPWR VGND sg13g2_decap_8
XFILLER_29_414 VPWR VGND sg13g2_fill_1
XFILLER_29_458 VPWR VGND sg13g2_decap_4
XFILLER_44_406 VPWR VGND sg13g2_decap_8
XFILLER_24_130 VPWR VGND sg13g2_decap_8
XFILLER_12_347 VPWR VGND sg13g2_decap_8
XFILLER_21_892 VPWR VGND sg13g2_fill_1
XFILLER_21_870 VPWR VGND sg13g2_fill_2
XFILLER_4_546 VPWR VGND sg13g2_decap_8
XFILLER_21_74 VPWR VGND sg13g2_decap_8
XFILLER_48_745 VPWR VGND sg13g2_fill_2
XFILLER_48_723 VPWR VGND sg13g2_fill_2
XFILLER_47_266 VPWR VGND sg13g2_decap_8
XFILLER_35_406 VPWR VGND sg13g2_decap_8
XFILLER_44_940 VPWR VGND sg13g2_fill_2
XFILLER_15_130 VPWR VGND sg13g2_decap_8
XFILLER_43_483 VPWR VGND sg13g2_decap_4
X_1810_ net225 VPWR _0715_ VGND state\[67\] net201 sg13g2_o21ai_1
XFILLER_30_144 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
X_1741_ VPWR VGND _0663_ net99 _0662_ _0199_ _0305_ net55 sg13g2_a221oi_1
X_1672_ VGND VPWR net119 daisychain\[31\] _0612_ net30 sg13g2_a21oi_1
XFILLER_8_885 VPWR VGND sg13g2_fill_1
XFILLER_7_98 VPWR VGND sg13g2_decap_8
X_2224_ _0983_ net126 state\[85\] VPWR VGND sg13g2_nand2_1
XFILLER_39_723 VPWR VGND sg13g2_decap_8
X_2155_ VGND VPWR _0665_ _0948_ _0434_ net93 sg13g2_a21oi_1
XFILLER_38_266 VPWR VGND sg13g2_decap_8
XFILLER_26_417 VPWR VGND sg13g2_decap_8
X_2086_ _0914_ net120 state\[16\] VPWR VGND sg13g2_nand2_1
XFILLER_34_483 VPWR VGND sg13g2_decap_8
XFILLER_22_612 VPWR VGND sg13g2_decap_8
XFILLER_21_144 VPWR VGND sg13g2_decap_8
X_1939_ net180 _0254_ _0811_ _0812_ VPWR VGND sg13g2_a21o_1
XFILLER_29_200 VPWR VGND sg13g2_decap_8
XFILLER_18_918 VPWR VGND sg13g2_fill_1
XFILLER_17_406 VPWR VGND sg13g2_decap_8
XFILLER_44_203 VPWR VGND sg13g2_decap_8
XFILLER_29_277 VPWR VGND sg13g2_decap_8
XFILLER_16_74 VPWR VGND sg13g2_decap_8
XFILLER_12_144 VPWR VGND sg13g2_decap_8
XFILLER_9_616 VPWR VGND sg13g2_fill_2
XFILLER_9_605 VPWR VGND sg13g2_decap_8
XFILLER_9_627 VPWR VGND sg13g2_fill_1
XFILLER_8_137 VPWR VGND sg13g2_decap_8
XFILLER_32_95 VPWR VGND sg13g2_decap_8
XFILLER_4_354 VPWR VGND sg13g2_decap_8
X_2501__233 VPWR VGND net232 sg13g2_tiehi
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_48_542 VPWR VGND sg13g2_fill_2
XFILLER_35_203 VPWR VGND sg13g2_decap_8
XFILLER_16_450 VPWR VGND sg13g2_decap_8
XFILLER_43_280 VPWR VGND sg13g2_decap_8
X_2842_ daisychain\[124\] net20 VPWR VGND sg13g2_buf_1
XFILLER_31_475 VPWR VGND sg13g2_fill_1
X_1724_ VGND VPWR net141 daisychain\[44\] _0651_ net50 sg13g2_a21oi_1
X_1655_ net165 _0176_ _0598_ _0599_ VPWR VGND sg13g2_a21o_1
X_1586_ net206 VPWR _0547_ VGND state\[11\] net162 sg13g2_o21ai_1
XFILLER_39_520 VPWR VGND sg13g2_decap_4
X_2207_ VGND VPWR _0743_ _0974_ _0460_ net106 sg13g2_a21oi_1
X_2138_ _0940_ net138 state\[42\] VPWR VGND sg13g2_nand2_1
XFILLER_26_214 VPWR VGND sg13g2_decap_8
X_2069_ VGND VPWR _0536_ _0905_ _0391_ net70 sg13g2_a21oi_1
XFILLER_41_217 VPWR VGND sg13g2_decap_8
XFILLER_23_932 VPWR VGND sg13g2_fill_1
XFILLER_34_291 VPWR VGND sg13g2_decap_8
XFILLER_23_954 VPWR VGND sg13g2_decap_8
XFILLER_22_431 VPWR VGND sg13g2_decap_8
XFILLER_10_626 VPWR VGND sg13g2_fill_1
XFILLER_22_486 VPWR VGND sg13g2_fill_1
XFILLER_10_648 VPWR VGND sg13g2_decap_8
XFILLER_2_836 VPWR VGND sg13g2_decap_8
XFILLER_1_357 VPWR VGND sg13g2_decap_8
X_2420__264 VPWR VGND net263 sg13g2_tiehi
XFILLER_17_203 VPWR VGND sg13g2_decap_8
XFILLER_33_707 VPWR VGND sg13g2_decap_4
XFILLER_27_84 VPWR VGND sg13g2_decap_8
XFILLER_32_228 VPWR VGND sg13g2_decap_8
XFILLER_26_770 VPWR VGND sg13g2_fill_2
XFILLER_13_431 VPWR VGND sg13g2_decap_8
XFILLER_25_291 VPWR VGND sg13g2_decap_8
XFILLER_13_486 VPWR VGND sg13g2_decap_8
XFILLER_9_424 VPWR VGND sg13g2_decap_8
XFILLER_40_294 VPWR VGND sg13g2_decap_8
XFILLER_4_151 VPWR VGND sg13g2_decap_8
X_1440_ VPWR _0254_ daisychain\[99\] VGND sg13g2_inv_1
XFILLER_5_696 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_decap_8
X_1371_ VPWR _0062_ state\[40\] VGND sg13g2_inv_1
XFILLER_4_88 VPWR VGND sg13g2_decap_8
XFILLER_49_895 VPWR VGND sg13g2_fill_1
XFILLER_48_350 VPWR VGND sg13g2_decap_8
XFILLER_36_545 VPWR VGND sg13g2_fill_1
XFILLER_23_228 VPWR VGND sg13g2_decap_8
XFILLER_16_291 VPWR VGND sg13g2_decap_8
X_1707_ net187 _0191_ _0637_ _0638_ VPWR VGND sg13g2_a21o_1
X_1638_ net223 VPWR _0586_ VGND state\[24\] net195 sg13g2_o21ai_1
X_1569_ VPWR VGND _0534_ net70 _0533_ _0222_ _0262_ net25 sg13g2_a221oi_1
XFILLER_48_28 VPWR VGND sg13g2_decap_8
XFILLER_39_350 VPWR VGND sg13g2_decap_8
XFILLER_27_545 VPWR VGND sg13g2_decap_8
XFILLER_27_578 VPWR VGND sg13g2_decap_8
XFILLER_14_228 VPWR VGND sg13g2_decap_8
Xfanout43 net48 net43 VPWR VGND sg13g2_buf_1
Xfanout54 net55 net54 VPWR VGND sg13g2_buf_1
Xfanout65 net67 net65 VPWR VGND sg13g2_buf_1
Xfanout32 net33 net32 VPWR VGND sg13g2_buf_1
XFILLER_23_784 VPWR VGND sg13g2_decap_4
Xfanout76 net77 net76 VPWR VGND sg13g2_buf_1
Xfanout87 net90 net87 VPWR VGND sg13g2_buf_1
Xfanout98 net101 net98 VPWR VGND sg13g2_buf_1
XFILLER_10_445 VPWR VGND sg13g2_decap_8
XFILLER_13_53 VPWR VGND sg13g2_decap_8
X_2565__355 VPWR VGND net354 sg13g2_tiehi
XFILLER_6_438 VPWR VGND sg13g2_decap_8
XFILLER_2_655 VPWR VGND sg13g2_decap_8
XFILLER_1_154 VPWR VGND sg13g2_decap_8
X_2322__460 VPWR VGND net459 sg13g2_tiehi
XFILLER_18_501 VPWR VGND sg13g2_fill_2
XFILLER_49_158 VPWR VGND sg13g2_decap_8
XFILLER_46_898 VPWR VGND sg13g2_fill_2
XFILLER_45_364 VPWR VGND sg13g2_decap_8
XFILLER_33_537 VPWR VGND sg13g2_fill_2
XFILLER_9_221 VPWR VGND sg13g2_decap_8
XFILLER_9_298 VPWR VGND sg13g2_decap_8
X_2541_ net378 VGND VPWR _0487_ state\[103\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2472_ net348 VGND VPWR _0418_ state\[34\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_1423_ VPWR _0146_ daisychain\[116\] VGND sg13g2_inv_1
X_1354_ VPWR _0080_ state\[57\] VGND sg13g2_inv_1
X_1285_ VPWR _0029_ state\[126\] VGND sg13g2_inv_1
XFILLER_36_364 VPWR VGND sg13g2_decap_8
Xclkload7 clkload7/Y clknet_leaf_13_clk VPWR VGND sg13g2_inv_2
Xfanout222 net228 net222 VPWR VGND sg13g2_buf_1
Xfanout211 net212 net211 VPWR VGND sg13g2_buf_1
Xfanout200 net203 net200 VPWR VGND sg13g2_buf_1
XFILLER_8_1024 VPWR VGND sg13g2_decap_4
XFILLER_8_1002 VPWR VGND sg13g2_fill_1
XFILLER_15_504 VPWR VGND sg13g2_fill_2
XFILLER_42_301 VPWR VGND sg13g2_decap_8
XFILLER_27_364 VPWR VGND sg13g2_decap_8
XFILLER_43_868 VPWR VGND sg13g2_decap_8
XFILLER_42_378 VPWR VGND sg13g2_decap_8
XFILLER_30_529 VPWR VGND sg13g2_decap_8
XFILLER_24_74 VPWR VGND sg13g2_decap_8
XFILLER_10_242 VPWR VGND sg13g2_decap_8
XFILLER_7_725 VPWR VGND sg13g2_decap_4
XFILLER_6_235 VPWR VGND sg13g2_decap_8
XFILLER_7_769 VPWR VGND sg13g2_decap_8
XFILLER_40_84 VPWR VGND sg13g2_decap_8
XFILLER_2_452 VPWR VGND sg13g2_decap_8
XFILLER_49_60 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_19_810 VPWR VGND sg13g2_decap_8
XFILLER_19_854 VPWR VGND sg13g2_decap_4
XFILLER_18_375 VPWR VGND sg13g2_decap_4
XFILLER_45_161 VPWR VGND sg13g2_decap_8
XFILLER_33_312 VPWR VGND sg13g2_decap_8
X_1972_ VGND VPWR net131 daisychain\[106\] _0837_ net44 sg13g2_a21oi_1
XFILLER_33_389 VPWR VGND sg13g2_decap_8
XdigitalenH.g\[0\].u.inv1 VPWR digitalenH.g\[0\].u.OUTN net7 VGND sg13g2_inv_1
X_2524_ net310 VGND VPWR _0470_ state\[86\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_46_0 VPWR VGND sg13g2_decap_8
X_2455_ net416 VGND VPWR _0401_ state\[17\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2386_ net331 VGND VPWR _0332_ daisychain\[76\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1406_ VPWR _0083_ state\[5\] VGND sg13g2_inv_1
X_1337_ VPWR _0099_ state\[74\] VGND sg13g2_inv_1
XFILLER_37_673 VPWR VGND sg13g2_fill_1
XFILLER_36_161 VPWR VGND sg13g2_decap_8
XFILLER_24_312 VPWR VGND sg13g2_decap_8
XFILLER_12_507 VPWR VGND sg13g2_decap_8
XFILLER_24_389 VPWR VGND sg13g2_decap_8
XFILLER_10_32 VPWR VGND sg13g2_decap_8
XFILLER_3_249 VPWR VGND sg13g2_decap_8
XFILLER_0_901 VPWR VGND sg13g2_decap_8
XFILLER_0_912 VPWR VGND sg13g2_decap_8
XFILLER_19_74 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_decap_8
XFILLER_43_610 VPWR VGND sg13g2_decap_8
XFILLER_34_109 VPWR VGND sg13g2_decap_8
XFILLER_27_161 VPWR VGND sg13g2_decap_8
XFILLER_15_312 VPWR VGND sg13g2_decap_8
XFILLER_43_676 VPWR VGND sg13g2_decap_4
XFILLER_35_84 VPWR VGND sg13g2_decap_8
XFILLER_15_389 VPWR VGND sg13g2_decap_8
XFILLER_43_698 VPWR VGND sg13g2_fill_2
XFILLER_42_175 VPWR VGND sg13g2_decap_8
XFILLER_30_326 VPWR VGND sg13g2_decap_8
XFILLER_7_511 VPWR VGND sg13g2_decap_8
XFILLER_7_588 VPWR VGND sg13g2_decap_8
X_2240_ _0991_ net150 state\[93\] VPWR VGND sg13g2_nand2_1
XFILLER_18_4 VPWR VGND sg13g2_decap_8
X_2171_ VGND VPWR _0689_ _0956_ _0442_ net97 sg13g2_a21oi_1
X_2474__341 VPWR VGND net340 sg13g2_tiehi
XFILLER_19_651 VPWR VGND sg13g2_fill_2
XFILLER_25_109 VPWR VGND sg13g2_decap_8
XFILLER_18_172 VPWR VGND sg13g2_decap_8
XFILLER_34_676 VPWR VGND sg13g2_decap_4
XFILLER_33_186 VPWR VGND sg13g2_decap_8
XFILLER_21_326 VPWR VGND sg13g2_decap_8
X_1955_ net181 _0132_ _0823_ _0824_ VPWR VGND sg13g2_a21o_1
XFILLER_30_860 VPWR VGND sg13g2_fill_1
X_1886_ net212 VPWR _0772_ VGND state\[86\] net174 sg13g2_o21ai_1
X_2507_ net446 VGND VPWR _0453_ state\[69\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2438_ net483 VGND VPWR _0384_ state\[0\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2369_ net365 VGND VPWR _0315_ daisychain\[59\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_16_109 VPWR VGND sg13g2_decap_8
X_2453__425 VPWR VGND net424 sg13g2_tiehi
XFILLER_12_326 VPWR VGND sg13g2_decap_8
XFILLER_24_186 VPWR VGND sg13g2_decap_8
XFILLER_8_319 VPWR VGND sg13g2_decap_8
XANTENNA_60 VPWR VGND daisychain\[126\] sg13g2_antennanp
XFILLER_4_525 VPWR VGND sg13g2_decap_8
XFILLER_21_53 VPWR VGND sg13g2_decap_8
XFILLER_0_720 VPWR VGND sg13g2_decap_4
XFILLER_43_1000 VPWR VGND sg13g2_fill_2
XFILLER_0_775 VPWR VGND sg13g2_fill_2
XFILLER_0_786 VPWR VGND sg13g2_decap_8
XFILLER_47_245 VPWR VGND sg13g2_decap_8
XFILLER_43_462 VPWR VGND sg13g2_fill_2
XFILLER_15_186 VPWR VGND sg13g2_decap_8
XFILLER_16_698 VPWR VGND sg13g2_decap_4
X_2430__244 VPWR VGND net243 sg13g2_tiehi
XFILLER_44_996 VPWR VGND sg13g2_fill_1
XFILLER_31_668 VPWR VGND sg13g2_decap_8
XFILLER_30_123 VPWR VGND sg13g2_decap_8
X_1740_ VGND VPWR net145 daisychain\[48\] _0663_ net55 sg13g2_a21oi_1
XFILLER_8_864 VPWR VGND sg13g2_fill_1
XFILLER_8_842 VPWR VGND sg13g2_fill_1
X_1671_ net167 _0181_ _0610_ _0611_ VPWR VGND sg13g2_a21o_1
XFILLER_7_77 VPWR VGND sg13g2_decap_8
XFILLER_7_385 VPWR VGND sg13g2_decap_8
XFILLER_3_580 VPWR VGND sg13g2_decap_8
X_2223_ VGND VPWR _0767_ _0982_ _0468_ net79 sg13g2_a21oi_1
X_2154_ _0948_ net139 state\[50\] VPWR VGND sg13g2_nand2_1
XFILLER_38_245 VPWR VGND sg13g2_decap_8
X_2085_ VGND VPWR _0560_ _0913_ _0399_ net77 sg13g2_a21oi_1
XFILLER_19_492 VPWR VGND sg13g2_decap_8
XFILLER_21_123 VPWR VGND sg13g2_decap_8
X_1938_ net214 VPWR _0811_ VGND state\[99\] net178 sg13g2_o21ai_1
X_1869_ VPWR VGND _0759_ net105 _0758_ _0235_ _0337_ net60 sg13g2_a221oi_1
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_1006 VPWR VGND sg13g2_fill_2
XFILLER_1_539 VPWR VGND sg13g2_decap_8
XFILLER_29_256 VPWR VGND sg13g2_decap_8
XFILLER_16_53 VPWR VGND sg13g2_decap_8
XFILLER_44_259 VPWR VGND sg13g2_decap_8
XFILLER_26_963 VPWR VGND sg13g2_decap_8
XFILLER_12_123 VPWR VGND sg13g2_decap_8
XFILLER_8_116 VPWR VGND sg13g2_decap_8
XFILLER_32_74 VPWR VGND sg13g2_decap_8
XFILLER_4_333 VPWR VGND sg13g2_decap_8
XFILLER_35_259 VPWR VGND sg13g2_decap_8
XFILLER_31_410 VPWR VGND sg13g2_decap_8
X_2332__440 VPWR VGND net439 sg13g2_tiehi
X_2841_ daisychain\[123\] net19 VPWR VGND sg13g2_buf_1
XFILLER_12_690 VPWR VGND sg13g2_decap_8
X_1723_ net185 _0195_ _0649_ _0650_ VPWR VGND sg13g2_a21o_1
XFILLER_7_182 VPWR VGND sg13g2_decap_8
X_1654_ net207 VPWR _0598_ VGND state\[28\] net165 sg13g2_o21ai_1
X_1585_ VPWR VGND _0546_ net74 _0545_ _0139_ _0266_ net28 sg13g2_a221oi_1
XFILLER_39_510 VPWR VGND sg13g2_decap_4
X_2206_ _0974_ net154 state\[76\] VPWR VGND sg13g2_nand2_1
XFILLER_39_532 VPWR VGND sg13g2_fill_1
XFILLER_2_1019 VPWR VGND sg13g2_decap_8
X_2137_ VGND VPWR _0638_ _0939_ _0425_ net92 sg13g2_a21oi_1
X_2068_ _0905_ net114 state\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_34_270 VPWR VGND sg13g2_decap_8
XFILLER_23_911 VPWR VGND sg13g2_decap_8
XFILLER_22_410 VPWR VGND sg13g2_decap_8
XFILLER_1_336 VPWR VGND sg13g2_decap_8
XFILLER_18_749 VPWR VGND sg13g2_decap_8
XFILLER_45_524 VPWR VGND sg13g2_decap_8
XFILLER_27_63 VPWR VGND sg13g2_decap_8
XFILLER_17_259 VPWR VGND sg13g2_decap_8
XFILLER_45_568 VPWR VGND sg13g2_decap_8
XFILLER_13_410 VPWR VGND sg13g2_decap_8
XFILLER_32_207 VPWR VGND sg13g2_decap_8
XFILLER_25_270 VPWR VGND sg13g2_decap_8
XFILLER_9_403 VPWR VGND sg13g2_decap_8
XFILLER_43_84 VPWR VGND sg13g2_decap_8
XFILLER_40_273 VPWR VGND sg13g2_decap_8
XFILLER_5_675 VPWR VGND sg13g2_decap_8
XFILLER_4_130 VPWR VGND sg13g2_decap_8
X_1370_ VPWR _0063_ state\[41\] VGND sg13g2_inv_1
XFILLER_4_67 VPWR VGND sg13g2_decap_8
XFILLER_49_863 VPWR VGND sg13g2_fill_2
XFILLER_23_207 VPWR VGND sg13g2_decap_8
XFILLER_16_270 VPWR VGND sg13g2_decap_8
XFILLER_31_284 VPWR VGND sg13g2_decap_8
X_1706_ net218 VPWR _0637_ VGND state\[41\] net186 sg13g2_o21ai_1
X_1637_ VPWR VGND _0585_ net102 _0584_ _0171_ _0279_ net57 sg13g2_a221oi_1
X_1568_ VGND VPWR net114 daisychain\[5\] _0534_ net25 sg13g2_a21oi_1
X_1499_ VPWR _0190_ daisychain\[40\] VGND sg13g2_inv_1
XFILLER_27_535 VPWR VGND sg13g2_decap_4
XFILLER_14_207 VPWR VGND sg13g2_decap_8
Xfanout44 net48 net44 VPWR VGND sg13g2_buf_1
Xfanout55 net56 net55 VPWR VGND sg13g2_buf_1
Xfanout33 net68 net33 VPWR VGND sg13g2_buf_1
XFILLER_10_424 VPWR VGND sg13g2_decap_8
XFILLER_13_32 VPWR VGND sg13g2_decap_8
Xfanout66 net67 net66 VPWR VGND sg13g2_buf_1
Xfanout77 net78 net77 VPWR VGND sg13g2_buf_1
Xfanout88 net90 net88 VPWR VGND sg13g2_buf_1
Xfanout99 net101 net99 VPWR VGND sg13g2_buf_1
XFILLER_22_284 VPWR VGND sg13g2_decap_8
XFILLER_6_417 VPWR VGND sg13g2_decap_8
XFILLER_2_634 VPWR VGND sg13g2_decap_8
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_49_137 VPWR VGND sg13g2_decap_8
XFILLER_38_84 VPWR VGND sg13g2_decap_8
XFILLER_46_866 VPWR VGND sg13g2_decap_4
XFILLER_45_343 VPWR VGND sg13g2_decap_8
XFILLER_9_200 VPWR VGND sg13g2_decap_8
XFILLER_13_284 VPWR VGND sg13g2_decap_8
XFILLER_9_277 VPWR VGND sg13g2_decap_8
X_2540_ net394 VGND VPWR _0486_ state\[102\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2471_ net352 VGND VPWR _0417_ state\[33\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_1422_ VPWR _0147_ daisychain\[117\] VGND sg13g2_inv_1
XFILLER_5_494 VPWR VGND sg13g2_decap_8
X_1353_ VPWR _0081_ state\[58\] VGND sg13g2_inv_1
X_1284_ VPWR _1026_ net211 VGND sg13g2_inv_1
XFILLER_49_693 VPWR VGND sg13g2_decap_8
XFILLER_36_343 VPWR VGND sg13g2_decap_8
XFILLER_24_549 VPWR VGND sg13g2_decap_4
X_2449__441 VPWR VGND net440 sg13g2_tiehi
Xclkload8 clknet_leaf_14_clk clkload8/Y VPWR VGND sg13g2_inv_4
Xfanout223 net227 net223 VPWR VGND sg13g2_buf_1
Xfanout212 net217 net212 VPWR VGND sg13g2_buf_1
Xfanout201 net203 net201 VPWR VGND sg13g2_buf_1
XFILLER_8_1014 VPWR VGND sg13g2_fill_1
XFILLER_28_811 VPWR VGND sg13g2_decap_8
XFILLER_27_343 VPWR VGND sg13g2_decap_8
XFILLER_42_357 VPWR VGND sg13g2_decap_8
XFILLER_30_519 VPWR VGND sg13g2_fill_2
XFILLER_30_508 VPWR VGND sg13g2_fill_2
XFILLER_24_53 VPWR VGND sg13g2_decap_8
XFILLER_10_221 VPWR VGND sg13g2_decap_8
XFILLER_6_214 VPWR VGND sg13g2_decap_8
XFILLER_10_298 VPWR VGND sg13g2_decap_8
XFILLER_40_63 VPWR VGND sg13g2_decap_8
XFILLER_3_921 VPWR VGND sg13g2_fill_2
XFILLER_2_431 VPWR VGND sg13g2_decap_8
XFILLER_38_619 VPWR VGND sg13g2_decap_4
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_18_354 VPWR VGND sg13g2_decap_8
XFILLER_45_140 VPWR VGND sg13g2_decap_8
XFILLER_19_888 VPWR VGND sg13g2_decap_4
XFILLER_33_368 VPWR VGND sg13g2_decap_8
X_1971_ net179 _0136_ _0835_ _0836_ VPWR VGND sg13g2_a21o_1
X_2523_ net318 VGND VPWR _0469_ state\[85\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XdigitalenH.g\[0\].u.inv2 VPWR digitalenH.g\[0\].u.OUTP digitalenH.g\[0\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_5_291 VPWR VGND sg13g2_decap_8
X_2454_ net420 VGND VPWR _0400_ state\[16\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2385_ net333 VGND VPWR _0331_ daisychain\[75\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_1405_ VPWR _0094_ state\[6\] VGND sg13g2_inv_1
XFILLER_39_0 VPWR VGND sg13g2_decap_8
X_1336_ VPWR _0100_ state\[75\] VGND sg13g2_inv_1
Xinput1 rst_n net1 VPWR VGND sg13g2_buf_1
XFILLER_37_685 VPWR VGND sg13g2_decap_4
XFILLER_37_663 VPWR VGND sg13g2_fill_2
XFILLER_36_140 VPWR VGND sg13g2_decap_8
XFILLER_24_368 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_decap_8
XFILLER_3_228 VPWR VGND sg13g2_decap_8
XFILLER_10_88 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_19_53 VPWR VGND sg13g2_decap_8
XFILLER_43_600 VPWR VGND sg13g2_fill_1
XFILLER_27_140 VPWR VGND sg13g2_decap_8
XFILLER_15_368 VPWR VGND sg13g2_decap_8
XFILLER_42_154 VPWR VGND sg13g2_decap_8
XFILLER_35_63 VPWR VGND sg13g2_decap_8
XFILLER_30_305 VPWR VGND sg13g2_decap_8
XFILLER_11_574 VPWR VGND sg13g2_decap_8
XFILLER_11_585 VPWR VGND sg13g2_fill_2
XFILLER_7_567 VPWR VGND sg13g2_decap_8
X_2170_ _0956_ net144 state\[58\] VPWR VGND sg13g2_nand2_1
XFILLER_20_1012 VPWR VGND sg13g2_decap_8
XFILLER_18_151 VPWR VGND sg13g2_decap_8
XFILLER_47_961 VPWR VGND sg13g2_decap_8
XFILLER_34_633 VPWR VGND sg13g2_decap_8
XFILLER_34_611 VPWR VGND sg13g2_decap_8
X_2515__383 VPWR VGND net382 sg13g2_tiehi
XFILLER_22_817 VPWR VGND sg13g2_fill_2
XFILLER_33_165 VPWR VGND sg13g2_decap_8
XFILLER_21_305 VPWR VGND sg13g2_decap_8
X_1954_ net216 VPWR _0823_ VGND state\[103\] net179 sg13g2_o21ai_1
X_1885_ VPWR VGND _0771_ net82 _0770_ _0239_ _0341_ net37 sg13g2_a221oi_1
X_2481__313 VPWR VGND net312 sg13g2_tiehi
X_2342__420 VPWR VGND net419 sg13g2_tiehi
X_2506_ net454 VGND VPWR _0452_ state\[68\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2437_ net229 VGND VPWR _0383_ daisychain\[127\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2368_ net367 VGND VPWR _0314_ daisychain\[58\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_2299_ VGND VPWR _0881_ _1020_ _0506_ net70 sg13g2_a21oi_1
X_1319_ VPWR _0119_ state\[92\] VGND sg13g2_inv_1
XFILLER_25_622 VPWR VGND sg13g2_decap_8
XFILLER_40_603 VPWR VGND sg13g2_fill_2
XFILLER_12_305 VPWR VGND sg13g2_decap_8
XFILLER_24_165 VPWR VGND sg13g2_decap_8
XANTENNA_50 VPWR VGND daisychain\[2\] sg13g2_antennanp
XANTENNA_61 VPWR VGND daisychain\[126\] sg13g2_antennanp
XFILLER_20_382 VPWR VGND sg13g2_decap_8
XFILLER_4_504 VPWR VGND sg13g2_decap_8
XFILLER_21_32 VPWR VGND sg13g2_decap_8
X_2527__287 VPWR VGND net286 sg13g2_tiehi
XFILLER_47_224 VPWR VGND sg13g2_decap_8
X_2319__466 VPWR VGND net465 sg13g2_tiehi
XFILLER_46_84 VPWR VGND sg13g2_decap_8
XFILLER_43_441 VPWR VGND sg13g2_decap_8
XFILLER_15_165 VPWR VGND sg13g2_decap_8
XFILLER_31_603 VPWR VGND sg13g2_decap_8
XFILLER_30_102 VPWR VGND sg13g2_decap_8
XFILLER_8_821 VPWR VGND sg13g2_fill_1
XFILLER_30_179 VPWR VGND sg13g2_decap_8
XFILLER_11_382 VPWR VGND sg13g2_decap_8
X_1670_ net208 VPWR _0610_ VGND state\[32\] net167 sg13g2_o21ai_1
XFILLER_8_898 VPWR VGND sg13g2_fill_1
XFILLER_7_56 VPWR VGND sg13g2_decap_8
XFILLER_7_364 VPWR VGND sg13g2_decap_8
XFILLER_30_4 VPWR VGND sg13g2_decap_8
X_2222_ _0982_ net123 state\[84\] VPWR VGND sg13g2_nand2_1
X_2153_ VGND VPWR _0662_ _0947_ _0433_ net97 sg13g2_a21oi_1
XFILLER_38_224 VPWR VGND sg13g2_decap_8
X_2084_ _0913_ net120 state\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_34_463 VPWR VGND sg13g2_decap_8
XFILLER_21_102 VPWR VGND sg13g2_decap_8
XFILLER_21_179 VPWR VGND sg13g2_decap_8
X_1937_ VPWR VGND _0810_ net84 _0809_ _0253_ _0354_ net41 sg13g2_a221oi_1
XFILLER_30_691 VPWR VGND sg13g2_decap_8
X_1868_ VGND VPWR net151 daisychain\[80\] _0759_ net60 sg13g2_a21oi_1
X_1799_ net199 _0216_ _0706_ _0707_ VPWR VGND sg13g2_a21o_1
XFILLER_1_518 VPWR VGND sg13g2_decap_8
XFILLER_18_909 VPWR VGND sg13g2_fill_2
XFILLER_29_235 VPWR VGND sg13g2_decap_8
XFILLER_44_238 VPWR VGND sg13g2_decap_8
XFILLER_26_942 VPWR VGND sg13g2_fill_2
XFILLER_16_32 VPWR VGND sg13g2_decap_8
XFILLER_12_102 VPWR VGND sg13g2_decap_8
XFILLER_13_658 VPWR VGND sg13g2_decap_8
XFILLER_12_179 VPWR VGND sg13g2_decap_8
XFILLER_32_53 VPWR VGND sg13g2_decap_8
XFILLER_21_680 VPWR VGND sg13g2_decap_4
XFILLER_4_312 VPWR VGND sg13g2_decap_8
XFILLER_4_389 VPWR VGND sg13g2_decap_8
XFILLER_48_511 VPWR VGND sg13g2_decap_8
XFILLER_0_595 VPWR VGND sg13g2_decap_8
XFILLER_48_544 VPWR VGND sg13g2_fill_1
XFILLER_35_238 VPWR VGND sg13g2_decap_8
XFILLER_16_474 VPWR VGND sg13g2_decap_4
XFILLER_44_794 VPWR VGND sg13g2_fill_2
XFILLER_44_783 VPWR VGND sg13g2_decap_8
XFILLER_32_923 VPWR VGND sg13g2_fill_1
X_2840_ daisychain\[122\] net18 VPWR VGND sg13g2_buf_1
XFILLER_32_945 VPWR VGND sg13g2_fill_1
X_1722_ net219 VPWR _0649_ VGND state\[45\] net185 sg13g2_o21ai_1
X_1653_ VPWR VGND _0597_ net76 _0596_ _0175_ _0283_ net30 sg13g2_a221oi_1
XFILLER_7_161 VPWR VGND sg13g2_decap_8
X_1584_ VGND VPWR net117 daisychain\[9\] _0546_ net28 sg13g2_a21oi_1
XFILLER_4_890 VPWR VGND sg13g2_fill_2
X_2205_ VGND VPWR _0740_ _0973_ _0459_ net106 sg13g2_a21oi_1
X_2136_ _0939_ net138 state\[41\] VPWR VGND sg13g2_nand2_1
X_2067_ VGND VPWR _0533_ _0904_ _0390_ net70 sg13g2_a21oi_1
XFILLER_42_709 VPWR VGND sg13g2_decap_8
XFILLER_26_249 VPWR VGND sg13g2_decap_8
XFILLER_23_978 VPWR VGND sg13g2_decap_8
XFILLER_5_109 VPWR VGND sg13g2_decap_8
XFILLER_1_315 VPWR VGND sg13g2_decap_8
XFILLER_49_319 VPWR VGND sg13g2_decap_8
XFILLER_27_42 VPWR VGND sg13g2_decap_8
XFILLER_17_238 VPWR VGND sg13g2_decap_8
XFILLER_26_794 VPWR VGND sg13g2_decap_4
XFILLER_43_63 VPWR VGND sg13g2_decap_8
XFILLER_40_252 VPWR VGND sg13g2_decap_8
XFILLER_9_459 VPWR VGND sg13g2_decap_8
XFILLER_5_632 VPWR VGND sg13g2_decap_4
XFILLER_4_46 VPWR VGND sg13g2_decap_8
XFILLER_4_186 VPWR VGND sg13g2_decap_8
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_48_385 VPWR VGND sg13g2_decap_8
XFILLER_32_742 VPWR VGND sg13g2_decap_8
XFILLER_32_720 VPWR VGND sg13g2_decap_8
XFILLER_32_753 VPWR VGND sg13g2_decap_8
XFILLER_32_797 VPWR VGND sg13g2_fill_1
XFILLER_31_263 VPWR VGND sg13g2_decap_8
XFILLER_20_948 VPWR VGND sg13g2_decap_8
X_1705_ VPWR VGND _0636_ net103 _0635_ _0190_ _0296_ net58 sg13g2_a221oi_1
XFILLER_8_481 VPWR VGND sg13g2_decap_8
X_1636_ VGND VPWR net148 daisychain\[22\] _0585_ net57 sg13g2_a21oi_1
X_1567_ net166 _0222_ _0532_ _0533_ VPWR VGND sg13g2_a21o_1
X_1498_ VPWR _0191_ daisychain\[41\] VGND sg13g2_inv_1
XFILLER_39_385 VPWR VGND sg13g2_decap_8
X_2119_ VGND VPWR _0611_ _0930_ _0416_ net76 sg13g2_a21oi_1
Xfanout45 net48 net45 VPWR VGND sg13g2_buf_1
Xfanout56 net68 net56 VPWR VGND sg13g2_buf_1
Xfanout34 net36 net34 VPWR VGND sg13g2_buf_1
XFILLER_10_403 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_decap_8
Xfanout67 net68 net67 VPWR VGND sg13g2_buf_1
Xfanout78 net112 net78 VPWR VGND sg13g2_buf_1
Xfanout89 net90 net89 VPWR VGND sg13g2_buf_1
XFILLER_22_263 VPWR VGND sg13g2_decap_8
XFILLER_7_919 VPWR VGND sg13g2_decap_8
XFILLER_13_88 VPWR VGND sg13g2_decap_8
XFILLER_2_613 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_49_116 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_38_63 VPWR VGND sg13g2_decap_8
XFILLER_18_525 VPWR VGND sg13g2_decap_8
XFILLER_46_834 VPWR VGND sg13g2_decap_8
XFILLER_45_322 VPWR VGND sg13g2_decap_8
XFILLER_33_506 VPWR VGND sg13g2_fill_1
XFILLER_45_399 VPWR VGND sg13g2_decap_8
XFILLER_33_539 VPWR VGND sg13g2_fill_1
XFILLER_41_561 VPWR VGND sg13g2_decap_8
XFILLER_13_263 VPWR VGND sg13g2_decap_8
XFILLER_9_256 VPWR VGND sg13g2_decap_8
XFILLER_6_963 VPWR VGND sg13g2_fill_1
XFILLER_6_952 VPWR VGND sg13g2_decap_8
X_2470_ net356 VGND VPWR _0416_ state\[32\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_5_473 VPWR VGND sg13g2_decap_8
X_1421_ VPWR _0148_ daisychain\[118\] VGND sg13g2_inv_1
X_1352_ VPWR _0082_ state\[59\] VGND sg13g2_inv_1
X_1283_ VPWR _0030_ state\[127\] VGND sg13g2_inv_1
XFILLER_49_672 VPWR VGND sg13g2_fill_2
XFILLER_48_182 VPWR VGND sg13g2_decap_8
XFILLER_36_322 VPWR VGND sg13g2_decap_8
XFILLER_36_399 VPWR VGND sg13g2_decap_8
Xclkload9 clkload9/Y clknet_leaf_16_clk VPWR VGND sg13g2_inv_8
X_1619_ net175 _0166_ _0571_ _0572_ VPWR VGND sg13g2_a21o_1
Xfanout213 net216 net213 VPWR VGND sg13g2_buf_1
Xfanout202 net203 net202 VPWR VGND sg13g2_buf_1
Xfanout224 net227 net224 VPWR VGND sg13g2_buf_1
X_2456__413 VPWR VGND net412 sg13g2_tiehi
XFILLER_46_119 VPWR VGND sg13g2_decap_8
XFILLER_39_182 VPWR VGND sg13g2_decap_8
XFILLER_27_322 VPWR VGND sg13g2_decap_8
XFILLER_15_506 VPWR VGND sg13g2_fill_1
X_2352__400 VPWR VGND net399 sg13g2_tiehi
XFILLER_42_336 VPWR VGND sg13g2_decap_8
XFILLER_27_399 VPWR VGND sg13g2_decap_8
XFILLER_24_32 VPWR VGND sg13g2_decap_8
XFILLER_10_200 VPWR VGND sg13g2_decap_8
XFILLER_10_277 VPWR VGND sg13g2_decap_8
XFILLER_40_42 VPWR VGND sg13g2_decap_8
XFILLER_3_900 VPWR VGND sg13g2_fill_1
XFILLER_3_955 VPWR VGND sg13g2_decap_8
XFILLER_2_410 VPWR VGND sg13g2_decap_8
XFILLER_2_487 VPWR VGND sg13g2_decap_8
XFILLER_49_95 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_19_801 VPWR VGND sg13g2_fill_1
XFILLER_18_333 VPWR VGND sg13g2_decap_8
XFILLER_19_867 VPWR VGND sg13g2_fill_2
XFILLER_18_399 VPWR VGND sg13g2_decap_8
XFILLER_45_196 VPWR VGND sg13g2_decap_8
X_1970_ net215 VPWR _0835_ VGND state\[107\] net179 sg13g2_o21ai_1
XFILLER_33_347 VPWR VGND sg13g2_decap_8
X_2329__446 VPWR VGND net445 sg13g2_tiehi
X_2522_ net326 VGND VPWR _0468_ state\[84\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_6_771 VPWR VGND sg13g2_fill_1
XFILLER_5_270 VPWR VGND sg13g2_decap_8
X_2453_ net424 VGND VPWR _0399_ state\[15\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2384_ net335 VGND VPWR _0330_ daisychain\[74\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1404_ VPWR _0105_ state\[7\] VGND sg13g2_inv_1
X_1335_ VPWR _0101_ state\[76\] VGND sg13g2_inv_1
Xinput2 ui_in[0] net2 VPWR VGND sg13g2_buf_1
XFILLER_49_480 VPWR VGND sg13g2_decap_8
XFILLER_37_620 VPWR VGND sg13g2_decap_8
XFILLER_25_826 VPWR VGND sg13g2_fill_1
XFILLER_36_196 VPWR VGND sg13g2_decap_8
XFILLER_25_859 VPWR VGND sg13g2_fill_2
XFILLER_24_347 VPWR VGND sg13g2_decap_8
XFILLER_3_207 VPWR VGND sg13g2_decap_8
XFILLER_10_67 VPWR VGND sg13g2_decap_8
XFILLER_0_958 VPWR VGND sg13g2_decap_8
XFILLER_0_969 VPWR VGND sg13g2_fill_1
XFILLER_48_918 VPWR VGND sg13g2_fill_2
XFILLER_19_32 VPWR VGND sg13g2_decap_8
XFILLER_47_406 VPWR VGND sg13g2_decap_8
XFILLER_28_642 VPWR VGND sg13g2_fill_1
XFILLER_28_631 VPWR VGND sg13g2_decap_8
XFILLER_35_42 VPWR VGND sg13g2_decap_8
XFILLER_15_347 VPWR VGND sg13g2_decap_8
XFILLER_42_133 VPWR VGND sg13g2_decap_8
XFILLER_31_807 VPWR VGND sg13g2_fill_1
XFILLER_27_196 VPWR VGND sg13g2_decap_8
XFILLER_24_881 VPWR VGND sg13g2_fill_2
XFILLER_11_564 VPWR VGND sg13g2_fill_1
XFILLER_7_546 VPWR VGND sg13g2_decap_8
XFILLER_3_752 VPWR VGND sg13g2_decap_8
XFILLER_2_284 VPWR VGND sg13g2_decap_8
XFILLER_38_406 VPWR VGND sg13g2_decap_4
XFILLER_18_130 VPWR VGND sg13g2_decap_8
XFILLER_19_675 VPWR VGND sg13g2_decap_4
XFILLER_46_483 VPWR VGND sg13g2_decap_8
XFILLER_33_144 VPWR VGND sg13g2_decap_8
X_1953_ VPWR VGND _0822_ net104 _0821_ _0131_ _0358_ net61 sg13g2_a221oi_1
X_1884_ VGND VPWR net126 daisychain\[84\] _0771_ net37 sg13g2_a21oi_1
X_2505_ net462 VGND VPWR _0451_ state\[67\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2436_ net231 VGND VPWR _0382_ daisychain\[126\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2367_ net369 VGND VPWR _0313_ daisychain\[57\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_5_1018 VPWR VGND sg13g2_decap_8
X_2298_ _1020_ net114 state\[122\] VPWR VGND sg13g2_nand2_1
X_1318_ VPWR _0120_ state\[93\] VGND sg13g2_inv_1
XFILLER_37_483 VPWR VGND sg13g2_decap_8
XFILLER_25_645 VPWR VGND sg13g2_decap_8
XFILLER_24_144 VPWR VGND sg13g2_decap_8
XFILLER_40_659 VPWR VGND sg13g2_decap_8
XFILLER_40_637 VPWR VGND sg13g2_fill_2
XFILLER_21_840 VPWR VGND sg13g2_decap_8
XANTENNA_40 VPWR VGND daisychain\[104\] sg13g2_antennanp
XANTENNA_51 VPWR VGND daisychain\[37\] sg13g2_antennanp
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_20_361 VPWR VGND sg13g2_decap_8
XFILLER_21_88 VPWR VGND sg13g2_decap_8
XFILLER_0_733 VPWR VGND sg13g2_fill_2
XFILLER_43_1002 VPWR VGND sg13g2_fill_1
XFILLER_47_203 VPWR VGND sg13g2_decap_8
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_15_144 VPWR VGND sg13g2_decap_8
XFILLER_43_420 VPWR VGND sg13g2_decap_8
XFILLER_43_464 VPWR VGND sg13g2_fill_1
XFILLER_31_648 VPWR VGND sg13g2_fill_1
XFILLER_31_637 VPWR VGND sg13g2_decap_8
XFILLER_30_158 VPWR VGND sg13g2_decap_8
XFILLER_11_361 VPWR VGND sg13g2_decap_8
XFILLER_8_855 VPWR VGND sg13g2_fill_1
XFILLER_7_35 VPWR VGND sg13g2_decap_8
XFILLER_8_877 VPWR VGND sg13g2_fill_1
XFILLER_7_343 VPWR VGND sg13g2_decap_8
X_2221_ VGND VPWR _0764_ _0981_ _0467_ net79 sg13g2_a21oi_1
XFILLER_39_704 VPWR VGND sg13g2_decap_8
XFILLER_38_203 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_decap_8
X_2152_ _0947_ net144 state\[49\] VPWR VGND sg13g2_nand2_1
XFILLER_39_737 VPWR VGND sg13g2_fill_2
X_2083_ VGND VPWR _0557_ _0912_ _0398_ net73 sg13g2_a21oi_1
XFILLER_47_770 VPWR VGND sg13g2_fill_1
XFILLER_46_280 VPWR VGND sg13g2_decap_8
XFILLER_34_442 VPWR VGND sg13g2_decap_8
XFILLER_22_626 VPWR VGND sg13g2_fill_1
XFILLER_34_497 VPWR VGND sg13g2_decap_8
XFILLER_21_158 VPWR VGND sg13g2_decap_8
X_1936_ VGND VPWR net128 daisychain\[97\] _0810_ net41 sg13g2_a21oi_1
X_1867_ net197 _0235_ _0757_ _0758_ VPWR VGND sg13g2_a21o_1
X_1798_ net225 VPWR _0706_ VGND state\[64\] net199 sg13g2_o21ai_1
XFILLER_27_1019 VPWR VGND sg13g2_decap_8
X_2419_ net265 VGND VPWR _0365_ daisychain\[109\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_29_214 VPWR VGND sg13g2_decap_8
XFILLER_16_11 VPWR VGND sg13g2_decap_8
XFILLER_45_729 VPWR VGND sg13g2_fill_1
XFILLER_44_217 VPWR VGND sg13g2_decap_8
XFILLER_26_932 VPWR VGND sg13g2_fill_2
XFILLER_26_921 VPWR VGND sg13g2_decap_8
XFILLER_37_280 VPWR VGND sg13g2_decap_8
XFILLER_25_442 VPWR VGND sg13g2_fill_1
XFILLER_25_431 VPWR VGND sg13g2_decap_8
XFILLER_16_88 VPWR VGND sg13g2_decap_8
XFILLER_40_445 VPWR VGND sg13g2_decap_8
XFILLER_12_158 VPWR VGND sg13g2_decap_8
XFILLER_40_456 VPWR VGND sg13g2_fill_2
XFILLER_32_32 VPWR VGND sg13g2_decap_8
XFILLER_4_368 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_decap_8
X_2360__384 VPWR VGND net383 sg13g2_tiehi
XFILLER_35_217 VPWR VGND sg13g2_decap_8
XFILLER_28_291 VPWR VGND sg13g2_decap_8
XFILLER_16_464 VPWR VGND sg13g2_decap_4
XFILLER_43_294 VPWR VGND sg13g2_decap_8
XFILLER_31_445 VPWR VGND sg13g2_decap_8
X_1721_ VPWR VGND _0648_ net94 _0647_ _0194_ _0300_ net50 sg13g2_a221oi_1
XFILLER_8_652 VPWR VGND sg13g2_decap_4
XFILLER_7_140 VPWR VGND sg13g2_decap_8
X_1652_ VGND VPWR net119 daisychain\[26\] _0597_ net30 sg13g2_a21oi_1
X_1583_ net164 _0139_ _0544_ _0545_ VPWR VGND sg13g2_a21o_1
X_2406__292 VPWR VGND net291 sg13g2_tiehi
X_2204_ _0973_ net154 state\[75\] VPWR VGND sg13g2_nand2_1
X_2135_ VGND VPWR _0635_ _0938_ _0424_ net95 sg13g2_a21oi_1
XFILLER_26_228 VPWR VGND sg13g2_decap_8
XFILLER_19_291 VPWR VGND sg13g2_decap_8
X_2066_ _0904_ net114 state\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_22_445 VPWR VGND sg13g2_decap_8
X_1919_ net180 _0249_ _0796_ _0797_ VPWR VGND sg13g2_a21o_1
XFILLER_17_217 VPWR VGND sg13g2_decap_8
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_27_98 VPWR VGND sg13g2_decap_8
XFILLER_13_445 VPWR VGND sg13g2_decap_8
XFILLER_13_456 VPWR VGND sg13g2_fill_1
XFILLER_13_467 VPWR VGND sg13g2_fill_1
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_40_231 VPWR VGND sg13g2_decap_8
XFILLER_9_438 VPWR VGND sg13g2_decap_8
XFILLER_22_990 VPWR VGND sg13g2_fill_1
XFILLER_5_611 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_4_165 VPWR VGND sg13g2_decap_8
XFILLER_49_810 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_49_843 VPWR VGND sg13g2_decap_8
XFILLER_48_364 VPWR VGND sg13g2_decap_8
XFILLER_32_776 VPWR VGND sg13g2_fill_1
XFILLER_31_242 VPWR VGND sg13g2_decap_8
X_1704_ VGND VPWR net149 daisychain\[39\] _0636_ net58 sg13g2_a21oi_1
XFILLER_8_460 VPWR VGND sg13g2_decap_8
X_1635_ net194 _0171_ _0583_ _0584_ VPWR VGND sg13g2_a21o_1
X_1566_ net207 VPWR _0532_ VGND state\[6\] net166 sg13g2_o21ai_1
X_1497_ VPWR _0192_ daisychain\[42\] VGND sg13g2_inv_1
X_2339__426 VPWR VGND net425 sg13g2_tiehi
XFILLER_39_364 VPWR VGND sg13g2_decap_8
X_2118_ _0930_ net119 state\[32\] VPWR VGND sg13g2_nand2_1
X_2049_ VPWR VGND _0894_ net69 _0893_ _0157_ _0382_ net24 sg13g2_a221oi_1
Xfanout35 net40 net35 VPWR VGND sg13g2_buf_1
Xfanout46 net47 net46 VPWR VGND sg13g2_buf_1
Xfanout24 net26 net24 VPWR VGND sg13g2_buf_1
XFILLER_22_242 VPWR VGND sg13g2_decap_8
Xfanout57 net67 net57 VPWR VGND sg13g2_buf_1
Xfanout68 _0515_ net68 VPWR VGND sg13g2_buf_1
Xfanout79 net81 net79 VPWR VGND sg13g2_buf_1
XFILLER_10_459 VPWR VGND sg13g2_decap_8
XFILLER_13_67 VPWR VGND sg13g2_decap_8
XFILLER_2_669 VPWR VGND sg13g2_decap_4
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_38_42 VPWR VGND sg13g2_decap_8
XFILLER_45_301 VPWR VGND sg13g2_decap_8
XFILLER_45_378 VPWR VGND sg13g2_decap_8
XFILLER_14_710 VPWR VGND sg13g2_fill_2
XFILLER_14_732 VPWR VGND sg13g2_decap_8
XFILLER_13_242 VPWR VGND sg13g2_decap_8
XFILLER_9_235 VPWR VGND sg13g2_decap_8
XFILLER_41_595 VPWR VGND sg13g2_decap_8
XFILLER_5_452 VPWR VGND sg13g2_decap_8
X_1420_ VPWR _0149_ daisychain\[119\] VGND sg13g2_inv_1
X_1351_ VPWR _0084_ state\[60\] VGND sg13g2_inv_1
XFILLER_23_1000 VPWR VGND sg13g2_fill_2
XFILLER_48_161 VPWR VGND sg13g2_decap_8
XFILLER_36_301 VPWR VGND sg13g2_decap_8
XFILLER_36_378 VPWR VGND sg13g2_decap_8
XFILLER_17_570 VPWR VGND sg13g2_decap_8
XFILLER_24_529 VPWR VGND sg13g2_fill_2
X_2484__301 VPWR VGND net300 sg13g2_tiehi
XFILLER_20_735 VPWR VGND sg13g2_decap_4
XFILLER_30_1015 VPWR VGND sg13g2_decap_8
XFILLER_20_779 VPWR VGND sg13g2_fill_2
X_1618_ net213 VPWR _0571_ VGND state\[19\] net175 sg13g2_o21ai_1
Xfanout214 net216 net214 VPWR VGND sg13g2_buf_1
Xfanout203 net204 net203 VPWR VGND sg13g2_buf_1
Xfanout225 net227 net225 VPWR VGND sg13g2_buf_1
X_1549_ VPWR VGND _0519_ net80 _0518_ _0167_ _0257_ net34 sg13g2_a221oi_1
XFILLER_39_161 VPWR VGND sg13g2_decap_8
XFILLER_27_301 VPWR VGND sg13g2_decap_8
XFILLER_43_827 VPWR VGND sg13g2_decap_4
XFILLER_27_378 VPWR VGND sg13g2_decap_8
XFILLER_42_315 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_11_724 VPWR VGND sg13g2_decap_8
XFILLER_24_88 VPWR VGND sg13g2_decap_8
XFILLER_10_256 VPWR VGND sg13g2_decap_8
XFILLER_6_249 VPWR VGND sg13g2_decap_8
XFILLER_40_21 VPWR VGND sg13g2_decap_8
XFILLER_40_98 VPWR VGND sg13g2_decap_8
XFILLER_3_923 VPWR VGND sg13g2_fill_1
XFILLER_2_466 VPWR VGND sg13g2_decap_8
XFILLER_49_74 VPWR VGND sg13g2_decap_8
XFILLER_19_824 VPWR VGND sg13g2_fill_2
XFILLER_18_312 VPWR VGND sg13g2_decap_8
XFILLER_46_654 VPWR VGND sg13g2_fill_2
XFILLER_45_175 VPWR VGND sg13g2_decap_8
XFILLER_33_326 VPWR VGND sg13g2_decap_8
XFILLER_41_392 VPWR VGND sg13g2_decap_8
X_2521_ net334 VGND VPWR _0467_ state\[83\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2452_ net428 VGND VPWR _0398_ state\[14\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2383_ net337 VGND VPWR _0329_ daisychain\[73\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1403_ VPWR _0116_ state\[8\] VGND sg13g2_inv_1
X_1334_ VPWR _0102_ state\[77\] VGND sg13g2_inv_1
XFILLER_28_109 VPWR VGND sg13g2_decap_8
Xinput3 ui_in[1] net3 VPWR VGND sg13g2_buf_1
XFILLER_37_643 VPWR VGND sg13g2_decap_8
XFILLER_36_175 VPWR VGND sg13g2_decap_8
XFILLER_24_326 VPWR VGND sg13g2_decap_8
XFILLER_10_46 VPWR VGND sg13g2_decap_8
XFILLER_0_926 VPWR VGND sg13g2_decap_4
XFILLER_19_11 VPWR VGND sg13g2_decap_8
XFILLER_19_109 VPWR VGND sg13g2_decap_8
XFILLER_19_88 VPWR VGND sg13g2_decap_8
XFILLER_15_326 VPWR VGND sg13g2_decap_8
XFILLER_43_624 VPWR VGND sg13g2_decap_8
XFILLER_42_112 VPWR VGND sg13g2_decap_8
XFILLER_35_21 VPWR VGND sg13g2_decap_8
XFILLER_27_175 VPWR VGND sg13g2_decap_8
XFILLER_43_668 VPWR VGND sg13g2_decap_4
XFILLER_35_98 VPWR VGND sg13g2_decap_8
XFILLER_42_189 VPWR VGND sg13g2_decap_8
XFILLER_24_893 VPWR VGND sg13g2_fill_2
XFILLER_11_543 VPWR VGND sg13g2_decap_8
XFILLER_11_554 VPWR VGND sg13g2_fill_1
XFILLER_7_525 VPWR VGND sg13g2_decap_8
XFILLER_3_720 VPWR VGND sg13g2_decap_8
XFILLER_2_263 VPWR VGND sg13g2_decap_8
XFILLER_18_186 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_8
XFILLER_34_602 VPWR VGND sg13g2_decap_4
XFILLER_33_123 VPWR VGND sg13g2_decap_8
X_2370__364 VPWR VGND net363 sg13g2_tiehi
XFILLER_22_819 VPWR VGND sg13g2_fill_1
X_1952_ VGND VPWR net150 daisychain\[101\] _0822_ net61 sg13g2_a21oi_1
X_1883_ net173 _0239_ _0769_ _0770_ VPWR VGND sg13g2_a21o_1
X_2504_ net470 VGND VPWR _0450_ state\[66\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_44_0 VPWR VGND sg13g2_decap_8
X_2435_ net233 VGND VPWR _0381_ daisychain\[125\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2366_ net371 VGND VPWR _0312_ daisychain\[56\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2297_ VGND VPWR _0878_ _1019_ _0505_ net69 sg13g2_a21oi_1
X_1317_ VPWR _0121_ state\[94\] VGND sg13g2_inv_1
XFILLER_37_462 VPWR VGND sg13g2_decap_8
XFILLER_24_123 VPWR VGND sg13g2_decap_8
X_2416__272 VPWR VGND net271 sg13g2_tiehi
XFILLER_40_616 VPWR VGND sg13g2_fill_2
XANTENNA_30 VPWR VGND _0200_ sg13g2_antennanp
XANTENNA_41 VPWR VGND daisychain\[114\] sg13g2_antennanp
XFILLER_20_340 VPWR VGND sg13g2_decap_8
XANTENNA_52 VPWR VGND daisychain\[41\] sg13g2_antennanp
XFILLER_21_885 VPWR VGND sg13g2_decap_8
XFILLER_4_539 VPWR VGND sg13g2_decap_8
XFILLER_21_67 VPWR VGND sg13g2_decap_8
XFILLER_43_1025 VPWR VGND sg13g2_decap_4
XFILLER_29_941 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_15_123 VPWR VGND sg13g2_decap_8
XFILLER_16_646 VPWR VGND sg13g2_fill_1
XFILLER_43_476 VPWR VGND sg13g2_decap_8
XFILLER_43_498 VPWR VGND sg13g2_decap_8
XFILLER_30_137 VPWR VGND sg13g2_decap_8
XFILLER_11_340 VPWR VGND sg13g2_decap_8
XFILLER_8_812 VPWR VGND sg13g2_fill_1
XFILLER_8_801 VPWR VGND sg13g2_fill_1
XFILLER_8_834 VPWR VGND sg13g2_fill_1
XFILLER_7_322 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_8_889 VPWR VGND sg13g2_fill_2
XFILLER_7_399 VPWR VGND sg13g2_decap_8
X_2220_ _0981_ net123 state\[83\] VPWR VGND sg13g2_nand2_1
XFILLER_3_594 VPWR VGND sg13g2_decap_8
XFILLER_16_4 VPWR VGND sg13g2_decap_8
X_2151_ VGND VPWR _0659_ _0946_ _0432_ net99 sg13g2_a21oi_1
X_2082_ _0912_ net116 state\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_38_259 VPWR VGND sg13g2_decap_8
XFILLER_34_410 VPWR VGND sg13g2_decap_8
XFILLER_34_476 VPWR VGND sg13g2_decap_8
X_1935_ net176 _0253_ _0808_ _0809_ VPWR VGND sg13g2_a21o_1
XFILLER_21_137 VPWR VGND sg13g2_decap_8
XFILLER_30_671 VPWR VGND sg13g2_decap_4
X_1866_ net224 VPWR _0757_ VGND state\[81\] net197 sg13g2_o21ai_1
X_1797_ VPWR VGND _0705_ net107 _0704_ _0215_ _0319_ net63 sg13g2_a221oi_1
X_2418_ net267 VGND VPWR _0364_ daisychain\[108\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2349_ net405 VGND VPWR _0295_ daisychain\[39\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_26_944 VPWR VGND sg13g2_fill_1
XFILLER_25_410 VPWR VGND sg13g2_decap_8
XFILLER_16_67 VPWR VGND sg13g2_decap_8
XFILLER_13_638 VPWR VGND sg13g2_decap_8
XFILLER_13_649 VPWR VGND sg13g2_decap_4
XFILLER_40_413 VPWR VGND sg13g2_fill_2
XFILLER_12_137 VPWR VGND sg13g2_decap_8
XFILLER_32_11 VPWR VGND sg13g2_decap_8
X_2349__406 VPWR VGND net405 sg13g2_tiehi
XFILLER_32_88 VPWR VGND sg13g2_decap_8
XFILLER_21_693 VPWR VGND sg13g2_decap_8
XFILLER_4_347 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_48_535 VPWR VGND sg13g2_decap_8
XFILLER_29_771 VPWR VGND sg13g2_decap_8
XFILLER_16_410 VPWR VGND sg13g2_decap_8
XFILLER_44_741 VPWR VGND sg13g2_decap_8
XFILLER_28_270 VPWR VGND sg13g2_decap_8
XFILLER_43_273 VPWR VGND sg13g2_decap_8
XFILLER_31_468 VPWR VGND sg13g2_decap_8
XFILLER_12_671 VPWR VGND sg13g2_fill_1
XFILLER_8_631 VPWR VGND sg13g2_decap_8
X_1720_ VGND VPWR net141 daisychain\[43\] _0648_ net50 sg13g2_a21oi_1
X_1651_ net167 _0175_ _0595_ _0596_ VPWR VGND sg13g2_a21o_1
XdacH daisychain\[64\] _0216_ daisychain\[65\] _0217_ daisychain\[66\] _0218_ daisychain\[67\]
+ _0219_ daisychain\[68\] _0220_ daisychain\[69\] _0221_ daisychain\[70\] _0223_ daisychain\[71\]
+ _0224_ daisychain\[72\] _0225_ digitalenH.g\[2\].u.OUTP digitalenH.g\[2\].u.OUTN
+ daisychain\[73\] _0226_ daisychain\[74\] _0227_ daisychain\[75\] _0228_ daisychain\[76\]
+ _0229_ daisychain\[77\] _0230_ daisychain\[78\] _0231_ daisychain\[79\] _0232_ daisychain\[80\]
+ _0234_ daisychain\[81\] _0235_ daisychain\[82\] _0236_ daisychain\[83\] _0237_ daisychain\[84\]
+ _0238_ daisychain\[85\] _0239_ daisychain\[86\] _0240_ daisychain\[87\] _0241_ daisychain\[88\]
+ _0242_ daisychain\[89\] _0243_ daisychain\[90\] _0245_ daisychain\[91\] _0246_ daisychain\[92\]
+ _0247_ daisychain\[93\] _0248_ daisychain\[94\] _0249_ daisychain\[95\] _0250_ daisychain\[96\]
+ _0251_ daisychain\[97\] _0252_ daisychain\[98\] _0253_ daisychain\[99\] _0254_ daisychain\[100\]
+ _0129_ daisychain\[101\] _0130_ daisychain\[102\] _0131_ daisychain\[103\] _0132_
+ daisychain\[104\] _0133_ daisychain\[105\] _0134_ daisychain\[106\] _0135_ daisychain\[107\]
+ _0136_ daisychain\[108\] _0137_ daisychain\[109\] _0138_ daisychain\[110\] _0140_
+ daisychain\[111\] _0141_ daisychain\[112\] _0142_ daisychain\[113\] _0143_ daisychain\[114\]
+ _0144_ daisychain\[115\] _0145_ daisychain\[116\] _0146_ daisychain\[117\] _0147_
+ daisychain\[118\] _0148_ daisychain\[119\] _0149_ daisychain\[120\] _0151_ daisychain\[121\]
+ _0152_ daisychain\[122\] _0153_ digitalenH.g\[3\].u.OUTP digitalenH.g\[3\].u.OUTN
+ daisychain\[123\] _0154_ daisychain\[124\] _0155_ daisychain\[125\] _0156_ daisychain\[126\]
+ _0157_ daisychain\[127\] _0158_ daisychain\[0\] _0128_ daisychain\[1\] _0167_ daisychain\[2\]
+ _0178_ daisychain\[3\] _0189_ daisychain\[4\] _0200_ daisychain\[5\] _0211_ daisychain\[6\]
+ digitalenH.g\[0\].u.OUTP digitalenH.g\[0\].u.OUTN _0222_ daisychain\[7\] _0233_
+ daisychain\[8\] _0244_ daisychain\[9\] _0255_ daisychain\[10\] _0139_ daisychain\[11\]
+ _0150_ daisychain\[12\] _0159_ daisychain\[13\] _0160_ daisychain\[14\] _0161_ daisychain\[15\]
+ _0162_ daisychain\[16\] _0163_ daisychain\[17\] _0164_ daisychain\[18\] _0165_ daisychain\[19\]
+ _0166_ daisychain\[20\] _0168_ daisychain\[21\] _0169_ daisychain\[22\] _0170_ daisychain\[23\]
+ _0171_ daisychain\[24\] _0172_ daisychain\[25\] _0173_ daisychain\[26\] _0174_ daisychain\[27\]
+ _0175_ daisychain\[28\] _0176_ daisychain\[29\] _0177_ daisychain\[30\] _0179_ daisychain\[31\]
+ _0180_ daisychain\[33\] _0182_ daisychain\[32\] _0181_ daisychain\[34\] _0183_ daisychain\[35\]
+ _0184_ daisychain\[36\] _0185_ daisychain\[37\] _0186_ daisychain\[38\] _0187_ daisychain\[39\]
+ _0188_ daisychain\[40\] _0190_ daisychain\[41\] _0191_ daisychain\[42\] _0192_ daisychain\[43\]
+ _0193_ daisychain\[44\] _0194_ daisychain\[45\] _0195_ daisychain\[46\] _0196_ daisychain\[47\]
+ _0197_ daisychain\[48\] _0198_ daisychain\[49\] _0199_ daisychain\[50\] _0201_ daisychain\[51\]
+ _0202_ daisychain\[52\] _0203_ daisychain\[53\] _0204_ daisychain\[54\] _0205_ daisychain\[55\]
+ _0206_ daisychain\[56\] _0207_ daisychain\[57\] _0208_ daisychain\[58\] _0209_ daisychain\[59\]
+ _0210_ daisychain\[60\] _0212_ daisychain\[61\] _0213_ daisychain\[62\] _0214_ daisychain\[63\]
+ _0215_ digitalenH.g\[1\].u.OUTP digitalenH.g\[1\].u.OUTN VGND VPWR dac128module
XFILLER_7_196 VPWR VGND sg13g2_decap_8
X_1582_ net206 VPWR _0544_ VGND state\[10\] net164 sg13g2_o21ai_1
X_2203_ VGND VPWR _0737_ _0972_ _0458_ net106 sg13g2_a21oi_1
XFILLER_39_524 VPWR VGND sg13g2_fill_1
X_2134_ _0938_ net141 state\[40\] VPWR VGND sg13g2_nand2_1
XFILLER_26_207 VPWR VGND sg13g2_decap_8
XFILLER_19_270 VPWR VGND sg13g2_decap_8
X_2065_ VGND VPWR _0530_ _0903_ _0389_ net77 sg13g2_a21oi_1
XFILLER_47_590 VPWR VGND sg13g2_decap_8
XFILLER_23_925 VPWR VGND sg13g2_decap_8
XFILLER_23_903 VPWR VGND sg13g2_fill_2
XFILLER_34_284 VPWR VGND sg13g2_decap_8
XFILLER_23_947 VPWR VGND sg13g2_decap_8
XFILLER_22_424 VPWR VGND sg13g2_decap_8
XFILLER_10_619 VPWR VGND sg13g2_decap_8
XFILLER_31_991 VPWR VGND sg13g2_decap_8
X_1918_ net215 VPWR _0796_ VGND state\[94\] net180 sg13g2_o21ai_1
X_1849_ VPWR VGND _0744_ net106 _0743_ _0229_ _0332_ net62 sg13g2_a221oi_1
XFILLER_2_829 VPWR VGND sg13g2_decap_8
X_2459__401 VPWR VGND net400 sg13g2_tiehi
XFILLER_45_538 VPWR VGND sg13g2_decap_8
XFILLER_27_77 VPWR VGND sg13g2_decap_8
XFILLER_13_424 VPWR VGND sg13g2_decap_8
XFILLER_43_21 VPWR VGND sg13g2_decap_8
XFILLER_41_733 VPWR VGND sg13g2_fill_2
XFILLER_40_210 VPWR VGND sg13g2_decap_8
XFILLER_25_284 VPWR VGND sg13g2_decap_8
XFILLER_9_417 VPWR VGND sg13g2_decap_8
XFILLER_13_479 VPWR VGND sg13g2_decap_8
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_40_287 VPWR VGND sg13g2_decap_8
XFILLER_4_144 VPWR VGND sg13g2_decap_8
XFILLER_49_1020 VPWR VGND sg13g2_decap_8
XFILLER_1_840 VPWR VGND sg13g2_fill_2
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_48_343 VPWR VGND sg13g2_decap_8
XFILLER_49_888 VPWR VGND sg13g2_decap_8
XFILLER_16_284 VPWR VGND sg13g2_decap_8
XFILLER_44_593 VPWR VGND sg13g2_decap_8
XFILLER_31_221 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_11_clk clknet_2_3__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
XFILLER_31_298 VPWR VGND sg13g2_decap_8
X_1703_ net195 _0190_ _0634_ _0635_ VPWR VGND sg13g2_a21o_1
X_1634_ net223 VPWR _0583_ VGND state\[23\] net194 sg13g2_o21ai_1
XdigitalenH.g\[3\].u.inv1 VPWR digitalenH.g\[3\].u.OUTN net7 VGND sg13g2_inv_1
X_1565_ VPWR VGND _0531_ net75 _0530_ _0211_ _0261_ net29 sg13g2_a221oi_1
X_1496_ VPWR _0193_ daisychain\[43\] VGND sg13g2_inv_1
XFILLER_39_343 VPWR VGND sg13g2_decap_8
X_2117_ VGND VPWR _0608_ _0929_ _0415_ net73 sg13g2_a21oi_1
X_2048_ VGND VPWR net113 daisychain\[125\] _0894_ net24 sg13g2_a21oi_1
XFILLER_35_560 VPWR VGND sg13g2_fill_2
XFILLER_23_711 VPWR VGND sg13g2_fill_2
Xfanout36 net40 net36 VPWR VGND sg13g2_buf_1
Xfanout47 net48 net47 VPWR VGND sg13g2_buf_1
Xfanout25 net26 net25 VPWR VGND sg13g2_buf_1
X_2530__263 VPWR VGND net262 sg13g2_tiehi
XFILLER_22_221 VPWR VGND sg13g2_decap_8
Xfanout58 net67 net58 VPWR VGND sg13g2_buf_1
Xfanout69 net72 net69 VPWR VGND sg13g2_buf_1
XFILLER_23_777 VPWR VGND sg13g2_decap_8
XFILLER_10_438 VPWR VGND sg13g2_decap_8
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_22_298 VPWR VGND sg13g2_decap_8
XFILLER_2_648 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_38_21 VPWR VGND sg13g2_decap_8
XFILLER_38_98 VPWR VGND sg13g2_decap_8
XFILLER_45_357 VPWR VGND sg13g2_decap_8
XFILLER_13_221 VPWR VGND sg13g2_decap_8
XFILLER_9_214 VPWR VGND sg13g2_decap_8
XFILLER_13_298 VPWR VGND sg13g2_decap_8
XFILLER_6_932 VPWR VGND sg13g2_decap_4
XFILLER_5_431 VPWR VGND sg13g2_decap_8
XFILLER_6_998 VPWR VGND sg13g2_fill_1
XFILLER_6_987 VPWR VGND sg13g2_fill_2
XFILLER_48_7 VPWR VGND sg13g2_decap_8
X_1350_ VPWR _0085_ state\[61\] VGND sg13g2_inv_1
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_49_674 VPWR VGND sg13g2_fill_1
XFILLER_49_663 VPWR VGND sg13g2_decap_4
XFILLER_48_140 VPWR VGND sg13g2_decap_8
XFILLER_36_357 VPWR VGND sg13g2_decap_8
XFILLER_32_585 VPWR VGND sg13g2_fill_2
XFILLER_20_747 VPWR VGND sg13g2_decap_4
XFILLER_8_291 VPWR VGND sg13g2_decap_8
X_1617_ VPWR VGND _0570_ net85 _0569_ _0165_ _0274_ net42 sg13g2_a221oi_1
X_2380__344 VPWR VGND net343 sg13g2_tiehi
Xfanout204 net5 net204 VPWR VGND sg13g2_buf_1
XFILLER_8_1006 VPWR VGND sg13g2_fill_2
Xfanout226 net227 net226 VPWR VGND sg13g2_buf_1
Xfanout215 net216 net215 VPWR VGND sg13g2_buf_1
X_1548_ VGND VPWR net124 daisychain\[0\] _0519_ net34 sg13g2_a21oi_1
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
X_1479_ VPWR _0212_ daisychain\[60\] VGND sg13g2_inv_1
XFILLER_39_140 VPWR VGND sg13g2_decap_8
XFILLER_28_825 VPWR VGND sg13g2_fill_2
XFILLER_27_357 VPWR VGND sg13g2_decap_8
XFILLER_24_67 VPWR VGND sg13g2_decap_8
XFILLER_10_235 VPWR VGND sg13g2_decap_8
XFILLER_7_729 VPWR VGND sg13g2_fill_1
XFILLER_7_718 VPWR VGND sg13g2_fill_2
XFILLER_6_228 VPWR VGND sg13g2_decap_8
XFILLER_40_77 VPWR VGND sg13g2_decap_8
X_2426__252 VPWR VGND net251 sg13g2_tiehi
XFILLER_2_445 VPWR VGND sg13g2_decap_8
XFILLER_49_53 VPWR VGND sg13g2_decap_8
XFILLER_46_622 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_19_858 VPWR VGND sg13g2_fill_2
XFILLER_18_368 VPWR VGND sg13g2_decap_8
XFILLER_45_154 VPWR VGND sg13g2_decap_8
XFILLER_18_379 VPWR VGND sg13g2_fill_2
XFILLER_33_305 VPWR VGND sg13g2_decap_8
XFILLER_14_574 VPWR VGND sg13g2_decap_4
XFILLER_41_371 VPWR VGND sg13g2_decap_8
X_2520_ net342 VGND VPWR _0466_ state\[82\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_6_762 VPWR VGND sg13g2_decap_8
X_2451_ net432 VGND VPWR _0397_ state\[13\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1402_ VPWR _0127_ state\[9\] VGND sg13g2_inv_1
X_2382_ net339 VGND VPWR _0328_ daisychain\[72\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1333_ VPWR _0103_ state\[78\] VGND sg13g2_inv_1
XFILLER_37_600 VPWR VGND sg13g2_fill_1
Xinput4 ui_in[2] net4 VPWR VGND sg13g2_buf_1
Xclkbuf_2_1__f_clk clknet_2_1__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_37_699 VPWR VGND sg13g2_fill_1
XFILLER_36_154 VPWR VGND sg13g2_decap_8
XFILLER_24_305 VPWR VGND sg13g2_decap_8
XFILLER_32_382 VPWR VGND sg13g2_decap_8
XFILLER_20_511 VPWR VGND sg13g2_fill_1
XFILLER_10_25 VPWR VGND sg13g2_decap_8
XFILLER_28_611 VPWR VGND sg13g2_fill_1
XFILLER_19_67 VPWR VGND sg13g2_decap_8
XFILLER_28_666 VPWR VGND sg13g2_fill_1
XFILLER_15_305 VPWR VGND sg13g2_decap_8
XFILLER_27_154 VPWR VGND sg13g2_decap_8
XFILLER_42_168 VPWR VGND sg13g2_decap_8
XFILLER_35_77 VPWR VGND sg13g2_decap_8
XFILLER_30_319 VPWR VGND sg13g2_decap_8
XFILLER_24_883 VPWR VGND sg13g2_fill_1
XFILLER_11_522 VPWR VGND sg13g2_decap_8
XFILLER_23_382 VPWR VGND sg13g2_decap_8
XFILLER_7_504 VPWR VGND sg13g2_decap_8
XFILLER_3_798 VPWR VGND sg13g2_fill_1
XFILLER_2_242 VPWR VGND sg13g2_decap_8
XFILLER_19_622 VPWR VGND sg13g2_fill_2
XFILLER_46_441 VPWR VGND sg13g2_decap_8
XFILLER_20_1026 VPWR VGND sg13g2_fill_2
XFILLER_18_165 VPWR VGND sg13g2_decap_8
XFILLER_34_625 VPWR VGND sg13g2_fill_1
XFILLER_33_102 VPWR VGND sg13g2_decap_8
XFILLER_34_669 VPWR VGND sg13g2_decap_8
XFILLER_34_647 VPWR VGND sg13g2_decap_4
XFILLER_33_179 VPWR VGND sg13g2_decap_8
XFILLER_21_319 VPWR VGND sg13g2_decap_8
XFILLER_14_382 VPWR VGND sg13g2_decap_8
X_1951_ net196 _0131_ _0820_ _0821_ VPWR VGND sg13g2_a21o_1
X_1882_ net212 VPWR _0769_ VGND state\[85\] net173 sg13g2_o21ai_1
X_2503_ net478 VGND VPWR _0449_ state\[65\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_6_592 VPWR VGND sg13g2_decap_8
X_2434_ net235 VGND VPWR _0380_ daisychain\[124\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2365_ net373 VGND VPWR _0311_ daisychain\[55\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
X_1316_ VPWR _0122_ state\[95\] VGND sg13g2_inv_1
X_2296_ _1019_ net113 state\[121\] VPWR VGND sg13g2_nand2_1
XFILLER_37_441 VPWR VGND sg13g2_decap_8
XFILLER_2_81 VPWR VGND sg13g2_decap_8
XFILLER_24_102 VPWR VGND sg13g2_decap_8
XFILLER_12_319 VPWR VGND sg13g2_decap_8
XFILLER_40_639 VPWR VGND sg13g2_fill_1
XFILLER_24_179 VPWR VGND sg13g2_decap_8
XFILLER_21_831 VPWR VGND sg13g2_fill_1
XANTENNA_20 VPWR VGND _0129_ sg13g2_antennanp
XANTENNA_31 VPWR VGND _0200_ sg13g2_antennanp
XANTENNA_42 VPWR VGND daisychain\[11\] sg13g2_antennanp
XANTENNA_53 VPWR VGND daisychain\[41\] sg13g2_antennanp
XFILLER_21_897 VPWR VGND sg13g2_fill_2
XFILLER_21_46 VPWR VGND sg13g2_decap_8
XFILLER_20_396 VPWR VGND sg13g2_decap_8
XFILLER_4_518 VPWR VGND sg13g2_decap_8
XFILLER_0_713 VPWR VGND sg13g2_fill_2
XFILLER_0_724 VPWR VGND sg13g2_fill_1
XFILLER_0_768 VPWR VGND sg13g2_decap_8
XFILLER_47_238 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_15_102 VPWR VGND sg13g2_decap_8
XFILLER_46_98 VPWR VGND sg13g2_decap_8
XFILLER_28_496 VPWR VGND sg13g2_decap_8
XFILLER_16_669 VPWR VGND sg13g2_decap_8
XFILLER_43_455 VPWR VGND sg13g2_decap_8
XFILLER_15_179 VPWR VGND sg13g2_decap_8
XFILLER_30_116 VPWR VGND sg13g2_decap_8
XFILLER_8_846 VPWR VGND sg13g2_fill_2
XFILLER_7_301 VPWR VGND sg13g2_decap_8
XFILLER_11_396 VPWR VGND sg13g2_decap_8
XFILLER_8_868 VPWR VGND sg13g2_fill_1
XFILLER_7_378 VPWR VGND sg13g2_decap_8
XFILLER_3_573 VPWR VGND sg13g2_decap_8
X_2150_ _0946_ net145 state\[48\] VPWR VGND sg13g2_nand2_1
X_2081_ VGND VPWR _0554_ _0911_ _0397_ net92 sg13g2_a21oi_1
XFILLER_38_238 VPWR VGND sg13g2_decap_8
XFILLER_47_761 VPWR VGND sg13g2_fill_1
XFILLER_19_452 VPWR VGND sg13g2_decap_8
XFILLER_21_116 VPWR VGND sg13g2_decap_8
X_1934_ net213 VPWR _0808_ VGND state\[98\] net175 sg13g2_o21ai_1
X_1865_ VPWR VGND _0756_ net104 _0755_ _0234_ _0336_ net59 sg13g2_a221oi_1
X_1796_ VGND VPWR net153 daisychain\[62\] _0705_ net63 sg13g2_a21oi_1
X_2417_ net269 VGND VPWR _0363_ daisychain\[107\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2348_ net407 VGND VPWR _0294_ daisychain\[38\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2279_ VGND VPWR _0851_ _1010_ _0496_ net80 sg13g2_a21oi_1
XFILLER_29_249 VPWR VGND sg13g2_decap_8
XFILLER_26_956 VPWR VGND sg13g2_decap_8
XFILLER_16_46 VPWR VGND sg13g2_decap_8
XFILLER_12_116 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_decap_8
XFILLER_40_469 VPWR VGND sg13g2_decap_8
XFILLER_21_650 VPWR VGND sg13g2_fill_2
XFILLER_32_67 VPWR VGND sg13g2_decap_8
XFILLER_20_193 VPWR VGND sg13g2_decap_8
XFILLER_4_326 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_48_525 VPWR VGND sg13g2_decap_4
XFILLER_29_761 VPWR VGND sg13g2_decap_4
XFILLER_43_252 VPWR VGND sg13g2_decap_8
XFILLER_32_915 VPWR VGND sg13g2_decap_4
XFILLER_31_403 VPWR VGND sg13g2_decap_8
XFILLER_11_193 VPWR VGND sg13g2_decap_8
X_1650_ net208 VPWR _0595_ VGND state\[27\] net167 sg13g2_o21ai_1
XFILLER_7_175 VPWR VGND sg13g2_decap_8
X_1581_ VPWR VGND _0543_ net74 _0542_ _0255_ _0265_ net28 sg13g2_a221oi_1
X_2202_ _0972_ net154 state\[74\] VPWR VGND sg13g2_nand2_1
XFILLER_39_503 VPWR VGND sg13g2_decap_8
X_2133_ VGND VPWR _0632_ _0937_ _0423_ net103 sg13g2_a21oi_1
XFILLER_39_558 VPWR VGND sg13g2_decap_8
XFILLER_39_547 VPWR VGND sg13g2_fill_1
X_2064_ _0903_ net121 state\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_34_263 VPWR VGND sg13g2_decap_8
XFILLER_22_403 VPWR VGND sg13g2_decap_8
X_1917_ VPWR VGND _0795_ net104 _0794_ _0248_ _0349_ net59 sg13g2_a221oi_1
X_1848_ VGND VPWR net154 daisychain\[75\] _0744_ net64 sg13g2_a21oi_1
X_1779_ net189 _0210_ _0691_ _0692_ VPWR VGND sg13g2_a21o_1
XFILLER_1_329 VPWR VGND sg13g2_decap_8
XFILLER_45_517 VPWR VGND sg13g2_decap_8
X_2390__324 VPWR VGND net323 sg13g2_tiehi
XFILLER_27_56 VPWR VGND sg13g2_decap_8
XFILLER_13_403 VPWR VGND sg13g2_decap_8
XFILLER_25_263 VPWR VGND sg13g2_decap_8
XFILLER_43_77 VPWR VGND sg13g2_decap_8
XFILLER_40_266 VPWR VGND sg13g2_decap_8
XFILLER_22_981 VPWR VGND sg13g2_decap_8
X_2507__447 VPWR VGND net446 sg13g2_tiehi
XFILLER_4_123 VPWR VGND sg13g2_decap_8
XFILLER_5_668 VPWR VGND sg13g2_decap_8
XFILLER_48_322 VPWR VGND sg13g2_decap_8
X_2436__232 VPWR VGND net231 sg13g2_tiehi
XFILLER_48_399 VPWR VGND sg13g2_decap_8
XFILLER_16_263 VPWR VGND sg13g2_decap_8
XFILLER_32_712 VPWR VGND sg13g2_decap_4
XFILLER_31_200 VPWR VGND sg13g2_decap_8
XFILLER_32_767 VPWR VGND sg13g2_decap_4
XFILLER_20_907 VPWR VGND sg13g2_fill_1
XFILLER_32_789 VPWR VGND sg13g2_decap_4
XFILLER_31_277 VPWR VGND sg13g2_decap_8
X_1702_ net220 VPWR _0634_ VGND state\[40\] net187 sg13g2_o21ai_1
X_1633_ VPWR VGND _0582_ net102 _0581_ _0170_ _0278_ net57 sg13g2_a221oi_1
XFILLER_8_495 VPWR VGND sg13g2_decap_8
XdigitalenH.g\[3\].u.inv2 VPWR digitalenH.g\[3\].u.OUTP digitalenH.g\[3\].u.OUTN VGND
+ sg13g2_inv_1
X_1564_ VGND VPWR net128 daisychain\[4\] _0531_ net41 sg13g2_a21oi_1
X_1495_ VPWR _0194_ daisychain\[44\] VGND sg13g2_inv_1
XFILLER_4_690 VPWR VGND sg13g2_decap_8
XFILLER_39_322 VPWR VGND sg13g2_decap_8
XFILLER_27_506 VPWR VGND sg13g2_decap_4
X_2116_ _0929_ net122 state\[31\] VPWR VGND sg13g2_nand2_1
XFILLER_39_399 VPWR VGND sg13g2_decap_8
XFILLER_27_539 VPWR VGND sg13g2_fill_2
X_2047_ net159 _0157_ _0892_ _0893_ VPWR VGND sg13g2_a21o_1
XFILLER_22_200 VPWR VGND sg13g2_decap_8
Xfanout37 net39 net37 VPWR VGND sg13g2_buf_1
Xfanout26 net33 net26 VPWR VGND sg13g2_buf_1
XFILLER_10_417 VPWR VGND sg13g2_decap_8
Xfanout48 net68 net48 VPWR VGND sg13g2_buf_1
Xfanout59 net61 net59 VPWR VGND sg13g2_buf_1
XFILLER_22_277 VPWR VGND sg13g2_decap_8
XFILLER_13_25 VPWR VGND sg13g2_decap_8
XFILLER_2_627 VPWR VGND sg13g2_decap_8
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_38_77 VPWR VGND sg13g2_decap_8
XFILLER_18_539 VPWR VGND sg13g2_fill_1
XFILLER_46_859 VPWR VGND sg13g2_decap_8
XFILLER_45_336 VPWR VGND sg13g2_decap_8
XFILLER_13_200 VPWR VGND sg13g2_decap_8
XFILLER_13_277 VPWR VGND sg13g2_decap_8
XFILLER_6_900 VPWR VGND sg13g2_decap_8
XFILLER_5_410 VPWR VGND sg13g2_decap_8
XFILLER_5_487 VPWR VGND sg13g2_decap_8
XFILLER_49_642 VPWR VGND sg13g2_fill_2
XFILLER_1_693 VPWR VGND sg13g2_fill_2
XFILLER_49_686 VPWR VGND sg13g2_decap_8
XFILLER_36_336 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_17_550 VPWR VGND sg13g2_decap_8
XFILLER_8_270 VPWR VGND sg13g2_decap_8
X_1616_ VGND VPWR net129 daisychain\[17\] _0570_ net42 sg13g2_a21oi_1
Xfanout205 net210 net205 VPWR VGND sg13g2_buf_1
XFILLER_5_81 VPWR VGND sg13g2_decap_8
Xfanout227 net228 net227 VPWR VGND sg13g2_buf_1
Xfanout216 net217 net216 VPWR VGND sg13g2_buf_1
X_1547_ net170 _0167_ _0517_ _0518_ VPWR VGND sg13g2_a21o_1
X_1478_ VPWR _0213_ daisychain\[61\] VGND sg13g2_inv_1
XFILLER_39_196 VPWR VGND sg13g2_decap_8
XFILLER_27_336 VPWR VGND sg13g2_decap_8
XFILLER_24_46 VPWR VGND sg13g2_decap_8
XFILLER_10_214 VPWR VGND sg13g2_decap_8
XFILLER_6_207 VPWR VGND sg13g2_decap_8
XFILLER_40_56 VPWR VGND sg13g2_decap_8
XFILLER_3_914 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_3_969 VPWR VGND sg13g2_decap_4
XFILLER_2_424 VPWR VGND sg13g2_decap_8
XFILLER_49_32 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_19_826 VPWR VGND sg13g2_fill_1
XFILLER_18_347 VPWR VGND sg13g2_decap_8
XFILLER_46_667 VPWR VGND sg13g2_decap_8
XFILLER_46_656 VPWR VGND sg13g2_fill_1
XFILLER_45_133 VPWR VGND sg13g2_decap_8
XFILLER_42_862 VPWR VGND sg13g2_decap_8
XFILLER_42_851 VPWR VGND sg13g2_decap_4
XFILLER_41_350 VPWR VGND sg13g2_decap_8
X_2450_ net436 VGND VPWR _0396_ state\[12\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_1401_ VPWR _0011_ state\[10\] VGND sg13g2_inv_1
XFILLER_5_284 VPWR VGND sg13g2_decap_8
X_2381_ net341 VGND VPWR _0327_ daisychain\[71\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2559__451 VPWR VGND net450 sg13g2_tiehi
X_1332_ VPWR _0104_ state\[79\] VGND sg13g2_inv_1
XFILLER_1_490 VPWR VGND sg13g2_decap_8
Xinput5 ui_in[3] net5 VPWR VGND sg13g2_buf_1
XFILLER_49_494 VPWR VGND sg13g2_decap_8
XFILLER_36_133 VPWR VGND sg13g2_decap_8
XFILLER_37_689 VPWR VGND sg13g2_fill_1
XFILLER_37_678 VPWR VGND sg13g2_fill_2
XFILLER_32_361 VPWR VGND sg13g2_decap_8
XFILLER_20_578 VPWR VGND sg13g2_decap_8
XFILLER_19_46 VPWR VGND sg13g2_decap_8
XFILLER_27_133 VPWR VGND sg13g2_decap_8
XFILLER_35_56 VPWR VGND sg13g2_decap_8
XFILLER_42_147 VPWR VGND sg13g2_decap_8
XFILLER_11_501 VPWR VGND sg13g2_decap_8
XFILLER_24_895 VPWR VGND sg13g2_fill_1
XFILLER_23_361 VPWR VGND sg13g2_decap_8
XFILLER_2_221 VPWR VGND sg13g2_decap_8
XFILLER_3_777 VPWR VGND sg13g2_fill_2
XFILLER_2_298 VPWR VGND sg13g2_decap_8
XFILLER_47_932 VPWR VGND sg13g2_fill_2
XFILLER_46_420 VPWR VGND sg13g2_decap_8
XFILLER_18_144 VPWR VGND sg13g2_decap_8
XFILLER_47_998 VPWR VGND sg13g2_fill_2
XFILLER_33_158 VPWR VGND sg13g2_decap_8
XFILLER_14_361 VPWR VGND sg13g2_decap_8
X_1950_ net224 VPWR _0820_ VGND state\[102\] net196 sg13g2_o21ai_1
X_1881_ VPWR VGND _0768_ net79 _0767_ _0238_ _0340_ net35 sg13g2_a221oi_1
X_2502_ net VGND VPWR _0448_ state\[64\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_6_571 VPWR VGND sg13g2_decap_8
X_2433_ net237 VGND VPWR _0379_ daisychain\[123\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2364_ net375 VGND VPWR _0310_ daisychain\[54\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1315_ VPWR _0123_ state\[96\] VGND sg13g2_inv_1
X_2295_ VGND VPWR _0875_ _1018_ _0504_ net83 sg13g2_a21oi_1
XFILLER_2_60 VPWR VGND sg13g2_decap_8
XFILLER_49_291 VPWR VGND sg13g2_decap_8
XFILLER_37_420 VPWR VGND sg13g2_fill_2
XFILLER_25_659 VPWR VGND sg13g2_decap_8
XFILLER_40_618 VPWR VGND sg13g2_fill_1
XFILLER_24_158 VPWR VGND sg13g2_decap_8
XFILLER_40_629 VPWR VGND sg13g2_decap_4
XFILLER_21_821 VPWR VGND sg13g2_fill_2
XANTENNA_10 VPWR VGND _0163_ sg13g2_antennanp
XANTENNA_21 VPWR VGND _0133_ sg13g2_antennanp
XANTENNA_32 VPWR VGND _0233_ sg13g2_antennanp
XANTENNA_43 VPWR VGND daisychain\[11\] sg13g2_antennanp
XANTENNA_54 VPWR VGND daisychain\[42\] sg13g2_antennanp
XFILLER_20_375 VPWR VGND sg13g2_decap_8
XFILLER_21_25 VPWR VGND sg13g2_decap_8
XFILLER_47_217 VPWR VGND sg13g2_decap_8
XFILLER_29_921 VPWR VGND sg13g2_fill_2
XFILLER_29_910 VPWR VGND sg13g2_decap_8
XFILLER_28_442 VPWR VGND sg13g2_decap_8
XFILLER_46_77 VPWR VGND sg13g2_decap_8
XFILLER_29_976 VPWR VGND sg13g2_fill_2
XFILLER_28_453 VPWR VGND sg13g2_fill_2
XFILLER_43_434 VPWR VGND sg13g2_decap_8
XFILLER_15_158 VPWR VGND sg13g2_decap_8
XFILLER_11_375 VPWR VGND sg13g2_decap_8
XFILLER_8_825 VPWR VGND sg13g2_fill_1
XFILLER_7_49 VPWR VGND sg13g2_decap_8
XFILLER_7_357 VPWR VGND sg13g2_decap_8
XFILLER_3_552 VPWR VGND sg13g2_decap_8
XFILLER_39_718 VPWR VGND sg13g2_fill_2
XFILLER_38_217 VPWR VGND sg13g2_decap_8
X_2080_ _0911_ net138 state\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_19_431 VPWR VGND sg13g2_fill_2
XFILLER_19_420 VPWR VGND sg13g2_decap_8
XFILLER_46_294 VPWR VGND sg13g2_decap_8
XFILLER_34_456 VPWR VGND sg13g2_decap_8
XFILLER_15_692 VPWR VGND sg13g2_decap_8
X_1933_ VPWR VGND _0807_ net84 _0806_ _0252_ _0353_ net41 sg13g2_a221oi_1
X_1864_ VGND VPWR net150 daisychain\[79\] _0756_ net59 sg13g2_a21oi_1
X_1795_ net193 _0215_ _0703_ _0704_ VPWR VGND sg13g2_a21o_1
XFILLER_7_891 VPWR VGND sg13g2_decap_8
X_2416_ net271 VGND VPWR _0362_ daisychain\[106\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2347_ net409 VGND VPWR _0293_ daisychain\[37\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2278_ _1010_ net124 state\[112\] VPWR VGND sg13g2_nand2_1
XFILLER_29_228 VPWR VGND sg13g2_decap_8
XFILLER_16_25 VPWR VGND sg13g2_decap_8
XFILLER_37_294 VPWR VGND sg13g2_decap_8
XFILLER_32_46 VPWR VGND sg13g2_decap_8
XFILLER_21_673 VPWR VGND sg13g2_decap_8
XFILLER_21_684 VPWR VGND sg13g2_fill_2
XFILLER_20_172 VPWR VGND sg13g2_decap_8
XFILLER_5_828 VPWR VGND sg13g2_decap_4
XFILLER_4_305 VPWR VGND sg13g2_decap_8
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_decap_8
XFILLER_48_504 VPWR VGND sg13g2_decap_8
XFILLER_29_751 VPWR VGND sg13g2_decap_4
XFILLER_43_231 VPWR VGND sg13g2_decap_8
XFILLER_16_478 VPWR VGND sg13g2_fill_2
XFILLER_32_949 VPWR VGND sg13g2_fill_1
XFILLER_31_459 VPWR VGND sg13g2_decap_4
XFILLER_11_172 VPWR VGND sg13g2_decap_8
XFILLER_8_688 VPWR VGND sg13g2_fill_1
XFILLER_7_154 VPWR VGND sg13g2_decap_8
X_1580_ VGND VPWR net117 daisychain\[8\] _0543_ net28 sg13g2_a21oi_1
XFILLER_4_883 VPWR VGND sg13g2_decap_8
XFILLER_3_382 VPWR VGND sg13g2_decap_8
XFILLER_26_1022 VPWR VGND sg13g2_decap_8
X_2201_ VGND VPWR _0734_ _0971_ _0457_ net109 sg13g2_a21oi_1
XFILLER_21_4 VPWR VGND sg13g2_decap_8
X_2132_ _0937_ net149 state\[39\] VPWR VGND sg13g2_nand2_1
X_2063_ VGND VPWR _0527_ _0902_ _0388_ net77 sg13g2_a21oi_1
XFILLER_34_242 VPWR VGND sg13g2_decap_8
XFILLER_23_905 VPWR VGND sg13g2_fill_1
X_1916_ VGND VPWR net150 daisychain\[92\] _0795_ net59 sg13g2_a21oi_1
X_1847_ net199 _0229_ _0742_ _0743_ VPWR VGND sg13g2_a21o_1
XFILLER_8_81 VPWR VGND sg13g2_decap_8
X_1778_ net221 VPWR _0691_ VGND state\[59\] net189 sg13g2_o21ai_1
XFILLER_1_308 VPWR VGND sg13g2_decap_8
XFILLER_27_35 VPWR VGND sg13g2_decap_8
XFILLER_25_242 VPWR VGND sg13g2_decap_8
XFILLER_26_798 VPWR VGND sg13g2_fill_1
XFILLER_26_787 VPWR VGND sg13g2_decap_8
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_41_735 VPWR VGND sg13g2_fill_1
XFILLER_40_245 VPWR VGND sg13g2_decap_8
XFILLER_5_636 VPWR VGND sg13g2_fill_1
XFILLER_5_625 VPWR VGND sg13g2_decap_8
XFILLER_4_102 VPWR VGND sg13g2_decap_8
XFILLER_4_39 VPWR VGND sg13g2_decap_8
XFILLER_4_179 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_49_857 VPWR VGND sg13g2_fill_2
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_36_507 VPWR VGND sg13g2_decap_8
XFILLER_17_732 VPWR VGND sg13g2_decap_4
XFILLER_16_242 VPWR VGND sg13g2_decap_8
XFILLER_31_256 VPWR VGND sg13g2_decap_8
X_1701_ VPWR VGND _0633_ net103 _0632_ _0188_ _0295_ net58 sg13g2_a221oi_1
X_1632_ VGND VPWR net148 daisychain\[21\] _0582_ net57 sg13g2_a21oi_1
XFILLER_8_474 VPWR VGND sg13g2_decap_8
X_1563_ net166 _0211_ _0529_ _0530_ VPWR VGND sg13g2_a21o_1
X_1494_ VPWR _0195_ daisychain\[45\] VGND sg13g2_inv_1
XFILLER_39_301 VPWR VGND sg13g2_decap_8
X_2115_ VGND VPWR _0605_ _0928_ _0414_ net77 sg13g2_a21oi_1
XFILLER_39_378 VPWR VGND sg13g2_decap_8
X_2046_ net205 VPWR _0892_ VGND state\[126\] net159 sg13g2_o21ai_1
XFILLER_35_562 VPWR VGND sg13g2_fill_1
Xfanout38 net40 net38 VPWR VGND sg13g2_buf_1
Xfanout27 net28 net27 VPWR VGND sg13g2_buf_1
XFILLER_23_746 VPWR VGND sg13g2_fill_2
Xfanout49 net51 net49 VPWR VGND sg13g2_buf_1
XFILLER_22_256 VPWR VGND sg13g2_decap_8
XFILLER_2_606 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_49_109 VPWR VGND sg13g2_decap_8
XFILLER_38_56 VPWR VGND sg13g2_decap_8
XFILLER_18_518 VPWR VGND sg13g2_decap_8
XFILLER_46_827 VPWR VGND sg13g2_decap_8
XFILLER_45_315 VPWR VGND sg13g2_decap_8
XFILLER_13_256 VPWR VGND sg13g2_decap_8
XFILLER_9_249 VPWR VGND sg13g2_decap_8
XFILLER_5_466 VPWR VGND sg13g2_decap_8
X_2403__298 VPWR VGND net297 sg13g2_tiehi
XFILLER_1_672 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_36_315 VPWR VGND sg13g2_decap_8
XFILLER_44_392 VPWR VGND sg13g2_decap_8
XFILLER_32_587 VPWR VGND sg13g2_fill_1
X_1615_ net177 _0165_ _0568_ _0569_ VPWR VGND sg13g2_a21o_1
X_1546_ net211 VPWR _0517_ VGND state\[1\] net170 sg13g2_o21ai_1
XFILLER_5_60 VPWR VGND sg13g2_decap_8
Xfanout228 net4 net228 VPWR VGND sg13g2_buf_1
Xfanout217 net228 net217 VPWR VGND sg13g2_buf_1
Xfanout206 net209 net206 VPWR VGND sg13g2_buf_1
X_1477_ VPWR _0214_ daisychain\[62\] VGND sg13g2_inv_1
XFILLER_39_175 VPWR VGND sg13g2_decap_8
XFILLER_28_827 VPWR VGND sg13g2_fill_1
XFILLER_27_315 VPWR VGND sg13g2_decap_8
X_2029_ VPWR VGND _0879_ net69 _0878_ _0152_ _0377_ net24 sg13g2_a221oi_1
XFILLER_42_329 VPWR VGND sg13g2_decap_8
XFILLER_35_392 VPWR VGND sg13g2_decap_8
XFILLER_23_532 VPWR VGND sg13g2_fill_1
XFILLER_23_521 VPWR VGND sg13g2_fill_2
XFILLER_24_25 VPWR VGND sg13g2_decap_8
XFILLER_11_738 VPWR VGND sg13g2_fill_1
XFILLER_40_35 VPWR VGND sg13g2_decap_8
XFILLER_2_403 VPWR VGND sg13g2_decap_8
XFILLER_49_11 VPWR VGND sg13g2_decap_8
XFILLER_49_88 VPWR VGND sg13g2_decap_8
XFILLER_18_326 VPWR VGND sg13g2_decap_8
XFILLER_45_112 VPWR VGND sg13g2_decap_8
XFILLER_45_189 VPWR VGND sg13g2_decap_8
XFILLER_6_797 VPWR VGND sg13g2_decap_8
XFILLER_5_263 VPWR VGND sg13g2_decap_8
X_1400_ VPWR _0022_ state\[11\] VGND sg13g2_inv_1
X_2380_ net343 VGND VPWR _0326_ daisychain\[70\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1331_ VPWR _0106_ state\[80\] VGND sg13g2_inv_1
XFILLER_2_981 VPWR VGND sg13g2_decap_8
Xinput6 ui_in[4] net6 VPWR VGND sg13g2_buf_1
XFILLER_49_473 VPWR VGND sg13g2_decap_8
XFILLER_37_613 VPWR VGND sg13g2_decap_8
XFILLER_36_112 VPWR VGND sg13g2_decap_8
XFILLER_25_819 VPWR VGND sg13g2_decap_8
XFILLER_36_189 VPWR VGND sg13g2_decap_8
XFILLER_17_392 VPWR VGND sg13g2_decap_8
XFILLER_32_340 VPWR VGND sg13g2_decap_8
X_1529_ VPWR _0139_ daisychain\[10\] VGND sg13g2_inv_1
XFILLER_19_25 VPWR VGND sg13g2_decap_8
XFILLER_28_624 VPWR VGND sg13g2_decap_8
XFILLER_27_112 VPWR VGND sg13g2_decap_8
X_2356__392 VPWR VGND net391 sg13g2_tiehi
XFILLER_43_638 VPWR VGND sg13g2_fill_2
XFILLER_42_126 VPWR VGND sg13g2_decap_8
XFILLER_35_35 VPWR VGND sg13g2_decap_8
XFILLER_27_189 VPWR VGND sg13g2_decap_8
XFILLER_23_340 VPWR VGND sg13g2_decap_8
XFILLER_7_539 VPWR VGND sg13g2_decap_8
XFILLER_3_734 VPWR VGND sg13g2_decap_4
XFILLER_2_200 VPWR VGND sg13g2_decap_8
XFILLER_2_277 VPWR VGND sg13g2_decap_8
XFILLER_18_123 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
X_2554__371 VPWR VGND net370 sg13g2_tiehi
XFILLER_46_476 VPWR VGND sg13g2_decap_8
XFILLER_19_668 VPWR VGND sg13g2_decap_8
X_2550__235 VPWR VGND net234 sg13g2_tiehi
XFILLER_14_340 VPWR VGND sg13g2_decap_8
XFILLER_33_137 VPWR VGND sg13g2_decap_8
X_1880_ VGND VPWR net123 daisychain\[83\] _0768_ net35 sg13g2_a21oi_1
XFILLER_42_693 VPWR VGND sg13g2_fill_2
X_2501_ net232 VGND VPWR _0447_ state\[63\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_6_550 VPWR VGND sg13g2_decap_8
X_2432_ net239 VGND VPWR _0378_ daisychain\[122\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_2363_ net377 VGND VPWR _0309_ daisychain\[53\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1314_ VPWR _0124_ state\[97\] VGND sg13g2_inv_1
X_2294_ _1018_ net127 state\[120\] VPWR VGND sg13g2_nand2_1
XFILLER_49_270 VPWR VGND sg13g2_decap_8
XFILLER_37_476 VPWR VGND sg13g2_decap_8
XFILLER_24_137 VPWR VGND sg13g2_decap_8
XANTENNA_11 VPWR VGND _0175_ sg13g2_antennanp
XANTENNA_22 VPWR VGND _0136_ sg13g2_antennanp
XFILLER_21_866 VPWR VGND sg13g2_decap_4
XFILLER_21_855 VPWR VGND sg13g2_fill_2
XANTENNA_33 VPWR VGND _0234_ sg13g2_antennanp
XANTENNA_44 VPWR VGND daisychain\[11\] sg13g2_antennanp
XANTENNA_55 VPWR VGND daisychain\[79\] sg13g2_antennanp
XFILLER_20_354 VPWR VGND sg13g2_decap_8
XFILLER_48_719 VPWR VGND sg13g2_decap_4
XFILLER_28_410 VPWR VGND sg13g2_decap_8
XFILLER_46_56 VPWR VGND sg13g2_decap_8
XFILLER_28_476 VPWR VGND sg13g2_decap_8
XFILLER_44_936 VPWR VGND sg13g2_decap_4
XFILLER_43_413 VPWR VGND sg13g2_decap_8
XFILLER_15_137 VPWR VGND sg13g2_decap_8
XFILLER_24_660 VPWR VGND sg13g2_fill_2
XFILLER_11_354 VPWR VGND sg13g2_decap_8
X_2545__315 VPWR VGND net314 sg13g2_tiehi
XFILLER_7_28 VPWR VGND sg13g2_decap_8
XFILLER_8_859 VPWR VGND sg13g2_fill_2
XFILLER_7_336 VPWR VGND sg13g2_decap_8
XFILLER_11_81 VPWR VGND sg13g2_decap_8
XFILLER_3_531 VPWR VGND sg13g2_decap_8
XFILLER_19_410 VPWR VGND sg13g2_decap_4
XFILLER_47_752 VPWR VGND sg13g2_decap_8
XFILLER_46_273 VPWR VGND sg13g2_decap_8
XFILLER_34_424 VPWR VGND sg13g2_decap_4
XFILLER_22_619 VPWR VGND sg13g2_decap_8
X_1932_ VGND VPWR net128 daisychain\[96\] _0807_ net41 sg13g2_a21oi_1
XFILLER_30_641 VPWR VGND sg13g2_fill_1
X_1863_ net194 _0234_ _0754_ _0755_ VPWR VGND sg13g2_a21o_1
X_1794_ net222 VPWR _0703_ VGND state\[63\] net192 sg13g2_o21ai_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
X_2415_ net273 VGND VPWR _0361_ daisychain\[105\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2346_ net411 VGND VPWR _0292_ daisychain\[36\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_29_207 VPWR VGND sg13g2_decap_8
X_2277_ VGND VPWR _0848_ _1009_ _0495_ net80 sg13g2_a21oi_1
XFILLER_37_273 VPWR VGND sg13g2_decap_8
XFILLER_25_424 VPWR VGND sg13g2_decap_8
XFILLER_40_427 VPWR VGND sg13g2_fill_2
XFILLER_40_438 VPWR VGND sg13g2_decap_8
XFILLER_32_25 VPWR VGND sg13g2_decap_8
XFILLER_21_652 VPWR VGND sg13g2_fill_1
XFILLER_20_151 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_16_424 VPWR VGND sg13g2_decap_8
XFILLER_44_711 VPWR VGND sg13g2_fill_1
XFILLER_43_210 VPWR VGND sg13g2_decap_8
XFILLER_29_785 VPWR VGND sg13g2_decap_4
XFILLER_28_284 VPWR VGND sg13g2_decap_8
XFILLER_16_435 VPWR VGND sg13g2_fill_2
XFILLER_16_457 VPWR VGND sg13g2_decap_8
XFILLER_16_468 VPWR VGND sg13g2_fill_1
XFILLER_43_287 VPWR VGND sg13g2_decap_8
XFILLER_31_427 VPWR VGND sg13g2_fill_2
XFILLER_11_151 VPWR VGND sg13g2_decap_8
XFILLER_8_645 VPWR VGND sg13g2_decap_8
XFILLER_7_133 VPWR VGND sg13g2_decap_8
XFILLER_3_361 VPWR VGND sg13g2_decap_8
X_2200_ _0971_ net156 state\[73\] VPWR VGND sg13g2_nand2_1
XFILLER_14_4 VPWR VGND sg13g2_decap_8
X_2131_ VGND VPWR _0629_ _0936_ _0422_ net92 sg13g2_a21oi_1
X_2062_ _0902_ net118 state\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_19_284 VPWR VGND sg13g2_decap_8
XFILLER_35_733 VPWR VGND sg13g2_fill_2
XFILLER_34_221 VPWR VGND sg13g2_decap_8
XFILLER_34_298 VPWR VGND sg13g2_decap_8
XFILLER_22_438 VPWR VGND sg13g2_decap_8
X_1915_ net196 _0248_ _0793_ _0794_ VPWR VGND sg13g2_a21o_1
X_2413__278 VPWR VGND net277 sg13g2_tiehi
Xclkbuf_leaf_14_clk clknet_2_2__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
XFILLER_8_60 VPWR VGND sg13g2_decap_8
XFILLER_30_471 VPWR VGND sg13g2_decap_4
X_1846_ net225 VPWR _0742_ VGND state\[76\] net199 sg13g2_o21ai_1
X_1777_ VPWR VGND _0690_ net97 _0689_ _0209_ _0314_ net56 sg13g2_a221oi_1
X_2329_ net445 VGND VPWR _0275_ daisychain\[19\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_26_766 VPWR VGND sg13g2_decap_4
XFILLER_25_221 VPWR VGND sg13g2_decap_8
XFILLER_13_438 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
XFILLER_40_224 VPWR VGND sg13g2_decap_8
XFILLER_25_298 VPWR VGND sg13g2_decap_8
XFILLER_21_482 VPWR VGND sg13g2_fill_2
XFILLER_5_604 VPWR VGND sg13g2_decap_8
XFILLER_4_158 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_1_810 VPWR VGND sg13g2_fill_2
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_49_803 VPWR VGND sg13g2_decap_8
XFILLER_49_836 VPWR VGND sg13g2_decap_8
XFILLER_1_898 VPWR VGND sg13g2_decap_4
X_2553__403 VPWR VGND net402 sg13g2_tiehi
XFILLER_48_357 VPWR VGND sg13g2_decap_8
XFILLER_16_221 VPWR VGND sg13g2_decap_8
XFILLER_17_91 VPWR VGND sg13g2_decap_8
XFILLER_16_298 VPWR VGND sg13g2_decap_8
XFILLER_31_235 VPWR VGND sg13g2_decap_8
XFILLER_8_431 VPWR VGND sg13g2_decap_8
XFILLER_12_493 VPWR VGND sg13g2_decap_8
X_1700_ VGND VPWR net149 daisychain\[38\] _0633_ net58 sg13g2_a21oi_1
XFILLER_8_453 VPWR VGND sg13g2_decap_8
X_1631_ net194 _0170_ _0580_ _0581_ VPWR VGND sg13g2_a21o_1
X_1562_ net207 VPWR _0529_ VGND state\[5\] net165 sg13g2_o21ai_1
X_1493_ VPWR _0196_ daisychain\[46\] VGND sg13g2_inv_1
Xclkbuf_leaf_3_clk clknet_2_1__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_2114_ _0928_ net120 state\[30\] VPWR VGND sg13g2_nand2_1
XFILLER_39_357 VPWR VGND sg13g2_decap_8
X_2045_ VPWR VGND _0891_ net69 _0890_ _0156_ _0381_ net24 sg13g2_a221oi_1
XFILLER_35_530 VPWR VGND sg13g2_decap_4
Xfanout28 net33 net28 VPWR VGND sg13g2_buf_1
X_2315__474 VPWR VGND net473 sg13g2_tiehi
Xfanout39 net40 net39 VPWR VGND sg13g2_buf_1
XFILLER_22_235 VPWR VGND sg13g2_decap_8
X_1829_ VPWR VGND _0729_ net105 _0728_ _0224_ _0327_ net60 sg13g2_a221oi_1
XFILLER_38_35 VPWR VGND sg13g2_decap_8
XFILLER_46_806 VPWR VGND sg13g2_fill_1
XFILLER_14_703 VPWR VGND sg13g2_fill_2
XFILLER_14_725 VPWR VGND sg13g2_decap_8
XFILLER_13_235 VPWR VGND sg13g2_decap_8
XFILLER_9_228 VPWR VGND sg13g2_decap_8
X_2366__372 VPWR VGND net371 sg13g2_tiehi
XFILLER_5_445 VPWR VGND sg13g2_decap_8
XFILLER_1_651 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_1_695 VPWR VGND sg13g2_fill_1
XFILLER_49_644 VPWR VGND sg13g2_fill_1
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_45_850 VPWR VGND sg13g2_fill_2
XFILLER_17_596 VPWR VGND sg13g2_decap_4
XFILLER_44_371 VPWR VGND sg13g2_decap_8
XFILLER_32_555 VPWR VGND sg13g2_fill_2
XFILLER_20_739 VPWR VGND sg13g2_fill_1
X_1614_ net213 VPWR _0568_ VGND state\[18\] net177 sg13g2_o21ai_1
X_1545_ VPWR VGND _0514_ net79 _0516_ _0128_ _0256_ net35 sg13g2_a221oi_1
Xfanout218 net220 net218 VPWR VGND sg13g2_buf_1
Xfanout207 net209 net207 VPWR VGND sg13g2_buf_1
X_1476_ VPWR _0215_ daisychain\[63\] VGND sg13g2_inv_1
XFILLER_39_154 VPWR VGND sg13g2_decap_8
X_2028_ VGND VPWR net113 daisychain\[120\] _0879_ net24 sg13g2_a21oi_1
XFILLER_42_308 VPWR VGND sg13g2_decap_8
XFILLER_35_371 VPWR VGND sg13g2_decap_8
XFILLER_23_500 VPWR VGND sg13g2_fill_2
XFILLER_10_249 VPWR VGND sg13g2_decap_8
XFILLER_40_14 VPWR VGND sg13g2_decap_8
XFILLER_2_459 VPWR VGND sg13g2_decap_8
XFILLER_49_67 VPWR VGND sg13g2_decap_8
XFILLER_18_305 VPWR VGND sg13g2_decap_8
XFILLER_19_817 VPWR VGND sg13g2_decap_8
XFILLER_46_636 VPWR VGND sg13g2_fill_2
XFILLER_45_168 VPWR VGND sg13g2_decap_8
XFILLER_33_319 VPWR VGND sg13g2_decap_8
XFILLER_26_382 VPWR VGND sg13g2_decap_8
XFILLER_14_566 VPWR VGND sg13g2_decap_4
XFILLER_41_385 VPWR VGND sg13g2_decap_8
XFILLER_14_81 VPWR VGND sg13g2_decap_8
XFILLER_5_242 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
X_1330_ VPWR _0107_ state\[81\] VGND sg13g2_inv_1
XFILLER_2_960 VPWR VGND sg13g2_fill_1
Xinput7 ui_in[5] net7 VPWR VGND sg13g2_buf_1
X_2555__339 VPWR VGND net338 sg13g2_tiehi
XFILLER_49_452 VPWR VGND sg13g2_decap_8
XFILLER_36_168 VPWR VGND sg13g2_decap_8
XFILLER_17_371 VPWR VGND sg13g2_decap_8
XFILLER_24_319 VPWR VGND sg13g2_decap_8
XFILLER_32_396 VPWR VGND sg13g2_decap_8
XFILLER_10_39 VPWR VGND sg13g2_decap_8
XFILLER_0_919 VPWR VGND sg13g2_decap_8
X_1528_ VPWR _0150_ daisychain\[11\] VGND sg13g2_inv_1
X_1459_ VPWR _0234_ daisychain\[80\] VGND sg13g2_inv_1
XFILLER_43_617 VPWR VGND sg13g2_decap_8
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_27_168 VPWR VGND sg13g2_decap_8
XFILLER_15_319 VPWR VGND sg13g2_decap_8
XFILLER_42_105 VPWR VGND sg13g2_decap_8
X_2510__423 VPWR VGND net422 sg13g2_tiehi
XFILLER_11_536 VPWR VGND sg13g2_decap_8
XFILLER_23_396 VPWR VGND sg13g2_decap_8
XFILLER_7_518 VPWR VGND sg13g2_decap_8
XFILLER_3_713 VPWR VGND sg13g2_decap_8
XFILLER_2_256 VPWR VGND sg13g2_decap_8
XFILLER_47_901 VPWR VGND sg13g2_decap_8
XFILLER_18_102 VPWR VGND sg13g2_decap_8
XFILLER_19_658 VPWR VGND sg13g2_fill_1
XFILLER_19_647 VPWR VGND sg13g2_decap_4
XFILLER_46_455 VPWR VGND sg13g2_decap_8
XFILLER_34_606 VPWR VGND sg13g2_fill_1
XFILLER_18_179 VPWR VGND sg13g2_decap_8
XFILLER_33_116 VPWR VGND sg13g2_decap_8
XFILLER_42_661 VPWR VGND sg13g2_decap_4
XFILLER_14_396 VPWR VGND sg13g2_decap_8
XFILLER_41_182 VPWR VGND sg13g2_decap_8
X_2500_ net236 VGND VPWR _0446_ state\[62\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_2431_ net241 VGND VPWR _0377_ daisychain\[121\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_2522__327 VPWR VGND net326 sg13g2_tiehi
X_2362_ net379 VGND VPWR _0308_ daisychain\[52\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2293_ VGND VPWR _0872_ _1017_ _0503_ net82 sg13g2_a21oi_1
X_1313_ VPWR _0125_ state\[98\] VGND sg13g2_inv_1
XFILLER_37_422 VPWR VGND sg13g2_fill_1
XFILLER_2_95 VPWR VGND sg13g2_decap_8
XFILLER_37_455 VPWR VGND sg13g2_decap_8
XFILLER_24_116 VPWR VGND sg13g2_decap_8
XFILLER_18_691 VPWR VGND sg13g2_fill_1
XANTENNA_12 VPWR VGND _0249_ sg13g2_antennanp
XANTENNA_23 VPWR VGND _0138_ sg13g2_antennanp
XFILLER_32_193 VPWR VGND sg13g2_decap_8
XFILLER_20_333 VPWR VGND sg13g2_decap_8
XANTENNA_34 VPWR VGND _0243_ sg13g2_antennanp
XANTENNA_45 VPWR VGND daisychain\[126\] sg13g2_antennanp
XANTENNA_56 VPWR VGND daisychain\[88\] sg13g2_antennanp
X_2423__258 VPWR VGND net257 sg13g2_tiehi
XFILLER_43_1018 VPWR VGND sg13g2_decap_8
XFILLER_29_934 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_29_978 VPWR VGND sg13g2_fill_1
XFILLER_15_116 VPWR VGND sg13g2_decap_8
XFILLER_16_639 VPWR VGND sg13g2_decap_8
XFILLER_43_469 VPWR VGND sg13g2_decap_8
XFILLER_8_805 VPWR VGND sg13g2_fill_1
XFILLER_11_333 VPWR VGND sg13g2_decap_8
XFILLER_8_838 VPWR VGND sg13g2_fill_1
XFILLER_8_816 VPWR VGND sg13g2_fill_2
XFILLER_7_315 VPWR VGND sg13g2_decap_8
XFILLER_23_193 VPWR VGND sg13g2_decap_8
XFILLER_11_60 VPWR VGND sg13g2_decap_8
XFILLER_3_510 VPWR VGND sg13g2_decap_8
XFILLER_3_587 VPWR VGND sg13g2_decap_8
XFILLER_47_742 VPWR VGND sg13g2_decap_8
XFILLER_19_466 VPWR VGND sg13g2_fill_2
XFILLER_46_252 VPWR VGND sg13g2_decap_8
XFILLER_34_403 VPWR VGND sg13g2_decap_8
XFILLER_19_499 VPWR VGND sg13g2_decap_4
XFILLER_15_661 VPWR VGND sg13g2_decap_8
X_1931_ net175 _0252_ _0805_ _0806_ VPWR VGND sg13g2_a21o_1
XFILLER_14_193 VPWR VGND sg13g2_decap_8
X_1862_ net223 VPWR _0754_ VGND state\[80\] net194 sg13g2_o21ai_1
XFILLER_30_664 VPWR VGND sg13g2_decap_8
XFILLER_30_675 VPWR VGND sg13g2_fill_1
X_1793_ VPWR VGND _0702_ net100 _0701_ _0214_ _0318_ net54 sg13g2_a221oi_1
X_2414_ net275 VGND VPWR _0360_ daisychain\[104\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_35_0 VPWR VGND sg13g2_decap_8
X_2345_ net413 VGND VPWR _0291_ daisychain\[35\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2276_ _1009_ net124 state\[111\] VPWR VGND sg13g2_nand2_1
XFILLER_37_252 VPWR VGND sg13g2_decap_8
XFILLER_25_403 VPWR VGND sg13g2_decap_8
XFILLER_40_406 VPWR VGND sg13g2_decap_8
XFILLER_21_664 VPWR VGND sg13g2_fill_1
XFILLER_20_130 VPWR VGND sg13g2_decap_8
X_2325__454 VPWR VGND net453 sg13g2_tiehi
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_16_403 VPWR VGND sg13g2_decap_8
XFILLER_28_263 VPWR VGND sg13g2_decap_8
XFILLER_43_266 VPWR VGND sg13g2_decap_8
XFILLER_31_417 VPWR VGND sg13g2_fill_2
XFILLER_11_130 VPWR VGND sg13g2_decap_8
XFILLER_12_697 VPWR VGND sg13g2_decap_4
XFILLER_8_624 VPWR VGND sg13g2_decap_8
XFILLER_7_112 VPWR VGND sg13g2_decap_8
XdacL state\[64\] _0088_ state\[65\] _0089_ state\[66\] _0090_ state\[67\] _0091_
+ state\[68\] _0092_ state\[69\] _0093_ state\[70\] _0095_ state\[71\] _0096_ state\[72\]
+ _0097_ digitalenL.g\[2\].u.OUTP digitalenL.g\[2\].u.OUTN state\[73\] _0098_ state\[74\]
+ _0099_ state\[75\] _0100_ state\[76\] _0101_ state\[77\] _0102_ state\[78\] _0103_
+ state\[79\] _0104_ state\[80\] _0106_ state\[81\] _0107_ state\[82\] _0108_ state\[83\]
+ _0109_ state\[84\] _0110_ state\[85\] _0111_ state\[86\] _0112_ state\[87\] _0113_
+ state\[88\] _0114_ state\[89\] _0115_ state\[90\] _0117_ state\[91\] _0118_ state\[92\]
+ _0119_ state\[93\] _0120_ state\[94\] _0121_ state\[95\] _0122_ state\[96\] _0123_
+ state\[97\] _0124_ state\[98\] _0125_ state\[99\] _0126_ state\[100\] _0001_ state\[101\]
+ _0002_ state\[102\] _0003_ state\[103\] _0004_ state\[104\] _0005_ state\[105\]
+ _0006_ state\[106\] _0007_ state\[107\] _0008_ state\[108\] _0009_ state\[109\]
+ _0010_ state\[110\] _0012_ state\[111\] _0013_ state\[112\] _0014_ state\[113\]
+ _0015_ state\[114\] _0016_ state\[115\] _0017_ state\[116\] _0018_ state\[117\]
+ _0019_ state\[118\] _0020_ state\[119\] _0021_ state\[120\] _0023_ state\[121\]
+ _0024_ state\[122\] _0025_ digitalenL.g\[3\].u.OUTP digitalenL.g\[3\].u.OUTN state\[123\]
+ _0026_ state\[124\] _0027_ state\[125\] _0028_ state\[126\] _0029_ state\[127\]
+ _0030_ state\[0\] _0000_ state\[1\] _0039_ state\[2\] _0050_ state\[3\] _0061_ state\[4\]
+ _0072_ state\[5\] _0083_ state\[6\] digitalenL.g\[0\].u.OUTP digitalenL.g\[0\].u.OUTN
+ _0094_ state\[7\] _0105_ state\[8\] _0116_ state\[9\] _0127_ state\[10\] _0011_
+ state\[11\] _0022_ state\[12\] _0031_ state\[13\] _0032_ state\[14\] _0033_ state\[15\]
+ _0034_ state\[16\] _0035_ state\[17\] _0036_ state\[18\] _0037_ state\[19\] _0038_
+ state\[20\] _0040_ state\[21\] _0041_ state\[22\] _0042_ state\[23\] _0043_ state\[24\]
+ _0044_ state\[25\] _0045_ state\[26\] _0046_ state\[27\] _0047_ state\[28\] _0048_
+ state\[29\] _0049_ state\[30\] _0051_ state\[31\] _0052_ state\[33\] _0054_ state\[32\]
+ _0053_ state\[34\] _0055_ state\[35\] _0056_ state\[36\] _0057_ state\[37\] _0058_
+ state\[38\] _0059_ state\[39\] _0060_ state\[40\] _0062_ state\[41\] _0063_ state\[42\]
+ _0064_ state\[43\] _0065_ state\[44\] _0066_ state\[45\] _0067_ state\[46\] _0068_
+ state\[47\] _0069_ state\[48\] _0070_ state\[49\] _0071_ state\[50\] _0073_ state\[51\]
+ _0074_ state\[52\] _0075_ state\[53\] _0076_ state\[54\] _0077_ state\[55\] _0078_
+ state\[56\] _0079_ state\[57\] _0080_ state\[58\] _0081_ state\[59\] _0082_ state\[60\]
+ _0084_ state\[61\] _0085_ state\[62\] _0086_ state\[63\] _0087_ digitalenL.g\[1\].u.OUTP
+ digitalenL.g\[1\].u.OUTN VGND VPWR dac128module
XFILLER_7_189 VPWR VGND sg13g2_decap_8
XFILLER_22_81 VPWR VGND sg13g2_decap_8
XFILLER_4_830 VPWR VGND sg13g2_decap_8
XFILLER_4_896 VPWR VGND sg13g2_decap_8
XFILLER_3_340 VPWR VGND sg13g2_decap_8
X_2130_ _0936_ net138 state\[38\] VPWR VGND sg13g2_nand2_1
XFILLER_39_528 VPWR VGND sg13g2_decap_4
X_2061_ VGND VPWR _0524_ _0901_ _0387_ net71 sg13g2_a21oi_1
X_2376__352 VPWR VGND net351 sg13g2_tiehi
XFILLER_19_263 VPWR VGND sg13g2_decap_8
XFILLER_47_572 VPWR VGND sg13g2_decap_4
XFILLER_34_200 VPWR VGND sg13g2_decap_8
XFILLER_23_918 VPWR VGND sg13g2_decap_4
XFILLER_22_417 VPWR VGND sg13g2_decap_8
XFILLER_34_277 VPWR VGND sg13g2_decap_8
X_1914_ net224 VPWR _0793_ VGND state\[93\] net196 sg13g2_o21ai_1
X_1845_ VPWR VGND _0741_ net106 _0740_ _0228_ _0331_ net62 sg13g2_a221oi_1
X_1776_ VGND VPWR net144 daisychain\[57\] _0690_ net56 sg13g2_a21oi_1
X_2328_ net447 VGND VPWR _0274_ daisychain\[18\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2259_ VGND VPWR _0821_ _1000_ _0486_ net90 sg13g2_a21oi_1
XFILLER_26_723 VPWR VGND sg13g2_fill_1
XFILLER_26_701 VPWR VGND sg13g2_decap_4
XFILLER_25_200 VPWR VGND sg13g2_decap_8
XFILLER_38_594 VPWR VGND sg13g2_decap_8
XFILLER_43_14 VPWR VGND sg13g2_decap_8
XFILLER_13_417 VPWR VGND sg13g2_decap_8
XFILLER_40_203 VPWR VGND sg13g2_decap_8
XFILLER_25_277 VPWR VGND sg13g2_decap_8
XFILLER_22_951 VPWR VGND sg13g2_decap_8
XFILLER_4_137 VPWR VGND sg13g2_decap_8
XFILLER_49_1013 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_48_336 VPWR VGND sg13g2_decap_8
XFILLER_16_200 VPWR VGND sg13g2_decap_8
XFILLER_17_70 VPWR VGND sg13g2_decap_8
XFILLER_16_277 VPWR VGND sg13g2_decap_8
XFILLER_31_214 VPWR VGND sg13g2_decap_8
XFILLER_12_472 VPWR VGND sg13g2_decap_8
XFILLER_8_410 VPWR VGND sg13g2_decap_8
X_1630_ net223 VPWR _0580_ VGND state\[22\] net194 sg13g2_o21ai_1
X_1561_ VPWR VGND _0528_ net84 _0527_ _0200_ _0260_ net41 sg13g2_a221oi_1
X_1492_ VPWR _0197_ daisychain\[47\] VGND sg13g2_inv_1
X_2113_ VGND VPWR _0602_ _0927_ _0413_ net77 sg13g2_a21oi_1
XFILLER_39_336 VPWR VGND sg13g2_decap_8
X_2044_ VGND VPWR net113 daisychain\[124\] _0891_ net24 sg13g2_a21oi_1
XFILLER_35_553 VPWR VGND sg13g2_decap_8
XFILLER_23_704 VPWR VGND sg13g2_decap_8
Xfanout29 net32 net29 VPWR VGND sg13g2_buf_1
XFILLER_23_726 VPWR VGND sg13g2_fill_2
XFILLER_22_214 VPWR VGND sg13g2_decap_8
XFILLER_13_39 VPWR VGND sg13g2_decap_8
XFILLER_30_291 VPWR VGND sg13g2_decap_8
X_1828_ VGND VPWR net151 daisychain\[70\] _0729_ net60 sg13g2_a21oi_1
X_1759_ net192 _0205_ _0676_ _0677_ VPWR VGND sg13g2_a21o_1
XFILLER_38_14 VPWR VGND sg13g2_decap_8
XFILLER_13_214 VPWR VGND sg13g2_decap_8
XFILLER_9_207 VPWR VGND sg13g2_decap_8
XFILLER_41_589 VPWR VGND sg13g2_fill_2
XFILLER_22_781 VPWR VGND sg13g2_fill_2
XFILLER_21_291 VPWR VGND sg13g2_decap_8
XFILLER_6_925 VPWR VGND sg13g2_decap_8
XFILLER_5_424 VPWR VGND sg13g2_decap_8
XFILLER_1_630 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_49_623 VPWR VGND sg13g2_decap_4
XFILLER_49_667 VPWR VGND sg13g2_fill_1
XFILLER_49_656 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_44_350 VPWR VGND sg13g2_decap_8
XFILLER_12_291 VPWR VGND sg13g2_decap_8
X_2525__303 VPWR VGND net302 sg13g2_tiehi
XFILLER_8_284 VPWR VGND sg13g2_decap_8
X_1613_ VPWR VGND _0567_ net102 _0566_ _0164_ _0273_ net57 sg13g2_a221oi_1
X_1544_ VGND VPWR net123 net2 _0516_ net35 sg13g2_a21oi_1
Xfanout219 net220 net219 VPWR VGND sg13g2_buf_1
Xfanout208 net209 net208 VPWR VGND sg13g2_buf_1
XFILLER_5_95 VPWR VGND sg13g2_decap_8
XFILLER_4_490 VPWR VGND sg13g2_decap_8
X_1475_ VPWR _0216_ daisychain\[64\] VGND sg13g2_inv_1
XFILLER_39_133 VPWR VGND sg13g2_decap_8
XFILLER_28_818 VPWR VGND sg13g2_decap_8
X_2027_ net159 _0152_ _0877_ _0878_ VPWR VGND sg13g2_a21o_1
XFILLER_35_350 VPWR VGND sg13g2_decap_8
XFILLER_10_228 VPWR VGND sg13g2_decap_8
XFILLER_2_438 VPWR VGND sg13g2_decap_8
XFILLER_49_46 VPWR VGND sg13g2_decap_8
XFILLER_46_1027 VPWR VGND sg13g2_fill_2
XFILLER_45_147 VPWR VGND sg13g2_decap_8
X_2433__238 VPWR VGND net237 sg13g2_tiehi
XFILLER_26_361 VPWR VGND sg13g2_decap_8
XFILLER_14_578 VPWR VGND sg13g2_fill_2
XFILLER_41_364 VPWR VGND sg13g2_decap_8
XFILLER_14_60 VPWR VGND sg13g2_decap_8
XFILLER_6_733 VPWR VGND sg13g2_decap_4
XFILLER_5_221 VPWR VGND sg13g2_decap_8
XFILLER_6_755 VPWR VGND sg13g2_decap_8
XFILLER_5_298 VPWR VGND sg13g2_decap_8
XFILLER_30_81 VPWR VGND sg13g2_decap_8
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_49_431 VPWR VGND sg13g2_decap_8
XFILLER_18_851 VPWR VGND sg13g2_fill_1
XdigitalenL.g\[1\].u.inv1 VPWR digitalenL.g\[1\].u.OUTN net6 VGND sg13g2_inv_1
XFILLER_36_147 VPWR VGND sg13g2_decap_8
XFILLER_17_350 VPWR VGND sg13g2_decap_8
XFILLER_45_670 VPWR VGND sg13g2_decap_4
XFILLER_32_375 VPWR VGND sg13g2_decap_8
XFILLER_10_18 VPWR VGND sg13g2_decap_8
X_1527_ VPWR _0159_ daisychain\[12\] VGND sg13g2_inv_1
X_1458_ VPWR _0235_ daisychain\[81\] VGND sg13g2_inv_1
X_1389_ VPWR _0042_ state\[22\] VGND sg13g2_inv_1
XFILLER_28_648 VPWR VGND sg13g2_fill_2
XFILLER_28_659 VPWR VGND sg13g2_decap_8
XFILLER_27_147 VPWR VGND sg13g2_decap_8
XFILLER_11_515 VPWR VGND sg13g2_decap_8
XFILLER_23_375 VPWR VGND sg13g2_decap_8
XFILLER_3_703 VPWR VGND sg13g2_fill_2
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_2_235 VPWR VGND sg13g2_decap_8
XFILLER_47_913 VPWR VGND sg13g2_decap_8
XFILLER_46_434 VPWR VGND sg13g2_decap_8
XFILLER_20_1019 VPWR VGND sg13g2_decap_8
XFILLER_18_158 VPWR VGND sg13g2_decap_8
XFILLER_47_968 VPWR VGND sg13g2_decap_4
X_2335__434 VPWR VGND net433 sg13g2_tiehi
XFILLER_34_618 VPWR VGND sg13g2_decap_8
XFILLER_42_640 VPWR VGND sg13g2_decap_8
XFILLER_25_81 VPWR VGND sg13g2_decap_8
XFILLER_14_375 VPWR VGND sg13g2_decap_8
XFILLER_42_695 VPWR VGND sg13g2_fill_1
XFILLER_41_161 VPWR VGND sg13g2_decap_8
XFILLER_30_824 VPWR VGND sg13g2_decap_4
XFILLER_41_91 VPWR VGND sg13g2_decap_8
X_2430_ net243 VGND VPWR _0376_ daisychain\[120\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_6_585 VPWR VGND sg13g2_decap_8
X_2361_ net381 VGND VPWR _0307_ daisychain\[51\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2292_ _1017_ net126 state\[119\] VPWR VGND sg13g2_nand2_1
X_1312_ VPWR _0126_ state\[99\] VGND sg13g2_inv_1
XFILLER_2_791 VPWR VGND sg13g2_fill_1
XFILLER_37_434 VPWR VGND sg13g2_decap_8
XFILLER_2_74 VPWR VGND sg13g2_decap_8
XFILLER_25_607 VPWR VGND sg13g2_fill_2
XFILLER_25_629 VPWR VGND sg13g2_decap_4
XFILLER_33_673 VPWR VGND sg13g2_fill_2
XFILLER_21_802 VPWR VGND sg13g2_fill_2
XANTENNA_13 VPWR VGND _0249_ sg13g2_antennanp
XFILLER_32_172 VPWR VGND sg13g2_decap_8
XFILLER_20_312 VPWR VGND sg13g2_decap_8
XANTENNA_24 VPWR VGND _0140_ sg13g2_antennanp
XANTENNA_35 VPWR VGND _0243_ sg13g2_antennanp
XANTENNA_46 VPWR VGND daisychain\[127\] sg13g2_antennanp
XANTENNA_57 VPWR VGND _0187_ sg13g2_antennanp
X_2386__332 VPWR VGND net331 sg13g2_tiehi
XFILLER_20_389 VPWR VGND sg13g2_decap_8
XFILLER_21_39 VPWR VGND sg13g2_decap_8
X_2559_ net450 VGND VPWR _0505_ state\[121\] clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_43_448 VPWR VGND sg13g2_decap_8
XFILLER_30_109 VPWR VGND sg13g2_decap_8
XFILLER_11_312 VPWR VGND sg13g2_decap_8
XFILLER_23_172 VPWR VGND sg13g2_decap_8
XFILLER_11_389 VPWR VGND sg13g2_decap_8
XFILLER_3_566 VPWR VGND sg13g2_decap_8
XFILLER_46_231 VPWR VGND sg13g2_decap_8
XFILLER_47_776 VPWR VGND sg13g2_fill_2
XFILLER_36_91 VPWR VGND sg13g2_decap_8
XFILLER_43_971 VPWR VGND sg13g2_fill_2
XFILLER_21_109 VPWR VGND sg13g2_decap_8
XFILLER_14_172 VPWR VGND sg13g2_decap_8
X_1930_ net213 VPWR _0805_ VGND state\[97\] net175 sg13g2_o21ai_1
X_1861_ VPWR VGND _0753_ net104 _0752_ _0232_ _0335_ net59 sg13g2_a221oi_1
XFILLER_30_698 VPWR VGND sg13g2_decap_4
X_1792_ VGND VPWR net146 daisychain\[61\] _0702_ net54 sg13g2_a21oi_1
X_2485__297 VPWR VGND net296 sg13g2_tiehi
XFILLER_7_850 VPWR VGND sg13g2_fill_1
XFILLER_6_382 VPWR VGND sg13g2_decap_8
X_2413_ net277 VGND VPWR _0359_ daisychain\[103\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2344_ net415 VGND VPWR _0290_ daisychain\[34\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2275_ VGND VPWR _0845_ _1008_ _0494_ net84 sg13g2_a21oi_1
XFILLER_37_231 VPWR VGND sg13g2_decap_8
XFILLER_16_39 VPWR VGND sg13g2_decap_8
XFILLER_26_949 VPWR VGND sg13g2_decap_8
XFILLER_12_109 VPWR VGND sg13g2_decap_8
XFILLER_21_643 VPWR VGND sg13g2_decap_8
XFILLER_20_186 VPWR VGND sg13g2_decap_8
XFILLER_4_319 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_48_518 VPWR VGND sg13g2_decap_8
XFILLER_48_529 VPWR VGND sg13g2_fill_2
XFILLER_29_765 VPWR VGND sg13g2_fill_1
XFILLER_28_242 VPWR VGND sg13g2_decap_8
XFILLER_43_245 VPWR VGND sg13g2_decap_8
XFILLER_32_919 VPWR VGND sg13g2_fill_1
XFILLER_31_429 VPWR VGND sg13g2_fill_1
XFILLER_12_676 VPWR VGND sg13g2_fill_2
XFILLER_11_186 VPWR VGND sg13g2_decap_8
XFILLER_22_60 VPWR VGND sg13g2_decap_8
XFILLER_7_168 VPWR VGND sg13g2_decap_8
XFILLER_4_864 VPWR VGND sg13g2_decap_4
XFILLER_3_396 VPWR VGND sg13g2_decap_8
XFILLER_26_1003 VPWR VGND sg13g2_decap_4
X_2060_ _0901_ net115 state\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_19_242 VPWR VGND sg13g2_decap_8
XFILLER_35_702 VPWR VGND sg13g2_decap_4
XFILLER_35_735 VPWR VGND sg13g2_fill_1
XFILLER_34_256 VPWR VGND sg13g2_decap_8
X_1913_ VPWR VGND _0792_ net105 _0791_ _0247_ _0348_ net61 sg13g2_a221oi_1
XFILLER_30_462 VPWR VGND sg13g2_fill_1
XFILLER_30_451 VPWR VGND sg13g2_decap_8
X_1844_ VGND VPWR net154 daisychain\[74\] _0741_ net64 sg13g2_a21oi_1
X_1775_ net188 _0209_ _0688_ _0689_ VPWR VGND sg13g2_a21o_1
XFILLER_8_95 VPWR VGND sg13g2_decap_8
X_2327_ net449 VGND VPWR _0273_ daisychain\[17\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2258_ _1000_ net134 state\[102\] VPWR VGND sg13g2_nand2_1
XFILLER_27_49 VPWR VGND sg13g2_decap_8
X_2189_ VGND VPWR _0716_ _0965_ _0451_ net109 sg13g2_a21oi_1
XFILLER_26_735 VPWR VGND sg13g2_fill_2
XFILLER_41_716 VPWR VGND sg13g2_decap_4
XFILLER_25_256 VPWR VGND sg13g2_decap_8
XFILLER_40_259 VPWR VGND sg13g2_decap_8
XFILLER_21_451 VPWR VGND sg13g2_decap_8
XFILLER_21_484 VPWR VGND sg13g2_fill_1
XFILLER_4_116 VPWR VGND sg13g2_decap_8
XFILLER_1_812 VPWR VGND sg13g2_fill_1
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_48_315 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_16_256 VPWR VGND sg13g2_decap_8
XFILLER_32_716 VPWR VGND sg13g2_fill_1
XFILLER_32_705 VPWR VGND sg13g2_decap_8
XFILLER_32_749 VPWR VGND sg13g2_fill_1
XFILLER_32_727 VPWR VGND sg13g2_fill_2
XFILLER_12_451 VPWR VGND sg13g2_decap_8
X_2412__280 VPWR VGND net279 sg13g2_tiehi
XFILLER_33_81 VPWR VGND sg13g2_decap_8
XFILLER_8_488 VPWR VGND sg13g2_decap_8
X_1560_ VGND VPWR net128 daisychain\[3\] _0528_ net41 sg13g2_a21oi_1
XFILLER_4_650 VPWR VGND sg13g2_fill_2
X_1491_ VPWR _0198_ daisychain\[48\] VGND sg13g2_inv_1
XFILLER_4_672 VPWR VGND sg13g2_fill_2
XFILLER_3_193 VPWR VGND sg13g2_decap_8
XFILLER_39_315 VPWR VGND sg13g2_decap_8
X_2112_ _0927_ net121 state\[29\] VPWR VGND sg13g2_nand2_1
X_2043_ net159 _0156_ _0889_ _0890_ VPWR VGND sg13g2_a21o_1
XFILLER_47_392 VPWR VGND sg13g2_decap_8
XFILLER_13_18 VPWR VGND sg13g2_decap_8
XFILLER_30_270 VPWR VGND sg13g2_decap_8
X_1827_ net197 _0224_ _0727_ _0728_ VPWR VGND sg13g2_a21o_1
X_1758_ net222 VPWR _0676_ VGND state\[54\] net192 sg13g2_o21ai_1
X_1689_ VPWR VGND _0624_ net94 _0623_ _0185_ _0292_ net49 sg13g2_a221oi_1
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_45_329 VPWR VGND sg13g2_decap_8
XFILLER_38_392 VPWR VGND sg13g2_decap_8
XFILLER_21_270 VPWR VGND sg13g2_decap_8
XFILLER_5_403 VPWR VGND sg13g2_decap_8
XFILLER_6_959 VPWR VGND sg13g2_decap_4
XFILLER_1_686 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
XFILLER_49_679 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_45_830 VPWR VGND sg13g2_decap_8
XFILLER_36_329 VPWR VGND sg13g2_decap_8
XFILLER_28_81 VPWR VGND sg13g2_decap_8
XFILLER_17_532 VPWR VGND sg13g2_fill_1
XFILLER_17_565 VPWR VGND sg13g2_fill_1
XFILLER_32_524 VPWR VGND sg13g2_decap_4
XFILLER_32_557 VPWR VGND sg13g2_fill_1
XFILLER_44_91 VPWR VGND sg13g2_decap_8
XFILLER_12_270 VPWR VGND sg13g2_decap_8
XFILLER_8_263 VPWR VGND sg13g2_decap_8
X_1612_ VGND VPWR net148 daisychain\[16\] _0567_ net57 sg13g2_a21oi_1
X_2345__414 VPWR VGND net413 sg13g2_tiehi
X_1543_ net211 net3 _0515_ VPWR VGND sg13g2_nor2_1
Xfanout209 net210 net209 VPWR VGND sg13g2_buf_1
X_1474_ VPWR _0217_ daisychain\[65\] VGND sg13g2_inv_1
XFILLER_5_74 VPWR VGND sg13g2_decap_8
XFILLER_39_112 VPWR VGND sg13g2_decap_8
XFILLER_48_690 VPWR VGND sg13g2_fill_2
XFILLER_39_189 VPWR VGND sg13g2_decap_8
XFILLER_27_329 VPWR VGND sg13g2_decap_8
X_2026_ net205 VPWR _0877_ VGND state\[121\] net159 sg13g2_o21ai_1
XFILLER_23_502 VPWR VGND sg13g2_fill_1
XFILLER_24_39 VPWR VGND sg13g2_decap_8
XFILLER_10_207 VPWR VGND sg13g2_decap_8
XFILLER_40_49 VPWR VGND sg13g2_decap_8
XFILLER_2_417 VPWR VGND sg13g2_decap_8
XFILLER_49_25 VPWR VGND sg13g2_decap_8
X_2396__312 VPWR VGND net311 sg13g2_tiehi
XFILLER_45_126 VPWR VGND sg13g2_decap_8
XFILLER_26_340 VPWR VGND sg13g2_decap_8
XFILLER_27_885 VPWR VGND sg13g2_fill_2
XFILLER_14_557 VPWR VGND sg13g2_decap_4
XFILLER_42_888 VPWR VGND sg13g2_fill_1
XFILLER_41_343 VPWR VGND sg13g2_decap_8
XFILLER_5_200 VPWR VGND sg13g2_decap_8
XFILLER_5_277 VPWR VGND sg13g2_decap_8
XFILLER_30_60 VPWR VGND sg13g2_decap_8
XFILLER_2_951 VPWR VGND sg13g2_decap_8
XFILLER_2_995 VPWR VGND sg13g2_fill_2
XFILLER_7_1011 VPWR VGND sg13g2_decap_8
XFILLER_49_410 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_39_91 VPWR VGND sg13g2_decap_8
XFILLER_18_830 VPWR VGND sg13g2_fill_1
XFILLER_49_487 VPWR VGND sg13g2_decap_8
XFILLER_37_627 VPWR VGND sg13g2_decap_8
XFILLER_36_126 VPWR VGND sg13g2_decap_8
XdigitalenL.g\[1\].u.inv2 VPWR digitalenL.g\[1\].u.OUTP digitalenL.g\[1\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_32_354 VPWR VGND sg13g2_decap_8
XFILLER_9_550 VPWR VGND sg13g2_decap_8
X_1526_ VPWR _0160_ daisychain\[13\] VGND sg13g2_inv_1
X_1457_ VPWR _0236_ daisychain\[82\] VGND sg13g2_inv_1
XFILLER_19_39 VPWR VGND sg13g2_decap_8
X_1388_ VPWR _0043_ state\[23\] VGND sg13g2_inv_1
XFILLER_28_638 VPWR VGND sg13g2_decap_4
XFILLER_27_126 VPWR VGND sg13g2_decap_8
XFILLER_35_49 VPWR VGND sg13g2_decap_8
X_2009_ VPWR VGND _0864_ net88 _0863_ _0146_ _0372_ net45 sg13g2_a221oi_1
XFILLER_23_354 VPWR VGND sg13g2_decap_8
XFILLER_2_214 VPWR VGND sg13g2_decap_8
XFILLER_47_925 VPWR VGND sg13g2_decap_8
XFILLER_46_413 VPWR VGND sg13g2_decap_8
XFILLER_18_137 VPWR VGND sg13g2_decap_8
XFILLER_14_354 VPWR VGND sg13g2_decap_8
XFILLER_42_652 VPWR VGND sg13g2_fill_1
XFILLER_41_140 VPWR VGND sg13g2_decap_8
XFILLER_25_60 VPWR VGND sg13g2_decap_8
XFILLER_10_593 VPWR VGND sg13g2_fill_2
X_2561__323 VPWR VGND net322 sg13g2_tiehi
XFILLER_41_70 VPWR VGND sg13g2_decap_8
XFILLER_6_564 VPWR VGND sg13g2_decap_8
X_2360_ net383 VGND VPWR _0306_ daisychain\[50\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2291_ VGND VPWR _0869_ _1016_ _0502_ net91 sg13g2_a21oi_1
X_1311_ VPWR _0001_ state\[100\] VGND sg13g2_inv_1
XFILLER_2_53 VPWR VGND sg13g2_decap_8
XFILLER_1_280 VPWR VGND sg13g2_decap_8
XFILLER_49_284 VPWR VGND sg13g2_decap_8
XFILLER_37_413 VPWR VGND sg13g2_decap_8
XFILLER_46_980 VPWR VGND sg13g2_fill_1
XANTENNA_14 VPWR VGND daisychain\[110\] sg13g2_antennanp
XFILLER_32_151 VPWR VGND sg13g2_decap_8
XFILLER_21_847 VPWR VGND sg13g2_fill_1
XANTENNA_25 VPWR VGND _0140_ sg13g2_antennanp
XANTENNA_36 VPWR VGND _0250_ sg13g2_antennanp
XANTENNA_47 VPWR VGND daisychain\[15\] sg13g2_antennanp
XANTENNA_58 VPWR VGND daisychain\[100\] sg13g2_antennanp
XFILLER_21_18 VPWR VGND sg13g2_decap_8
XFILLER_20_368 VPWR VGND sg13g2_decap_8
XFILLER_0_729 VPWR VGND sg13g2_decap_4
X_2558_ net242 VGND VPWR _0504_ state\[120\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2489_ net280 VGND VPWR _0435_ state\[51\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1509_ VPWR _0179_ daisychain\[30\] VGND sg13g2_inv_1
XFILLER_29_903 VPWR VGND sg13g2_decap_8
XFILLER_28_424 VPWR VGND sg13g2_decap_8
XFILLER_29_969 VPWR VGND sg13g2_decap_8
XFILLER_28_435 VPWR VGND sg13g2_decap_8
XFILLER_43_427 VPWR VGND sg13g2_decap_8
X_2514__391 VPWR VGND net390 sg13g2_tiehi
XFILLER_23_151 VPWR VGND sg13g2_decap_8
XFILLER_8_829 VPWR VGND sg13g2_fill_2
XFILLER_11_368 VPWR VGND sg13g2_decap_8
XFILLER_3_545 VPWR VGND sg13g2_decap_8
XFILLER_11_95 VPWR VGND sg13g2_decap_8
XFILLER_47_766 VPWR VGND sg13g2_decap_4
XFILLER_46_210 VPWR VGND sg13g2_decap_8
XFILLER_19_446 VPWR VGND sg13g2_fill_2
XFILLER_15_630 VPWR VGND sg13g2_decap_8
XFILLER_46_287 VPWR VGND sg13g2_decap_8
XFILLER_36_70 VPWR VGND sg13g2_decap_8
XFILLER_34_449 VPWR VGND sg13g2_decap_8
XFILLER_27_490 VPWR VGND sg13g2_fill_2
XFILLER_15_641 VPWR VGND sg13g2_fill_2
XFILLER_14_151 VPWR VGND sg13g2_decap_8
XFILLER_15_685 VPWR VGND sg13g2_decap_8
X_1860_ VGND VPWR net150 daisychain\[78\] _0753_ net59 sg13g2_a21oi_1
X_1791_ net190 _0214_ _0700_ _0701_ VPWR VGND sg13g2_a21o_1
XFILLER_7_884 VPWR VGND sg13g2_decap_8
XFILLER_7_862 VPWR VGND sg13g2_decap_8
XFILLER_6_361 VPWR VGND sg13g2_decap_8
X_2526__295 VPWR VGND net294 sg13g2_tiehi
X_2412_ net279 VGND VPWR _0358_ daisychain\[102\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2343_ net417 VGND VPWR _0289_ daisychain\[33\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2422__260 VPWR VGND net259 sg13g2_tiehi
X_2274_ _1008_ net128 state\[110\] VPWR VGND sg13g2_nand2_1
XFILLER_42_1020 VPWR VGND sg13g2_decap_8
XFILLER_38_733 VPWR VGND sg13g2_decap_4
XFILLER_37_210 VPWR VGND sg13g2_decap_8
X_2492__269 VPWR VGND net268 sg13g2_tiehi
XFILLER_26_928 VPWR VGND sg13g2_decap_4
XFILLER_16_18 VPWR VGND sg13g2_decap_8
XFILLER_37_287 VPWR VGND sg13g2_decap_8
XFILLER_25_438 VPWR VGND sg13g2_decap_4
XFILLER_18_490 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_17_clk clknet_2_2__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
X_2353__398 VPWR VGND net397 sg13g2_tiehi
XFILLER_33_460 VPWR VGND sg13g2_decap_8
XFILLER_32_39 VPWR VGND sg13g2_decap_8
XFILLER_20_165 VPWR VGND sg13g2_decap_8
X_1989_ VPWR VGND _0849_ net80 _0848_ _0141_ _0367_ net34 sg13g2_a221oi_1
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_29_755 VPWR VGND sg13g2_fill_1
XFILLER_29_744 VPWR VGND sg13g2_decap_8
XFILLER_28_221 VPWR VGND sg13g2_decap_8
XFILLER_43_224 VPWR VGND sg13g2_decap_8
XFILLER_28_298 VPWR VGND sg13g2_decap_8
XFILLER_12_611 VPWR VGND sg13g2_decap_4
XFILLER_12_633 VPWR VGND sg13g2_decap_8
XFILLER_11_165 VPWR VGND sg13g2_decap_8
X_2549__251 VPWR VGND net250 sg13g2_tiehi
XFILLER_7_147 VPWR VGND sg13g2_decap_8
XFILLER_3_375 VPWR VGND sg13g2_decap_8
XFILLER_26_1015 VPWR VGND sg13g2_decap_8
XFILLER_19_221 VPWR VGND sg13g2_decap_8
XFILLER_47_91 VPWR VGND sg13g2_decap_8
XFILLER_19_298 VPWR VGND sg13g2_decap_8
XFILLER_34_235 VPWR VGND sg13g2_decap_8
XFILLER_43_780 VPWR VGND sg13g2_fill_1
X_1912_ VGND VPWR net151 daisychain\[91\] _0792_ net61 sg13g2_a21oi_1
XFILLER_31_953 VPWR VGND sg13g2_fill_1
X_1843_ net199 _0228_ _0739_ _0740_ VPWR VGND sg13g2_a21o_1
XFILLER_8_74 VPWR VGND sg13g2_decap_8
X_1774_ net221 VPWR _0688_ VGND state\[58\] net188 sg13g2_o21ai_1
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
XFILLER_40_0 VPWR VGND sg13g2_decap_8
X_2326_ net451 VGND VPWR _0272_ daisychain\[16\] clknet_leaf_8_clk sg13g2_dfrbpq_1
X_2257_ VGND VPWR _0818_ _0999_ _0485_ net89 sg13g2_a21oi_1
XFILLER_27_28 VPWR VGND sg13g2_decap_8
X_2188_ _0965_ net156 state\[67\] VPWR VGND sg13g2_nand2_1
XFILLER_25_235 VPWR VGND sg13g2_decap_8
XFILLER_43_49 VPWR VGND sg13g2_decap_8
XFILLER_40_238 VPWR VGND sg13g2_decap_8
XFILLER_5_618 VPWR VGND sg13g2_decap_8
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
XFILLER_49_817 VPWR VGND sg13g2_fill_2
XFILLER_17_725 VPWR VGND sg13g2_decap_8
XFILLER_16_235 VPWR VGND sg13g2_decap_8
XFILLER_25_780 VPWR VGND sg13g2_decap_8
XFILLER_12_430 VPWR VGND sg13g2_decap_8
XFILLER_31_249 VPWR VGND sg13g2_decap_8
XFILLER_25_791 VPWR VGND sg13g2_fill_2
XFILLER_33_60 VPWR VGND sg13g2_decap_8
XFILLER_8_467 VPWR VGND sg13g2_decap_8
X_1490_ VPWR _0199_ daisychain\[49\] VGND sg13g2_inv_1
XFILLER_3_172 VPWR VGND sg13g2_decap_8
XFILLER_0_890 VPWR VGND sg13g2_decap_4
XFILLER_12_4 VPWR VGND sg13g2_decap_8
X_2111_ VGND VPWR _0599_ _0926_ _0412_ net75 sg13g2_a21oi_1
X_2042_ net205 VPWR _0889_ VGND state\[125\] net159 sg13g2_o21ai_1
XFILLER_47_371 VPWR VGND sg13g2_decap_8
XFILLER_23_728 VPWR VGND sg13g2_fill_1
XFILLER_22_249 VPWR VGND sg13g2_decap_8
X_1826_ net224 VPWR _0727_ VGND state\[71\] net197 sg13g2_o21ai_1
X_1757_ VPWR VGND _0675_ net99 _0674_ _0204_ _0309_ net53 sg13g2_a221oi_1
X_1688_ VGND VPWR net140 daisychain\[35\] _0624_ net49 sg13g2_a21oi_1
X_2309_ VGND VPWR _0896_ _1025_ _0511_ net72 sg13g2_a21oi_1
XFILLER_38_49 VPWR VGND sg13g2_decap_8
XFILLER_45_308 VPWR VGND sg13g2_decap_8
XFILLER_38_371 VPWR VGND sg13g2_decap_8
XFILLER_26_511 VPWR VGND sg13g2_fill_2
XFILLER_13_249 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_490 VPWR VGND uio_oe[6] sg13g2_tiehi
XFILLER_5_459 VPWR VGND sg13g2_decap_8
XFILLER_49_603 VPWR VGND sg13g2_fill_2
XFILLER_1_665 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_36_308 VPWR VGND sg13g2_decap_8
XFILLER_29_382 VPWR VGND sg13g2_decap_8
XFILLER_28_60 VPWR VGND sg13g2_decap_8
XFILLER_17_577 VPWR VGND sg13g2_fill_2
XFILLER_45_875 VPWR VGND sg13g2_decap_4
XFILLER_44_70 VPWR VGND sg13g2_decap_8
XFILLER_44_385 VPWR VGND sg13g2_decap_8
XFILLER_9_732 VPWR VGND sg13g2_fill_1
XFILLER_8_242 VPWR VGND sg13g2_decap_8
X_1611_ net187 _0164_ _0565_ _0566_ VPWR VGND sg13g2_a21o_1
X_1542_ net170 _0128_ _0513_ _0514_ VPWR VGND sg13g2_a21o_1
XFILLER_5_53 VPWR VGND sg13g2_decap_8
XFILLER_4_470 VPWR VGND sg13g2_fill_2
X_1473_ VPWR _0218_ daisychain\[66\] VGND sg13g2_inv_1
XFILLER_39_168 VPWR VGND sg13g2_decap_8
XFILLER_27_308 VPWR VGND sg13g2_decap_8
X_2025_ VPWR VGND _0876_ net83 _0875_ _0151_ _0376_ net38 sg13g2_a221oi_1
XFILLER_23_514 VPWR VGND sg13g2_decap_8
XFILLER_35_385 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_8
XFILLER_40_28 VPWR VGND sg13g2_decap_8
X_1809_ VPWR VGND _0714_ net107 _0713_ _0218_ _0322_ net63 sg13g2_a221oi_1
XFILLER_18_319 VPWR VGND sg13g2_decap_8
XFILLER_45_105 VPWR VGND sg13g2_decap_8
XFILLER_42_801 VPWR VGND sg13g2_fill_1
XFILLER_27_897 VPWR VGND sg13g2_fill_1
XFILLER_41_322 VPWR VGND sg13g2_decap_8
XFILLER_26_396 VPWR VGND sg13g2_decap_8
XFILLER_42_878 VPWR VGND sg13g2_fill_1
XFILLER_41_399 VPWR VGND sg13g2_decap_8
XFILLER_22_580 VPWR VGND sg13g2_decap_8
XFILLER_14_95 VPWR VGND sg13g2_decap_8
XFILLER_22_591 VPWR VGND sg13g2_fill_1
XFILLER_5_256 VPWR VGND sg13g2_decap_8
XFILLER_2_930 VPWR VGND sg13g2_fill_1
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_49_466 VPWR VGND sg13g2_decap_8
XFILLER_39_70 VPWR VGND sg13g2_decap_8
XFILLER_36_105 VPWR VGND sg13g2_decap_8
XFILLER_18_842 VPWR VGND sg13g2_fill_2
XFILLER_17_385 VPWR VGND sg13g2_decap_8
XFILLER_44_182 VPWR VGND sg13g2_decap_8
XFILLER_32_333 VPWR VGND sg13g2_decap_8
X_2488__285 VPWR VGND net284 sg13g2_tiehi
X_2529__271 VPWR VGND net270 sg13g2_tiehi
X_1525_ VPWR _0161_ daisychain\[14\] VGND sg13g2_inv_1
XFILLER_19_18 VPWR VGND sg13g2_decap_8
X_1456_ VPWR _0237_ daisychain\[83\] VGND sg13g2_inv_1
X_1387_ VPWR _0044_ state\[24\] VGND sg13g2_inv_1
XFILLER_28_617 VPWR VGND sg13g2_fill_2
XFILLER_27_105 VPWR VGND sg13g2_decap_8
XFILLER_35_28 VPWR VGND sg13g2_decap_8
X_2008_ VGND VPWR net132 daisychain\[115\] _0864_ net45 sg13g2_a21oi_1
X_2432__240 VPWR VGND net239 sg13g2_tiehi
XFILLER_42_119 VPWR VGND sg13g2_decap_8
XFILLER_35_182 VPWR VGND sg13g2_decap_8
XFILLER_23_333 VPWR VGND sg13g2_decap_8
X_2467__369 VPWR VGND net368 sg13g2_tiehi
XFILLER_3_727 VPWR VGND sg13g2_decap_8
XFILLER_3_705 VPWR VGND sg13g2_fill_1
X_2363__378 VPWR VGND net377 sg13g2_tiehi
XFILLER_3_738 VPWR VGND sg13g2_fill_1
XFILLER_18_116 VPWR VGND sg13g2_decap_8
XFILLER_46_469 VPWR VGND sg13g2_decap_8
XFILLER_14_333 VPWR VGND sg13g2_decap_8
XFILLER_26_193 VPWR VGND sg13g2_decap_8
XFILLER_41_196 VPWR VGND sg13g2_decap_8
XFILLER_10_550 VPWR VGND sg13g2_decap_8
XFILLER_6_543 VPWR VGND sg13g2_decap_8
X_2409__286 VPWR VGND net285 sg13g2_tiehi
Xheichips25_pudding VPWR VGND uio_oe[0] sg13g2_tiehi
XFILLER_44_7 VPWR VGND sg13g2_decap_8
XFILLER_29_1024 VPWR VGND sg13g2_decap_4
X_2290_ _1016_ net127 state\[118\] VPWR VGND sg13g2_nand2_1
X_1310_ VPWR _0002_ state\[101\] VGND sg13g2_inv_1
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_49_263 VPWR VGND sg13g2_decap_8
XFILLER_37_469 VPWR VGND sg13g2_decap_8
XFILLER_17_182 VPWR VGND sg13g2_decap_8
XFILLER_33_642 VPWR VGND sg13g2_decap_8
XFILLER_32_130 VPWR VGND sg13g2_decap_8
XANTENNA_15 VPWR VGND daisychain\[110\] sg13g2_antennanp
XANTENNA_26 VPWR VGND _0166_ sg13g2_antennanp
XANTENNA_37 VPWR VGND _0251_ sg13g2_antennanp
XANTENNA_48 VPWR VGND daisychain\[29\] sg13g2_antennanp
XFILLER_20_347 VPWR VGND sg13g2_decap_8
XANTENNA_59 VPWR VGND daisychain\[126\] sg13g2_antennanp
X_2557_ net274 VGND VPWR _0503_ state\[119\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2488_ net284 VGND VPWR _0434_ state\[50\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1508_ VPWR _0180_ daisychain\[31\] VGND sg13g2_inv_1
X_1439_ VPWR _0129_ daisychain\[100\] VGND sg13g2_inv_1
XFILLER_29_948 VPWR VGND sg13g2_fill_2
XFILLER_28_403 VPWR VGND sg13g2_decap_8
XFILLER_46_49 VPWR VGND sg13g2_decap_8
XFILLER_44_929 VPWR VGND sg13g2_decap_8
XFILLER_43_406 VPWR VGND sg13g2_decap_8
XFILLER_23_130 VPWR VGND sg13g2_decap_8
XFILLER_11_347 VPWR VGND sg13g2_decap_8
XFILLER_7_329 VPWR VGND sg13g2_decap_8
XFILLER_11_74 VPWR VGND sg13g2_decap_8
XFILLER_3_524 VPWR VGND sg13g2_decap_8
XFILLER_47_701 VPWR VGND sg13g2_fill_2
XFILLER_19_414 VPWR VGND sg13g2_fill_2
XFILLER_19_403 VPWR VGND sg13g2_decap_8
XFILLER_46_266 VPWR VGND sg13g2_decap_8
XFILLER_34_428 VPWR VGND sg13g2_fill_2
XFILLER_34_417 VPWR VGND sg13g2_decap_8
XFILLER_14_130 VPWR VGND sg13g2_decap_8
XFILLER_43_973 VPWR VGND sg13g2_fill_1
XFILLER_15_675 VPWR VGND sg13g2_fill_2
XFILLER_43_984 VPWR VGND sg13g2_fill_1
XFILLER_42_450 VPWR VGND sg13g2_decap_4
XFILLER_30_601 VPWR VGND sg13g2_decap_8
X_1790_ net222 VPWR _0700_ VGND state\[62\] net190 sg13g2_o21ai_1
X_2563__419 VPWR VGND net418 sg13g2_tiehi
XFILLER_6_340 VPWR VGND sg13g2_decap_8
X_2411_ net281 VGND VPWR _0357_ daisychain\[101\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2342_ net419 VGND VPWR _0288_ daisychain\[32\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2273_ VGND VPWR _0842_ _1007_ _0493_ net86 sg13g2_a21oi_1
XFILLER_37_266 VPWR VGND sg13g2_decap_8
XFILLER_25_417 VPWR VGND sg13g2_decap_8
XFILLER_32_18 VPWR VGND sg13g2_decap_8
XFILLER_20_144 VPWR VGND sg13g2_decap_8
X_1988_ VGND VPWR net128 daisychain\[110\] _0849_ net43 sg13g2_a21oi_1
XFILLER_28_200 VPWR VGND sg13g2_decap_8
Xclkbuf_2_2__f_clk clknet_2_2__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_44_704 VPWR VGND sg13g2_decap_8
XFILLER_29_789 VPWR VGND sg13g2_fill_1
XFILLER_29_778 VPWR VGND sg13g2_decap_8
XFILLER_16_417 VPWR VGND sg13g2_decap_8
XFILLER_44_748 VPWR VGND sg13g2_decap_4
XFILLER_43_203 VPWR VGND sg13g2_decap_8
XFILLER_28_277 VPWR VGND sg13g2_decap_8
XFILLER_25_995 VPWR VGND sg13g2_fill_2
XFILLER_11_144 VPWR VGND sg13g2_decap_8
XFILLER_8_638 VPWR VGND sg13g2_decap_8
XFILLER_8_605 VPWR VGND sg13g2_decap_4
XFILLER_7_126 VPWR VGND sg13g2_decap_8
XFILLER_22_95 VPWR VGND sg13g2_decap_8
XFILLER_3_354 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_19_200 VPWR VGND sg13g2_decap_8
Xfanout190 net191 net190 VPWR VGND sg13g2_buf_1
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_19_277 VPWR VGND sg13g2_decap_8
XFILLER_47_597 VPWR VGND sg13g2_decap_8
XFILLER_35_726 VPWR VGND sg13g2_decap_8
XFILLER_34_214 VPWR VGND sg13g2_decap_8
XFILLER_31_921 VPWR VGND sg13g2_fill_2
X_1911_ net197 _0247_ _0790_ _0791_ VPWR VGND sg13g2_a21o_1
XFILLER_42_280 VPWR VGND sg13g2_decap_8
X_1842_ net225 VPWR _0739_ VGND state\[75\] net199 sg13g2_o21ai_1
XFILLER_8_53 VPWR VGND sg13g2_decap_8
XFILLER_31_998 VPWR VGND sg13g2_fill_2
XFILLER_30_475 VPWR VGND sg13g2_fill_2
X_1773_ VPWR VGND _0687_ net97 _0686_ _0208_ _0313_ net56 sg13g2_a221oi_1
XFILLER_7_660 VPWR VGND sg13g2_fill_1
XFILLER_7_693 VPWR VGND sg13g2_fill_1
XFILLER_7_682 VPWR VGND sg13g2_decap_8
X_2325_ net453 VGND VPWR _0271_ daisychain\[15\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2256_ _0999_ net133 state\[101\] VPWR VGND sg13g2_nand2_1
X_2187_ VGND VPWR _0713_ _0964_ _0450_ net107 sg13g2_a21oi_1
XFILLER_38_575 VPWR VGND sg13g2_fill_2
XFILLER_26_737 VPWR VGND sg13g2_fill_1
XFILLER_25_214 VPWR VGND sg13g2_decap_8
XFILLER_26_759 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
XFILLER_40_217 VPWR VGND sg13g2_decap_8
XFILLER_22_921 VPWR VGND sg13g2_decap_4
XFILLER_21_431 VPWR VGND sg13g2_decap_8
XFILLER_33_291 VPWR VGND sg13g2_decap_8
XFILLER_21_475 VPWR VGND sg13g2_decap_8
XFILLER_49_1027 VPWR VGND sg13g2_fill_2
XFILLER_1_869 VPWR VGND sg13g2_fill_2
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_16_214 VPWR VGND sg13g2_decap_8
XFILLER_17_84 VPWR VGND sg13g2_decap_8
XFILLER_32_729 VPWR VGND sg13g2_fill_1
XFILLER_31_228 VPWR VGND sg13g2_decap_8
XFILLER_24_291 VPWR VGND sg13g2_decap_8
XFILLER_12_486 VPWR VGND sg13g2_decap_8
XFILLER_8_446 VPWR VGND sg13g2_decap_8
XFILLER_8_424 VPWR VGND sg13g2_decap_8
XFILLER_4_652 VPWR VGND sg13g2_fill_1
XFILLER_4_630 VPWR VGND sg13g2_decap_8
XFILLER_3_151 VPWR VGND sg13g2_decap_8
XFILLER_0_880 VPWR VGND sg13g2_fill_1
X_2110_ _0926_ net118 state\[28\] VPWR VGND sg13g2_nand2_1
X_2041_ VPWR VGND _0888_ net71 _0887_ _0155_ _0380_ net24 sg13g2_a221oi_1
XFILLER_47_350 VPWR VGND sg13g2_decap_8
XFILLER_35_523 VPWR VGND sg13g2_decap_8
XFILLER_35_545 VPWR VGND sg13g2_fill_2
XFILLER_35_534 VPWR VGND sg13g2_fill_2
XFILLER_22_228 VPWR VGND sg13g2_decap_8
XFILLER_15_291 VPWR VGND sg13g2_decap_8
XFILLER_31_751 VPWR VGND sg13g2_decap_8
X_1825_ VPWR VGND _0726_ net108 _0725_ _0223_ _0326_ net65 sg13g2_a221oi_1
X_1756_ VGND VPWR net145 daisychain\[52\] _0675_ net53 sg13g2_a21oi_1
XFILLER_7_490 VPWR VGND sg13g2_decap_8
X_1687_ net186 _0185_ _0622_ _0623_ VPWR VGND sg13g2_a21o_1
X_2308_ _1025_ state\[127\] net115 VPWR VGND sg13g2_nand2_1
XFILLER_38_28 VPWR VGND sg13g2_decap_8
X_2239_ VGND VPWR _0791_ _0990_ _0476_ net105 sg13g2_a21oi_1
XFILLER_38_350 VPWR VGND sg13g2_decap_8
XFILLER_13_228 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_491 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_22_773 VPWR VGND sg13g2_fill_2
XFILLER_5_438 VPWR VGND sg13g2_decap_8
X_2546__299 VPWR VGND net298 sg13g2_tiehi
XFILLER_1_644 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_29_361 VPWR VGND sg13g2_decap_8
X_2373__358 VPWR VGND net357 sg13g2_tiehi
XFILLER_17_589 VPWR VGND sg13g2_fill_2
XFILLER_44_364 VPWR VGND sg13g2_decap_8
XFILLER_8_221 VPWR VGND sg13g2_decap_8
X_1610_ net220 VPWR _0565_ VGND state\[17\] net187 sg13g2_o21ai_1
XFILLER_8_298 VPWR VGND sg13g2_decap_8
X_1541_ net211 VPWR _0513_ VGND state\[0\] net170 sg13g2_o21ai_1
XFILLER_5_32 VPWR VGND sg13g2_decap_8
X_1472_ VPWR _0219_ daisychain\[67\] VGND sg13g2_inv_1
X_2460__397 VPWR VGND net396 sg13g2_tiehi
XFILLER_39_147 VPWR VGND sg13g2_decap_8
X_2024_ VGND VPWR net127 daisychain\[119\] _0876_ net38 sg13g2_a21oi_1
X_2419__266 VPWR VGND net265 sg13g2_tiehi
XFILLER_35_364 VPWR VGND sg13g2_decap_8
X_1808_ VGND VPWR net157 daisychain\[65\] _0714_ net64 sg13g2_a21oi_1
X_1739_ net192 _0199_ _0661_ _0662_ VPWR VGND sg13g2_a21o_1
XFILLER_46_629 VPWR VGND sg13g2_decap_8
XFILLER_14_504 VPWR VGND sg13g2_decap_4
XFILLER_27_887 VPWR VGND sg13g2_fill_1
XFILLER_41_301 VPWR VGND sg13g2_decap_8
XFILLER_26_375 VPWR VGND sg13g2_decap_8
XFILLER_41_378 VPWR VGND sg13g2_decap_8
XFILLER_10_721 VPWR VGND sg13g2_decap_8
XFILLER_10_732 VPWR VGND sg13g2_fill_1
XFILLER_14_74 VPWR VGND sg13g2_decap_8
XFILLER_6_769 VPWR VGND sg13g2_fill_2
XFILLER_5_235 VPWR VGND sg13g2_decap_8
XFILLER_30_95 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_49_445 VPWR VGND sg13g2_decap_8
XFILLER_18_821 VPWR VGND sg13g2_fill_2
XFILLER_17_364 VPWR VGND sg13g2_decap_8
XFILLER_44_161 VPWR VGND sg13g2_decap_8
XFILLER_32_312 VPWR VGND sg13g2_decap_8
XFILLER_32_389 VPWR VGND sg13g2_decap_8
XFILLER_13_592 VPWR VGND sg13g2_fill_2
X_1524_ VPWR _0162_ daisychain\[15\] VGND sg13g2_inv_1
X_1455_ VPWR _0238_ daisychain\[84\] VGND sg13g2_inv_1
X_2495__257 VPWR VGND net256 sg13g2_tiehi
X_1386_ VPWR _0045_ state\[25\] VGND sg13g2_inv_1
X_2007_ net182 _0146_ _0862_ _0863_ VPWR VGND sg13g2_a21o_1
XFILLER_35_161 VPWR VGND sg13g2_decap_8
XFILLER_24_846 VPWR VGND sg13g2_decap_4
XFILLER_23_312 VPWR VGND sg13g2_decap_8
XFILLER_11_529 VPWR VGND sg13g2_decap_8
XFILLER_23_389 VPWR VGND sg13g2_decap_8
XFILLER_2_249 VPWR VGND sg13g2_decap_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
XFILLER_33_109 VPWR VGND sg13g2_decap_8
XFILLER_14_312 VPWR VGND sg13g2_decap_8
XFILLER_26_172 VPWR VGND sg13g2_decap_8
XFILLER_42_665 VPWR VGND sg13g2_fill_1
XFILLER_14_389 VPWR VGND sg13g2_decap_8
XFILLER_41_175 VPWR VGND sg13g2_decap_8
XFILLER_25_95 VPWR VGND sg13g2_decap_8
XFILLER_10_595 VPWR VGND sg13g2_fill_1
XFILLER_6_522 VPWR VGND sg13g2_decap_8
XFILLER_6_599 VPWR VGND sg13g2_fill_2
XFILLER_2_750 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_49_242 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_37_448 VPWR VGND sg13g2_decap_8
XFILLER_2_88 VPWR VGND sg13g2_decap_8
XFILLER_17_161 VPWR VGND sg13g2_decap_8
XFILLER_18_684 VPWR VGND sg13g2_fill_2
XFILLER_24_109 VPWR VGND sg13g2_decap_8
XANTENNA_16 VPWR VGND daisychain\[113\] sg13g2_antennanp
XANTENNA_27 VPWR VGND _0179_ sg13g2_antennanp
XANTENNA_38 VPWR VGND _0253_ sg13g2_antennanp
XFILLER_32_186 VPWR VGND sg13g2_decap_8
XFILLER_20_326 VPWR VGND sg13g2_decap_8
XANTENNA_49 VPWR VGND daisychain\[29\] sg13g2_antennanp
XFILLER_9_382 VPWR VGND sg13g2_decap_8
XFILLER_0_709 VPWR VGND sg13g2_decap_4
X_2556_ net306 VGND VPWR _0502_ state\[118\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2487_ net288 VGND VPWR _0433_ state\[49\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1507_ VPWR _0181_ daisychain\[32\] VGND sg13g2_inv_1
X_1438_ VPWR _0130_ daisychain\[101\] VGND sg13g2_inv_1
X_1369_ VPWR _0064_ state\[42\] VGND sg13g2_inv_1
XFILLER_46_28 VPWR VGND sg13g2_decap_8
XFILLER_15_109 VPWR VGND sg13g2_decap_8
XFILLER_24_698 VPWR VGND sg13g2_decap_8
XFILLER_11_326 VPWR VGND sg13g2_decap_8
XFILLER_23_186 VPWR VGND sg13g2_decap_8
XFILLER_7_308 VPWR VGND sg13g2_decap_8
XFILLER_3_503 VPWR VGND sg13g2_decap_8
XFILLER_11_53 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_47_735 VPWR VGND sg13g2_fill_2
XFILLER_46_245 VPWR VGND sg13g2_decap_8
XFILLER_19_459 VPWR VGND sg13g2_decap_8
XFILLER_15_654 VPWR VGND sg13g2_fill_2
XFILLER_14_186 VPWR VGND sg13g2_decap_8
XFILLER_30_646 VPWR VGND sg13g2_fill_2
XFILLER_7_820 VPWR VGND sg13g2_fill_1
X_2410_ net283 VGND VPWR _0356_ daisychain\[100\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_6_396 VPWR VGND sg13g2_decap_8
X_2341_ net421 VGND VPWR _0287_ daisychain\[31\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2272_ _1007_ net130 state\[109\] VPWR VGND sg13g2_nand2_1
XFILLER_37_245 VPWR VGND sg13g2_decap_8
XFILLER_20_123 VPWR VGND sg13g2_decap_8
X_1987_ net175 _0141_ _0847_ _0848_ VPWR VGND sg13g2_a21o_1
X_2544__331 VPWR VGND net330 sg13g2_tiehi
X_2539_ net410 VGND VPWR _0485_ state\[101\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_0_539 VPWR VGND sg13g2_decap_8
X_2401__302 VPWR VGND net301 sg13g2_tiehi
XFILLER_28_256 VPWR VGND sg13g2_decap_8
XFILLER_43_259 VPWR VGND sg13g2_decap_8
XFILLER_24_451 VPWR VGND sg13g2_fill_2
XFILLER_11_123 VPWR VGND sg13g2_decap_8
XFILLER_7_105 VPWR VGND sg13g2_decap_8
XFILLER_22_74 VPWR VGND sg13g2_decap_8
XFILLER_4_823 VPWR VGND sg13g2_decap_8
XFILLER_3_333 VPWR VGND sg13g2_decap_8
Xfanout191 net193 net191 VPWR VGND sg13g2_buf_1
Xfanout180 net182 net180 VPWR VGND sg13g2_buf_1
XFILLER_19_256 VPWR VGND sg13g2_decap_8
XFILLER_47_565 VPWR VGND sg13g2_decap_8
XFILLER_28_790 VPWR VGND sg13g2_decap_8
XFILLER_43_760 VPWR VGND sg13g2_fill_1
X_1910_ net224 VPWR _0790_ VGND state\[92\] net197 sg13g2_o21ai_1
XFILLER_30_410 VPWR VGND sg13g2_decap_8
X_1841_ VPWR VGND _0738_ net106 _0737_ _0227_ _0330_ net62 sg13g2_a221oi_1
XFILLER_8_32 VPWR VGND sg13g2_decap_8
X_1772_ VGND VPWR net145 daisychain\[56\] _0687_ net53 sg13g2_a21oi_1
X_2383__338 VPWR VGND net337 sg13g2_tiehi
XFILLER_6_193 VPWR VGND sg13g2_decap_8
X_2324_ net455 VGND VPWR _0270_ daisychain\[14\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2539__411 VPWR VGND net410 sg13g2_tiehi
X_2255_ VGND VPWR _0815_ _0998_ _0484_ net89 sg13g2_a21oi_1
X_2186_ _0964_ net153 state\[66\] VPWR VGND sg13g2_nand2_1
XFILLER_26_716 VPWR VGND sg13g2_decap_8
XFILLER_33_270 VPWR VGND sg13g2_decap_8
XFILLER_22_944 VPWR VGND sg13g2_decap_8
XFILLER_21_410 VPWR VGND sg13g2_decap_8
XFILLER_22_988 VPWR VGND sg13g2_fill_2
X_2429__246 VPWR VGND net245 sg13g2_tiehi
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_49_819 VPWR VGND sg13g2_fill_1
XFILLER_48_329 VPWR VGND sg13g2_decap_8
XFILLER_17_63 VPWR VGND sg13g2_decap_8
XFILLER_31_207 VPWR VGND sg13g2_decap_8
XFILLER_25_771 VPWR VGND sg13g2_decap_4
XFILLER_12_410 VPWR VGND sg13g2_fill_2
XFILLER_24_270 VPWR VGND sg13g2_decap_8
XFILLER_8_403 VPWR VGND sg13g2_decap_8
XFILLER_12_465 VPWR VGND sg13g2_decap_8
XFILLER_33_95 VPWR VGND sg13g2_decap_8
XFILLER_3_130 VPWR VGND sg13g2_decap_8
XFILLER_4_697 VPWR VGND sg13g2_decap_4
XFILLER_0_870 VPWR VGND sg13g2_decap_4
XFILLER_39_329 VPWR VGND sg13g2_decap_8
X_2040_ VGND VPWR net113 daisychain\[123\] _0888_ net24 sg13g2_a21oi_1
XFILLER_48_852 VPWR VGND sg13g2_fill_2
XFILLER_48_885 VPWR VGND sg13g2_decap_4
XFILLER_35_513 VPWR VGND sg13g2_decap_4
XFILLER_22_207 VPWR VGND sg13g2_decap_8
XFILLER_15_270 VPWR VGND sg13g2_decap_8
X_1824_ VGND VPWR net155 daisychain\[69\] _0726_ net65 sg13g2_a21oi_1
XFILLER_30_284 VPWR VGND sg13g2_decap_8
X_1755_ net189 _0204_ _0673_ _0674_ VPWR VGND sg13g2_a21o_1
X_1686_ net209 VPWR _0622_ VGND state\[36\] net163 sg13g2_o21ai_1
X_2307_ VGND VPWR _0893_ _1024_ _0510_ net69 sg13g2_a21oi_1
X_2238_ _0990_ net151 state\[92\] VPWR VGND sg13g2_nand2_1
X_2169_ VGND VPWR _0686_ _0955_ _0441_ net97 sg13g2_a21oi_1
XFILLER_13_207 VPWR VGND sg13g2_decap_8
XFILLER_41_527 VPWR VGND sg13g2_decap_8
XFILLER_6_907 VPWR VGND sg13g2_fill_2
XFILLER_21_284 VPWR VGND sg13g2_decap_8
XFILLER_5_417 VPWR VGND sg13g2_decap_8
XFILLER_1_623 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_49_616 VPWR VGND sg13g2_decap_8
XFILLER_49_649 VPWR VGND sg13g2_decap_8
XFILLER_49_627 VPWR VGND sg13g2_fill_2
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_29_340 VPWR VGND sg13g2_decap_8
XFILLER_28_95 VPWR VGND sg13g2_decap_8
XFILLER_17_557 VPWR VGND sg13g2_fill_2
XFILLER_17_579 VPWR VGND sg13g2_fill_1
XFILLER_44_343 VPWR VGND sg13g2_decap_8
XFILLER_8_200 VPWR VGND sg13g2_decap_8
XFILLER_12_284 VPWR VGND sg13g2_decap_8
XFILLER_8_277 VPWR VGND sg13g2_decap_8
X_1540_ VPWR _0512_ net1 VGND sg13g2_inv_1
XFILLER_5_11 VPWR VGND sg13g2_decap_8
X_1471_ VPWR _0220_ daisychain\[68\] VGND sg13g2_inv_1
XFILLER_5_88 VPWR VGND sg13g2_decap_8
XFILLER_4_483 VPWR VGND sg13g2_decap_8
XFILLER_39_126 VPWR VGND sg13g2_decap_8
X_2023_ net174 _0151_ _0874_ _0875_ VPWR VGND sg13g2_a21o_1
XFILLER_35_343 VPWR VGND sg13g2_decap_8
XFILLER_23_538 VPWR VGND sg13g2_decap_8
XFILLER_31_560 VPWR VGND sg13g2_fill_2
X_1807_ net200 _0218_ _0712_ _0713_ VPWR VGND sg13g2_a21o_1
X_1738_ net221 VPWR _0661_ VGND state\[49\] net188 sg13g2_o21ai_1
X_1669_ VPWR VGND _0609_ net77 _0608_ _0180_ _0287_ net31 sg13g2_a221oi_1
XFILLER_49_39 VPWR VGND sg13g2_decap_8
XFILLER_26_354 VPWR VGND sg13g2_decap_8
XFILLER_42_858 VPWR VGND sg13g2_fill_1
XFILLER_41_357 VPWR VGND sg13g2_decap_8
XFILLER_14_53 VPWR VGND sg13g2_decap_8
XFILLER_6_726 VPWR VGND sg13g2_decap_8
XFILLER_6_748 VPWR VGND sg13g2_decap_8
XFILLER_6_737 VPWR VGND sg13g2_fill_2
XFILLER_5_214 VPWR VGND sg13g2_decap_8
XFILLER_30_74 VPWR VGND sg13g2_decap_8
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_7_1025 VPWR VGND sg13g2_decap_4
XFILLER_49_424 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_17_343 VPWR VGND sg13g2_decap_8
XFILLER_18_855 VPWR VGND sg13g2_fill_1
XFILLER_45_663 VPWR VGND sg13g2_decap_8
XFILLER_44_140 VPWR VGND sg13g2_decap_8
XFILLER_45_674 VPWR VGND sg13g2_fill_1
XFILLER_32_368 VPWR VGND sg13g2_decap_8
XFILLER_9_575 VPWR VGND sg13g2_fill_2
X_1523_ VPWR _0163_ daisychain\[16\] VGND sg13g2_inv_1
X_1454_ VPWR _0239_ daisychain\[85\] VGND sg13g2_inv_1
XFILLER_4_291 VPWR VGND sg13g2_decap_8
X_2503__479 VPWR VGND net478 sg13g2_tiehi
X_1385_ VPWR _0046_ state\[26\] VGND sg13g2_inv_1
XFILLER_49_991 VPWR VGND sg13g2_decap_8
XFILLER_48_490 VPWR VGND sg13g2_decap_8
X_2006_ net215 VPWR _0862_ VGND state\[116\] net182 sg13g2_o21ai_1
XFILLER_35_140 VPWR VGND sg13g2_decap_8
XFILLER_11_508 VPWR VGND sg13g2_decap_8
XFILLER_23_368 VPWR VGND sg13g2_decap_8
X_2839_ daisychain\[121\] net17 VPWR VGND sg13g2_buf_1
XFILLER_2_228 VPWR VGND sg13g2_decap_8
XFILLER_46_427 VPWR VGND sg13g2_decap_8
XFILLER_26_151 VPWR VGND sg13g2_decap_8
XFILLER_42_633 VPWR VGND sg13g2_decap_8
XFILLER_14_368 VPWR VGND sg13g2_decap_8
XFILLER_41_154 VPWR VGND sg13g2_decap_8
XFILLER_30_817 VPWR VGND sg13g2_decap_8
XFILLER_25_74 VPWR VGND sg13g2_decap_8
XFILLER_6_501 VPWR VGND sg13g2_decap_8
X_2311__482 VPWR VGND net481 sg13g2_tiehi
XFILLER_41_84 VPWR VGND sg13g2_decap_8
XFILLER_6_578 VPWR VGND sg13g2_decap_8
XFILLER_2_784 VPWR VGND sg13g2_decap_8
XFILLER_49_221 VPWR VGND sg13g2_decap_8
XFILLER_1_294 VPWR VGND sg13g2_decap_8
XFILLER_2_67 VPWR VGND sg13g2_decap_8
XFILLER_49_298 VPWR VGND sg13g2_decap_8
XFILLER_37_427 VPWR VGND sg13g2_decap_8
XFILLER_46_950 VPWR VGND sg13g2_fill_2
XFILLER_17_140 VPWR VGND sg13g2_decap_8
XFILLER_46_994 VPWR VGND sg13g2_decap_4
XFILLER_33_655 VPWR VGND sg13g2_fill_1
XFILLER_32_165 VPWR VGND sg13g2_decap_8
XFILLER_21_817 VPWR VGND sg13g2_decap_4
XFILLER_20_305 VPWR VGND sg13g2_decap_8
XANTENNA_17 VPWR VGND daisychain\[27\] sg13g2_antennanp
XANTENNA_28 VPWR VGND _0179_ sg13g2_antennanp
XANTENNA_39 VPWR VGND _0253_ sg13g2_antennanp
XFILLER_9_361 VPWR VGND sg13g2_decap_8
X_2555_ net338 VGND VPWR _0501_ state\[117\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2362__380 VPWR VGND net379 sg13g2_tiehi
X_2486_ net292 VGND VPWR _0432_ state\[48\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1506_ VPWR _0182_ daisychain\[33\] VGND sg13g2_inv_1
X_1437_ VPWR _0131_ daisychain\[102\] VGND sg13g2_inv_1
X_1368_ VPWR _0065_ state\[43\] VGND sg13g2_inv_1
XFILLER_29_917 VPWR VGND sg13g2_decap_4
X_2393__318 VPWR VGND net317 sg13g2_tiehi
XFILLER_28_449 VPWR VGND sg13g2_decap_4
X_2438__484 VPWR VGND net483 sg13g2_tiehi
X_1299_ VPWR _0014_ state\[112\] VGND sg13g2_inv_1
XFILLER_11_305 VPWR VGND sg13g2_decap_8
XFILLER_24_666 VPWR VGND sg13g2_fill_1
XFILLER_23_165 VPWR VGND sg13g2_decap_8
XFILLER_11_32 VPWR VGND sg13g2_decap_8
XFILLER_3_559 VPWR VGND sg13g2_decap_8
XFILLER_47_703 VPWR VGND sg13g2_fill_1
XFILLER_46_224 VPWR VGND sg13g2_decap_8
XFILLER_19_427 VPWR VGND sg13g2_decap_4
XFILLER_15_600 VPWR VGND sg13g2_decap_4
XFILLER_36_84 VPWR VGND sg13g2_decap_8
XFILLER_15_677 VPWR VGND sg13g2_fill_1
XFILLER_14_165 VPWR VGND sg13g2_decap_8
XFILLER_7_832 VPWR VGND sg13g2_decap_8
XFILLER_10_382 VPWR VGND sg13g2_decap_8
XFILLER_7_876 VPWR VGND sg13g2_decap_4
XFILLER_7_898 VPWR VGND sg13g2_decap_8
XFILLER_6_375 VPWR VGND sg13g2_decap_8
X_2340_ net423 VGND VPWR _0286_ daisychain\[30\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2271_ VGND VPWR _0839_ _1006_ _0492_ net86 sg13g2_a21oi_1
XFILLER_2_592 VPWR VGND sg13g2_decap_8
XFILLER_28_4 VPWR VGND sg13g2_decap_8
XFILLER_37_224 VPWR VGND sg13g2_decap_8
XFILLER_19_994 VPWR VGND sg13g2_fill_1
XFILLER_46_791 VPWR VGND sg13g2_decap_8
XFILLER_21_636 VPWR VGND sg13g2_decap_8
XFILLER_20_102 VPWR VGND sg13g2_decap_8
X_1986_ net213 VPWR _0847_ VGND state\[111\] net170 sg13g2_o21ai_1
XFILLER_20_179 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_9_clk clknet_2_3__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
XFILLER_0_518 VPWR VGND sg13g2_decap_8
X_2538_ net426 VGND VPWR _0484_ state\[100\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2469_ net360 VGND VPWR _0415_ state\[31\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_28_235 VPWR VGND sg13g2_decap_8
XFILLER_44_717 VPWR VGND sg13g2_decap_4
XFILLER_43_238 VPWR VGND sg13g2_decap_8
XFILLER_11_102 VPWR VGND sg13g2_decap_8
XFILLER_11_179 VPWR VGND sg13g2_decap_8
XFILLER_22_53 VPWR VGND sg13g2_decap_8
XFILLER_3_312 VPWR VGND sg13g2_decap_8
XFILLER_4_868 VPWR VGND sg13g2_fill_2
XFILLER_4_857 VPWR VGND sg13g2_decap_8
XFILLER_4_846 VPWR VGND sg13g2_decap_4
XFILLER_3_389 VPWR VGND sg13g2_decap_8
XFILLER_26_1007 VPWR VGND sg13g2_fill_1
Xfanout192 net193 net192 VPWR VGND sg13g2_buf_1
Xfanout181 net182 net181 VPWR VGND sg13g2_buf_1
Xfanout170 net172 net170 VPWR VGND sg13g2_buf_1
XFILLER_19_235 VPWR VGND sg13g2_decap_8
XFILLER_35_706 VPWR VGND sg13g2_fill_2
XFILLER_34_249 VPWR VGND sg13g2_decap_8
XFILLER_15_452 VPWR VGND sg13g2_decap_4
XFILLER_15_496 VPWR VGND sg13g2_decap_4
X_1840_ VGND VPWR net154 daisychain\[73\] _0738_ net62 sg13g2_a21oi_1
XFILLER_8_11 VPWR VGND sg13g2_decap_8
XFILLER_30_444 VPWR VGND sg13g2_decap_8
X_1771_ net191 _0208_ _0685_ _0686_ VPWR VGND sg13g2_a21o_1
XFILLER_8_88 VPWR VGND sg13g2_decap_8
X_2463__385 VPWR VGND net384 sg13g2_tiehi
XFILLER_6_172 VPWR VGND sg13g2_decap_8
X_2323_ net457 VGND VPWR _0269_ daisychain\[13\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2254_ _0998_ net133 state\[100\] VPWR VGND sg13g2_nand2_1
X_2185_ VGND VPWR _0710_ _0963_ _0449_ net107 sg13g2_a21oi_1
XFILLER_26_728 VPWR VGND sg13g2_decap_8
XFILLER_25_249 VPWR VGND sg13g2_decap_8
XFILLER_41_709 VPWR VGND sg13g2_decap_8
X_1969_ VPWR VGND _0834_ net87 _0833_ _0135_ _0362_ net45 sg13g2_a221oi_1
XFILLER_4_109 VPWR VGND sg13g2_decap_8
X_2442__469 VPWR VGND net468 sg13g2_tiehi
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_17_42 VPWR VGND sg13g2_decap_8
XFILLER_16_249 VPWR VGND sg13g2_decap_8
XFILLER_12_444 VPWR VGND sg13g2_decap_8
XFILLER_33_74 VPWR VGND sg13g2_decap_8
XFILLER_4_665 VPWR VGND sg13g2_decap_8
XFILLER_3_186 VPWR VGND sg13g2_decap_8
XFILLER_39_308 VPWR VGND sg13g2_decap_8
XFILLER_47_385 VPWR VGND sg13g2_decap_8
XFILLER_35_547 VPWR VGND sg13g2_fill_1
XFILLER_31_764 VPWR VGND sg13g2_fill_2
XFILLER_30_263 VPWR VGND sg13g2_decap_8
X_1823_ net201 _0223_ _0724_ _0725_ VPWR VGND sg13g2_a21o_1
X_1754_ net221 VPWR _0673_ VGND state\[53\] net189 sg13g2_o21ai_1
XFILLER_8_993 VPWR VGND sg13g2_fill_2
XFILLER_8_960 VPWR VGND sg13g2_fill_1
X_1685_ VPWR VGND _0621_ net92 _0620_ _0184_ _0291_ net52 sg13g2_a221oi_1
X_2506__455 VPWR VGND net454 sg13g2_tiehi
X_2541__379 VPWR VGND net378 sg13g2_tiehi
X_2498__245 VPWR VGND net244 sg13g2_tiehi
X_2306_ _1024_ net113 state\[126\] VPWR VGND sg13g2_nand2_1
X_2237_ VGND VPWR _0788_ _0989_ _0475_ net103 sg13g2_a21oi_1
X_2168_ _0955_ net143 state\[57\] VPWR VGND sg13g2_nand2_1
XFILLER_38_385 VPWR VGND sg13g2_decap_8
X_2099_ VGND VPWR _0581_ _0920_ _0406_ net102 sg13g2_a21oi_1
XFILLER_22_775 VPWR VGND sg13g2_fill_1
XFILLER_21_263 VPWR VGND sg13g2_decap_8
XFILLER_1_602 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
X_2477__329 VPWR VGND net328 sg13g2_tiehi
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_1_679 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
X_2518__359 VPWR VGND net358 sg13g2_tiehi
XFILLER_28_74 VPWR VGND sg13g2_decap_8
XFILLER_45_823 VPWR VGND sg13g2_fill_2
XFILLER_44_322 VPWR VGND sg13g2_decap_8
XFILLER_29_396 VPWR VGND sg13g2_decap_8
XFILLER_44_399 VPWR VGND sg13g2_decap_8
XFILLER_9_702 VPWR VGND sg13g2_fill_1
XFILLER_44_84 VPWR VGND sg13g2_decap_8
XFILLER_12_263 VPWR VGND sg13g2_decap_8
XFILLER_40_594 VPWR VGND sg13g2_fill_2
XFILLER_8_256 VPWR VGND sg13g2_decap_8
X_1470_ VPWR _0221_ daisychain\[69\] VGND sg13g2_inv_1
XFILLER_5_67 VPWR VGND sg13g2_decap_8
XFILLER_39_105 VPWR VGND sg13g2_decap_8
X_2321__462 VPWR VGND net461 sg13g2_tiehi
XFILLER_10_4 VPWR VGND sg13g2_decap_8
X_2022_ net217 VPWR _0874_ VGND state\[120\] net174 sg13g2_o21ai_1
X_2536__459 VPWR VGND net458 sg13g2_tiehi
XFILLER_47_182 VPWR VGND sg13g2_decap_8
XFILLER_35_322 VPWR VGND sg13g2_decap_8
XFILLER_35_399 VPWR VGND sg13g2_decap_8
XFILLER_16_591 VPWR VGND sg13g2_fill_1
X_1806_ net225 VPWR _0712_ VGND state\[66\] net200 sg13g2_o21ai_1
X_1737_ VPWR VGND _0660_ net106 _0659_ _0198_ _0304_ net62 sg13g2_a221oi_1
X_1668_ VGND VPWR net120 daisychain\[30\] _0609_ net31 sg13g2_a21oi_1
XFILLER_49_18 VPWR VGND sg13g2_decap_8
X_1599_ net162 _0161_ _0556_ _0557_ VPWR VGND sg13g2_a21o_1
XFILLER_45_119 VPWR VGND sg13g2_decap_8
XFILLER_38_182 VPWR VGND sg13g2_decap_8
XFILLER_27_878 VPWR VGND sg13g2_decap_8
XFILLER_26_333 VPWR VGND sg13g2_decap_8
X_2372__360 VPWR VGND net359 sg13g2_tiehi
XFILLER_42_815 VPWR VGND sg13g2_decap_8
XFILLER_41_336 VPWR VGND sg13g2_decap_8
XFILLER_14_32 VPWR VGND sg13g2_decap_8
XFILLER_22_550 VPWR VGND sg13g2_fill_2
XFILLER_30_53 VPWR VGND sg13g2_decap_8
XFILLER_49_403 VPWR VGND sg13g2_decap_8
XFILLER_2_988 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
XFILLER_39_84 VPWR VGND sg13g2_decap_8
XFILLER_18_801 VPWR VGND sg13g2_fill_1
XFILLER_17_322 VPWR VGND sg13g2_decap_8
XFILLER_18_834 VPWR VGND sg13g2_fill_1
XFILLER_36_119 VPWR VGND sg13g2_decap_8
XFILLER_29_193 VPWR VGND sg13g2_decap_8
XFILLER_17_399 VPWR VGND sg13g2_decap_8
XFILLER_44_196 VPWR VGND sg13g2_decap_8
XFILLER_32_347 VPWR VGND sg13g2_decap_8
XFILLER_20_509 VPWR VGND sg13g2_fill_2
XFILLER_13_594 VPWR VGND sg13g2_fill_1
XFILLER_9_543 VPWR VGND sg13g2_decap_8
X_1522_ VPWR _0164_ daisychain\[17\] VGND sg13g2_inv_1
X_1453_ VPWR _0240_ daisychain\[86\] VGND sg13g2_inv_1
XFILLER_4_270 VPWR VGND sg13g2_decap_8
X_1384_ VPWR _0047_ state\[27\] VGND sg13g2_inv_1
XFILLER_28_609 VPWR VGND sg13g2_fill_2
XFILLER_27_119 VPWR VGND sg13g2_decap_8
X_2005_ VPWR VGND _0861_ net87 _0860_ _0145_ _0371_ net44 sg13g2_a221oi_1
XFILLER_35_196 VPWR VGND sg13g2_decap_8
XFILLER_23_347 VPWR VGND sg13g2_decap_8
X_2838_ daisychain\[120\] net16 VPWR VGND sg13g2_buf_1
XFILLER_2_207 VPWR VGND sg13g2_decap_8
XFILLER_46_406 VPWR VGND sg13g2_decap_8
XFILLER_39_491 VPWR VGND sg13g2_decap_4
XFILLER_26_130 VPWR VGND sg13g2_decap_8
XFILLER_27_664 VPWR VGND sg13g2_decap_8
XFILLER_14_347 VPWR VGND sg13g2_decap_8
XFILLER_25_53 VPWR VGND sg13g2_decap_8
XFILLER_41_133 VPWR VGND sg13g2_decap_8
XFILLER_41_63 VPWR VGND sg13g2_decap_8
XFILLER_6_557 VPWR VGND sg13g2_decap_8
XFILLER_2_774 VPWR VGND sg13g2_decap_4
XFILLER_49_200 VPWR VGND sg13g2_decap_8
XFILLER_1_273 VPWR VGND sg13g2_decap_8
XFILLER_37_406 VPWR VGND sg13g2_decap_8
XFILLER_2_46 VPWR VGND sg13g2_decap_8
XFILLER_49_277 VPWR VGND sg13g2_decap_8
XFILLER_18_686 VPWR VGND sg13g2_fill_1
XFILLER_17_196 VPWR VGND sg13g2_decap_8
XFILLER_33_667 VPWR VGND sg13g2_fill_2
XFILLER_32_144 VPWR VGND sg13g2_decap_8
XANTENNA_18 VPWR VGND daisychain\[27\] sg13g2_antennanp
XANTENNA_29 VPWR VGND _0190_ sg13g2_antennanp
XFILLER_9_340 VPWR VGND sg13g2_decap_8
X_2554_ net370 VGND VPWR _0500_ state\[116\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_1505_ VPWR _0183_ daisychain\[34\] VGND sg13g2_inv_1
XFILLER_5_590 VPWR VGND sg13g2_decap_8
X_2485_ net296 VGND VPWR _0431_ state\[47\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1436_ VPWR _0132_ daisychain\[103\] VGND sg13g2_inv_1
X_1367_ VPWR _0066_ state\[44\] VGND sg13g2_inv_1
XFILLER_28_417 VPWR VGND sg13g2_decap_8
X_1298_ VPWR _0015_ state\[113\] VGND sg13g2_inv_1
XFILLER_36_472 VPWR VGND sg13g2_decap_8
XFILLER_23_144 VPWR VGND sg13g2_decap_8
XFILLER_11_11 VPWR VGND sg13g2_decap_8
XFILLER_11_88 VPWR VGND sg13g2_decap_8
XFILLER_3_538 VPWR VGND sg13g2_decap_8
XFILLER_46_203 VPWR VGND sg13g2_decap_8
XFILLER_47_759 VPWR VGND sg13g2_fill_2
XFILLER_36_63 VPWR VGND sg13g2_decap_8
XFILLER_28_995 VPWR VGND sg13g2_decap_8
XFILLER_28_973 VPWR VGND sg13g2_decap_8
XFILLER_27_450 VPWR VGND sg13g2_fill_1
XFILLER_15_623 VPWR VGND sg13g2_fill_2
XFILLER_42_420 VPWR VGND sg13g2_fill_1
XFILLER_27_483 VPWR VGND sg13g2_decap_8
XFILLER_14_144 VPWR VGND sg13g2_decap_8
XFILLER_30_648 VPWR VGND sg13g2_fill_1
XFILLER_10_361 VPWR VGND sg13g2_decap_8
XFILLER_7_855 VPWR VGND sg13g2_decap_8
XFILLER_6_354 VPWR VGND sg13g2_decap_8
XFILLER_42_7 VPWR VGND sg13g2_decap_8
X_2270_ _1006_ net130 state\[108\] VPWR VGND sg13g2_nand2_1
XFILLER_2_571 VPWR VGND sg13g2_decap_8
XFILLER_38_737 VPWR VGND sg13g2_fill_2
XFILLER_37_203 VPWR VGND sg13g2_decap_8
XFILLER_18_483 VPWR VGND sg13g2_decap_8
XFILLER_45_280 VPWR VGND sg13g2_decap_8
X_1985_ VPWR VGND _0846_ net84 _0845_ _0140_ _0366_ net43 sg13g2_a221oi_1
XFILLER_20_158 VPWR VGND sg13g2_decap_8
X_2509__431 VPWR VGND net430 sg13g2_tiehi
X_2537_ net442 VGND VPWR _0483_ state\[99\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2468_ net364 VGND VPWR _0414_ state\[30\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_1419_ VPWR _0151_ daisychain\[120\] VGND sg13g2_inv_1
X_2399_ net305 VGND VPWR _0345_ daisychain\[89\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_28_214 VPWR VGND sg13g2_decap_8
XFILLER_43_217 VPWR VGND sg13g2_decap_8
XFILLER_36_280 VPWR VGND sg13g2_decap_8
XFILLER_25_976 VPWR VGND sg13g2_fill_2
XFILLER_24_453 VPWR VGND sg13g2_fill_1
XFILLER_24_431 VPWR VGND sg13g2_fill_2
XFILLER_12_615 VPWR VGND sg13g2_fill_2
XFILLER_12_626 VPWR VGND sg13g2_decap_8
XFILLER_24_497 VPWR VGND sg13g2_fill_1
XFILLER_24_486 VPWR VGND sg13g2_decap_8
XFILLER_11_158 VPWR VGND sg13g2_decap_8
XFILLER_22_32 VPWR VGND sg13g2_decap_8
XFILLER_3_368 VPWR VGND sg13g2_decap_8
XFILLER_19_214 VPWR VGND sg13g2_decap_8
Xfanout182 net183 net182 VPWR VGND sg13g2_buf_1
Xfanout171 net172 net171 VPWR VGND sg13g2_buf_1
Xfanout160 net161 net160 VPWR VGND sg13g2_buf_1
XFILLER_47_523 VPWR VGND sg13g2_fill_2
Xfanout193 net204 net193 VPWR VGND sg13g2_buf_1
XFILLER_47_84 VPWR VGND sg13g2_decap_8
X_2491__273 VPWR VGND net272 sg13g2_tiehi
XFILLER_34_228 VPWR VGND sg13g2_decap_8
XFILLER_27_280 VPWR VGND sg13g2_decap_8
XFILLER_15_431 VPWR VGND sg13g2_decap_8
XFILLER_43_784 VPWR VGND sg13g2_decap_4
XFILLER_42_294 VPWR VGND sg13g2_decap_8
XFILLER_31_957 VPWR VGND sg13g2_fill_2
X_1770_ net221 VPWR _0685_ VGND state\[57\] net188 sg13g2_o21ai_1
XFILLER_8_67 VPWR VGND sg13g2_decap_8
XFILLER_6_151 VPWR VGND sg13g2_decap_8
X_2322_ net459 VGND VPWR _0268_ daisychain\[12\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_2253_ VGND VPWR _0812_ _0997_ _0483_ net86 sg13g2_a21oi_1
X_2184_ _0963_ net153 state\[65\] VPWR VGND sg13g2_nand2_1
XFILLER_25_228 VPWR VGND sg13g2_decap_8
XFILLER_19_792 VPWR VGND sg13g2_decap_8
XFILLER_18_291 VPWR VGND sg13g2_decap_8
X_2470__357 VPWR VGND net356 sg13g2_tiehi
X_2331__442 VPWR VGND net441 sg13g2_tiehi
XFILLER_21_445 VPWR VGND sg13g2_fill_2
X_1968_ VGND VPWR net131 daisychain\[105\] _0834_ net45 sg13g2_a21oi_1
X_1899_ net178 _0243_ _0781_ _0782_ VPWR VGND sg13g2_a21o_1
XFILLER_17_21 VPWR VGND sg13g2_decap_8
XFILLER_17_718 VPWR VGND sg13g2_decap_8
XFILLER_44_515 VPWR VGND sg13g2_fill_2
XFILLER_16_228 VPWR VGND sg13g2_decap_8
XFILLER_17_98 VPWR VGND sg13g2_decap_8
XFILLER_12_423 VPWR VGND sg13g2_decap_8
XFILLER_40_732 VPWR VGND sg13g2_fill_2
XFILLER_33_53 VPWR VGND sg13g2_decap_8
XFILLER_32_1001 VPWR VGND sg13g2_fill_1
XFILLER_8_438 VPWR VGND sg13g2_decap_4
X_2382__340 VPWR VGND net339 sg13g2_tiehi
XFILLER_3_165 VPWR VGND sg13g2_decap_8
XFILLER_47_364 VPWR VGND sg13g2_decap_8
X_1822_ net226 VPWR _0724_ VGND state\[70\] net201 sg13g2_o21ai_1
XFILLER_30_242 VPWR VGND sg13g2_decap_8
X_1753_ VPWR VGND _0672_ net99 _0671_ _0203_ _0308_ net55 sg13g2_a221oi_1
XFILLER_8_972 VPWR VGND sg13g2_fill_2
X_1684_ VGND VPWR net116 daisychain\[34\] _0621_ net28 sg13g2_a21oi_1
X_2305_ VGND VPWR _0890_ _1023_ _0509_ net69 sg13g2_a21oi_1
X_2236_ _0989_ net149 state\[91\] VPWR VGND sg13g2_nand2_1
X_2359__386 VPWR VGND net385 sg13g2_tiehi
XFILLER_38_364 VPWR VGND sg13g2_decap_8
XFILLER_26_504 VPWR VGND sg13g2_decap_8
X_2167_ VGND VPWR _0683_ _0954_ _0440_ net98 sg13g2_a21oi_1
X_2098_ _0920_ net148 state\[22\] VPWR VGND sg13g2_nand2_1
XFILLER_21_242 VPWR VGND sg13g2_decap_8
XFILLER_1_658 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_28_53 VPWR VGND sg13g2_decap_8
XFILLER_45_846 VPWR VGND sg13g2_decap_4
XFILLER_44_301 VPWR VGND sg13g2_decap_8
XFILLER_29_375 VPWR VGND sg13g2_decap_8
XFILLER_17_559 VPWR VGND sg13g2_fill_1
XFILLER_45_879 VPWR VGND sg13g2_fill_1
XFILLER_45_868 VPWR VGND sg13g2_decap_8
XFILLER_44_378 VPWR VGND sg13g2_decap_8
XFILLER_44_63 VPWR VGND sg13g2_decap_8
XFILLER_12_242 VPWR VGND sg13g2_decap_8
XFILLER_9_725 VPWR VGND sg13g2_decap_8
XFILLER_40_551 VPWR VGND sg13g2_decap_8
XFILLER_8_235 VPWR VGND sg13g2_decap_8
XFILLER_5_931 VPWR VGND sg13g2_fill_2
XFILLER_5_46 VPWR VGND sg13g2_decap_8
XFILLER_4_452 VPWR VGND sg13g2_decap_8
X_2021_ VPWR VGND _0873_ net82 _0872_ _0149_ _0375_ net37 sg13g2_a221oi_1
XFILLER_47_161 VPWR VGND sg13g2_decap_8
XFILLER_35_301 VPWR VGND sg13g2_decap_8
XFILLER_35_378 VPWR VGND sg13g2_decap_8
XFILLER_23_507 VPWR VGND sg13g2_decap_8
XFILLER_31_562 VPWR VGND sg13g2_fill_1
X_1805_ VPWR VGND _0711_ net107 _0710_ _0217_ _0321_ net63 sg13g2_a221oi_1
X_1736_ VGND VPWR net154 daisychain\[47\] _0660_ net62 sg13g2_a21oi_1
X_1667_ net163 _0180_ _0607_ _0608_ VPWR VGND sg13g2_a21o_1
X_1598_ net206 VPWR _0556_ VGND state\[14\] net162 sg13g2_o21ai_1
X_2219_ VGND VPWR _0761_ _0980_ _0466_ net79 sg13g2_a21oi_1
XFILLER_38_161 VPWR VGND sg13g2_decap_8
XFILLER_26_312 VPWR VGND sg13g2_decap_8
XFILLER_41_315 VPWR VGND sg13g2_decap_8
XFILLER_26_389 VPWR VGND sg13g2_decap_8
XFILLER_14_11 VPWR VGND sg13g2_decap_8
XFILLER_22_573 VPWR VGND sg13g2_decap_8
XFILLER_14_88 VPWR VGND sg13g2_decap_8
XFILLER_30_32 VPWR VGND sg13g2_decap_8
XFILLER_5_249 VPWR VGND sg13g2_decap_8
XFILLER_2_912 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_39_63 VPWR VGND sg13g2_decap_8
XFILLER_49_459 VPWR VGND sg13g2_decap_8
XFILLER_17_301 VPWR VGND sg13g2_decap_8
XFILLER_18_813 VPWR VGND sg13g2_fill_1
XFILLER_29_172 VPWR VGND sg13g2_decap_8
XFILLER_17_378 VPWR VGND sg13g2_decap_8
XFILLER_44_175 VPWR VGND sg13g2_decap_8
XFILLER_32_326 VPWR VGND sg13g2_decap_8
XFILLER_26_890 VPWR VGND sg13g2_decap_4
XFILLER_9_522 VPWR VGND sg13g2_decap_8
XFILLER_9_577 VPWR VGND sg13g2_fill_1
XFILLER_40_392 VPWR VGND sg13g2_decap_8
X_1521_ VPWR _0165_ daisychain\[18\] VGND sg13g2_inv_1
XFILLER_5_772 VPWR VGND sg13g2_fill_2
XFILLER_5_761 VPWR VGND sg13g2_decap_8
X_1452_ VPWR _0241_ daisychain\[87\] VGND sg13g2_inv_1
XFILLER_45_1022 VPWR VGND sg13g2_decap_8
X_1383_ VPWR _0048_ state\[28\] VGND sg13g2_inv_1
X_2004_ VGND VPWR net131 daisychain\[114\] _0861_ net37 sg13g2_a21oi_1
XFILLER_36_676 VPWR VGND sg13g2_fill_2
XFILLER_35_175 VPWR VGND sg13g2_decap_8
XFILLER_23_326 VPWR VGND sg13g2_decap_8
X_2837_ state\[127\] net15 VPWR VGND sg13g2_buf_1
X_1719_ net185 _0194_ _0646_ _0647_ VPWR VGND sg13g2_a21o_1
XFILLER_47_908 VPWR VGND sg13g2_fill_2
XFILLER_18_109 VPWR VGND sg13g2_decap_8
XFILLER_14_326 VPWR VGND sg13g2_decap_8
XFILLER_41_112 VPWR VGND sg13g2_decap_8
XFILLER_26_186 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_decap_8
XFILLER_41_189 VPWR VGND sg13g2_decap_8
XFILLER_10_543 VPWR VGND sg13g2_decap_8
XFILLER_6_536 VPWR VGND sg13g2_decap_8
XFILLER_41_42 VPWR VGND sg13g2_decap_8
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_1_252 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_49_256 VPWR VGND sg13g2_decap_8
XFILLER_18_654 VPWR VGND sg13g2_decap_4
XFILLER_33_613 VPWR VGND sg13g2_fill_2
XFILLER_17_175 VPWR VGND sg13g2_decap_8
XFILLER_32_123 VPWR VGND sg13g2_decap_8
XANTENNA_19 VPWR VGND daisychain\[9\] sg13g2_antennanp
X_2466__373 VPWR VGND net372 sg13g2_tiehi
XFILLER_9_396 VPWR VGND sg13g2_decap_8
X_2553_ net402 VGND VPWR _0499_ state\[115\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_1504_ VPWR _0184_ daisychain\[35\] VGND sg13g2_inv_1
X_2484_ net300 VGND VPWR _0430_ state\[46\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1435_ VPWR _0133_ daisychain\[104\] VGND sg13g2_inv_1
X_1366_ VPWR _0067_ state\[45\] VGND sg13g2_inv_1
X_1297_ VPWR _0016_ state\[114\] VGND sg13g2_inv_1
XFILLER_36_451 VPWR VGND sg13g2_decap_8
XFILLER_23_123 VPWR VGND sg13g2_decap_8
XFILLER_20_841 VPWR VGND sg13g2_decap_4
XFILLER_11_67 VPWR VGND sg13g2_decap_8
X_2445__457 VPWR VGND net456 sg13g2_tiehi
XFILLER_3_517 VPWR VGND sg13g2_decap_8
X_2341__422 VPWR VGND net421 sg13g2_tiehi
XFILLER_46_259 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_decap_8
XFILLER_14_123 VPWR VGND sg13g2_decap_8
XFILLER_15_668 VPWR VGND sg13g2_decap_8
XFILLER_42_443 VPWR VGND sg13g2_decap_8
XFILLER_23_690 VPWR VGND sg13g2_fill_2
XFILLER_10_340 VPWR VGND sg13g2_decap_8
XFILLER_6_333 VPWR VGND sg13g2_decap_8
XFILLER_2_550 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_decap_8
X_2392__320 VPWR VGND net319 sg13g2_tiehi
XFILLER_37_259 VPWR VGND sg13g2_decap_8
X_2318__468 VPWR VGND net467 sg13g2_tiehi
XFILLER_33_410 VPWR VGND sg13g2_decap_8
X_1984_ VGND VPWR net128 daisychain\[109\] _0846_ net43 sg13g2_a21oi_1
XFILLER_20_137 VPWR VGND sg13g2_decap_8
XFILLER_9_193 VPWR VGND sg13g2_decap_8
X_2536_ net458 VGND VPWR _0482_ state\[98\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2467_ net368 VGND VPWR _0413_ state\[29\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_1418_ VPWR _0152_ daisychain\[121\] VGND sg13g2_inv_1
X_2398_ net307 VGND VPWR _0344_ daisychain\[88\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_29_705 VPWR VGND sg13g2_decap_4
X_1349_ VPWR _0086_ state\[62\] VGND sg13g2_inv_1
XFILLER_24_410 VPWR VGND sg13g2_decap_8
XFILLER_25_988 VPWR VGND sg13g2_decap_8
XFILLER_11_137 VPWR VGND sg13g2_decap_8
XdigitalenH.g\[2\].u.inv1 VPWR digitalenH.g\[2\].u.OUTN net7 VGND sg13g2_inv_1
XFILLER_8_609 VPWR VGND sg13g2_fill_2
XFILLER_7_119 VPWR VGND sg13g2_decap_8
XFILLER_22_11 VPWR VGND sg13g2_decap_8
X_2369__366 VPWR VGND net365 sg13g2_tiehi
XFILLER_22_88 VPWR VGND sg13g2_decap_8
XFILLER_3_347 VPWR VGND sg13g2_decap_8
Xfanout183 net204 net183 VPWR VGND sg13g2_buf_1
Xfanout172 net183 net172 VPWR VGND sg13g2_buf_1
Xfanout161 net169 net161 VPWR VGND sg13g2_buf_1
Xfanout150 net152 net150 VPWR VGND sg13g2_buf_1
Xfanout194 net195 net194 VPWR VGND sg13g2_buf_1
XFILLER_47_63 VPWR VGND sg13g2_decap_8
XFILLER_34_207 VPWR VGND sg13g2_decap_8
XFILLER_15_410 VPWR VGND sg13g2_decap_8
XFILLER_42_273 VPWR VGND sg13g2_decap_8
XFILLER_8_46 VPWR VGND sg13g2_decap_8
XFILLER_6_130 VPWR VGND sg13g2_decap_8
X_2321_ net461 VGND VPWR _0267_ daisychain\[11\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2252_ _0997_ net130 state\[99\] VPWR VGND sg13g2_nand2_1
X_2500__237 VPWR VGND net236 sg13g2_tiehi
XFILLER_33_4 VPWR VGND sg13g2_decap_8
X_2183_ VGND VPWR _0707_ _0962_ _0448_ net107 sg13g2_a21oi_1
XFILLER_18_270 VPWR VGND sg13g2_decap_8
XFILLER_25_207 VPWR VGND sg13g2_decap_8
XFILLER_22_925 VPWR VGND sg13g2_fill_1
XFILLER_33_284 VPWR VGND sg13g2_decap_8
XFILLER_22_958 VPWR VGND sg13g2_fill_1
XFILLER_21_424 VPWR VGND sg13g2_decap_8
XFILLER_21_468 VPWR VGND sg13g2_decap_8
X_1967_ net182 _0135_ _0832_ _0833_ VPWR VGND sg13g2_a21o_1
X_1898_ net214 VPWR _0781_ VGND state\[89\] net178 sg13g2_o21ai_1
X_2519_ net350 VGND VPWR _0465_ state\[81\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_29_579 VPWR VGND sg13g2_fill_2
XFILLER_16_207 VPWR VGND sg13g2_decap_8
XFILLER_17_77 VPWR VGND sg13g2_decap_8
XFILLER_33_32 VPWR VGND sg13g2_decap_8
XFILLER_24_284 VPWR VGND sg13g2_decap_8
XFILLER_12_479 VPWR VGND sg13g2_decap_8
XFILLER_8_417 VPWR VGND sg13g2_decap_8
XFILLER_32_1024 VPWR VGND sg13g2_decap_4
XFILLER_4_623 VPWR VGND sg13g2_decap_8
XFILLER_3_144 VPWR VGND sg13g2_decap_8
XFILLER_0_851 VPWR VGND sg13g2_fill_2
XFILLER_47_343 VPWR VGND sg13g2_decap_8
XFILLER_28_590 VPWR VGND sg13g2_fill_2
XFILLER_15_284 VPWR VGND sg13g2_decap_8
XFILLER_31_744 VPWR VGND sg13g2_fill_2
XFILLER_30_221 VPWR VGND sg13g2_decap_8
X_1821_ VPWR VGND _0723_ net109 _0722_ _0221_ _0325_ net66 sg13g2_a221oi_1
XFILLER_31_766 VPWR VGND sg13g2_fill_1
XFILLER_30_298 VPWR VGND sg13g2_decap_8
X_1752_ VGND VPWR net145 daisychain\[51\] _0672_ net55 sg13g2_a21oi_1
Xclkbuf_leaf_10_clk clknet_2_3__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
X_1683_ net184 _0184_ _0619_ _0620_ VPWR VGND sg13g2_a21o_1
XFILLER_7_483 VPWR VGND sg13g2_decap_8
X_2304_ _1023_ net113 state\[125\] VPWR VGND sg13g2_nand2_1
X_2235_ VGND VPWR _0785_ _0988_ _0474_ net103 sg13g2_a21oi_1
X_2166_ _0954_ net143 state\[56\] VPWR VGND sg13g2_nand2_1
XFILLER_38_343 VPWR VGND sg13g2_decap_8
X_2097_ VGND VPWR _0578_ _0919_ _0405_ net75 sg13g2_a21oi_1
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_21_221 VPWR VGND sg13g2_decap_8
XFILLER_21_298 VPWR VGND sg13g2_decap_8
XFILLER_1_637 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_28_32 VPWR VGND sg13g2_decap_8
XFILLER_29_354 VPWR VGND sg13g2_decap_8
XFILLER_45_825 VPWR VGND sg13g2_fill_1
XFILLER_44_357 VPWR VGND sg13g2_decap_8
XFILLER_44_42 VPWR VGND sg13g2_decap_8
XFILLER_12_221 VPWR VGND sg13g2_decap_8
XFILLER_40_530 VPWR VGND sg13g2_fill_2
XFILLER_8_214 VPWR VGND sg13g2_decap_8
XFILLER_12_298 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_decap_8
XFILLER_4_431 VPWR VGND sg13g2_decap_8
XFILLER_4_497 VPWR VGND sg13g2_decap_8
X_2020_ VGND VPWR net126 daisychain\[118\] _0873_ net37 sg13g2_a21oi_1
XFILLER_47_140 VPWR VGND sg13g2_decap_8
XFILLER_35_357 VPWR VGND sg13g2_decap_8
X_1804_ VGND VPWR net153 daisychain\[64\] _0711_ net63 sg13g2_a21oi_1
X_1735_ net192 _0198_ _0658_ _0659_ VPWR VGND sg13g2_a21o_1
XFILLER_7_280 VPWR VGND sg13g2_decap_8
X_1666_ net206 VPWR _0607_ VGND state\[31\] net162 sg13g2_o21ai_1
X_1597_ VPWR VGND _0555_ net92 _0554_ _0160_ _0269_ net52 sg13g2_a221oi_1
XFILLER_39_663 VPWR VGND sg13g2_fill_1
X_2218_ _0980_ net123 state\[82\] VPWR VGND sg13g2_nand2_1
XFILLER_38_140 VPWR VGND sg13g2_decap_8
X_2149_ VGND VPWR _0656_ _0945_ _0431_ net93 sg13g2_a21oi_1
XFILLER_14_508 VPWR VGND sg13g2_fill_1
XFILLER_26_368 VPWR VGND sg13g2_decap_8
XFILLER_22_552 VPWR VGND sg13g2_fill_1
XFILLER_14_67 VPWR VGND sg13g2_decap_8
XFILLER_5_228 VPWR VGND sg13g2_decap_8
XFILLER_30_11 VPWR VGND sg13g2_decap_8
XFILLER_30_88 VPWR VGND sg13g2_decap_8
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_39_42 VPWR VGND sg13g2_decap_8
XFILLER_49_438 VPWR VGND sg13g2_decap_8
XFILLER_29_151 VPWR VGND sg13g2_decap_8
XFILLER_18_847 VPWR VGND sg13g2_fill_1
XFILLER_17_357 VPWR VGND sg13g2_decap_8
X_2351__402 VPWR VGND net401 sg13g2_tiehi
XFILLER_44_154 VPWR VGND sg13g2_decap_8
XFILLER_32_305 VPWR VGND sg13g2_decap_8
XFILLER_13_530 VPWR VGND sg13g2_fill_1
XFILLER_9_501 VPWR VGND sg13g2_decap_8
XFILLER_40_371 VPWR VGND sg13g2_decap_8
X_1520_ VPWR _0166_ daisychain\[19\] VGND sg13g2_inv_1
X_1451_ VPWR _0242_ daisychain\[88\] VGND sg13g2_inv_1
X_1382_ VPWR _0049_ state\[29\] VGND sg13g2_inv_1
X_2003_ net179 _0145_ _0859_ _0860_ VPWR VGND sg13g2_a21o_1
XFILLER_36_655 VPWR VGND sg13g2_fill_1
XFILLER_36_622 VPWR VGND sg13g2_fill_2
XFILLER_35_154 VPWR VGND sg13g2_decap_8
XFILLER_23_305 VPWR VGND sg13g2_decap_8
XFILLER_24_839 VPWR VGND sg13g2_decap_8
X_2836_ state\[126\] net14 VPWR VGND sg13g2_buf_1
XFILLER_31_382 VPWR VGND sg13g2_decap_8
X_1718_ net218 VPWR _0646_ VGND state\[44\] net185 sg13g2_o21ai_1
X_2328__448 VPWR VGND net447 sg13g2_tiehi
X_1649_ VPWR VGND _0594_ net76 _0593_ _0174_ _0282_ net30 sg13g2_a221oi_1
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_14_305 VPWR VGND sg13g2_decap_8
XFILLER_26_165 VPWR VGND sg13g2_decap_8
XFILLER_25_88 VPWR VGND sg13g2_decap_8
XFILLER_41_168 VPWR VGND sg13g2_decap_8
XFILLER_10_522 VPWR VGND sg13g2_decap_8
XFILLER_41_21 VPWR VGND sg13g2_decap_8
XFILLER_22_382 VPWR VGND sg13g2_decap_8
XFILLER_6_515 VPWR VGND sg13g2_decap_8
XFILLER_41_98 VPWR VGND sg13g2_decap_8
XFILLER_2_721 VPWR VGND sg13g2_decap_8
XFILLER_1_231 VPWR VGND sg13g2_decap_8
X_2379__346 VPWR VGND net345 sg13g2_tiehi
XFILLER_49_235 VPWR VGND sg13g2_decap_8
XFILLER_18_611 VPWR VGND sg13g2_decap_8
X_2494__261 VPWR VGND net260 sg13g2_tiehi
XFILLER_17_154 VPWR VGND sg13g2_decap_8
XFILLER_45_441 VPWR VGND sg13g2_decap_8
XFILLER_32_102 VPWR VGND sg13g2_decap_8
XFILLER_33_669 VPWR VGND sg13g2_fill_1
XFILLER_32_179 VPWR VGND sg13g2_decap_8
XFILLER_20_319 VPWR VGND sg13g2_decap_8
XFILLER_13_382 VPWR VGND sg13g2_decap_8
XFILLER_41_680 VPWR VGND sg13g2_fill_1
XFILLER_9_375 VPWR VGND sg13g2_decap_8
X_2552_ net434 VGND VPWR _0498_ state\[114\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_1503_ VPWR _0185_ daisychain\[36\] VGND sg13g2_inv_1
X_2483_ net304 VGND VPWR _0429_ state\[45\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1434_ VPWR _0134_ daisychain\[105\] VGND sg13g2_inv_1
X_1365_ VPWR _0068_ state\[46\] VGND sg13g2_inv_1
X_2473__345 VPWR VGND net344 sg13g2_tiehi
X_1296_ VPWR _0017_ state\[115\] VGND sg13g2_inv_1
XFILLER_49_780 VPWR VGND sg13g2_fill_2
XFILLER_23_102 VPWR VGND sg13g2_decap_8
XFILLER_11_319 VPWR VGND sg13g2_decap_8
XFILLER_23_179 VPWR VGND sg13g2_decap_8
XFILLER_32_680 VPWR VGND sg13g2_fill_1
XFILLER_11_46 VPWR VGND sg13g2_decap_8
X_2521__335 VPWR VGND net334 sg13g2_tiehi
XFILLER_46_238 VPWR VGND sg13g2_decap_8
XFILLER_36_21 VPWR VGND sg13g2_decap_8
X_2452__429 VPWR VGND net428 sg13g2_tiehi
XFILLER_27_441 VPWR VGND sg13g2_decap_8
XFILLER_14_102 VPWR VGND sg13g2_decap_8
XFILLER_15_647 VPWR VGND sg13g2_fill_2
XFILLER_43_978 VPWR VGND sg13g2_fill_1
XFILLER_36_98 VPWR VGND sg13g2_decap_8
XFILLER_14_179 VPWR VGND sg13g2_decap_8
XFILLER_30_639 VPWR VGND sg13g2_fill_2
XFILLER_7_813 VPWR VGND sg13g2_decap_8
XFILLER_7_846 VPWR VGND sg13g2_decap_4
XFILLER_6_312 VPWR VGND sg13g2_decap_8
XFILLER_10_396 VPWR VGND sg13g2_decap_8
XFILLER_6_389 VPWR VGND sg13g2_decap_8
XFILLER_37_238 VPWR VGND sg13g2_decap_8
X_2533__239 VPWR VGND net238 sg13g2_tiehi
XFILLER_18_463 VPWR VGND sg13g2_fill_2
XFILLER_21_617 VPWR VGND sg13g2_fill_2
X_1983_ net176 _0140_ _0844_ _0845_ VPWR VGND sg13g2_a21o_1
XFILLER_20_116 VPWR VGND sg13g2_decap_8
XFILLER_9_172 VPWR VGND sg13g2_decap_8
X_2535_ net474 VGND VPWR _0481_ state\[97\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2466_ net372 VGND VPWR _0412_ state\[28\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_1417_ VPWR _0153_ daisychain\[122\] VGND sg13g2_inv_1
X_2397_ net309 VGND VPWR _0343_ daisychain\[87\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_1348_ VPWR _0087_ state\[63\] VGND sg13g2_inv_1
XFILLER_3_1020 VPWR VGND sg13g2_decap_8
XFILLER_28_249 VPWR VGND sg13g2_decap_8
XFILLER_25_978 VPWR VGND sg13g2_fill_1
XFILLER_24_444 VPWR VGND sg13g2_decap_8
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_11_116 VPWR VGND sg13g2_decap_8
XdigitalenH.g\[2\].u.inv2 VPWR digitalenH.g\[2\].u.OUTP digitalenH.g\[2\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_22_67 VPWR VGND sg13g2_decap_8
XFILLER_3_326 VPWR VGND sg13g2_decap_8
Xfanout140 net142 net140 VPWR VGND sg13g2_buf_1
Xfanout173 net174 net173 VPWR VGND sg13g2_buf_1
Xfanout162 net164 net162 VPWR VGND sg13g2_buf_1
Xfanout151 net152 net151 VPWR VGND sg13g2_buf_1
Xfanout195 net198 net195 VPWR VGND sg13g2_buf_1
Xfanout184 net186 net184 VPWR VGND sg13g2_buf_1
XFILLER_47_525 VPWR VGND sg13g2_fill_1
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_19_249 VPWR VGND sg13g2_decap_8
XFILLER_28_783 VPWR VGND sg13g2_decap_8
XFILLER_43_731 VPWR VGND sg13g2_fill_2
XFILLER_15_477 VPWR VGND sg13g2_decap_4
XFILLER_42_252 VPWR VGND sg13g2_decap_8
XFILLER_30_403 VPWR VGND sg13g2_decap_8
XFILLER_31_959 VPWR VGND sg13g2_fill_1
XFILLER_30_425 VPWR VGND sg13g2_fill_2
XFILLER_8_25 VPWR VGND sg13g2_decap_8
XFILLER_30_458 VPWR VGND sg13g2_decap_4
XFILLER_11_694 VPWR VGND sg13g2_decap_4
XFILLER_10_193 VPWR VGND sg13g2_decap_8
XFILLER_7_698 VPWR VGND sg13g2_decap_4
XFILLER_6_186 VPWR VGND sg13g2_decap_8
X_2320_ net463 VGND VPWR _0266_ daisychain\[10\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2251_ VGND VPWR _0809_ _0996_ _0482_ net86 sg13g2_a21oi_1
XFILLER_26_4 VPWR VGND sg13g2_decap_8
X_2182_ _0962_ net153 state\[64\] VPWR VGND sg13g2_nand2_1
XFILLER_19_761 VPWR VGND sg13g2_decap_8
XFILLER_33_263 VPWR VGND sg13g2_decap_8
XFILLER_21_403 VPWR VGND sg13g2_decap_8
X_1966_ net215 VPWR _0832_ VGND state\[106\] net179 sg13g2_o21ai_1
XFILLER_21_458 VPWR VGND sg13g2_fill_2
X_1897_ VPWR VGND _0780_ net83 _0779_ _0242_ _0344_ net38 sg13g2_a221oi_1
X_2518_ net358 VGND VPWR _0464_ state\[80\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_0_329 VPWR VGND sg13g2_decap_8
X_2405__294 VPWR VGND net293 sg13g2_tiehi
X_2449_ net440 VGND VPWR _0395_ state\[11\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_17_56 VPWR VGND sg13g2_decap_8
XFILLER_12_403 VPWR VGND sg13g2_decap_8
XFILLER_24_263 VPWR VGND sg13g2_decap_8
XFILLER_33_11 VPWR VGND sg13g2_decap_8
XFILLER_12_458 VPWR VGND sg13g2_decap_8
XFILLER_33_88 VPWR VGND sg13g2_decap_8
XFILLER_20_480 VPWR VGND sg13g2_fill_2
XFILLER_4_602 VPWR VGND sg13g2_decap_8
XFILLER_3_123 VPWR VGND sg13g2_decap_8
XFILLER_0_830 VPWR VGND sg13g2_decap_8
XFILLER_0_863 VPWR VGND sg13g2_decap_8
XFILLER_0_874 VPWR VGND sg13g2_fill_2
XFILLER_47_322 VPWR VGND sg13g2_decap_8
XFILLER_48_889 VPWR VGND sg13g2_fill_2
XFILLER_35_517 VPWR VGND sg13g2_fill_2
XFILLER_47_399 VPWR VGND sg13g2_decap_8
XFILLER_15_263 VPWR VGND sg13g2_decap_8
XFILLER_30_200 VPWR VGND sg13g2_decap_8
X_1820_ VGND VPWR net156 daisychain\[68\] _0723_ net66 sg13g2_a21oi_1
XFILLER_30_277 VPWR VGND sg13g2_decap_8
XFILLER_11_480 VPWR VGND sg13g2_decap_8
X_1751_ net188 _0203_ _0670_ _0671_ VPWR VGND sg13g2_a21o_1
XFILLER_8_952 VPWR VGND sg13g2_fill_1
X_1682_ net218 VPWR _0619_ VGND state\[35\] net162 sg13g2_o21ai_1
XFILLER_8_985 VPWR VGND sg13g2_fill_1
XFILLER_7_462 VPWR VGND sg13g2_decap_8
X_2303_ VGND VPWR _0887_ _1022_ _0508_ net69 sg13g2_a21oi_1
X_2234_ _0988_ net148 state\[90\] VPWR VGND sg13g2_nand2_1
XFILLER_38_322 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
X_2165_ VGND VPWR _0680_ _0953_ _0439_ net100 sg13g2_a21oi_1
XFILLER_0_1001 VPWR VGND sg13g2_fill_2
XFILLER_0_1012 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
X_2096_ _0919_ net118 state\[21\] VPWR VGND sg13g2_nand2_1
XFILLER_38_399 VPWR VGND sg13g2_decap_8
XFILLER_34_594 VPWR VGND sg13g2_decap_4
XFILLER_21_200 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_485 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_21_277 VPWR VGND sg13g2_decap_8
X_1949_ VPWR VGND _0819_ net89 _0818_ _0130_ _0357_ net47 sg13g2_a221oi_1
XFILLER_1_616 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_49_609 VPWR VGND sg13g2_decap_8
XFILLER_48_119 VPWR VGND sg13g2_decap_8
XFILLER_28_11 VPWR VGND sg13g2_decap_8
XFILLER_29_333 VPWR VGND sg13g2_decap_8
X_2338__428 VPWR VGND net427 sg13g2_tiehi
XFILLER_28_88 VPWR VGND sg13g2_decap_8
XFILLER_44_336 VPWR VGND sg13g2_decap_8
XFILLER_44_21 VPWR VGND sg13g2_decap_8
XFILLER_25_550 VPWR VGND sg13g2_decap_8
XFILLER_12_200 VPWR VGND sg13g2_decap_8
XFILLER_25_572 VPWR VGND sg13g2_decap_4
XFILLER_44_98 VPWR VGND sg13g2_decap_8
XFILLER_12_277 VPWR VGND sg13g2_decap_8
XFILLER_5_900 VPWR VGND sg13g2_decap_4
XFILLER_4_410 VPWR VGND sg13g2_decap_8
XFILLER_4_476 VPWR VGND sg13g2_decap_8
XFILLER_39_119 VPWR VGND sg13g2_decap_8
XFILLER_0_693 VPWR VGND sg13g2_decap_8
XFILLER_47_196 VPWR VGND sg13g2_decap_8
XFILLER_35_336 VPWR VGND sg13g2_decap_8
X_2389__326 VPWR VGND net325 sg13g2_tiehi
XFILLER_31_553 VPWR VGND sg13g2_decap_8
X_2469__361 VPWR VGND net360 sg13g2_tiehi
X_1803_ net200 _0217_ _0709_ _0710_ VPWR VGND sg13g2_a21o_1
X_1734_ net222 VPWR _0658_ VGND state\[48\] net192 sg13g2_o21ai_1
XFILLER_8_771 VPWR VGND sg13g2_fill_1
XFILLER_8_760 VPWR VGND sg13g2_fill_2
X_1665_ VPWR VGND _0606_ net76 _0605_ _0179_ _0286_ net31 sg13g2_a221oi_1
X_1596_ VGND VPWR net138 daisychain\[12\] _0555_ net52 sg13g2_a21oi_1
X_2217_ VGND VPWR _0758_ _0979_ _0465_ net105 sg13g2_a21oi_1
XFILLER_39_675 VPWR VGND sg13g2_decap_4
X_2148_ _0945_ net139 state\[47\] VPWR VGND sg13g2_nand2_1
XFILLER_38_196 VPWR VGND sg13g2_decap_8
XFILLER_27_859 VPWR VGND sg13g2_fill_2
XFILLER_26_347 VPWR VGND sg13g2_decap_8
X_2079_ VGND VPWR _0551_ _0910_ _0396_ net73 sg13g2_a21oi_1
XFILLER_14_46 VPWR VGND sg13g2_decap_8
X_2448__445 VPWR VGND net444 sg13g2_tiehi
XFILLER_5_207 VPWR VGND sg13g2_decap_8
X_2524__311 VPWR VGND net310 sg13g2_tiehi
XFILLER_30_67 VPWR VGND sg13g2_decap_8
XFILLER_2_958 VPWR VGND sg13g2_fill_2
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_39_21 VPWR VGND sg13g2_decap_8
XFILLER_7_1018 VPWR VGND sg13g2_decap_8
XFILLER_49_417 VPWR VGND sg13g2_decap_8
XFILLER_39_98 VPWR VGND sg13g2_decap_8
XFILLER_29_130 VPWR VGND sg13g2_decap_8
XFILLER_18_826 VPWR VGND sg13g2_fill_1
XFILLER_45_601 VPWR VGND sg13g2_decap_4
XFILLER_17_336 VPWR VGND sg13g2_decap_8
XFILLER_18_859 VPWR VGND sg13g2_fill_1
XFILLER_45_656 VPWR VGND sg13g2_fill_2
XFILLER_44_133 VPWR VGND sg13g2_decap_8
XFILLER_40_350 VPWR VGND sg13g2_decap_8
XFILLER_9_568 VPWR VGND sg13g2_decap_8
XFILLER_9_557 VPWR VGND sg13g2_decap_8
X_1450_ VPWR _0243_ daisychain\[89\] VGND sg13g2_inv_1
XFILLER_4_284 VPWR VGND sg13g2_decap_8
XFILLER_45_1002 VPWR VGND sg13g2_decap_4
X_1381_ VPWR _0051_ state\[30\] VGND sg13g2_inv_1
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_49_984 VPWR VGND sg13g2_decap_8
X_2002_ net215 VPWR _0859_ VGND state\[115\] net179 sg13g2_o21ai_1
XFILLER_48_483 VPWR VGND sg13g2_decap_8
XFILLER_35_133 VPWR VGND sg13g2_decap_8
XFILLER_31_361 VPWR VGND sg13g2_decap_8
X_2835_ state\[125\] net13 VPWR VGND sg13g2_buf_1
X_1717_ VPWR VGND _0645_ net94 _0644_ _0193_ _0299_ net50 sg13g2_a221oi_1
X_1648_ VGND VPWR net119 daisychain\[25\] _0594_ net30 sg13g2_a21oi_1
X_1579_ net164 _0255_ _0541_ _0542_ VPWR VGND sg13g2_a21o_1
XFILLER_26_144 VPWR VGND sg13g2_decap_8
XFILLER_42_626 VPWR VGND sg13g2_decap_8
XFILLER_41_147 VPWR VGND sg13g2_decap_8
XFILLER_25_67 VPWR VGND sg13g2_decap_8
XFILLER_10_501 VPWR VGND sg13g2_decap_8
XFILLER_22_361 VPWR VGND sg13g2_decap_8
XFILLER_41_77 VPWR VGND sg13g2_decap_8
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_49_214 VPWR VGND sg13g2_decap_8
XFILLER_1_287 VPWR VGND sg13g2_decap_8
XFILLER_46_943 VPWR VGND sg13g2_decap_8
XFILLER_45_420 VPWR VGND sg13g2_decap_8
XFILLER_17_133 VPWR VGND sg13g2_decap_8
XFILLER_46_976 VPWR VGND sg13g2_fill_1
XFILLER_46_965 VPWR VGND sg13g2_fill_1
XFILLER_46_998 VPWR VGND sg13g2_fill_2
XFILLER_13_361 VPWR VGND sg13g2_decap_8
XFILLER_32_158 VPWR VGND sg13g2_decap_8
XFILLER_9_354 VPWR VGND sg13g2_decap_8
X_2551_ net466 VGND VPWR _0497_ state\[113\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_2482_ net308 VGND VPWR _0428_ state\[44\] clknet_leaf_15_clk sg13g2_dfrbpq_1
X_1502_ VPWR _0186_ daisychain\[37\] VGND sg13g2_inv_1
X_1433_ VPWR _0135_ daisychain\[106\] VGND sg13g2_inv_1
X_1364_ VPWR _0069_ state\[47\] VGND sg13g2_inv_1
X_1295_ VPWR _0018_ state\[116\] VGND sg13g2_inv_1
XFILLER_49_792 VPWR VGND sg13g2_fill_1
XFILLER_48_280 VPWR VGND sg13g2_decap_8
XFILLER_36_486 VPWR VGND sg13g2_fill_1
XFILLER_23_158 VPWR VGND sg13g2_decap_8
XFILLER_11_25 VPWR VGND sg13g2_decap_8
X_2480__317 VPWR VGND net316 sg13g2_tiehi
XFILLER_46_217 VPWR VGND sg13g2_decap_8
XFILLER_39_280 VPWR VGND sg13g2_decap_8
XFILLER_27_420 VPWR VGND sg13g2_decap_8
XFILLER_15_604 VPWR VGND sg13g2_fill_1
XFILLER_36_77 VPWR VGND sg13g2_decap_8
XFILLER_15_637 VPWR VGND sg13g2_decap_4
XFILLER_14_158 VPWR VGND sg13g2_decap_8
X_2415__274 VPWR VGND net273 sg13g2_tiehi
XFILLER_23_692 VPWR VGND sg13g2_fill_1
XFILLER_7_825 VPWR VGND sg13g2_decap_8
XFILLER_10_375 VPWR VGND sg13g2_decap_8
XFILLER_7_869 VPWR VGND sg13g2_decap_8
XFILLER_6_368 VPWR VGND sg13g2_decap_8
XFILLER_2_585 VPWR VGND sg13g2_decap_8
XFILLER_42_1027 VPWR VGND sg13g2_fill_2
XFILLER_37_217 VPWR VGND sg13g2_decap_8
XFILLER_18_420 VPWR VGND sg13g2_decap_8
XFILLER_19_954 VPWR VGND sg13g2_decap_8
XFILLER_46_784 VPWR VGND sg13g2_decap_8
XFILLER_18_497 VPWR VGND sg13g2_decap_4
XFILLER_45_294 VPWR VGND sg13g2_decap_8
XFILLER_33_467 VPWR VGND sg13g2_fill_1
XFILLER_14_692 VPWR VGND sg13g2_decap_8
X_1982_ net213 VPWR _0844_ VGND state\[110\] net175 sg13g2_o21ai_1
XFILLER_9_151 VPWR VGND sg13g2_decap_8
X_2534_ net230 VGND VPWR _0480_ state\[96\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_2465_ net376 VGND VPWR _0411_ state\[27\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2396_ net311 VGND VPWR _0342_ daisychain\[86\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_1416_ VPWR _0154_ daisychain\[123\] VGND sg13g2_inv_1
X_1347_ VPWR _0088_ state\[64\] VGND sg13g2_inv_1
XFILLER_3_81 VPWR VGND sg13g2_decap_8
XFILLER_29_718 VPWR VGND sg13g2_fill_1
XFILLER_28_228 VPWR VGND sg13g2_decap_8
XFILLER_36_294 VPWR VGND sg13g2_decap_8
XFILLER_22_46 VPWR VGND sg13g2_decap_8
XFILLER_3_305 VPWR VGND sg13g2_decap_8
Xfanout130 net136 net130 VPWR VGND sg13g2_buf_1
Xfanout174 net183 net174 VPWR VGND sg13g2_buf_1
Xfanout163 net164 net163 VPWR VGND sg13g2_buf_1
Xfanout152 net158 net152 VPWR VGND sg13g2_buf_1
Xfanout141 net142 net141 VPWR VGND sg13g2_buf_1
XFILLER_47_504 VPWR VGND sg13g2_decap_4
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_19_228 VPWR VGND sg13g2_decap_8
Xfanout196 net198 net196 VPWR VGND sg13g2_buf_1
Xfanout185 net186 net185 VPWR VGND sg13g2_buf_1
XFILLER_47_98 VPWR VGND sg13g2_decap_8
XFILLER_28_773 VPWR VGND sg13g2_fill_1
XFILLER_28_762 VPWR VGND sg13g2_decap_8
XFILLER_15_445 VPWR VGND sg13g2_decap_8
XFILLER_27_294 VPWR VGND sg13g2_decap_8
XFILLER_15_456 VPWR VGND sg13g2_fill_1
X_2317__470 VPWR VGND net469 sg13g2_tiehi
XFILLER_42_231 VPWR VGND sg13g2_decap_8
XFILLER_15_489 VPWR VGND sg13g2_decap_8
XFILLER_30_437 VPWR VGND sg13g2_decap_8
X_2348__408 VPWR VGND net407 sg13g2_tiehi
XFILLER_10_172 VPWR VGND sg13g2_decap_8
XFILLER_6_165 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_decap_8
X_2250_ _0996_ net130 state\[98\] VPWR VGND sg13g2_nand2_1
XFILLER_2_382 VPWR VGND sg13g2_decap_8
X_2181_ VGND VPWR _0704_ _0961_ _0447_ net100 sg13g2_a21oi_1
XFILLER_19_4 VPWR VGND sg13g2_decap_8
XFILLER_46_570 VPWR VGND sg13g2_fill_1
XFILLER_33_242 VPWR VGND sg13g2_decap_8
X_1965_ VPWR VGND _0831_ net89 _0830_ _0134_ _0361_ net47 sg13g2_a221oi_1
X_1896_ VGND VPWR net127 daisychain\[87\] _0780_ net38 sg13g2_a21oi_1
XFILLER_0_308 VPWR VGND sg13g2_decap_8
X_2399__306 VPWR VGND net305 sg13g2_tiehi
X_2517_ net366 VGND VPWR _0463_ state\[79\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_2448_ net444 VGND VPWR _0394_ state\[10\] clknet_leaf_18_clk sg13g2_dfrbpq_1
X_2379_ net345 VGND VPWR _0325_ daisychain\[69\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_17_35 VPWR VGND sg13g2_decap_8
XFILLER_24_242 VPWR VGND sg13g2_decap_8
XFILLER_12_437 VPWR VGND sg13g2_decap_8
XFILLER_25_787 VPWR VGND sg13g2_decap_4
XFILLER_33_67 VPWR VGND sg13g2_decap_8
XFILLER_3_102 VPWR VGND sg13g2_decap_8
XFILLER_4_658 VPWR VGND sg13g2_decap_8
XFILLER_3_179 VPWR VGND sg13g2_decap_8
XFILLER_0_853 VPWR VGND sg13g2_fill_1
XFILLER_47_301 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
XFILLER_15_242 VPWR VGND sg13g2_decap_8
XFILLER_43_562 VPWR VGND sg13g2_decap_8
XFILLER_43_540 VPWR VGND sg13g2_fill_2
XFILLER_31_746 VPWR VGND sg13g2_fill_1
X_1750_ net221 VPWR _0670_ VGND state\[52\] net188 sg13g2_o21ai_1
XFILLER_8_931 VPWR VGND sg13g2_fill_1
XFILLER_30_256 VPWR VGND sg13g2_decap_8
XFILLER_8_964 VPWR VGND sg13g2_fill_1
XFILLER_7_441 VPWR VGND sg13g2_decap_8
X_1681_ VPWR VGND _0618_ net74 _0617_ _0183_ _0290_ net28 sg13g2_a221oi_1
X_2302_ _1022_ net115 state\[124\] VPWR VGND sg13g2_nand2_1
X_2441__473 VPWR VGND net472 sg13g2_tiehi
X_2233_ VGND VPWR _0782_ _0987_ _0473_ net86 sg13g2_a21oi_1
XFILLER_38_301 VPWR VGND sg13g2_decap_8
X_2164_ _0953_ net146 state\[55\] VPWR VGND sg13g2_nand2_1
X_2552__435 VPWR VGND net434 sg13g2_tiehi
XFILLER_38_378 VPWR VGND sg13g2_decap_8
X_2095_ VGND VPWR _0575_ _0918_ _0404_ net75 sg13g2_a21oi_1
XFILLER_34_562 VPWR VGND sg13g2_decap_8
XFILLER_34_573 VPWR VGND sg13g2_fill_1
Xheichips25_pudding_486 VPWR VGND uio_oe[2] sg13g2_tiehi
XFILLER_21_256 VPWR VGND sg13g2_decap_8
X_1948_ VGND VPWR net133 daisychain\[100\] _0819_ net47 sg13g2_a21oi_1
X_1879_ net172 _0238_ _0766_ _0767_ VPWR VGND sg13g2_a21o_1
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_29_312 VPWR VGND sg13g2_decap_8
XFILLER_28_67 VPWR VGND sg13g2_decap_8
XFILLER_44_315 VPWR VGND sg13g2_decap_8
XFILLER_29_389 VPWR VGND sg13g2_decap_8
XFILLER_44_77 VPWR VGND sg13g2_decap_8
XFILLER_12_256 VPWR VGND sg13g2_decap_8
XFILLER_8_249 VPWR VGND sg13g2_decap_8
XFILLER_4_466 VPWR VGND sg13g2_decap_4
XFILLER_0_672 VPWR VGND sg13g2_decap_8
Xclkbuf_2_3__f_clk clknet_2_3__leaf_clk clknet_0_clk VPWR VGND sg13g2_buf_16
XFILLER_47_175 VPWR VGND sg13g2_decap_8
XFILLER_35_315 VPWR VGND sg13g2_decap_8
XFILLER_43_392 VPWR VGND sg13g2_decap_8
XFILLER_31_532 VPWR VGND sg13g2_decap_4
X_1802_ net225 VPWR _0709_ VGND state\[65\] net200 sg13g2_o21ai_1
X_1733_ VPWR VGND _0657_ net106 _0656_ _0197_ _0303_ net62 sg13g2_a221oi_1
XFILLER_8_783 VPWR VGND sg13g2_fill_1
X_1664_ VGND VPWR net119 daisychain\[29\] _0606_ net31 sg13g2_a21oi_1
X_1595_ net184 _0160_ _0553_ _0554_ VPWR VGND sg13g2_a21o_1
X_2216_ _0979_ net151 state\[81\] VPWR VGND sg13g2_nand2_1
X_2476__333 VPWR VGND net332 sg13g2_tiehi
XFILLER_22_1025 VPWR VGND sg13g2_decap_4
X_2147_ VGND VPWR _0653_ _0944_ _0430_ net93 sg13g2_a21oi_1
XFILLER_38_175 VPWR VGND sg13g2_decap_8
XFILLER_26_326 VPWR VGND sg13g2_decap_8
X_2078_ _0910_ net116 state\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_41_329 VPWR VGND sg13g2_decap_8
XFILLER_22_510 VPWR VGND sg13g2_decap_8
XFILLER_14_25 VPWR VGND sg13g2_decap_8
XFILLER_22_587 VPWR VGND sg13g2_decap_4
XFILLER_22_565 VPWR VGND sg13g2_fill_2
XFILLER_30_46 VPWR VGND sg13g2_decap_8
XFILLER_2_926 VPWR VGND sg13g2_decap_4
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_39_77 VPWR VGND sg13g2_decap_8
XFILLER_18_805 VPWR VGND sg13g2_fill_1
X_2455__417 VPWR VGND net416 sg13g2_tiehi
XFILLER_17_315 VPWR VGND sg13g2_decap_8
XFILLER_18_838 VPWR VGND sg13g2_fill_1
XFILLER_44_112 VPWR VGND sg13g2_decap_8
XFILLER_29_186 VPWR VGND sg13g2_decap_8
XFILLER_44_189 VPWR VGND sg13g2_decap_8
XFILLER_9_536 VPWR VGND sg13g2_decap_8
X_2425__254 VPWR VGND net253 sg13g2_tiehi
XFILLER_4_263 VPWR VGND sg13g2_decap_8
X_1380_ VPWR _0052_ state\[31\] VGND sg13g2_inv_1
X_2001_ VPWR VGND _0858_ net82 _0857_ _0144_ _0370_ net37 sg13g2_a221oi_1
XFILLER_48_462 VPWR VGND sg13g2_decap_8
XFILLER_35_112 VPWR VGND sg13g2_decap_8
XFILLER_24_819 VPWR VGND sg13g2_decap_8
XFILLER_35_189 VPWR VGND sg13g2_decap_8
XFILLER_32_852 VPWR VGND sg13g2_decap_4
XFILLER_32_874 VPWR VGND sg13g2_fill_2
XFILLER_31_340 VPWR VGND sg13g2_decap_8
X_2834_ state\[124\] net12 VPWR VGND sg13g2_buf_1
X_1716_ VGND VPWR net140 daisychain\[42\] _0645_ net50 sg13g2_a21oi_1
X_1647_ net167 _0174_ _0592_ _0593_ VPWR VGND sg13g2_a21o_1
XFILLER_6_81 VPWR VGND sg13g2_decap_8
X_1578_ net206 VPWR _0541_ VGND state\[9\] net164 sg13g2_o21ai_1
XFILLER_39_440 VPWR VGND sg13g2_decap_4
XFILLER_39_495 VPWR VGND sg13g2_fill_1
XFILLER_27_635 VPWR VGND sg13g2_decap_4
XFILLER_27_657 VPWR VGND sg13g2_decap_8
XFILLER_26_123 VPWR VGND sg13g2_decap_8
XFILLER_41_126 VPWR VGND sg13g2_decap_8
XFILLER_25_46 VPWR VGND sg13g2_decap_8
XFILLER_22_340 VPWR VGND sg13g2_decap_8
XFILLER_41_56 VPWR VGND sg13g2_decap_8
XFILLER_2_712 VPWR VGND sg13g2_decap_4
XFILLER_2_745 VPWR VGND sg13g2_fill_1
XFILLER_2_778 VPWR VGND sg13g2_fill_2
XFILLER_1_266 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_46_911 VPWR VGND sg13g2_decap_4
XFILLER_17_112 VPWR VGND sg13g2_decap_8
XFILLER_18_668 VPWR VGND sg13g2_decap_8
XFILLER_17_189 VPWR VGND sg13g2_decap_8
XFILLER_45_498 VPWR VGND sg13g2_decap_8
XFILLER_32_137 VPWR VGND sg13g2_decap_8
XFILLER_13_340 VPWR VGND sg13g2_decap_8
XFILLER_9_333 VPWR VGND sg13g2_decap_8
X_2550_ net234 VGND VPWR _0496_ state\[112\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2327__450 VPWR VGND net449 sg13g2_tiehi
X_2481_ net312 VGND VPWR _0427_ state\[43\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1501_ VPWR _0187_ daisychain\[38\] VGND sg13g2_inv_1
XFILLER_5_583 VPWR VGND sg13g2_decap_8
X_1432_ VPWR _0136_ daisychain\[107\] VGND sg13g2_inv_1
XFILLER_49_4 VPWR VGND sg13g2_decap_8
X_1363_ VPWR _0070_ state\[48\] VGND sg13g2_inv_1
X_1294_ VPWR _0019_ state\[117\] VGND sg13g2_inv_1
XFILLER_24_605 VPWR VGND sg13g2_fill_1
XFILLER_23_137 VPWR VGND sg13g2_decap_8
XFILLER_15_616 VPWR VGND sg13g2_decap_8
XFILLER_43_914 VPWR VGND sg13g2_fill_2
XFILLER_42_413 VPWR VGND sg13g2_decap_8
XFILLER_36_56 VPWR VGND sg13g2_decap_8
XFILLER_28_988 VPWR VGND sg13g2_decap_8
XFILLER_14_137 VPWR VGND sg13g2_decap_8
XFILLER_30_608 VPWR VGND sg13g2_decap_4
XFILLER_10_354 VPWR VGND sg13g2_decap_8
XFILLER_6_347 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_2_564 VPWR VGND sg13g2_decap_8
XFILLER_19_900 VPWR VGND sg13g2_decap_8
XFILLER_19_922 VPWR VGND sg13g2_decap_8
XFILLER_18_454 VPWR VGND sg13g2_fill_1
XFILLER_45_273 VPWR VGND sg13g2_decap_8
X_1981_ VPWR VGND _0843_ net87 _0842_ _0138_ _0365_ net44 sg13g2_a221oi_1
XFILLER_9_130 VPWR VGND sg13g2_decap_8
X_2533_ net238 VGND VPWR _0479_ state\[95\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_6_892 VPWR VGND sg13g2_fill_2
X_2464_ net380 VGND VPWR _0410_ state\[26\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_2395_ net313 VGND VPWR _0341_ daisychain\[85\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_1415_ VPWR _0155_ daisychain\[124\] VGND sg13g2_inv_1
X_1346_ VPWR _0089_ state\[65\] VGND sg13g2_inv_1
XFILLER_3_60 VPWR VGND sg13g2_decap_8
XFILLER_28_207 VPWR VGND sg13g2_decap_8
XFILLER_36_273 VPWR VGND sg13g2_decap_8
XFILLER_24_424 VPWR VGND sg13g2_decap_8
XFILLER_24_479 VPWR VGND sg13g2_decap_8
XFILLER_22_25 VPWR VGND sg13g2_decap_8
XFILLER_20_641 VPWR VGND sg13g2_decap_4
XFILLER_0_7 VPWR VGND sg13g2_decap_8
Xfanout131 net135 net131 VPWR VGND sg13g2_buf_1
Xfanout120 net121 net120 VPWR VGND sg13g2_buf_1
Xfanout164 net169 net164 VPWR VGND sg13g2_buf_1
Xfanout153 net157 net153 VPWR VGND sg13g2_buf_1
Xfanout142 net147 net142 VPWR VGND sg13g2_buf_1
XFILLER_19_207 VPWR VGND sg13g2_decap_8
Xfanout197 net198 net197 VPWR VGND sg13g2_buf_1
Xfanout186 net187 net186 VPWR VGND sg13g2_buf_1
Xfanout175 net178 net175 VPWR VGND sg13g2_buf_1
XFILLER_47_516 VPWR VGND sg13g2_decap_8
XFILLER_47_77 VPWR VGND sg13g2_decap_8
XFILLER_15_424 VPWR VGND sg13g2_decap_8
XFILLER_42_210 VPWR VGND sg13g2_decap_8
XFILLER_27_273 VPWR VGND sg13g2_decap_8
XFILLER_42_287 VPWR VGND sg13g2_decap_8
XFILLER_30_427 VPWR VGND sg13g2_fill_1
XFILLER_10_151 VPWR VGND sg13g2_decap_8
XFILLER_6_144 VPWR VGND sg13g2_decap_8
XFILLER_2_361 VPWR VGND sg13g2_decap_8
X_2180_ _0961_ net146 state\[63\] VPWR VGND sg13g2_nand2_1
XFILLER_19_785 VPWR VGND sg13g2_decap_8
XFILLER_18_284 VPWR VGND sg13g2_decap_8
XFILLER_33_221 VPWR VGND sg13g2_decap_8
XFILLER_14_490 VPWR VGND sg13g2_decap_8
X_1964_ VGND VPWR net133 daisychain\[104\] _0831_ net46 sg13g2_a21oi_1
Xclkbuf_leaf_13_clk clknet_2_2__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
XFILLER_33_298 VPWR VGND sg13g2_decap_8
XFILLER_21_438 VPWR VGND sg13g2_decap_8
XFILLER_30_983 VPWR VGND sg13g2_fill_1
XFILLER_30_972 VPWR VGND sg13g2_decap_8
X_1895_ net173 _0242_ _0778_ _0779_ VPWR VGND sg13g2_a21o_1
X_2516_ net374 VGND VPWR _0462_ state\[78\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2447_ net448 VGND VPWR _0393_ state\[9\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_2378_ net347 VGND VPWR _0324_ daisychain\[68\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_17_14 VPWR VGND sg13g2_decap_8
X_1329_ VPWR _0108_ state\[82\] VGND sg13g2_inv_1
XFILLER_44_508 VPWR VGND sg13g2_decap_8
XFILLER_37_571 VPWR VGND sg13g2_fill_2
XFILLER_24_221 VPWR VGND sg13g2_decap_8
XFILLER_12_416 VPWR VGND sg13g2_decap_8
XFILLER_40_725 VPWR VGND sg13g2_decap_8
XFILLER_33_46 VPWR VGND sg13g2_decap_8
XFILLER_24_298 VPWR VGND sg13g2_decap_8
XFILLER_21_983 VPWR VGND sg13g2_decap_8
XFILLER_4_637 VPWR VGND sg13g2_decap_4
XFILLER_3_158 VPWR VGND sg13g2_decap_8
XFILLER_47_357 VPWR VGND sg13g2_decap_8
XFILLER_15_221 VPWR VGND sg13g2_decap_8
XFILLER_31_714 VPWR VGND sg13g2_fill_2
XFILLER_15_298 VPWR VGND sg13g2_decap_8
XFILLER_31_758 VPWR VGND sg13g2_fill_2
XFILLER_30_235 VPWR VGND sg13g2_decap_8
XFILLER_8_910 VPWR VGND sg13g2_fill_1
XFILLER_8_943 VPWR VGND sg13g2_fill_1
XFILLER_7_420 VPWR VGND sg13g2_decap_8
X_1680_ VGND VPWR net117 daisychain\[33\] _0618_ net28 sg13g2_a21oi_1
XFILLER_8_998 VPWR VGND sg13g2_decap_4
XFILLER_7_497 VPWR VGND sg13g2_decap_8
XFILLER_48_1001 VPWR VGND sg13g2_fill_1
X_2301_ VGND VPWR _0884_ _1021_ _0507_ net70 sg13g2_a21oi_1
XFILLER_31_4 VPWR VGND sg13g2_decap_8
X_2232_ _0987_ net130 state\[89\] VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
X_2163_ VGND VPWR _0677_ _0952_ _0438_ net99 sg13g2_a21oi_1
XFILLER_38_357 VPWR VGND sg13g2_decap_8
X_2094_ _0918_ net118 state\[20\] VPWR VGND sg13g2_nand2_1
X_2435__234 VPWR VGND net233 sg13g2_tiehi
Xheichips25_pudding_487 VPWR VGND uio_oe[3] sg13g2_tiehi
XFILLER_21_235 VPWR VGND sg13g2_decap_8
XFILLER_9_81 VPWR VGND sg13g2_decap_8
X_1947_ net180 _0130_ _0817_ _0818_ VPWR VGND sg13g2_a21o_1
XFILLER_30_791 VPWR VGND sg13g2_decap_8
X_1878_ net211 VPWR _0766_ VGND state\[84\] net172 sg13g2_o21ai_1
XFILLER_28_46 VPWR VGND sg13g2_decap_8
XFILLER_29_368 VPWR VGND sg13g2_decap_8
XFILLER_44_56 VPWR VGND sg13g2_decap_8
XFILLER_12_235 VPWR VGND sg13g2_decap_8
XFILLER_13_736 VPWR VGND sg13g2_fill_2
XFILLER_9_707 VPWR VGND sg13g2_fill_2
XFILLER_8_228 VPWR VGND sg13g2_decap_8
XFILLER_40_599 VPWR VGND sg13g2_decap_4
XFILLER_21_791 VPWR VGND sg13g2_decap_8
XFILLER_5_39 VPWR VGND sg13g2_decap_8
XFILLER_4_445 VPWR VGND sg13g2_decap_8
X_2540__395 VPWR VGND net394 sg13g2_tiehi
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_47_154 VPWR VGND sg13g2_decap_8
XFILLER_16_530 VPWR VGND sg13g2_decap_4
XFILLER_44_850 VPWR VGND sg13g2_fill_1
XFILLER_43_371 VPWR VGND sg13g2_decap_8
X_1801_ VPWR VGND _0708_ net107 _0707_ _0216_ _0320_ net63 sg13g2_a221oi_1
X_1732_ VGND VPWR net154 daisychain\[46\] _0657_ net62 sg13g2_a21oi_1
XFILLER_8_762 VPWR VGND sg13g2_fill_1
X_1663_ net168 _0179_ _0604_ _0605_ VPWR VGND sg13g2_a21o_1
XFILLER_7_294 VPWR VGND sg13g2_decap_8
X_1594_ net218 VPWR _0553_ VGND state\[13\] net184 sg13g2_o21ai_1
X_2215_ VGND VPWR _0755_ _0978_ _0464_ net102 sg13g2_a21oi_1
XFILLER_38_154 VPWR VGND sg13g2_decap_8
X_2146_ _0944_ net139 state\[46\] VPWR VGND sg13g2_nand2_1
X_2337__430 VPWR VGND net429 sg13g2_tiehi
XFILLER_27_839 VPWR VGND sg13g2_fill_2
XFILLER_26_305 VPWR VGND sg13g2_decap_8
X_2077_ VGND VPWR _0548_ _0909_ _0395_ net73 sg13g2_a21oi_1
XFILLER_41_308 VPWR VGND sg13g2_decap_8
XFILLER_34_382 VPWR VGND sg13g2_decap_8
XFILLER_10_728 VPWR VGND sg13g2_decap_4
X_2483__305 VPWR VGND net304 sg13g2_tiehi
XFILLER_30_25 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_39_56 VPWR VGND sg13g2_decap_8
XFILLER_18_817 VPWR VGND sg13g2_fill_1
XFILLER_45_636 VPWR VGND sg13g2_fill_2
XFILLER_29_165 VPWR VGND sg13g2_decap_8
X_2535__475 VPWR VGND net474 sg13g2_tiehi
XFILLER_45_658 VPWR VGND sg13g2_fill_1
XFILLER_45_647 VPWR VGND sg13g2_fill_1
XFILLER_13_500 VPWR VGND sg13g2_decap_8
XFILLER_44_168 VPWR VGND sg13g2_decap_8
XFILLER_32_319 VPWR VGND sg13g2_decap_8
XFILLER_13_511 VPWR VGND sg13g2_decap_4
XFILLER_25_382 VPWR VGND sg13g2_decap_8
XFILLER_9_515 VPWR VGND sg13g2_decap_8
XFILLER_40_385 VPWR VGND sg13g2_decap_8
XFILLER_5_754 VPWR VGND sg13g2_decap_8
XFILLER_4_242 VPWR VGND sg13g2_decap_8
XFILLER_45_1015 VPWR VGND sg13g2_decap_8
X_2000_ VGND VPWR net126 daisychain\[113\] _0858_ net37 sg13g2_a21oi_1
XFILLER_49_964 VPWR VGND sg13g2_decap_4
XFILLER_48_441 VPWR VGND sg13g2_decap_8
XFILLER_35_168 VPWR VGND sg13g2_decap_8
XFILLER_23_319 VPWR VGND sg13g2_decap_8
XFILLER_16_382 VPWR VGND sg13g2_decap_8
XFILLER_32_842 VPWR VGND sg13g2_fill_1
X_2833_ state\[123\] net11 VPWR VGND sg13g2_buf_1
XFILLER_31_396 VPWR VGND sg13g2_decap_8
X_1715_ net185 _0193_ _0643_ _0644_ VPWR VGND sg13g2_a21o_1
XFILLER_6_60 VPWR VGND sg13g2_decap_8
X_1646_ net208 VPWR _0592_ VGND state\[26\] net167 sg13g2_o21ai_1
X_1577_ VPWR VGND _0540_ net70 _0539_ _0244_ _0264_ net33 sg13g2_a221oi_1
XFILLER_26_102 VPWR VGND sg13g2_decap_8
X_2129_ VGND VPWR _0626_ _0935_ _0421_ net92 sg13g2_a21oi_1
XFILLER_14_319 VPWR VGND sg13g2_decap_8
XFILLER_41_105 VPWR VGND sg13g2_decap_8
XFILLER_26_179 VPWR VGND sg13g2_decap_8
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_10_536 VPWR VGND sg13g2_decap_8
XFILLER_41_35 VPWR VGND sg13g2_decap_8
XFILLER_22_396 VPWR VGND sg13g2_decap_8
XFILLER_6_529 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_2_757 VPWR VGND sg13g2_fill_2
XFILLER_2_735 VPWR VGND sg13g2_fill_1
XFILLER_1_245 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_49_249 VPWR VGND sg13g2_decap_8
XFILLER_18_647 VPWR VGND sg13g2_decap_8
XFILLER_18_658 VPWR VGND sg13g2_fill_1
XFILLER_45_455 VPWR VGND sg13g2_decap_8
XFILLER_17_168 VPWR VGND sg13g2_decap_8
XFILLER_33_606 VPWR VGND sg13g2_decap_4
XFILLER_32_116 VPWR VGND sg13g2_decap_8
XFILLER_9_312 VPWR VGND sg13g2_decap_8
XFILLER_13_396 VPWR VGND sg13g2_decap_8
XFILLER_40_182 VPWR VGND sg13g2_decap_8
XFILLER_9_389 VPWR VGND sg13g2_decap_8
X_2480_ net316 VGND VPWR _0426_ state\[42\] clknet_leaf_16_clk sg13g2_dfrbpq_1
X_1500_ VPWR _0188_ daisychain\[39\] VGND sg13g2_inv_1
XFILLER_5_562 VPWR VGND sg13g2_decap_8
X_1431_ VPWR _0137_ daisychain\[108\] VGND sg13g2_inv_1
X_1362_ VPWR _0071_ state\[49\] VGND sg13g2_inv_1
X_1293_ VPWR _0020_ state\[118\] VGND sg13g2_inv_1
XFILLER_49_772 VPWR VGND sg13g2_decap_4
XFILLER_36_444 VPWR VGND sg13g2_decap_8
XFILLER_23_116 VPWR VGND sg13g2_decap_8
XFILLER_32_650 VPWR VGND sg13g2_fill_1
XFILLER_31_193 VPWR VGND sg13g2_decap_8
X_1629_ VPWR VGND _0579_ net75 _0578_ _0169_ _0277_ net29 sg13g2_a221oi_1
X_2560__387 VPWR VGND net386 sg13g2_tiehi
XFILLER_36_35 VPWR VGND sg13g2_decap_8
XFILLER_14_116 VPWR VGND sg13g2_decap_8
XFILLER_42_436 VPWR VGND sg13g2_decap_8
XFILLER_27_499 VPWR VGND sg13g2_decap_8
XFILLER_23_683 VPWR VGND sg13g2_fill_2
XFILLER_10_333 VPWR VGND sg13g2_decap_8
XFILLER_22_193 VPWR VGND sg13g2_decap_8
XFILLER_6_326 VPWR VGND sg13g2_decap_8
XFILLER_2_543 VPWR VGND sg13g2_decap_8
XFILLER_46_742 VPWR VGND sg13g2_decap_8
XFILLER_46_720 VPWR VGND sg13g2_fill_2
XFILLER_45_252 VPWR VGND sg13g2_decap_8
XFILLER_33_403 VPWR VGND sg13g2_decap_8
X_1980_ VGND VPWR net131 daisychain\[108\] _0843_ net44 sg13g2_a21oi_1
XFILLER_42_992 VPWR VGND sg13g2_fill_1
XFILLER_13_193 VPWR VGND sg13g2_decap_8
XFILLER_41_480 VPWR VGND sg13g2_fill_1
XFILLER_9_186 VPWR VGND sg13g2_decap_8
X_2532_ net246 VGND VPWR _0478_ state\[94\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_6_860 VPWR VGND sg13g2_fill_2
X_2444__461 VPWR VGND net460 sg13g2_tiehi
X_2463_ net384 VGND VPWR _0409_ state\[25\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_2394_ net315 VGND VPWR _0340_ daisychain\[84\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1414_ VPWR _0156_ daisychain\[125\] VGND sg13g2_inv_1
X_1345_ VPWR _0090_ state\[66\] VGND sg13g2_inv_1
XFILLER_36_252 VPWR VGND sg13g2_decap_8
XFILLER_25_915 VPWR VGND sg13g2_fill_2
XFILLER_24_403 VPWR VGND sg13g2_decap_8
XFILLER_20_697 VPWR VGND sg13g2_fill_2
Xfanout121 net122 net121 VPWR VGND sg13g2_buf_1
Xfanout110 net111 net110 VPWR VGND sg13g2_buf_1
Xfanout165 net168 net165 VPWR VGND sg13g2_buf_1
Xfanout154 net157 net154 VPWR VGND sg13g2_buf_1
Xfanout143 net144 net143 VPWR VGND sg13g2_buf_1
Xfanout132 net135 net132 VPWR VGND sg13g2_buf_1
Xfanout198 net204 net198 VPWR VGND sg13g2_buf_1
Xfanout187 net193 net187 VPWR VGND sg13g2_buf_1
Xfanout176 net178 net176 VPWR VGND sg13g2_buf_1
XFILLER_47_56 VPWR VGND sg13g2_decap_8
XFILLER_27_252 VPWR VGND sg13g2_decap_8
XFILLER_15_403 VPWR VGND sg13g2_decap_8
XFILLER_28_797 VPWR VGND sg13g2_decap_4
XFILLER_42_266 VPWR VGND sg13g2_decap_8
XFILLER_8_39 VPWR VGND sg13g2_decap_8
XFILLER_10_130 VPWR VGND sg13g2_decap_8
XFILLER_6_123 VPWR VGND sg13g2_decap_8
XFILLER_12_81 VPWR VGND sg13g2_decap_8
XFILLER_2_340 VPWR VGND sg13g2_decap_8
XFILLER_18_263 VPWR VGND sg13g2_decap_8
XFILLER_33_200 VPWR VGND sg13g2_decap_8
XFILLER_33_277 VPWR VGND sg13g2_decap_8
XFILLER_21_417 VPWR VGND sg13g2_decap_8
X_1963_ net181 _0134_ _0829_ _0830_ VPWR VGND sg13g2_a21o_1
X_1894_ net211 VPWR _0778_ VGND state\[88\] net170 sg13g2_o21ai_1
X_2515_ net382 VGND VPWR _0461_ state\[77\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2446_ net452 VGND VPWR _0392_ state\[8\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_2479__321 VPWR VGND net320 sg13g2_tiehi
X_2377_ net349 VGND VPWR _0323_ daisychain\[67\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_1328_ VPWR _0109_ state\[83\] VGND sg13g2_inv_1
XFILLER_24_200 VPWR VGND sg13g2_decap_8
XFILLER_40_737 VPWR VGND sg13g2_fill_2
XFILLER_33_25 VPWR VGND sg13g2_decap_8
XFILLER_24_277 VPWR VGND sg13g2_decap_8
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
X_2347__410 VPWR VGND net409 sg13g2_tiehi
XFILLER_4_616 VPWR VGND sg13g2_decap_8
XFILLER_3_137 VPWR VGND sg13g2_decap_8
XFILLER_0_800 VPWR VGND sg13g2_decap_8
XFILLER_0_844 VPWR VGND sg13g2_fill_2
X_2458__405 VPWR VGND net404 sg13g2_tiehi
XFILLER_48_848 VPWR VGND sg13g2_decap_4
XFILLER_47_336 VPWR VGND sg13g2_decap_8
XFILLER_15_200 VPWR VGND sg13g2_decap_8
XFILLER_15_277 VPWR VGND sg13g2_decap_8
XFILLER_31_726 VPWR VGND sg13g2_fill_2
XFILLER_30_214 VPWR VGND sg13g2_decap_8
XFILLER_11_494 VPWR VGND sg13g2_decap_8
XFILLER_8_977 VPWR VGND sg13g2_fill_2
XFILLER_7_476 VPWR VGND sg13g2_decap_8
X_2300_ _1021_ net114 state\[123\] VPWR VGND sg13g2_nand2_1
X_2231_ VGND VPWR _0779_ _0986_ _0472_ net81 sg13g2_a21oi_1
XFILLER_24_4 VPWR VGND sg13g2_decap_8
X_2162_ _0952_ net145 state\[54\] VPWR VGND sg13g2_nand2_1
XFILLER_38_336 VPWR VGND sg13g2_decap_8
X_2093_ VGND VPWR _0572_ _0917_ _0403_ net84 sg13g2_a21oi_1
XFILLER_0_1026 VPWR VGND sg13g2_fill_2
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_34_531 VPWR VGND sg13g2_decap_4
XFILLER_22_715 VPWR VGND sg13g2_decap_4
Xheichips25_pudding_488 VPWR VGND uio_oe[4] sg13g2_tiehi
XFILLER_21_214 VPWR VGND sg13g2_decap_8
XFILLER_9_60 VPWR VGND sg13g2_decap_8
X_1946_ net215 VPWR _0817_ VGND state\[101\] net181 sg13g2_o21ai_1
X_1877_ VPWR VGND _0765_ net79 _0764_ _0237_ _0339_ net35 sg13g2_a221oi_1
XdigitalenL.g\[0\].u.inv1 VPWR digitalenL.g\[0\].u.OUTN net6 VGND sg13g2_inv_1
X_2429_ net245 VGND VPWR _0375_ daisychain\[119\] clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_28_25 VPWR VGND sg13g2_decap_8
XFILLER_29_347 VPWR VGND sg13g2_decap_8
XFILLER_44_35 VPWR VGND sg13g2_decap_8
XFILLER_40_501 VPWR VGND sg13g2_fill_2
XFILLER_12_214 VPWR VGND sg13g2_decap_8
XFILLER_40_512 VPWR VGND sg13g2_decap_8
XFILLER_8_207 VPWR VGND sg13g2_decap_8
XFILLER_20_291 VPWR VGND sg13g2_decap_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_4_424 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_8
XFILLER_48_656 VPWR VGND sg13g2_decap_8
XFILLER_47_133 VPWR VGND sg13g2_decap_8
XFILLER_43_350 VPWR VGND sg13g2_decap_8
X_1800_ VGND VPWR net153 daisychain\[63\] _0708_ net63 sg13g2_a21oi_1
XFILLER_8_730 VPWR VGND sg13g2_decap_4
XFILLER_11_291 VPWR VGND sg13g2_decap_8
X_1731_ net187 _0197_ _0655_ _0656_ VPWR VGND sg13g2_a21o_1
X_1662_ net208 VPWR _0604_ VGND state\[30\] net168 sg13g2_o21ai_1
XFILLER_7_273 VPWR VGND sg13g2_decap_8
X_1593_ VPWR VGND _0552_ net73 _0551_ _0159_ _0268_ net27 sg13g2_a221oi_1
X_2214_ _0978_ net148 state\[80\] VPWR VGND sg13g2_nand2_1
XFILLER_39_634 VPWR VGND sg13g2_fill_2
X_2145_ VGND VPWR _0650_ _0943_ _0429_ net93 sg13g2_a21oi_1
XFILLER_38_133 VPWR VGND sg13g2_decap_8
X_2076_ _0909_ net116 state\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_34_361 VPWR VGND sg13g2_decap_8
XFILLER_22_567 VPWR VGND sg13g2_fill_1
X_1929_ VPWR VGND _0804_ net86 _0803_ _0251_ _0352_ net42 sg13g2_a221oi_1
XFILLER_2_906 VPWR VGND sg13g2_fill_1
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_39_35 VPWR VGND sg13g2_decap_8
XFILLER_29_144 VPWR VGND sg13g2_decap_8
XFILLER_44_147 VPWR VGND sg13g2_decap_8
XFILLER_25_361 VPWR VGND sg13g2_decap_8
XFILLER_40_364 VPWR VGND sg13g2_decap_8
XFILLER_5_722 VPWR VGND sg13g2_decap_8
XFILLER_5_711 VPWR VGND sg13g2_fill_2
XFILLER_4_221 VPWR VGND sg13g2_decap_8
XFILLER_4_298 VPWR VGND sg13g2_decap_8
XFILLER_20_81 VPWR VGND sg13g2_decap_8
XFILLER_49_932 VPWR VGND sg13g2_decap_8
XFILLER_49_921 VPWR VGND sg13g2_fill_2
XFILLER_48_420 VPWR VGND sg13g2_decap_8
XFILLER_49_998 VPWR VGND sg13g2_decap_8
XFILLER_48_497 VPWR VGND sg13g2_decap_8
XFILLER_35_147 VPWR VGND sg13g2_decap_8
XFILLER_16_361 VPWR VGND sg13g2_decap_8
X_2832_ state\[122\] net10 VPWR VGND sg13g2_buf_1
XFILLER_31_375 VPWR VGND sg13g2_decap_8
X_1714_ net218 VPWR _0643_ VGND state\[43\] net185 sg13g2_o21ai_1
XFILLER_8_593 VPWR VGND sg13g2_fill_1
X_1645_ VPWR VGND _0591_ net102 _0590_ _0173_ _0281_ net57 sg13g2_a221oi_1
X_1576_ VGND VPWR net114 daisychain\[7\] _0540_ net25 sg13g2_a21oi_1
X_2128_ _0935_ net138 state\[37\] VPWR VGND sg13g2_nand2_1
X_2059_ VGND VPWR _0521_ _0900_ _0386_ net71 sg13g2_a21oi_1
XFILLER_26_158 VPWR VGND sg13g2_decap_8
XFILLER_23_821 VPWR VGND sg13g2_fill_1
XFILLER_10_515 VPWR VGND sg13g2_decap_8
XFILLER_41_14 VPWR VGND sg13g2_decap_8
XFILLER_22_375 VPWR VGND sg13g2_decap_8
XFILLER_6_508 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_decap_8
XFILLER_49_228 VPWR VGND sg13g2_decap_8
XFILLER_18_604 VPWR VGND sg13g2_fill_2
XFILLER_45_434 VPWR VGND sg13g2_decap_8
XFILLER_17_147 VPWR VGND sg13g2_decap_8
XFILLER_33_618 VPWR VGND sg13g2_fill_1
X_2355__394 VPWR VGND net393 sg13g2_tiehi
XFILLER_45_489 VPWR VGND sg13g2_fill_1
XFILLER_13_375 VPWR VGND sg13g2_decap_8
XFILLER_15_81 VPWR VGND sg13g2_decap_8
XFILLER_41_673 VPWR VGND sg13g2_decap_8
XFILLER_40_161 VPWR VGND sg13g2_decap_8
XFILLER_9_368 VPWR VGND sg13g2_decap_8
XFILLER_5_541 VPWR VGND sg13g2_decap_8
X_1430_ VPWR _0138_ daisychain\[109\] VGND sg13g2_inv_1
X_1361_ VPWR _0073_ state\[50\] VGND sg13g2_inv_1
X_1292_ VPWR _0021_ state\[119\] VGND sg13g2_inv_1
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_31_172 VPWR VGND sg13g2_decap_8
XFILLER_11_39 VPWR VGND sg13g2_decap_8
X_1628_ VGND VPWR net118 daisychain\[20\] _0579_ net29 sg13g2_a21oi_1
X_1559_ net175 _0200_ _0526_ _0527_ VPWR VGND sg13g2_a21o_1
XFILLER_39_294 VPWR VGND sg13g2_decap_8
XFILLER_36_14 VPWR VGND sg13g2_decap_8
XFILLER_27_434 VPWR VGND sg13g2_decap_8
XFILLER_10_312 VPWR VGND sg13g2_decap_8
XFILLER_7_806 VPWR VGND sg13g2_decap_8
XFILLER_22_172 VPWR VGND sg13g2_decap_8
XFILLER_7_839 VPWR VGND sg13g2_decap_8
XFILLER_6_305 VPWR VGND sg13g2_decap_8
XFILLER_10_389 VPWR VGND sg13g2_decap_8
XFILLER_2_522 VPWR VGND sg13g2_decap_8
XFILLER_2_599 VPWR VGND sg13g2_decap_8
XFILLER_18_434 VPWR VGND sg13g2_decap_4
XFILLER_45_231 VPWR VGND sg13g2_decap_8
XFILLER_42_982 VPWR VGND sg13g2_decap_4
XFILLER_42_971 VPWR VGND sg13g2_fill_1
XFILLER_20_109 VPWR VGND sg13g2_decap_8
XFILLER_13_172 VPWR VGND sg13g2_decap_8
XFILLER_9_165 VPWR VGND sg13g2_decap_8
X_2531_ net254 VGND VPWR _0477_ state\[93\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_6_894 VPWR VGND sg13g2_fill_1
XFILLER_5_382 VPWR VGND sg13g2_decap_8
X_2462_ net388 VGND VPWR _0408_ state\[24\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2393_ net317 VGND VPWR _0339_ daisychain\[83\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1413_ VPWR _0157_ daisychain\[126\] VGND sg13g2_inv_1
X_1344_ VPWR _0091_ state\[67\] VGND sg13g2_inv_1
XFILLER_3_95 VPWR VGND sg13g2_decap_8
XFILLER_3_1013 VPWR VGND sg13g2_decap_8
XFILLER_36_231 VPWR VGND sg13g2_decap_8
X_2451__433 VPWR VGND net432 sg13g2_tiehi
XFILLER_24_437 VPWR VGND sg13g2_decap_8
XFILLER_11_109 VPWR VGND sg13g2_decap_8
XFILLER_32_470 VPWR VGND sg13g2_fill_2
XFILLER_20_676 VPWR VGND sg13g2_fill_2
XFILLER_20_687 VPWR VGND sg13g2_fill_1
XFILLER_3_319 VPWR VGND sg13g2_decap_8
Xfanout122 net137 net122 VPWR VGND sg13g2_buf_1
Xfanout111 net112 net111 VPWR VGND sg13g2_buf_1
Xfanout100 net101 net100 VPWR VGND sg13g2_buf_1
Xfanout155 net157 net155 VPWR VGND sg13g2_buf_1
Xfanout144 net147 net144 VPWR VGND sg13g2_buf_1
Xfanout133 net135 net133 VPWR VGND sg13g2_buf_1
Xfanout199 net203 net199 VPWR VGND sg13g2_buf_1
Xfanout188 net191 net188 VPWR VGND sg13g2_buf_1
Xfanout177 net178 net177 VPWR VGND sg13g2_buf_1
Xfanout166 net168 net166 VPWR VGND sg13g2_buf_1
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_27_231 VPWR VGND sg13g2_decap_8
XFILLER_42_245 VPWR VGND sg13g2_decap_8
XFILLER_8_18 VPWR VGND sg13g2_decap_8
XFILLER_11_654 VPWR VGND sg13g2_decap_4
XFILLER_10_186 VPWR VGND sg13g2_decap_8
XFILLER_6_102 VPWR VGND sg13g2_decap_8
XFILLER_12_60 VPWR VGND sg13g2_decap_8
XFILLER_6_179 VPWR VGND sg13g2_decap_8
XFILLER_2_396 VPWR VGND sg13g2_decap_8
XFILLER_19_710 VPWR VGND sg13g2_fill_1
XFILLER_18_242 VPWR VGND sg13g2_decap_8
XFILLER_46_540 VPWR VGND sg13g2_decap_8
XFILLER_34_702 VPWR VGND sg13g2_decap_4
XFILLER_34_735 VPWR VGND sg13g2_fill_1
XFILLER_33_256 VPWR VGND sg13g2_decap_8
X_1962_ net216 VPWR _0829_ VGND state\[105\] net181 sg13g2_o21ai_1
X_1893_ VPWR VGND _0777_ net83 _0776_ _0241_ _0343_ net38 sg13g2_a221oi_1
XFILLER_30_952 VPWR VGND sg13g2_decap_8
X_2514_ net390 VGND VPWR _0460_ state\[76\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_2445_ net456 VGND VPWR _0391_ state\[7\] clknet_leaf_0_clk sg13g2_dfrbpq_1
X_2376_ net351 VGND VPWR _0322_ daisychain\[66\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1327_ VPWR _0110_ state\[84\] VGND sg13g2_inv_1
XFILLER_37_551 VPWR VGND sg13g2_fill_2
XFILLER_17_49 VPWR VGND sg13g2_decap_8
XFILLER_24_256 VPWR VGND sg13g2_decap_8
XFILLER_3_116 VPWR VGND sg13g2_decap_8
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_16_702 VPWR VGND sg13g2_fill_2
XFILLER_16_724 VPWR VGND sg13g2_decap_4
XFILLER_43_521 VPWR VGND sg13g2_fill_1
XFILLER_15_256 VPWR VGND sg13g2_decap_8
XFILLER_31_716 VPWR VGND sg13g2_fill_1
XFILLER_8_923 VPWR VGND sg13g2_fill_1
XFILLER_11_473 VPWR VGND sg13g2_decap_8
XFILLER_8_956 VPWR VGND sg13g2_fill_1
XFILLER_23_81 VPWR VGND sg13g2_decap_8
XFILLER_8_989 VPWR VGND sg13g2_fill_1
XFILLER_7_455 VPWR VGND sg13g2_decap_8
XFILLER_3_650 VPWR VGND sg13g2_decap_8
X_2230_ _0986_ net125 state\[88\] VPWR VGND sg13g2_nand2_1
XFILLER_2_193 VPWR VGND sg13g2_decap_8
X_2161_ VGND VPWR _0674_ _0951_ _0437_ net98 sg13g2_a21oi_1
XFILLER_38_315 VPWR VGND sg13g2_decap_8
X_2092_ _0917_ net121 state\[19\] VPWR VGND sg13g2_nand2_1
XFILLER_19_562 VPWR VGND sg13g2_decap_4
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_46_392 VPWR VGND sg13g2_decap_8
Xheichips25_pudding_489 VPWR VGND uio_oe[5] sg13g2_tiehi
XFILLER_34_587 VPWR VGND sg13g2_decap_8
X_1945_ VPWR VGND _0816_ net89 _0815_ _0129_ _0356_ net46 sg13g2_a221oi_1
X_1876_ VGND VPWR net123 daisychain\[82\] _0765_ net35 sg13g2_a21oi_1
XdigitalenL.g\[0\].u.inv2 VPWR digitalenL.g\[0\].u.OUTP digitalenL.g\[0\].u.OUTN VGND
+ sg13g2_inv_1
XFILLER_1_609 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
X_2428_ net247 VGND VPWR _0374_ daisychain\[118\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2359_ net385 VGND VPWR _0305_ daisychain\[49\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_29_326 VPWR VGND sg13g2_decap_8
XFILLER_44_329 VPWR VGND sg13g2_decap_8
XFILLER_44_14 VPWR VGND sg13g2_decap_8
XFILLER_37_392 VPWR VGND sg13g2_decap_8
XFILLER_25_543 VPWR VGND sg13g2_decap_8
XFILLER_25_565 VPWR VGND sg13g2_decap_8
XFILLER_13_738 VPWR VGND sg13g2_fill_1
X_2314__476 VPWR VGND net475 sg13g2_tiehi
XFILLER_21_771 VPWR VGND sg13g2_fill_1
XFILLER_20_270 VPWR VGND sg13g2_decap_8
XFILLER_4_403 VPWR VGND sg13g2_decap_8
XFILLER_0_686 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_decap_8
XFILLER_35_329 VPWR VGND sg13g2_decap_8
XFILLER_29_860 VPWR VGND sg13g2_fill_1
XFILLER_18_81 VPWR VGND sg13g2_decap_8
XFILLER_31_546 VPWR VGND sg13g2_decap_8
XFILLER_11_270 VPWR VGND sg13g2_decap_8
X_1730_ net219 VPWR _0655_ VGND state\[47\] net185 sg13g2_o21ai_1
X_1661_ VPWR VGND _0603_ net75 _0602_ _0177_ _0285_ net32 sg13g2_a221oi_1
XFILLER_8_797 VPWR VGND sg13g2_fill_1
XFILLER_8_775 VPWR VGND sg13g2_fill_1
XFILLER_7_252 VPWR VGND sg13g2_decap_8
X_2365__374 VPWR VGND net373 sg13g2_tiehi
X_1592_ VGND VPWR net116 daisychain\[11\] _0552_ net27 sg13g2_a21oi_1
X_2213_ VGND VPWR _0752_ _0977_ _0463_ net104 sg13g2_a21oi_1
XFILLER_38_112 VPWR VGND sg13g2_decap_8
X_2144_ _0943_ net139 state\[45\] VPWR VGND sg13g2_nand2_1
XFILLER_39_668 VPWR VGND sg13g2_decap_8
XFILLER_39_679 VPWR VGND sg13g2_fill_2
X_2075_ VGND VPWR _0545_ _0908_ _0394_ net74 sg13g2_a21oi_1
XFILLER_47_690 VPWR VGND sg13g2_decap_8
XFILLER_38_189 VPWR VGND sg13g2_decap_8
XFILLER_34_340 VPWR VGND sg13g2_decap_8
XFILLER_14_39 VPWR VGND sg13g2_decap_8
X_1928_ VGND VPWR net129 daisychain\[95\] _0804_ net43 sg13g2_a21oi_1
X_1859_ net196 _0232_ _0751_ _0752_ VPWR VGND sg13g2_a21o_1
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_39_14 VPWR VGND sg13g2_decap_8
XFILLER_29_123 VPWR VGND sg13g2_decap_8
XFILLER_17_329 VPWR VGND sg13g2_decap_8
XFILLER_44_126 VPWR VGND sg13g2_decap_8
XFILLER_25_340 VPWR VGND sg13g2_decap_8
XFILLER_40_343 VPWR VGND sg13g2_decap_8
XFILLER_4_200 VPWR VGND sg13g2_decap_8
XFILLER_20_60 VPWR VGND sg13g2_decap_8
XFILLER_4_277 VPWR VGND sg13g2_decap_8
XFILLER_45_1006 VPWR VGND sg13g2_fill_2
XFILLER_49_900 VPWR VGND sg13g2_decap_8
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_48_476 VPWR VGND sg13g2_decap_8
XFILLER_35_126 VPWR VGND sg13g2_decap_8
XFILLER_16_340 VPWR VGND sg13g2_decap_8
X_2831_ state\[121\] net9 VPWR VGND sg13g2_buf_1
XFILLER_31_354 VPWR VGND sg13g2_decap_8
X_1713_ VPWR VGND _0642_ net94 _0641_ _0192_ _0298_ net51 sg13g2_a221oi_1
XFILLER_8_572 VPWR VGND sg13g2_decap_8
X_1644_ VGND VPWR net148 daisychain\[24\] _0591_ net57 sg13g2_a21oi_1
X_1575_ net169 _0244_ _0538_ _0539_ VPWR VGND sg13g2_a21o_1
XFILLER_6_95 VPWR VGND sg13g2_decap_8
X_2127_ VGND VPWR _0623_ _0934_ _0420_ net74 sg13g2_a21oi_1
XFILLER_26_137 VPWR VGND sg13g2_decap_8
X_2058_ _0900_ net115 state\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_22_354 VPWR VGND sg13g2_decap_8
XFILLER_1_203 VPWR VGND sg13g2_decap_8
XFILLER_2_759 VPWR VGND sg13g2_fill_1
XFILLER_49_207 VPWR VGND sg13g2_decap_8
XFILLER_17_126 VPWR VGND sg13g2_decap_8
XFILLER_46_969 VPWR VGND sg13g2_decap_8
XFILLER_45_413 VPWR VGND sg13g2_decap_8
XFILLER_13_354 VPWR VGND sg13g2_decap_8
XFILLER_15_60 VPWR VGND sg13g2_decap_8
XFILLER_40_140 VPWR VGND sg13g2_decap_8
XFILLER_9_347 VPWR VGND sg13g2_decap_8
XFILLER_5_520 VPWR VGND sg13g2_decap_8
XFILLER_31_81 VPWR VGND sg13g2_decap_8
XFILLER_5_597 VPWR VGND sg13g2_decap_8
X_1360_ VPWR _0074_ state\[51\] VGND sg13g2_inv_1
XFILLER_0_280 VPWR VGND sg13g2_decap_8
X_1291_ VPWR _0023_ state\[120\] VGND sg13g2_inv_1
XFILLER_49_752 VPWR VGND sg13g2_decap_8
XFILLER_49_785 VPWR VGND sg13g2_decap_8
XFILLER_49_763 VPWR VGND sg13g2_fill_1
XFILLER_48_273 VPWR VGND sg13g2_decap_8
XFILLER_36_413 VPWR VGND sg13g2_decap_4
XFILLER_36_479 VPWR VGND sg13g2_decap_8
XFILLER_31_151 VPWR VGND sg13g2_decap_8
XFILLER_11_18 VPWR VGND sg13g2_decap_8
X_1627_ net165 _0169_ _0577_ _0578_ VPWR VGND sg13g2_a21o_1
X_1558_ net207 VPWR _0526_ VGND state\[4\] net165 sg13g2_o21ai_1
X_1489_ VPWR _0201_ daisychain\[50\] VGND sg13g2_inv_1
XFILLER_39_273 VPWR VGND sg13g2_decap_8
XFILLER_27_413 VPWR VGND sg13g2_decap_8
XFILLER_22_151 VPWR VGND sg13g2_decap_8
XFILLER_10_368 VPWR VGND sg13g2_decap_8
XFILLER_2_501 VPWR VGND sg13g2_decap_8
XFILLER_2_578 VPWR VGND sg13g2_decap_8
XFILLER_46_700 VPWR VGND sg13g2_fill_2
XFILLER_18_413 VPWR VGND sg13g2_decap_8
XFILLER_45_210 VPWR VGND sg13g2_decap_8
XFILLER_19_947 VPWR VGND sg13g2_decap_8
XFILLER_19_936 VPWR VGND sg13g2_fill_1
XFILLER_45_287 VPWR VGND sg13g2_decap_8
XFILLER_14_630 VPWR VGND sg13g2_decap_8
XFILLER_26_81 VPWR VGND sg13g2_decap_8
XFILLER_13_151 VPWR VGND sg13g2_decap_8
XFILLER_14_685 VPWR VGND sg13g2_decap_8
XFILLER_9_144 VPWR VGND sg13g2_decap_8
XFILLER_42_91 VPWR VGND sg13g2_decap_8
X_2530_ net262 VGND VPWR _0476_ state\[92\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_2461_ net392 VGND VPWR _0407_ state\[23\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_5_361 VPWR VGND sg13g2_decap_8
X_1412_ VPWR _0158_ daisychain\[127\] VGND sg13g2_inv_1
X_2392_ net319 VGND VPWR _0338_ daisychain\[82\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_1343_ VPWR _0092_ state\[68\] VGND sg13g2_inv_1
XFILLER_3_74 VPWR VGND sg13g2_decap_8
XFILLER_49_571 VPWR VGND sg13g2_fill_2
XFILLER_36_210 VPWR VGND sg13g2_decap_8
XFILLER_36_287 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_16_clk clknet_2_2__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
XFILLER_32_482 VPWR VGND sg13g2_decap_8
XFILLER_22_39 VPWR VGND sg13g2_decap_8
XFILLER_20_699 VPWR VGND sg13g2_fill_1
Xfanout112 _0512_ net112 VPWR VGND sg13g2_buf_1
Xfanout101 net112 net101 VPWR VGND sg13g2_buf_1
Xfanout156 net157 net156 VPWR VGND sg13g2_buf_1
Xfanout145 net147 net145 VPWR VGND sg13g2_buf_1
Xfanout134 net135 net134 VPWR VGND sg13g2_buf_1
Xfanout123 net125 net123 VPWR VGND sg13g2_buf_1
Xfanout189 net191 net189 VPWR VGND sg13g2_buf_1
Xfanout178 net183 net178 VPWR VGND sg13g2_buf_1
Xfanout167 net168 net167 VPWR VGND sg13g2_buf_1
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_27_210 VPWR VGND sg13g2_decap_8
XFILLER_15_438 VPWR VGND sg13g2_decap_8
XFILLER_42_224 VPWR VGND sg13g2_decap_8
XFILLER_27_287 VPWR VGND sg13g2_decap_8
XFILLER_24_950 VPWR VGND sg13g2_decap_4
XFILLER_24_994 VPWR VGND sg13g2_decap_4
XFILLER_10_165 VPWR VGND sg13g2_decap_8
XFILLER_6_158 VPWR VGND sg13g2_decap_8
XFILLER_3_865 VPWR VGND sg13g2_fill_2
X_2324__456 VPWR VGND net455 sg13g2_tiehi
XFILLER_2_375 VPWR VGND sg13g2_decap_8
XFILLER_18_221 VPWR VGND sg13g2_decap_8
XFILLER_37_91 VPWR VGND sg13g2_decap_8
XFILLER_19_799 VPWR VGND sg13g2_fill_2
XFILLER_18_298 VPWR VGND sg13g2_decap_8
XFILLER_33_235 VPWR VGND sg13g2_decap_8
X_1961_ VPWR VGND _0828_ net89 _0827_ _0133_ _0360_ net46 sg13g2_a221oi_1
X_1892_ VGND VPWR net127 daisychain\[86\] _0777_ net38 sg13g2_a21oi_1
X_2513_ net398 VGND VPWR _0459_ state\[75\] clknet_leaf_12_clk sg13g2_dfrbpq_1
X_2444_ net460 VGND VPWR _0390_ state\[6\] clknet_leaf_0_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_5_clk clknet_2_1__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_2375_ net353 VGND VPWR _0321_ daisychain\[65\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_38_0 VPWR VGND sg13g2_decap_8
X_1326_ VPWR _0111_ state\[85\] VGND sg13g2_inv_1
XFILLER_17_28 VPWR VGND sg13g2_decap_8
X_2375__354 VPWR VGND net353 sg13g2_tiehi
XFILLER_24_235 VPWR VGND sg13g2_decap_8
X_2562__259 VPWR VGND net258 sg13g2_tiehi
XFILLER_0_846 VPWR VGND sg13g2_fill_1
XFILLER_15_235 VPWR VGND sg13g2_decap_8
XFILLER_43_533 VPWR VGND sg13g2_decap_8
XFILLER_8_902 VPWR VGND sg13g2_fill_1
XFILLER_30_249 VPWR VGND sg13g2_decap_8
XFILLER_11_452 VPWR VGND sg13g2_decap_8
XFILLER_8_935 VPWR VGND sg13g2_fill_1
XFILLER_23_60 VPWR VGND sg13g2_decap_8
XFILLER_8_968 VPWR VGND sg13g2_fill_1
XFILLER_7_434 VPWR VGND sg13g2_decap_8
XFILLER_2_172 VPWR VGND sg13g2_decap_8
X_2160_ _0951_ net143 state\[53\] VPWR VGND sg13g2_nand2_1
X_2091_ VGND VPWR _0569_ _0916_ _0402_ net85 sg13g2_a21oi_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_19_552 VPWR VGND sg13g2_decap_4
XFILLER_0_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_371 VPWR VGND sg13g2_decap_8
XFILLER_19_585 VPWR VGND sg13g2_decap_4
X_1944_ VGND VPWR net133 daisychain\[99\] _0816_ net46 sg13g2_a21oi_1
XFILLER_21_249 VPWR VGND sg13g2_decap_8
XFILLER_9_95 VPWR VGND sg13g2_decap_8
X_1875_ net172 _0237_ _0763_ _0764_ VPWR VGND sg13g2_a21o_1
XFILLER_7_990 VPWR VGND sg13g2_decap_8
X_2427_ net249 VGND VPWR _0373_ daisychain\[117\] clknet_leaf_4_clk sg13g2_dfrbpq_1
X_2358_ net387 VGND VPWR _0304_ daisychain\[48\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_29_305 VPWR VGND sg13g2_decap_8
X_2289_ VGND VPWR _0866_ _1015_ _0501_ net82 sg13g2_a21oi_1
X_1309_ VPWR _0003_ state\[102\] VGND sg13g2_inv_1
XFILLER_44_308 VPWR VGND sg13g2_decap_8
XFILLER_37_371 VPWR VGND sg13g2_decap_8
XFILLER_12_249 VPWR VGND sg13g2_decap_8
XFILLER_40_547 VPWR VGND sg13g2_fill_1
X_2505__463 VPWR VGND net462 sg13g2_tiehi
XFILLER_4_459 VPWR VGND sg13g2_decap_8
XFILLER_0_665 VPWR VGND sg13g2_decap_8
XFILLER_18_60 VPWR VGND sg13g2_decap_8
XFILLER_47_168 VPWR VGND sg13g2_decap_8
XFILLER_35_308 VPWR VGND sg13g2_decap_8
XFILLER_44_820 VPWR VGND sg13g2_fill_1
XFILLER_28_382 VPWR VGND sg13g2_decap_8
XFILLER_44_886 VPWR VGND sg13g2_fill_2
XFILLER_43_385 VPWR VGND sg13g2_decap_8
XFILLER_31_536 VPWR VGND sg13g2_fill_2
XFILLER_31_525 VPWR VGND sg13g2_decap_8
XFILLER_31_503 VPWR VGND sg13g2_fill_2
XFILLER_34_81 VPWR VGND sg13g2_decap_8
XFILLER_8_754 VPWR VGND sg13g2_fill_2
XFILLER_7_231 VPWR VGND sg13g2_decap_8
X_1660_ VGND VPWR net118 daisychain\[28\] _0603_ net29 sg13g2_a21oi_1
XFILLER_8_787 VPWR VGND sg13g2_decap_8
X_1591_ net162 _0159_ _0550_ _0551_ VPWR VGND sg13g2_a21o_1
XFILLER_4_982 VPWR VGND sg13g2_decap_8
X_2212_ _0977_ net150 state\[79\] VPWR VGND sg13g2_nand2_1
X_2143_ VGND VPWR _0647_ _0942_ _0428_ net93 sg13g2_a21oi_1
XFILLER_22_1018 VPWR VGND sg13g2_decap_8
XFILLER_38_168 VPWR VGND sg13g2_decap_8
XFILLER_26_319 VPWR VGND sg13g2_decap_8
XFILLER_19_382 VPWR VGND sg13g2_decap_8
X_2074_ _0908_ net117 state\[10\] VPWR VGND sg13g2_nand2_1
X_2517__367 VPWR VGND net366 sg13g2_tiehi
XFILLER_14_18 VPWR VGND sg13g2_decap_8
XFILLER_22_503 VPWR VGND sg13g2_decap_8
XFILLER_34_396 VPWR VGND sg13g2_decap_8
XFILLER_22_558 VPWR VGND sg13g2_fill_2
X_1927_ net177 _0251_ _0802_ _0803_ VPWR VGND sg13g2_a21o_1
XFILLER_30_591 VPWR VGND sg13g2_fill_1
X_1858_ net224 VPWR _0751_ VGND state\[79\] net196 sg13g2_o21ai_1
XFILLER_30_39 VPWR VGND sg13g2_decap_8
X_1789_ VPWR VGND _0699_ net100 _0698_ _0213_ _0317_ net54 sg13g2_a221oi_1
XFILLER_2_919 VPWR VGND sg13g2_decap_8
XFILLER_29_102 VPWR VGND sg13g2_decap_8
XFILLER_18_809 VPWR VGND sg13g2_fill_1
XFILLER_17_308 VPWR VGND sg13g2_decap_8
XFILLER_29_179 VPWR VGND sg13g2_decap_8
XFILLER_44_105 VPWR VGND sg13g2_decap_8
XFILLER_13_558 VPWR VGND sg13g2_decap_8
XFILLER_40_322 VPWR VGND sg13g2_decap_8
XFILLER_25_396 VPWR VGND sg13g2_decap_8
XFILLER_9_529 VPWR VGND sg13g2_decap_8
XFILLER_40_399 VPWR VGND sg13g2_decap_8
XFILLER_5_713 VPWR VGND sg13g2_fill_1
XFILLER_5_768 VPWR VGND sg13g2_decap_4
XFILLER_4_256 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_49_923 VPWR VGND sg13g2_fill_1
XFILLER_48_455 VPWR VGND sg13g2_decap_8
XFILLER_29_81 VPWR VGND sg13g2_decap_8
XFILLER_35_105 VPWR VGND sg13g2_decap_8
XFILLER_29_691 VPWR VGND sg13g2_decap_8
XFILLER_45_91 VPWR VGND sg13g2_decap_8
XFILLER_32_801 VPWR VGND sg13g2_fill_2
XFILLER_16_396 VPWR VGND sg13g2_decap_8
X_2830_ state\[120\] net8 VPWR VGND sg13g2_buf_1
XFILLER_43_182 VPWR VGND sg13g2_decap_8
XFILLER_31_333 VPWR VGND sg13g2_decap_8
X_1712_ VGND VPWR net140 daisychain\[41\] _0642_ net51 sg13g2_a21oi_1
XFILLER_8_551 VPWR VGND sg13g2_decap_8
XANTENNA_1 VPWR VGND _0131_ sg13g2_antennanp
X_1643_ net194 _0173_ _0589_ _0590_ VPWR VGND sg13g2_a21o_1
XFILLER_6_74 VPWR VGND sg13g2_decap_8
X_1574_ net206 VPWR _0538_ VGND state\[8\] net169 sg13g2_o21ai_1
XFILLER_6_1023 VPWR VGND sg13g2_decap_4
XFILLER_39_433 VPWR VGND sg13g2_decap_8
XFILLER_39_466 VPWR VGND sg13g2_decap_8
XFILLER_27_606 VPWR VGND sg13g2_fill_2
X_2126_ _0934_ net117 state\[36\] VPWR VGND sg13g2_nand2_1
X_2454__421 VPWR VGND net420 sg13g2_tiehi
XFILLER_27_639 VPWR VGND sg13g2_fill_1
XFILLER_26_116 VPWR VGND sg13g2_decap_8
X_2057_ VGND VPWR _0518_ _0899_ _0385_ net80 sg13g2_a21oi_1
XFILLER_41_119 VPWR VGND sg13g2_decap_8
XFILLER_35_683 VPWR VGND sg13g2_fill_1
XFILLER_25_39 VPWR VGND sg13g2_decap_8
XFILLER_23_812 VPWR VGND sg13g2_decap_8
XFILLER_23_801 VPWR VGND sg13g2_fill_2
XFILLER_34_193 VPWR VGND sg13g2_decap_8
XFILLER_22_333 VPWR VGND sg13g2_decap_8
XFILLER_41_49 VPWR VGND sg13g2_decap_8
XFILLER_2_716 VPWR VGND sg13g2_fill_1
XFILLER_1_259 VPWR VGND sg13g2_decap_8
XFILLER_46_915 VPWR VGND sg13g2_fill_2
XFILLER_46_904 VPWR VGND sg13g2_decap_8
XFILLER_17_105 VPWR VGND sg13g2_decap_8
XFILLER_46_937 VPWR VGND sg13g2_fill_2
XFILLER_26_672 VPWR VGND sg13g2_fill_2
XFILLER_13_333 VPWR VGND sg13g2_decap_8
XFILLER_26_694 VPWR VGND sg13g2_decap_8
XFILLER_25_193 VPWR VGND sg13g2_decap_8
XFILLER_41_686 VPWR VGND sg13g2_decap_8
XFILLER_9_326 VPWR VGND sg13g2_decap_8
XFILLER_40_196 VPWR VGND sg13g2_decap_8
XFILLER_31_60 VPWR VGND sg13g2_decap_8
XFILLER_5_576 VPWR VGND sg13g2_decap_8
X_1290_ VPWR _0024_ state\[121\] VGND sg13g2_inv_1
XFILLER_49_720 VPWR VGND sg13g2_decap_8
XFILLER_48_252 VPWR VGND sg13g2_decap_8
XFILLER_36_458 VPWR VGND sg13g2_fill_1
X_2334__436 VPWR VGND net435 sg13g2_tiehi
XFILLER_16_193 VPWR VGND sg13g2_decap_8
XFILLER_44_491 VPWR VGND sg13g2_decap_8
XFILLER_31_130 VPWR VGND sg13g2_decap_8
X_1626_ net207 VPWR _0577_ VGND state\[21\] net165 sg13g2_o21ai_1
X_1557_ VPWR VGND _0525_ net80 _0524_ _0189_ _0259_ net34 sg13g2_a221oi_1
X_1488_ VPWR _0202_ daisychain\[51\] VGND sg13g2_inv_1
XFILLER_39_252 VPWR VGND sg13g2_decap_8
XFILLER_15_609 VPWR VGND sg13g2_decap_8
X_2109_ VGND VPWR _0596_ _0925_ _0411_ net76 sg13g2_a21oi_1
XFILLER_36_49 VPWR VGND sg13g2_decap_8
XFILLER_42_406 VPWR VGND sg13g2_decap_8
XFILLER_35_480 VPWR VGND sg13g2_fill_1
XFILLER_23_631 VPWR VGND sg13g2_fill_2
XFILLER_23_620 VPWR VGND sg13g2_decap_8
XFILLER_23_653 VPWR VGND sg13g2_fill_2
XFILLER_22_130 VPWR VGND sg13g2_decap_8
XFILLER_23_697 VPWR VGND sg13g2_decap_8
XFILLER_10_347 VPWR VGND sg13g2_decap_8
X_2385__334 VPWR VGND net333 sg13g2_tiehi
XFILLER_2_557 VPWR VGND sg13g2_decap_8
XFILLER_18_447 VPWR VGND sg13g2_decap_8
XFILLER_46_756 VPWR VGND sg13g2_fill_1
XFILLER_45_266 VPWR VGND sg13g2_decap_8
XFILLER_33_417 VPWR VGND sg13g2_decap_4
XFILLER_26_60 VPWR VGND sg13g2_decap_8
XFILLER_13_130 VPWR VGND sg13g2_decap_8
XFILLER_9_123 VPWR VGND sg13g2_decap_8
XFILLER_42_70 VPWR VGND sg13g2_decap_8
XFILLER_5_340 VPWR VGND sg13g2_decap_8
X_2460_ net396 VGND VPWR _0406_ state\[22\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_1411_ VPWR _0000_ state\[0\] VGND sg13g2_inv_1
X_2391_ net321 VGND VPWR _0337_ daisychain\[81\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1342_ VPWR _0093_ state\[69\] VGND sg13g2_inv_1
XFILLER_3_53 VPWR VGND sg13g2_decap_8
XFILLER_36_266 VPWR VGND sg13g2_decap_8
XFILLER_24_417 VPWR VGND sg13g2_decap_8
XFILLER_32_472 VPWR VGND sg13g2_fill_1
XFILLER_22_18 VPWR VGND sg13g2_decap_8
X_1609_ VPWR VGND _0564_ net85 _0563_ _0163_ _0272_ net42 sg13g2_a221oi_1
Xfanout113 net115 net113 VPWR VGND sg13g2_buf_1
Xfanout102 net103 net102 VPWR VGND sg13g2_buf_1
Xfanout146 net147 net146 VPWR VGND sg13g2_buf_1
Xfanout135 net136 net135 VPWR VGND sg13g2_buf_1
Xfanout124 net125 net124 VPWR VGND sg13g2_buf_1
Xfanout179 net182 net179 VPWR VGND sg13g2_buf_1
Xfanout168 net169 net168 VPWR VGND sg13g2_buf_1
Xfanout157 net158 net157 VPWR VGND sg13g2_buf_1
XFILLER_28_701 VPWR VGND sg13g2_fill_2
XFILLER_15_417 VPWR VGND sg13g2_decap_8
XFILLER_42_203 VPWR VGND sg13g2_decap_8
XFILLER_27_266 VPWR VGND sg13g2_decap_8
XFILLER_23_483 VPWR VGND sg13g2_decap_4
XFILLER_10_144 VPWR VGND sg13g2_decap_8
XFILLER_6_137 VPWR VGND sg13g2_decap_8
XFILLER_12_95 VPWR VGND sg13g2_decap_8
XFILLER_3_833 VPWR VGND sg13g2_fill_1
XFILLER_2_354 VPWR VGND sg13g2_decap_8
XFILLER_18_200 VPWR VGND sg13g2_decap_8
XFILLER_18_277 VPWR VGND sg13g2_decap_8
XFILLER_37_70 VPWR VGND sg13g2_decap_8
XFILLER_33_214 VPWR VGND sg13g2_decap_8
X_1960_ VGND VPWR net133 daisychain\[103\] _0828_ net46 sg13g2_a21oi_1
XFILLER_30_921 VPWR VGND sg13g2_decap_4
X_1891_ net173 _0241_ _0775_ _0776_ VPWR VGND sg13g2_a21o_1
XFILLER_41_280 VPWR VGND sg13g2_decap_8
X_2512_ net406 VGND VPWR _0458_ state\[74\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_2443_ net464 VGND VPWR _0389_ state\[5\] clknet_leaf_1_clk sg13g2_dfrbpq_1
X_2374_ net355 VGND VPWR _0320_ daisychain\[64\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1325_ VPWR _0112_ state\[86\] VGND sg13g2_inv_1
XFILLER_37_564 VPWR VGND sg13g2_decap_8
XFILLER_25_737 VPWR VGND sg13g2_fill_1
XFILLER_24_214 VPWR VGND sg13g2_decap_8
XFILLER_33_39 VPWR VGND sg13g2_decap_8
XFILLER_21_910 VPWR VGND sg13g2_decap_8
XFILLER_32_291 VPWR VGND sg13g2_decap_8
XFILLER_20_431 VPWR VGND sg13g2_decap_8
XFILLER_0_814 VPWR VGND sg13g2_fill_2
XFILLER_15_214 VPWR VGND sg13g2_decap_8
XFILLER_43_512 VPWR VGND sg13g2_fill_1
XFILLER_30_228 VPWR VGND sg13g2_decap_8
XFILLER_11_431 VPWR VGND sg13g2_decap_8
XFILLER_8_914 VPWR VGND sg13g2_fill_2
XFILLER_23_291 VPWR VGND sg13g2_decap_8
XFILLER_8_947 VPWR VGND sg13g2_fill_2
XFILLER_7_413 VPWR VGND sg13g2_decap_8
XFILLER_3_696 VPWR VGND sg13g2_decap_8
XFILLER_2_151 VPWR VGND sg13g2_decap_8
X_2090_ _0916_ net129 state\[18\] VPWR VGND sg13g2_nand2_1
XFILLER_48_91 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_46_350 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_21_228 VPWR VGND sg13g2_decap_8
XFILLER_14_291 VPWR VGND sg13g2_decap_8
X_1943_ net180 _0129_ _0814_ _0815_ VPWR VGND sg13g2_a21o_1
X_2411__282 VPWR VGND net281 sg13g2_tiehi
XFILLER_9_74 VPWR VGND sg13g2_decap_8
XFILLER_30_784 VPWR VGND sg13g2_decap_8
X_1874_ net211 VPWR _0763_ VGND state\[83\] net172 sg13g2_o21ai_1
X_2426_ net251 VGND VPWR _0372_ daisychain\[116\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2357_ net389 VGND VPWR _0303_ daisychain\[47\] clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_28_39 VPWR VGND sg13g2_decap_8
X_2288_ _1015_ net136 state\[117\] VPWR VGND sg13g2_nand2_1
X_1308_ VPWR _0004_ state\[103\] VGND sg13g2_inv_1
XFILLER_37_350 VPWR VGND sg13g2_decap_8
XFILLER_25_523 VPWR VGND sg13g2_decap_8
XFILLER_44_49 VPWR VGND sg13g2_decap_8
XFILLER_13_729 VPWR VGND sg13g2_decap_8
XFILLER_40_526 VPWR VGND sg13g2_decap_4
XFILLER_12_228 VPWR VGND sg13g2_decap_8
XFILLER_21_762 VPWR VGND sg13g2_decap_8
XFILLER_4_438 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_decap_8
XFILLER_29_851 VPWR VGND sg13g2_decap_8
XFILLER_16_523 VPWR VGND sg13g2_decap_8
XFILLER_16_534 VPWR VGND sg13g2_fill_1
XFILLER_28_361 VPWR VGND sg13g2_decap_8
XFILLER_16_589 VPWR VGND sg13g2_fill_2
XFILLER_43_364 VPWR VGND sg13g2_decap_8
XFILLER_34_60 VPWR VGND sg13g2_decap_8
XFILLER_8_744 VPWR VGND sg13g2_decap_8
XFILLER_7_210 VPWR VGND sg13g2_decap_8
XFILLER_8_766 VPWR VGND sg13g2_fill_2
X_1590_ net206 VPWR _0550_ VGND state\[12\] net162 sg13g2_o21ai_1
XFILLER_7_287 VPWR VGND sg13g2_decap_8
XFILLER_3_482 VPWR VGND sg13g2_decap_8
X_2211_ VGND VPWR _0749_ _0976_ _0462_ net104 sg13g2_a21oi_1
XFILLER_22_4 VPWR VGND sg13g2_decap_8
X_2142_ _0942_ net139 state\[44\] VPWR VGND sg13g2_nand2_1
X_2073_ VGND VPWR _0542_ _0907_ _0393_ net74 sg13g2_a21oi_1
XFILLER_38_147 VPWR VGND sg13g2_decap_8
XFILLER_19_361 VPWR VGND sg13g2_decap_8
XFILLER_34_375 VPWR VGND sg13g2_decap_8
X_1926_ net214 VPWR _0802_ VGND state\[96\] net177 sg13g2_o21ai_1
X_1857_ VPWR VGND _0750_ net105 _0749_ _0231_ _0334_ net60 sg13g2_a221oi_1
XFILLER_30_18 VPWR VGND sg13g2_decap_8
X_2344__416 VPWR VGND net415 sg13g2_tiehi
X_1788_ VGND VPWR net146 daisychain\[60\] _0699_ net54 sg13g2_a21oi_1
X_2409_ net285 VGND VPWR _0355_ daisychain\[99\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_39_49 VPWR VGND sg13g2_decap_8
XFILLER_29_158 VPWR VGND sg13g2_decap_8
XFILLER_26_854 VPWR VGND sg13g2_decap_4
XFILLER_40_301 VPWR VGND sg13g2_decap_8
XFILLER_25_375 VPWR VGND sg13g2_decap_8
XFILLER_9_508 VPWR VGND sg13g2_decap_8
XFILLER_40_378 VPWR VGND sg13g2_decap_8
XFILLER_5_703 VPWR VGND sg13g2_fill_2
XFILLER_5_736 VPWR VGND sg13g2_fill_2
XFILLER_4_235 VPWR VGND sg13g2_decap_8
XFILLER_20_95 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
X_2395__314 VPWR VGND net313 sg13g2_tiehi
XFILLER_49_968 VPWR VGND sg13g2_fill_2
XFILLER_49_957 VPWR VGND sg13g2_decap_8
XFILLER_49_946 VPWR VGND sg13g2_decap_4
XFILLER_48_434 VPWR VGND sg13g2_decap_8
XFILLER_29_60 VPWR VGND sg13g2_decap_8
XFILLER_49_979 VPWR VGND sg13g2_fill_1
XFILLER_36_618 VPWR VGND sg13g2_decap_4
XFILLER_16_375 VPWR VGND sg13g2_decap_8
XFILLER_45_70 VPWR VGND sg13g2_decap_8
XFILLER_43_161 VPWR VGND sg13g2_decap_8
XFILLER_31_312 VPWR VGND sg13g2_decap_8
XFILLER_8_530 VPWR VGND sg13g2_decap_8
XFILLER_31_389 VPWR VGND sg13g2_decap_8
X_1711_ net184 _0192_ _0640_ _0641_ VPWR VGND sg13g2_a21o_1
XANTENNA_2 VPWR VGND _0144_ sg13g2_antennanp
X_1642_ net223 VPWR _0589_ VGND state\[25\] net194 sg13g2_o21ai_1
XFILLER_6_53 VPWR VGND sg13g2_decap_8
X_1573_ VPWR VGND _0537_ net70 _0536_ _0233_ _0263_ net26 sg13g2_a221oi_1
XFILLER_39_456 VPWR VGND sg13g2_fill_1
X_2125_ VGND VPWR _0620_ _0933_ _0419_ net92 sg13g2_a21oi_1
X_2056_ _0899_ net124 state\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_25_18 VPWR VGND sg13g2_decap_8
XFILLER_35_695 VPWR VGND sg13g2_decap_8
XFILLER_34_172 VPWR VGND sg13g2_decap_8
XFILLER_23_857 VPWR VGND sg13g2_decap_4
XFILLER_22_312 VPWR VGND sg13g2_decap_8
XFILLER_23_868 VPWR VGND sg13g2_decap_4
XFILLER_10_529 VPWR VGND sg13g2_decap_8
XFILLER_41_28 VPWR VGND sg13g2_decap_8
XFILLER_22_389 VPWR VGND sg13g2_decap_8
X_1909_ VPWR VGND _0789_ net105 _0788_ _0246_ _0347_ net60 sg13g2_a221oi_1
XFILLER_2_706 VPWR VGND sg13g2_fill_1
XFILLER_2_728 VPWR VGND sg13g2_decap_8
XFILLER_1_238 VPWR VGND sg13g2_decap_8
XFILLER_18_618 VPWR VGND sg13g2_fill_2
XFILLER_45_448 VPWR VGND sg13g2_decap_8
XFILLER_32_109 VPWR VGND sg13g2_decap_8
XFILLER_13_312 VPWR VGND sg13g2_decap_8
XFILLER_25_172 VPWR VGND sg13g2_decap_8
XFILLER_9_305 VPWR VGND sg13g2_decap_8
XFILLER_13_389 VPWR VGND sg13g2_decap_8
XFILLER_15_95 VPWR VGND sg13g2_decap_8
XFILLER_40_175 VPWR VGND sg13g2_decap_8
XFILLER_5_555 VPWR VGND sg13g2_decap_8
XFILLER_1_750 VPWR VGND sg13g2_fill_1
XFILLER_48_231 VPWR VGND sg13g2_decap_8
XFILLER_23_109 VPWR VGND sg13g2_decap_8
XFILLER_16_172 VPWR VGND sg13g2_decap_8
XFILLER_32_698 VPWR VGND sg13g2_decap_8
XFILLER_31_186 VPWR VGND sg13g2_decap_8
XFILLER_8_382 VPWR VGND sg13g2_decap_8
X_1625_ VPWR VGND _0576_ net75 _0575_ _0168_ _0276_ net29 sg13g2_a221oi_1
X_1556_ VGND VPWR net124 daisychain\[2\] _0525_ net34 sg13g2_a21oi_1
X_2558__243 VPWR VGND net242 sg13g2_tiehi
X_1487_ VPWR _0203_ daisychain\[52\] VGND sg13g2_inv_1
XFILLER_39_231 VPWR VGND sg13g2_decap_8
XFILLER_28_916 VPWR VGND sg13g2_fill_2
XFILLER_36_28 VPWR VGND sg13g2_decap_8
X_2108_ _0925_ net119 state\[27\] VPWR VGND sg13g2_nand2_1
XFILLER_27_448 VPWR VGND sg13g2_fill_2
XFILLER_14_109 VPWR VGND sg13g2_decap_8
X_2039_ net161 _0155_ _0886_ _0887_ VPWR VGND sg13g2_a21o_1
XFILLER_42_429 VPWR VGND sg13g2_decap_8
XFILLER_10_326 VPWR VGND sg13g2_decap_8
XFILLER_22_186 VPWR VGND sg13g2_decap_8
XFILLER_6_319 VPWR VGND sg13g2_decap_8
XFILLER_2_536 VPWR VGND sg13g2_decap_8
XFILLER_46_713 VPWR VGND sg13g2_fill_2
XFILLER_18_459 VPWR VGND sg13g2_decap_4
XFILLER_45_245 VPWR VGND sg13g2_decap_8
XFILLER_14_665 VPWR VGND sg13g2_fill_2
XFILLER_9_102 VPWR VGND sg13g2_decap_8
XFILLER_13_186 VPWR VGND sg13g2_decap_8
XFILLER_9_179 VPWR VGND sg13g2_decap_8
XFILLER_6_853 VPWR VGND sg13g2_decap_8
X_1410_ VPWR _0039_ state\[1\] VGND sg13g2_inv_1
XFILLER_5_396 VPWR VGND sg13g2_decap_8
X_2390_ net323 VGND VPWR _0336_ daisychain\[80\] clknet_leaf_9_clk sg13g2_dfrbpq_1
X_1341_ VPWR _0095_ state\[70\] VGND sg13g2_inv_1
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_3_1027 VPWR VGND sg13g2_fill_2
XFILLER_25_908 VPWR VGND sg13g2_decap_8
XFILLER_18_960 VPWR VGND sg13g2_fill_1
XFILLER_36_245 VPWR VGND sg13g2_decap_8
XFILLER_17_470 VPWR VGND sg13g2_fill_1
XFILLER_45_790 VPWR VGND sg13g2_fill_1
XFILLER_9_691 VPWR VGND sg13g2_decap_8
X_2564__291 VPWR VGND net290 sg13g2_tiehi
X_1608_ VGND VPWR net129 daisychain\[15\] _0564_ net42 sg13g2_a21oi_1
Xfanout103 net111 net103 VPWR VGND sg13g2_buf_1
X_2421__262 VPWR VGND net261 sg13g2_tiehi
Xfanout147 net158 net147 VPWR VGND sg13g2_buf_1
Xfanout136 net137 net136 VPWR VGND sg13g2_buf_1
Xfanout125 net136 net125 VPWR VGND sg13g2_buf_1
Xfanout114 net115 net114 VPWR VGND sg13g2_buf_1
XdigitalenL.g\[3\].u.inv1 VPWR digitalenL.g\[3\].u.OUTN net6 VGND sg13g2_inv_1
X_1539_ VPWR _0128_ daisychain\[0\] VGND sg13g2_inv_1
Xfanout169 net204 net169 VPWR VGND sg13g2_buf_1
Xfanout158 _1026_ net158 VPWR VGND sg13g2_buf_1
XFILLER_47_49 VPWR VGND sg13g2_decap_8
XFILLER_43_727 VPWR VGND sg13g2_decap_4
XFILLER_27_245 VPWR VGND sg13g2_decap_8
XFILLER_42_259 VPWR VGND sg13g2_decap_8
XFILLER_10_123 VPWR VGND sg13g2_decap_8
XFILLER_6_116 VPWR VGND sg13g2_decap_8
XFILLER_12_74 VPWR VGND sg13g2_decap_8
XFILLER_3_867 VPWR VGND sg13g2_fill_1
XFILLER_2_333 VPWR VGND sg13g2_decap_8
XFILLER_18_256 VPWR VGND sg13g2_decap_8
XFILLER_19_768 VPWR VGND sg13g2_fill_2
XFILLER_42_760 VPWR VGND sg13g2_decap_8
XFILLER_30_933 VPWR VGND sg13g2_fill_2
X_1890_ net212 VPWR _0775_ VGND state\[87\] net173 sg13g2_o21ai_1
XFILLER_42_793 VPWR VGND sg13g2_fill_1
XFILLER_30_988 VPWR VGND sg13g2_decap_8
X_2511_ net414 VGND VPWR _0457_ state\[73\] clknet_leaf_10_clk sg13g2_dfrbpq_1
X_2442_ net468 VGND VPWR _0388_ state\[4\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_5_193 VPWR VGND sg13g2_decap_8
X_2373_ net357 VGND VPWR _0319_ daisychain\[63\] clknet_leaf_11_clk sg13g2_dfrbpq_1
X_1324_ VPWR _0113_ state\[87\] VGND sg13g2_inv_1
XFILLER_33_18 VPWR VGND sg13g2_decap_8
XFILLER_32_270 VPWR VGND sg13g2_decap_8
XFILLER_20_410 VPWR VGND sg13g2_decap_8
XFILLER_20_476 VPWR VGND sg13g2_decap_4
XFILLER_4_609 VPWR VGND sg13g2_decap_8
XFILLER_0_837 VPWR VGND sg13g2_decap_8
XFILLER_47_329 VPWR VGND sg13g2_decap_8
XFILLER_30_207 VPWR VGND sg13g2_decap_8
XFILLER_11_410 VPWR VGND sg13g2_decap_8
XFILLER_23_270 VPWR VGND sg13g2_decap_8
XFILLER_11_487 VPWR VGND sg13g2_decap_8
XFILLER_23_95 VPWR VGND sg13g2_decap_8
XFILLER_7_469 VPWR VGND sg13g2_decap_8
XFILLER_3_664 VPWR VGND sg13g2_decap_4
XFILLER_2_130 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_17_7 VPWR VGND sg13g2_decap_8
XFILLER_38_329 VPWR VGND sg13g2_decap_8
XFILLER_0_1019 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_34_524 VPWR VGND sg13g2_decap_8
XFILLER_21_207 VPWR VGND sg13g2_decap_8
XFILLER_14_270 VPWR VGND sg13g2_decap_8
X_1942_ net215 VPWR _0814_ VGND state\[100\] net180 sg13g2_o21ai_1
XFILLER_9_53 VPWR VGND sg13g2_decap_8
XFILLER_30_741 VPWR VGND sg13g2_fill_1
X_1873_ VPWR VGND _0762_ net79 _0761_ _0236_ _0338_ net35 sg13g2_a221oi_1
XFILLER_6_480 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
X_2425_ net253 VGND VPWR _0371_ daisychain\[115\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2356_ net391 VGND VPWR _0302_ daisychain\[46\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_28_18 VPWR VGND sg13g2_decap_8
X_2287_ VGND VPWR _0863_ _1014_ _0500_ net88 sg13g2_a21oi_1
X_1307_ VPWR _0005_ state\[104\] VGND sg13g2_inv_1
XFILLER_44_28 VPWR VGND sg13g2_decap_8
XFILLER_12_207 VPWR VGND sg13g2_decap_8
XFILLER_21_785 VPWR VGND sg13g2_fill_2
XFILLER_20_284 VPWR VGND sg13g2_decap_8
XFILLER_4_417 VPWR VGND sg13g2_decap_8
XFILLER_0_623 VPWR VGND sg13g2_decap_8
XFILLER_47_126 VPWR VGND sg13g2_decap_8
XFILLER_28_340 VPWR VGND sg13g2_decap_8
XFILLER_18_95 VPWR VGND sg13g2_decap_8
XFILLER_29_885 VPWR VGND sg13g2_decap_4
XFILLER_43_343 VPWR VGND sg13g2_decap_8
XFILLER_44_888 VPWR VGND sg13g2_fill_1
XFILLER_12_730 VPWR VGND sg13g2_decap_8
XFILLER_11_284 VPWR VGND sg13g2_decap_8
XFILLER_8_756 VPWR VGND sg13g2_fill_1
XFILLER_8_734 VPWR VGND sg13g2_fill_2
XFILLER_8_723 VPWR VGND sg13g2_decap_8
XFILLER_7_266 VPWR VGND sg13g2_decap_8
XFILLER_4_973 VPWR VGND sg13g2_decap_4
XFILLER_3_461 VPWR VGND sg13g2_decap_8
X_2210_ _0976_ net150 state\[78\] VPWR VGND sg13g2_nand2_1
XFILLER_15_4 VPWR VGND sg13g2_decap_8
X_2141_ VGND VPWR _0644_ _0941_ _0427_ net93 sg13g2_a21oi_1
XFILLER_38_126 VPWR VGND sg13g2_decap_8
XFILLER_19_340 VPWR VGND sg13g2_decap_8
X_2072_ _0907_ net117 state\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_34_354 VPWR VGND sg13g2_decap_8
X_1925_ VPWR VGND _0801_ net85 _0800_ _0250_ _0351_ net43 sg13g2_a221oi_1
X_1856_ VGND VPWR net151 daisychain\[77\] _0750_ net60 sg13g2_a21oi_1
X_1787_ net190 _0213_ _0697_ _0698_ VPWR VGND sg13g2_a21o_1
XFILLER_39_28 VPWR VGND sg13g2_decap_8
X_2408_ net287 VGND VPWR _0354_ daisychain\[98\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_2339_ net425 VGND VPWR _0285_ daisychain\[29\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_29_137 VPWR VGND sg13g2_decap_8
XFILLER_26_822 VPWR VGND sg13g2_decap_8
XFILLER_25_354 VPWR VGND sg13g2_decap_8
XFILLER_40_357 VPWR VGND sg13g2_decap_8
XFILLER_4_214 VPWR VGND sg13g2_decap_8
XFILLER_20_74 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_49_914 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_48_413 VPWR VGND sg13g2_decap_8
XFILLER_16_354 VPWR VGND sg13g2_decap_8
XFILLER_43_140 VPWR VGND sg13g2_decap_8
XFILLER_31_368 VPWR VGND sg13g2_decap_8
XFILLER_12_582 VPWR VGND sg13g2_decap_8
XFILLER_12_593 VPWR VGND sg13g2_fill_1
X_1710_ net218 VPWR _0640_ VGND state\[42\] net184 sg13g2_o21ai_1
XANTENNA_3 VPWR VGND _0144_ sg13g2_antennanp
X_1641_ VPWR VGND _0588_ net103 _0587_ _0172_ _0280_ net58 sg13g2_a221oi_1
XFILLER_8_586 VPWR VGND sg13g2_decap_8
XFILLER_6_32 VPWR VGND sg13g2_decap_8
X_1572_ VGND VPWR net114 daisychain\[6\] _0537_ net25 sg13g2_a21oi_1
XFILLER_6_1003 VPWR VGND sg13g2_fill_1
XFILLER_3_291 VPWR VGND sg13g2_decap_8
X_2124_ _0933_ net138 state\[35\] VPWR VGND sg13g2_nand2_1
XFILLER_39_479 VPWR VGND sg13g2_decap_8
X_2055_ VGND VPWR _0514_ _0898_ _0384_ net79 sg13g2_a21oi_1
XFILLER_47_490 VPWR VGND sg13g2_decap_8
XFILLER_34_151 VPWR VGND sg13g2_decap_8
XFILLER_10_508 VPWR VGND sg13g2_decap_8
XFILLER_22_368 VPWR VGND sg13g2_decap_8
X_1908_ VGND VPWR net151 daisychain\[90\] _0789_ net60 sg13g2_a21oi_1
X_1839_ net199 _0227_ _0736_ _0737_ VPWR VGND sg13g2_a21o_1
XFILLER_1_217 VPWR VGND sg13g2_decap_8
XFILLER_45_427 VPWR VGND sg13g2_decap_8
XFILLER_25_151 VPWR VGND sg13g2_decap_8
X_2431__242 VPWR VGND net241 sg13g2_tiehi
XFILLER_13_368 VPWR VGND sg13g2_decap_8
XFILLER_15_74 VPWR VGND sg13g2_decap_8
XFILLER_40_154 VPWR VGND sg13g2_decap_8
XFILLER_5_501 VPWR VGND sg13g2_decap_8
XFILLER_5_534 VPWR VGND sg13g2_decap_8
XFILLER_31_95 VPWR VGND sg13g2_decap_8
XFILLER_49_700 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_45_983 VPWR VGND sg13g2_fill_1
XFILLER_16_151 VPWR VGND sg13g2_decap_8
XFILLER_44_471 VPWR VGND sg13g2_decap_8
XFILLER_31_165 VPWR VGND sg13g2_decap_8
XFILLER_8_361 VPWR VGND sg13g2_decap_8
X_1624_ VGND VPWR net118 daisychain\[19\] _0576_ net29 sg13g2_a21oi_1
X_2408__288 VPWR VGND net287 sg13g2_tiehi
X_1555_ net161 _0189_ _0523_ _0524_ VPWR VGND sg13g2_a21o_1
X_1486_ VPWR _0204_ daisychain\[53\] VGND sg13g2_inv_1
XFILLER_39_210 VPWR VGND sg13g2_decap_8
X_2107_ VGND VPWR _0593_ _0924_ _0410_ net76 sg13g2_a21oi_1
Xclkbuf_leaf_19_clk clknet_2_0__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_39_287 VPWR VGND sg13g2_decap_8
XFILLER_27_427 VPWR VGND sg13g2_decap_8
X_2038_ net210 VPWR _0886_ VGND state\[124\] net159 sg13g2_o21ai_1
XFILLER_23_655 VPWR VGND sg13g2_fill_1
XFILLER_10_305 VPWR VGND sg13g2_decap_8
XFILLER_22_165 VPWR VGND sg13g2_decap_8
XFILLER_2_515 VPWR VGND sg13g2_decap_8
XFILLER_18_427 VPWR VGND sg13g2_decap_8
XFILLER_18_438 VPWR VGND sg13g2_fill_2
XFILLER_45_224 VPWR VGND sg13g2_decap_8
XFILLER_14_611 VPWR VGND sg13g2_decap_8
XFILLER_42_975 VPWR VGND sg13g2_decap_8
XFILLER_26_95 VPWR VGND sg13g2_decap_8
XFILLER_13_165 VPWR VGND sg13g2_decap_8
XFILLER_14_677 VPWR VGND sg13g2_fill_2
XFILLER_14_699 VPWR VGND sg13g2_decap_4
XFILLER_42_986 VPWR VGND sg13g2_fill_1
XFILLER_9_158 VPWR VGND sg13g2_decap_8
XFILLER_6_843 VPWR VGND sg13g2_fill_1
XFILLER_5_375 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
X_2520__343 VPWR VGND net342 sg13g2_tiehi
X_1340_ VPWR _0096_ state\[71\] VGND sg13g2_inv_1
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_3_88 VPWR VGND sg13g2_decap_8
XFILLER_1_581 VPWR VGND sg13g2_decap_8
XFILLER_49_596 VPWR VGND sg13g2_decap_8
XFILLER_36_224 VPWR VGND sg13g2_decap_8
XFILLER_32_463 VPWR VGND sg13g2_decap_8
XFILLER_32_496 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_8_clk clknet_2_3__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_1607_ net177 _0163_ _0562_ _0563_ VPWR VGND sg13g2_a21o_1
Xfanout104 net111 net104 VPWR VGND sg13g2_buf_1
Xfanout137 net158 net137 VPWR VGND sg13g2_buf_1
Xfanout126 net127 net126 VPWR VGND sg13g2_buf_1
Xfanout115 net137 net115 VPWR VGND sg13g2_buf_1
XdigitalenL.g\[3\].u.inv2 VPWR digitalenL.g\[3\].u.OUTP digitalenL.g\[3\].u.OUTN VGND
+ sg13g2_inv_1
X_1538_ VPWR _0167_ daisychain\[1\] VGND sg13g2_inv_1
Xfanout159 net161 net159 VPWR VGND sg13g2_buf_1
Xfanout148 net152 net148 VPWR VGND sg13g2_buf_1
X_1469_ VPWR _0223_ daisychain\[70\] VGND sg13g2_inv_1
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_28_703 VPWR VGND sg13g2_fill_1
XFILLER_27_224 VPWR VGND sg13g2_decap_8
XFILLER_28_769 VPWR VGND sg13g2_decap_4
X_2532__247 VPWR VGND net246 sg13g2_tiehi
XFILLER_42_238 VPWR VGND sg13g2_decap_8
XFILLER_10_102 VPWR VGND sg13g2_decap_8
XFILLER_11_647 VPWR VGND sg13g2_decap_8
XFILLER_11_658 VPWR VGND sg13g2_fill_1
XFILLER_10_179 VPWR VGND sg13g2_decap_8
XFILLER_12_53 VPWR VGND sg13g2_decap_8
XFILLER_2_312 VPWR VGND sg13g2_decap_8
XFILLER_2_389 VPWR VGND sg13g2_decap_8
XFILLER_46_533 VPWR VGND sg13g2_decap_8
XFILLER_19_747 VPWR VGND sg13g2_fill_1
XFILLER_18_235 VPWR VGND sg13g2_decap_8
XFILLER_46_566 VPWR VGND sg13g2_decap_4
XFILLER_34_706 VPWR VGND sg13g2_fill_2
XFILLER_33_249 VPWR VGND sg13g2_decap_8
XFILLER_14_452 VPWR VGND sg13g2_decap_4
XFILLER_30_945 VPWR VGND sg13g2_decap_8
X_2510_ net422 VGND VPWR _0456_ state\[72\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_6_640 VPWR VGND sg13g2_decap_4
X_2441_ net472 VGND VPWR _0387_ state\[3\] clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_5_172 VPWR VGND sg13g2_decap_8
X_2372_ net359 VGND VPWR _0318_ daisychain\[62\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_1323_ VPWR _0114_ state\[88\] VGND sg13g2_inv_1
XFILLER_49_382 VPWR VGND sg13g2_decap_8
XFILLER_25_728 VPWR VGND sg13g2_fill_1
XFILLER_24_249 VPWR VGND sg13g2_decap_8
XFILLER_3_109 VPWR VGND sg13g2_decap_8
XFILLER_0_816 VPWR VGND sg13g2_fill_1
XFILLER_47_308 VPWR VGND sg13g2_decap_8
XFILLER_16_717 VPWR VGND sg13g2_decap_8
XFILLER_16_728 VPWR VGND sg13g2_fill_2
XFILLER_15_249 VPWR VGND sg13g2_decap_8
XFILLER_11_466 VPWR VGND sg13g2_decap_8
XFILLER_8_927 VPWR VGND sg13g2_fill_1
XFILLER_7_448 VPWR VGND sg13g2_decap_8
XFILLER_23_74 VPWR VGND sg13g2_decap_8
XFILLER_3_643 VPWR VGND sg13g2_decap_8
XFILLER_2_186 VPWR VGND sg13g2_decap_8
XFILLER_38_308 VPWR VGND sg13g2_decap_8
XFILLER_19_522 VPWR VGND sg13g2_fill_2
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_46_385 VPWR VGND sg13g2_decap_8
XFILLER_34_569 VPWR VGND sg13g2_fill_1
X_1941_ VPWR VGND _0813_ net89 _0812_ _0254_ _0355_ net46 sg13g2_a221oi_1
XFILLER_9_32 VPWR VGND sg13g2_decap_8
X_1872_ VGND VPWR net123 daisychain\[81\] _0762_ net35 sg13g2_a21oi_1
X_2424_ net255 VGND VPWR _0370_ daisychain\[114\] clknet_leaf_5_clk sg13g2_dfrbpq_1
X_2355_ net393 VGND VPWR _0301_ daisychain\[45\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
X_1306_ VPWR _0006_ state\[105\] VGND sg13g2_inv_1
XFILLER_29_319 VPWR VGND sg13g2_decap_8
X_2286_ _1014_ net132 state\[116\] VPWR VGND sg13g2_nand2_1
XFILLER_37_385 VPWR VGND sg13g2_decap_8
XFILLER_33_580 VPWR VGND sg13g2_decap_8
XFILLER_21_731 VPWR VGND sg13g2_decap_8
XFILLER_20_263 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_decap_8
XFILLER_0_679 VPWR VGND sg13g2_decap_8
XFILLER_48_628 VPWR VGND sg13g2_fill_1
XFILLER_47_105 VPWR VGND sg13g2_decap_8
XFILLER_18_74 VPWR VGND sg13g2_decap_8
XFILLER_43_322 VPWR VGND sg13g2_decap_8
XFILLER_28_396 VPWR VGND sg13g2_decap_8
XFILLER_43_399 VPWR VGND sg13g2_decap_8
XFILLER_34_95 VPWR VGND sg13g2_decap_8
XFILLER_11_263 VPWR VGND sg13g2_decap_8
XFILLER_8_779 VPWR VGND sg13g2_fill_1
XFILLER_7_245 VPWR VGND sg13g2_decap_8
XFILLER_4_963 VPWR VGND sg13g2_fill_1
XFILLER_4_952 VPWR VGND sg13g2_decap_8
XFILLER_4_996 VPWR VGND sg13g2_fill_1
XFILLER_3_440 VPWR VGND sg13g2_decap_8
X_2140_ _0941_ net138 state\[43\] VPWR VGND sg13g2_nand2_1
XFILLER_39_628 VPWR VGND sg13g2_fill_2
XFILLER_38_105 VPWR VGND sg13g2_decap_8
X_2071_ VGND VPWR _0539_ _0906_ _0392_ net78 sg13g2_a21oi_1
XFILLER_47_683 VPWR VGND sg13g2_decap_8
XFILLER_46_182 VPWR VGND sg13g2_decap_8
XFILLER_34_333 VPWR VGND sg13g2_decap_8
XFILLER_19_396 VPWR VGND sg13g2_decap_8
XFILLER_22_517 VPWR VGND sg13g2_fill_2
X_1924_ VGND VPWR net129 daisychain\[94\] _0801_ net42 sg13g2_a21oi_1
X_1855_ net196 _0231_ _0748_ _0749_ VPWR VGND sg13g2_a21o_1
X_1786_ net222 VPWR _0697_ VGND state\[61\] net190 sg13g2_o21ai_1
X_2407_ net289 VGND VPWR _0353_ daisychain\[97\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_2338_ net427 VGND VPWR _0284_ daisychain\[28\] clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_29_116 VPWR VGND sg13g2_decap_8
X_2269_ VGND VPWR _0836_ _1005_ _0491_ net88 sg13g2_a21oi_1
XFILLER_44_119 VPWR VGND sg13g2_decap_8
X_2418__268 VPWR VGND net267 sg13g2_tiehi
XFILLER_37_182 VPWR VGND sg13g2_decap_8
XFILLER_25_333 VPWR VGND sg13g2_decap_8
XFILLER_13_528 VPWR VGND sg13g2_fill_2
XFILLER_40_336 VPWR VGND sg13g2_decap_8
XFILLER_5_705 VPWR VGND sg13g2_fill_1
XFILLER_20_53 VPWR VGND sg13g2_decap_8
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_48_469 VPWR VGND sg13g2_decap_8
XFILLER_29_95 VPWR VGND sg13g2_decap_8
XFILLER_35_119 VPWR VGND sg13g2_decap_8
XFILLER_16_333 VPWR VGND sg13g2_decap_8
XFILLER_44_620 VPWR VGND sg13g2_fill_2
XFILLER_28_193 VPWR VGND sg13g2_decap_8
XFILLER_44_653 VPWR VGND sg13g2_fill_1
XFILLER_44_697 VPWR VGND sg13g2_decap_8
XFILLER_43_196 VPWR VGND sg13g2_decap_8
XFILLER_31_347 VPWR VGND sg13g2_decap_8
X_1640_ VGND VPWR net149 daisychain\[23\] _0588_ net58 sg13g2_a21oi_1
XFILLER_8_598 VPWR VGND sg13g2_decap_8
XFILLER_8_565 VPWR VGND sg13g2_decap_8
XFILLER_6_11 VPWR VGND sg13g2_decap_8
XANTENNA_4 VPWR VGND _0150_ sg13g2_antennanp
X_1571_ net160 _0233_ _0535_ _0536_ VPWR VGND sg13g2_a21o_1
XFILLER_6_88 VPWR VGND sg13g2_decap_8
XFILLER_4_782 VPWR VGND sg13g2_decap_8
XFILLER_3_270 VPWR VGND sg13g2_decap_8
X_2123_ VGND VPWR _0617_ _0932_ _0418_ net74 sg13g2_a21oi_1
X_2054_ _0898_ net123 state\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_19_193 VPWR VGND sg13g2_decap_8
XFILLER_34_130 VPWR VGND sg13g2_decap_8
XFILLER_22_347 VPWR VGND sg13g2_decap_8
X_1907_ net198 _0246_ _0787_ _0788_ VPWR VGND sg13g2_a21o_1
X_1838_ net225 VPWR _0736_ VGND state\[74\] net199 sg13g2_o21ai_1
X_1769_ VPWR VGND _0684_ net99 _0683_ _0207_ _0312_ net53 sg13g2_a221oi_1
XFILLER_45_406 VPWR VGND sg13g2_decap_8
XFILLER_17_119 VPWR VGND sg13g2_decap_8
XFILLER_38_480 VPWR VGND sg13g2_fill_1
XFILLER_25_130 VPWR VGND sg13g2_decap_8
XFILLER_13_347 VPWR VGND sg13g2_decap_8
XFILLER_15_53 VPWR VGND sg13g2_decap_8
XFILLER_40_133 VPWR VGND sg13g2_decap_8
XFILLER_5_513 VPWR VGND sg13g2_decap_8
XFILLER_31_74 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_49_745 VPWR VGND sg13g2_decap_8
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_36_406 VPWR VGND sg13g2_decap_8
XFILLER_17_620 VPWR VGND sg13g2_decap_4
XFILLER_29_480 VPWR VGND sg13g2_decap_8
XFILLER_16_130 VPWR VGND sg13g2_decap_8
XFILLER_45_962 VPWR VGND sg13g2_decap_8
XFILLER_45_995 VPWR VGND sg13g2_decap_8
XFILLER_32_678 VPWR VGND sg13g2_fill_2
XFILLER_31_144 VPWR VGND sg13g2_decap_8
XFILLER_8_340 VPWR VGND sg13g2_decap_8
X_2310__483 VPWR VGND net482 sg13g2_tiehi
X_1623_ net165 _0168_ _0574_ _0575_ VPWR VGND sg13g2_a21o_1
X_1554_ net205 VPWR _0523_ VGND state\[3\] net161 sg13g2_o21ai_1
X_1485_ VPWR _0205_ daisychain\[54\] VGND sg13g2_inv_1
.ends

