* Extracted by KLayout with SG13G2 LVS runset on : 27/08/2025 20:52

.SUBCKT PCSOURCE2U
M$1 \$2 \$5 \$10 \$2 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p PS=3.58u
+ PD=1.75u
M$2 \$10 \$1 \$6 \$2 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p PS=1.75u
+ PD=3.26u
.ENDS PCSOURCE2U
