VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DAC2U128OUT4IN
  CLASS BLOCK ;
  FOREIGN DAC2U128OUT4IN ;
  ORIGIN 0.310 0.200 ;
  SIZE 134.420 BY 26.590 ;
  PIN VbiasP[1]
    ANTENNAGATEAREA 478.500000 ;
    ANTENNADIFFAREA 5.010000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.900 14.950 1.080 19.950 ;
        RECT 2.530 14.950 3.080 19.950 ;
        RECT 4.530 14.950 5.080 19.950 ;
        RECT 6.530 14.950 7.080 19.950 ;
        RECT 8.530 14.950 9.080 19.950 ;
        RECT 10.530 14.950 11.080 19.950 ;
        RECT 12.530 14.950 13.080 19.950 ;
        RECT 14.530 14.950 15.080 19.950 ;
        RECT 16.530 14.950 17.080 19.950 ;
        RECT 18.530 14.950 19.080 19.950 ;
        RECT 20.530 14.950 21.080 19.950 ;
        RECT 22.530 14.950 23.080 19.950 ;
        RECT 24.530 14.950 25.080 19.950 ;
        RECT 26.530 14.950 27.080 19.950 ;
        RECT 28.530 14.950 29.080 19.950 ;
        RECT 30.530 14.950 31.080 19.950 ;
        RECT 32.530 14.950 33.080 19.950 ;
        RECT 34.530 14.950 35.080 19.950 ;
        RECT 36.530 14.950 37.080 19.950 ;
        RECT 38.530 14.950 39.080 19.950 ;
        RECT 40.530 14.950 41.080 19.950 ;
        RECT 42.530 14.950 43.080 19.950 ;
        RECT 44.530 14.950 45.080 19.950 ;
        RECT 46.530 14.950 47.080 19.950 ;
        RECT 48.530 14.950 49.080 19.950 ;
        RECT 50.530 14.950 51.080 19.950 ;
        RECT 52.530 14.950 53.080 19.950 ;
        RECT 54.530 14.950 55.080 19.950 ;
        RECT 56.530 14.950 57.080 19.950 ;
        RECT 58.530 14.950 59.080 19.950 ;
        RECT 60.530 14.950 61.080 19.950 ;
        RECT 62.530 14.950 63.080 19.950 ;
        RECT 64.530 14.950 65.080 19.950 ;
        RECT 66.530 14.950 67.080 19.950 ;
        RECT 68.530 14.950 69.080 19.950 ;
        RECT 70.530 14.950 71.080 19.950 ;
        RECT 72.530 14.950 73.080 19.950 ;
        RECT 74.530 14.950 75.080 19.950 ;
        RECT 76.530 14.950 77.080 19.950 ;
        RECT 78.530 14.950 79.080 19.950 ;
        RECT 80.530 14.950 81.080 19.950 ;
        RECT 82.530 14.950 83.080 19.950 ;
        RECT 84.530 14.950 85.080 19.950 ;
        RECT 86.530 14.950 87.080 19.950 ;
        RECT 88.530 14.950 89.080 19.950 ;
        RECT 90.530 14.950 91.080 19.950 ;
        RECT 92.530 14.950 93.080 19.950 ;
        RECT 94.530 14.950 95.080 19.950 ;
        RECT 96.530 14.950 97.080 19.950 ;
        RECT 98.530 14.950 99.080 19.950 ;
        RECT 100.530 14.950 101.080 19.950 ;
        RECT 102.530 14.950 103.080 19.950 ;
        RECT 104.530 14.950 105.080 19.950 ;
        RECT 106.530 14.950 107.080 19.950 ;
        RECT 108.530 14.950 109.080 19.950 ;
        RECT 110.530 14.950 111.080 19.950 ;
        RECT 112.530 14.950 113.080 19.950 ;
        RECT 114.530 14.950 115.080 19.950 ;
        RECT 116.530 14.950 117.080 19.950 ;
        RECT 118.530 14.950 119.080 19.950 ;
        RECT 120.530 14.950 121.080 19.950 ;
        RECT 122.530 14.950 123.080 19.950 ;
        RECT 124.530 14.950 125.080 19.950 ;
        RECT 126.530 14.950 127.080 19.950 ;
        RECT 128.530 14.950 129.080 19.950 ;
        RECT 130.530 14.950 131.080 19.950 ;
        RECT 132.530 14.950 132.900 19.950 ;
      LAYER Metal1 ;
        RECT 0.900 19.520 132.900 19.880 ;
        RECT 0.600 14.950 133.200 19.520 ;
        RECT 0.600 13.670 0.760 14.950 ;
        RECT 1.085 13.665 2.275 14.950 ;
        RECT 131.085 13.665 132.275 14.950 ;
        RECT 133.040 13.670 133.200 14.950 ;
    END
  END VbiasP[1]
  PIN Iout
    ANTENNADIFFAREA 66.047997 ;
    PORT
      LAYER Metal1 ;
        RECT 3.085 13.445 130.275 13.875 ;
        RECT 0.000 12.745 133.800 13.445 ;
        RECT 3.525 12.315 130.715 12.745 ;
    END
  END Iout
  PIN VbiasP[0]
    ANTENNAGATEAREA 478.500000 ;
    ANTENNADIFFAREA 5.010000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.900 6.240 1.270 11.240 ;
        RECT 2.720 6.240 3.270 11.240 ;
        RECT 4.720 6.240 5.270 11.240 ;
        RECT 6.720 6.240 7.270 11.240 ;
        RECT 8.720 6.240 9.270 11.240 ;
        RECT 10.720 6.240 11.270 11.240 ;
        RECT 12.720 6.240 13.270 11.240 ;
        RECT 14.720 6.240 15.270 11.240 ;
        RECT 16.720 6.240 17.270 11.240 ;
        RECT 18.720 6.240 19.270 11.240 ;
        RECT 20.720 6.240 21.270 11.240 ;
        RECT 22.720 6.240 23.270 11.240 ;
        RECT 24.720 6.240 25.270 11.240 ;
        RECT 26.720 6.240 27.270 11.240 ;
        RECT 28.720 6.240 29.270 11.240 ;
        RECT 30.720 6.240 31.270 11.240 ;
        RECT 32.720 6.240 33.270 11.240 ;
        RECT 34.720 6.240 35.270 11.240 ;
        RECT 36.720 6.240 37.270 11.240 ;
        RECT 38.720 6.240 39.270 11.240 ;
        RECT 40.720 6.240 41.270 11.240 ;
        RECT 42.720 6.240 43.270 11.240 ;
        RECT 44.720 6.240 45.270 11.240 ;
        RECT 46.720 6.240 47.270 11.240 ;
        RECT 48.720 6.240 49.270 11.240 ;
        RECT 50.720 6.240 51.270 11.240 ;
        RECT 52.720 6.240 53.270 11.240 ;
        RECT 54.720 6.240 55.270 11.240 ;
        RECT 56.720 6.240 57.270 11.240 ;
        RECT 58.720 6.240 59.270 11.240 ;
        RECT 60.720 6.240 61.270 11.240 ;
        RECT 62.720 6.240 63.270 11.240 ;
        RECT 64.720 6.240 65.270 11.240 ;
        RECT 66.720 6.240 67.270 11.240 ;
        RECT 68.720 6.240 69.270 11.240 ;
        RECT 70.720 6.240 71.270 11.240 ;
        RECT 72.720 6.240 73.270 11.240 ;
        RECT 74.720 6.240 75.270 11.240 ;
        RECT 76.720 6.240 77.270 11.240 ;
        RECT 78.720 6.240 79.270 11.240 ;
        RECT 80.720 6.240 81.270 11.240 ;
        RECT 82.720 6.240 83.270 11.240 ;
        RECT 84.720 6.240 85.270 11.240 ;
        RECT 86.720 6.240 87.270 11.240 ;
        RECT 88.720 6.240 89.270 11.240 ;
        RECT 90.720 6.240 91.270 11.240 ;
        RECT 92.720 6.240 93.270 11.240 ;
        RECT 94.720 6.240 95.270 11.240 ;
        RECT 96.720 6.240 97.270 11.240 ;
        RECT 98.720 6.240 99.270 11.240 ;
        RECT 100.720 6.240 101.270 11.240 ;
        RECT 102.720 6.240 103.270 11.240 ;
        RECT 104.720 6.240 105.270 11.240 ;
        RECT 106.720 6.240 107.270 11.240 ;
        RECT 108.720 6.240 109.270 11.240 ;
        RECT 110.720 6.240 111.270 11.240 ;
        RECT 112.720 6.240 113.270 11.240 ;
        RECT 114.720 6.240 115.270 11.240 ;
        RECT 116.720 6.240 117.270 11.240 ;
        RECT 118.720 6.240 119.270 11.240 ;
        RECT 120.720 6.240 121.270 11.240 ;
        RECT 122.720 6.240 123.270 11.240 ;
        RECT 124.720 6.240 125.270 11.240 ;
        RECT 126.720 6.240 127.270 11.240 ;
        RECT 128.720 6.240 129.270 11.240 ;
        RECT 130.720 6.240 131.270 11.240 ;
        RECT 132.720 6.240 132.900 11.240 ;
      LAYER Metal1 ;
        RECT 0.600 11.240 0.760 12.520 ;
        RECT 1.525 11.240 2.715 12.525 ;
        RECT 131.525 11.240 132.715 12.525 ;
        RECT 133.040 11.240 133.200 12.520 ;
        RECT 0.600 6.670 133.200 11.240 ;
        RECT 0.900 6.310 132.900 6.670 ;
    END
  END VbiasP[0]
  PIN ON[64]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 130.090 23.380 130.390 23.680 ;
        RECT 130.090 23.310 130.220 23.380 ;
        RECT 130.090 22.830 130.220 23.010 ;
      LAYER Metal1 ;
        RECT 130.030 23.470 130.320 23.760 ;
        RECT 130.160 23.400 130.320 23.470 ;
      LAYER Metal2 ;
        RECT 130.030 23.470 130.320 26.190 ;
    END
  END ON[64]
  PIN ONB[64]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 129.410 23.380 129.710 23.680 ;
        RECT 129.580 23.310 129.710 23.380 ;
        RECT 129.580 22.830 129.710 23.010 ;
      LAYER Metal1 ;
        RECT 129.480 23.470 129.770 23.760 ;
        RECT 129.480 23.400 129.640 23.470 ;
      LAYER Metal2 ;
        RECT 129.480 23.470 129.770 26.190 ;
    END
  END ONB[64]
  PIN ON[65]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 128.090 23.380 128.390 23.680 ;
        RECT 128.090 23.310 128.220 23.380 ;
        RECT 128.090 22.830 128.220 23.010 ;
      LAYER Metal1 ;
        RECT 128.030 23.470 128.320 23.760 ;
        RECT 128.160 23.400 128.320 23.470 ;
      LAYER Metal2 ;
        RECT 128.030 23.470 128.320 26.190 ;
    END
  END ON[65]
  PIN ONB[65]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 127.410 23.380 127.710 23.680 ;
        RECT 127.580 23.310 127.710 23.380 ;
        RECT 127.580 22.830 127.710 23.010 ;
      LAYER Metal1 ;
        RECT 127.480 23.470 127.770 23.760 ;
        RECT 127.480 23.400 127.640 23.470 ;
      LAYER Metal2 ;
        RECT 127.480 23.470 127.770 26.190 ;
    END
  END ONB[65]
  PIN ON[66]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 126.090 23.380 126.390 23.680 ;
        RECT 126.090 23.310 126.220 23.380 ;
        RECT 126.090 22.830 126.220 23.010 ;
      LAYER Metal1 ;
        RECT 126.030 23.470 126.320 23.760 ;
        RECT 126.160 23.400 126.320 23.470 ;
      LAYER Metal2 ;
        RECT 126.030 23.470 126.320 26.190 ;
    END
  END ON[66]
  PIN ONB[66]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 125.410 23.380 125.710 23.680 ;
        RECT 125.580 23.310 125.710 23.380 ;
        RECT 125.580 22.830 125.710 23.010 ;
      LAYER Metal1 ;
        RECT 125.480 23.470 125.770 23.760 ;
        RECT 125.480 23.400 125.640 23.470 ;
      LAYER Metal2 ;
        RECT 125.480 23.470 125.770 26.190 ;
    END
  END ONB[66]
  PIN ON[67]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 124.090 23.380 124.390 23.680 ;
        RECT 124.090 23.310 124.220 23.380 ;
        RECT 124.090 22.830 124.220 23.010 ;
      LAYER Metal1 ;
        RECT 124.030 23.470 124.320 23.760 ;
        RECT 124.160 23.400 124.320 23.470 ;
      LAYER Metal2 ;
        RECT 124.030 23.470 124.320 26.190 ;
    END
  END ON[67]
  PIN ONB[67]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 123.410 23.380 123.710 23.680 ;
        RECT 123.580 23.310 123.710 23.380 ;
        RECT 123.580 22.830 123.710 23.010 ;
      LAYER Metal1 ;
        RECT 123.480 23.470 123.770 23.760 ;
        RECT 123.480 23.400 123.640 23.470 ;
      LAYER Metal2 ;
        RECT 123.480 23.470 123.770 26.190 ;
    END
  END ONB[67]
  PIN ON[68]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 122.090 23.380 122.390 23.680 ;
        RECT 122.090 23.310 122.220 23.380 ;
        RECT 122.090 22.830 122.220 23.010 ;
      LAYER Metal1 ;
        RECT 122.030 23.470 122.320 23.760 ;
        RECT 122.160 23.400 122.320 23.470 ;
      LAYER Metal2 ;
        RECT 122.030 23.470 122.320 26.190 ;
    END
  END ON[68]
  PIN ONB[68]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 121.410 23.380 121.710 23.680 ;
        RECT 121.580 23.310 121.710 23.380 ;
        RECT 121.580 22.830 121.710 23.010 ;
      LAYER Metal1 ;
        RECT 121.480 23.470 121.770 23.760 ;
        RECT 121.480 23.400 121.640 23.470 ;
      LAYER Metal2 ;
        RECT 121.480 23.470 121.770 26.190 ;
    END
  END ONB[68]
  PIN ON[69]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 120.090 23.380 120.390 23.680 ;
        RECT 120.090 23.310 120.220 23.380 ;
        RECT 120.090 22.830 120.220 23.010 ;
      LAYER Metal1 ;
        RECT 120.030 23.470 120.320 23.760 ;
        RECT 120.160 23.400 120.320 23.470 ;
      LAYER Metal2 ;
        RECT 120.030 23.470 120.320 26.190 ;
    END
  END ON[69]
  PIN ONB[69]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 119.410 23.380 119.710 23.680 ;
        RECT 119.580 23.310 119.710 23.380 ;
        RECT 119.580 22.830 119.710 23.010 ;
      LAYER Metal1 ;
        RECT 119.480 23.470 119.770 23.760 ;
        RECT 119.480 23.400 119.640 23.470 ;
      LAYER Metal2 ;
        RECT 119.480 23.470 119.770 26.190 ;
    END
  END ONB[69]
  PIN ON[70]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 118.090 23.380 118.390 23.680 ;
        RECT 118.090 23.310 118.220 23.380 ;
        RECT 118.090 22.830 118.220 23.010 ;
      LAYER Metal1 ;
        RECT 118.030 23.470 118.320 23.760 ;
        RECT 118.160 23.400 118.320 23.470 ;
      LAYER Metal2 ;
        RECT 118.030 23.470 118.320 26.190 ;
    END
  END ON[70]
  PIN ONB[70]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 117.410 23.380 117.710 23.680 ;
        RECT 117.580 23.310 117.710 23.380 ;
        RECT 117.580 22.830 117.710 23.010 ;
      LAYER Metal1 ;
        RECT 117.480 23.470 117.770 23.760 ;
        RECT 117.480 23.400 117.640 23.470 ;
      LAYER Metal2 ;
        RECT 117.480 23.470 117.770 26.190 ;
    END
  END ONB[70]
  PIN ON[71]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 116.090 23.380 116.390 23.680 ;
        RECT 116.090 23.310 116.220 23.380 ;
        RECT 116.090 22.830 116.220 23.010 ;
      LAYER Metal1 ;
        RECT 116.030 23.470 116.320 23.760 ;
        RECT 116.160 23.400 116.320 23.470 ;
      LAYER Metal2 ;
        RECT 116.030 23.470 116.320 26.190 ;
    END
  END ON[71]
  PIN ONB[71]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 115.410 23.380 115.710 23.680 ;
        RECT 115.580 23.310 115.710 23.380 ;
        RECT 115.580 22.830 115.710 23.010 ;
      LAYER Metal1 ;
        RECT 115.480 23.470 115.770 23.760 ;
        RECT 115.480 23.400 115.640 23.470 ;
      LAYER Metal2 ;
        RECT 115.480 23.470 115.770 26.190 ;
    END
  END ONB[71]
  PIN ON[72]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 114.090 23.380 114.390 23.680 ;
        RECT 114.090 23.310 114.220 23.380 ;
        RECT 114.090 22.830 114.220 23.010 ;
      LAYER Metal1 ;
        RECT 114.030 23.470 114.320 23.760 ;
        RECT 114.160 23.400 114.320 23.470 ;
      LAYER Metal2 ;
        RECT 114.030 23.470 114.320 26.190 ;
    END
  END ON[72]
  PIN ONB[72]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 113.410 23.380 113.710 23.680 ;
        RECT 113.580 23.310 113.710 23.380 ;
        RECT 113.580 22.830 113.710 23.010 ;
      LAYER Metal1 ;
        RECT 113.480 23.470 113.770 23.760 ;
        RECT 113.480 23.400 113.640 23.470 ;
      LAYER Metal2 ;
        RECT 113.480 23.470 113.770 26.190 ;
    END
  END ONB[72]
  PIN ON[73]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 112.090 23.380 112.390 23.680 ;
        RECT 112.090 23.310 112.220 23.380 ;
        RECT 112.090 22.830 112.220 23.010 ;
      LAYER Metal1 ;
        RECT 112.030 23.470 112.320 23.760 ;
        RECT 112.160 23.400 112.320 23.470 ;
      LAYER Metal2 ;
        RECT 112.030 23.470 112.320 26.190 ;
    END
  END ON[73]
  PIN ONB[73]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 111.410 23.380 111.710 23.680 ;
        RECT 111.580 23.310 111.710 23.380 ;
        RECT 111.580 22.830 111.710 23.010 ;
      LAYER Metal1 ;
        RECT 111.480 23.470 111.770 23.760 ;
        RECT 111.480 23.400 111.640 23.470 ;
      LAYER Metal2 ;
        RECT 111.480 23.470 111.770 26.190 ;
    END
  END ONB[73]
  PIN ON[74]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 110.090 23.380 110.390 23.680 ;
        RECT 110.090 23.310 110.220 23.380 ;
        RECT 110.090 22.830 110.220 23.010 ;
      LAYER Metal1 ;
        RECT 110.030 23.470 110.320 23.760 ;
        RECT 110.160 23.400 110.320 23.470 ;
      LAYER Metal2 ;
        RECT 110.030 23.470 110.320 26.190 ;
    END
  END ON[74]
  PIN ONB[74]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 109.410 23.380 109.710 23.680 ;
        RECT 109.580 23.310 109.710 23.380 ;
        RECT 109.580 22.830 109.710 23.010 ;
      LAYER Metal1 ;
        RECT 109.480 23.470 109.770 23.760 ;
        RECT 109.480 23.400 109.640 23.470 ;
      LAYER Metal2 ;
        RECT 109.480 23.470 109.770 26.190 ;
    END
  END ONB[74]
  PIN ON[75]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 108.090 23.380 108.390 23.680 ;
        RECT 108.090 23.310 108.220 23.380 ;
        RECT 108.090 22.830 108.220 23.010 ;
      LAYER Metal1 ;
        RECT 108.030 23.470 108.320 23.760 ;
        RECT 108.160 23.400 108.320 23.470 ;
      LAYER Metal2 ;
        RECT 108.030 23.470 108.320 26.190 ;
    END
  END ON[75]
  PIN ONB[75]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 107.410 23.380 107.710 23.680 ;
        RECT 107.580 23.310 107.710 23.380 ;
        RECT 107.580 22.830 107.710 23.010 ;
      LAYER Metal1 ;
        RECT 107.480 23.470 107.770 23.760 ;
        RECT 107.480 23.400 107.640 23.470 ;
      LAYER Metal2 ;
        RECT 107.480 23.470 107.770 26.190 ;
    END
  END ONB[75]
  PIN ON[76]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 106.090 23.380 106.390 23.680 ;
        RECT 106.090 23.310 106.220 23.380 ;
        RECT 106.090 22.830 106.220 23.010 ;
      LAYER Metal1 ;
        RECT 106.030 23.470 106.320 23.760 ;
        RECT 106.160 23.400 106.320 23.470 ;
      LAYER Metal2 ;
        RECT 106.030 23.470 106.320 26.190 ;
    END
  END ON[76]
  PIN ONB[76]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 105.410 23.380 105.710 23.680 ;
        RECT 105.580 23.310 105.710 23.380 ;
        RECT 105.580 22.830 105.710 23.010 ;
      LAYER Metal1 ;
        RECT 105.480 23.470 105.770 23.760 ;
        RECT 105.480 23.400 105.640 23.470 ;
      LAYER Metal2 ;
        RECT 105.480 23.470 105.770 26.190 ;
    END
  END ONB[76]
  PIN ON[77]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 104.090 23.380 104.390 23.680 ;
        RECT 104.090 23.310 104.220 23.380 ;
        RECT 104.090 22.830 104.220 23.010 ;
      LAYER Metal1 ;
        RECT 104.030 23.470 104.320 23.760 ;
        RECT 104.160 23.400 104.320 23.470 ;
      LAYER Metal2 ;
        RECT 104.030 23.470 104.320 26.190 ;
    END
  END ON[77]
  PIN ONB[77]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 103.410 23.380 103.710 23.680 ;
        RECT 103.580 23.310 103.710 23.380 ;
        RECT 103.580 22.830 103.710 23.010 ;
      LAYER Metal1 ;
        RECT 103.480 23.470 103.770 23.760 ;
        RECT 103.480 23.400 103.640 23.470 ;
      LAYER Metal2 ;
        RECT 103.480 23.470 103.770 26.190 ;
    END
  END ONB[77]
  PIN ON[78]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 102.090 23.380 102.390 23.680 ;
        RECT 102.090 23.310 102.220 23.380 ;
        RECT 102.090 22.830 102.220 23.010 ;
      LAYER Metal1 ;
        RECT 102.030 23.470 102.320 23.760 ;
        RECT 102.160 23.400 102.320 23.470 ;
      LAYER Metal2 ;
        RECT 102.030 23.470 102.320 26.190 ;
    END
  END ON[78]
  PIN ONB[78]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 101.410 23.380 101.710 23.680 ;
        RECT 101.580 23.310 101.710 23.380 ;
        RECT 101.580 22.830 101.710 23.010 ;
      LAYER Metal1 ;
        RECT 101.480 23.470 101.770 23.760 ;
        RECT 101.480 23.400 101.640 23.470 ;
      LAYER Metal2 ;
        RECT 101.480 23.470 101.770 26.190 ;
    END
  END ONB[78]
  PIN ON[79]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 100.090 23.380 100.390 23.680 ;
        RECT 100.090 23.310 100.220 23.380 ;
        RECT 100.090 22.830 100.220 23.010 ;
      LAYER Metal1 ;
        RECT 100.030 23.470 100.320 23.760 ;
        RECT 100.160 23.400 100.320 23.470 ;
      LAYER Metal2 ;
        RECT 100.030 23.470 100.320 26.190 ;
    END
  END ON[79]
  PIN ONB[79]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 99.410 23.380 99.710 23.680 ;
        RECT 99.580 23.310 99.710 23.380 ;
        RECT 99.580 22.830 99.710 23.010 ;
      LAYER Metal1 ;
        RECT 99.480 23.470 99.770 23.760 ;
        RECT 99.480 23.400 99.640 23.470 ;
      LAYER Metal2 ;
        RECT 99.480 23.470 99.770 26.190 ;
    END
  END ONB[79]
  PIN ON[80]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 98.090 23.380 98.390 23.680 ;
        RECT 98.090 23.310 98.220 23.380 ;
        RECT 98.090 22.830 98.220 23.010 ;
      LAYER Metal1 ;
        RECT 98.030 23.470 98.320 23.760 ;
        RECT 98.160 23.400 98.320 23.470 ;
      LAYER Metal2 ;
        RECT 98.030 23.470 98.320 26.190 ;
    END
  END ON[80]
  PIN ONB[80]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 97.410 23.380 97.710 23.680 ;
        RECT 97.580 23.310 97.710 23.380 ;
        RECT 97.580 22.830 97.710 23.010 ;
      LAYER Metal1 ;
        RECT 97.480 23.470 97.770 23.760 ;
        RECT 97.480 23.400 97.640 23.470 ;
      LAYER Metal2 ;
        RECT 97.480 23.470 97.770 26.190 ;
    END
  END ONB[80]
  PIN ON[81]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 96.090 23.380 96.390 23.680 ;
        RECT 96.090 23.310 96.220 23.380 ;
        RECT 96.090 22.830 96.220 23.010 ;
      LAYER Metal1 ;
        RECT 96.030 23.470 96.320 23.760 ;
        RECT 96.160 23.400 96.320 23.470 ;
      LAYER Metal2 ;
        RECT 96.030 23.470 96.320 26.190 ;
    END
  END ON[81]
  PIN ONB[81]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 95.410 23.380 95.710 23.680 ;
        RECT 95.580 23.310 95.710 23.380 ;
        RECT 95.580 22.830 95.710 23.010 ;
      LAYER Metal1 ;
        RECT 95.480 23.470 95.770 23.760 ;
        RECT 95.480 23.400 95.640 23.470 ;
      LAYER Metal2 ;
        RECT 95.480 23.470 95.770 26.190 ;
    END
  END ONB[81]
  PIN ON[82]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 94.090 23.380 94.390 23.680 ;
        RECT 94.090 23.310 94.220 23.380 ;
        RECT 94.090 22.830 94.220 23.010 ;
      LAYER Metal1 ;
        RECT 94.030 23.470 94.320 23.760 ;
        RECT 94.160 23.400 94.320 23.470 ;
      LAYER Metal2 ;
        RECT 94.030 23.470 94.320 26.190 ;
    END
  END ON[82]
  PIN ONB[82]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 93.410 23.380 93.710 23.680 ;
        RECT 93.580 23.310 93.710 23.380 ;
        RECT 93.580 22.830 93.710 23.010 ;
      LAYER Metal1 ;
        RECT 93.480 23.470 93.770 23.760 ;
        RECT 93.480 23.400 93.640 23.470 ;
      LAYER Metal2 ;
        RECT 93.480 23.470 93.770 26.190 ;
    END
  END ONB[82]
  PIN ON[83]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 92.090 23.380 92.390 23.680 ;
        RECT 92.090 23.310 92.220 23.380 ;
        RECT 92.090 22.830 92.220 23.010 ;
      LAYER Metal1 ;
        RECT 92.030 23.470 92.320 23.760 ;
        RECT 92.160 23.400 92.320 23.470 ;
      LAYER Metal2 ;
        RECT 92.030 23.470 92.320 26.190 ;
    END
  END ON[83]
  PIN ONB[83]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 91.410 23.380 91.710 23.680 ;
        RECT 91.580 23.310 91.710 23.380 ;
        RECT 91.580 22.830 91.710 23.010 ;
      LAYER Metal1 ;
        RECT 91.480 23.470 91.770 23.760 ;
        RECT 91.480 23.400 91.640 23.470 ;
      LAYER Metal2 ;
        RECT 91.480 23.470 91.770 26.190 ;
    END
  END ONB[83]
  PIN ON[84]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 90.090 23.380 90.390 23.680 ;
        RECT 90.090 23.310 90.220 23.380 ;
        RECT 90.090 22.830 90.220 23.010 ;
      LAYER Metal1 ;
        RECT 90.030 23.470 90.320 23.760 ;
        RECT 90.160 23.400 90.320 23.470 ;
      LAYER Metal2 ;
        RECT 90.030 23.470 90.320 26.190 ;
    END
  END ON[84]
  PIN ONB[84]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 89.410 23.380 89.710 23.680 ;
        RECT 89.580 23.310 89.710 23.380 ;
        RECT 89.580 22.830 89.710 23.010 ;
      LAYER Metal1 ;
        RECT 89.480 23.470 89.770 23.760 ;
        RECT 89.480 23.400 89.640 23.470 ;
      LAYER Metal2 ;
        RECT 89.480 23.470 89.770 26.190 ;
    END
  END ONB[84]
  PIN ON[85]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 88.090 23.380 88.390 23.680 ;
        RECT 88.090 23.310 88.220 23.380 ;
        RECT 88.090 22.830 88.220 23.010 ;
      LAYER Metal1 ;
        RECT 88.030 23.470 88.320 23.760 ;
        RECT 88.160 23.400 88.320 23.470 ;
      LAYER Metal2 ;
        RECT 88.030 23.470 88.320 26.190 ;
    END
  END ON[85]
  PIN ONB[85]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 87.410 23.380 87.710 23.680 ;
        RECT 87.580 23.310 87.710 23.380 ;
        RECT 87.580 22.830 87.710 23.010 ;
      LAYER Metal1 ;
        RECT 87.480 23.470 87.770 23.760 ;
        RECT 87.480 23.400 87.640 23.470 ;
      LAYER Metal2 ;
        RECT 87.480 23.470 87.770 26.190 ;
    END
  END ONB[85]
  PIN ON[86]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 86.090 23.380 86.390 23.680 ;
        RECT 86.090 23.310 86.220 23.380 ;
        RECT 86.090 22.830 86.220 23.010 ;
      LAYER Metal1 ;
        RECT 86.030 23.470 86.320 23.760 ;
        RECT 86.160 23.400 86.320 23.470 ;
      LAYER Metal2 ;
        RECT 86.030 23.470 86.320 26.190 ;
    END
  END ON[86]
  PIN ONB[86]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 85.410 23.380 85.710 23.680 ;
        RECT 85.580 23.310 85.710 23.380 ;
        RECT 85.580 22.830 85.710 23.010 ;
      LAYER Metal1 ;
        RECT 85.480 23.470 85.770 23.760 ;
        RECT 85.480 23.400 85.640 23.470 ;
      LAYER Metal2 ;
        RECT 85.480 23.470 85.770 26.190 ;
    END
  END ONB[86]
  PIN ON[87]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 84.090 23.380 84.390 23.680 ;
        RECT 84.090 23.310 84.220 23.380 ;
        RECT 84.090 22.830 84.220 23.010 ;
      LAYER Metal1 ;
        RECT 84.030 23.470 84.320 23.760 ;
        RECT 84.160 23.400 84.320 23.470 ;
      LAYER Metal2 ;
        RECT 84.030 23.470 84.320 26.190 ;
    END
  END ON[87]
  PIN ONB[87]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 83.410 23.380 83.710 23.680 ;
        RECT 83.580 23.310 83.710 23.380 ;
        RECT 83.580 22.830 83.710 23.010 ;
      LAYER Metal1 ;
        RECT 83.480 23.470 83.770 23.760 ;
        RECT 83.480 23.400 83.640 23.470 ;
      LAYER Metal2 ;
        RECT 83.480 23.470 83.770 26.190 ;
    END
  END ONB[87]
  PIN ON[88]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 82.090 23.380 82.390 23.680 ;
        RECT 82.090 23.310 82.220 23.380 ;
        RECT 82.090 22.830 82.220 23.010 ;
      LAYER Metal1 ;
        RECT 82.030 23.470 82.320 23.760 ;
        RECT 82.160 23.400 82.320 23.470 ;
      LAYER Metal2 ;
        RECT 82.030 23.470 82.320 26.190 ;
    END
  END ON[88]
  PIN ONB[88]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 81.410 23.380 81.710 23.680 ;
        RECT 81.580 23.310 81.710 23.380 ;
        RECT 81.580 22.830 81.710 23.010 ;
      LAYER Metal1 ;
        RECT 81.480 23.470 81.770 23.760 ;
        RECT 81.480 23.400 81.640 23.470 ;
      LAYER Metal2 ;
        RECT 81.480 23.470 81.770 26.190 ;
    END
  END ONB[88]
  PIN ON[89]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 80.090 23.380 80.390 23.680 ;
        RECT 80.090 23.310 80.220 23.380 ;
        RECT 80.090 22.830 80.220 23.010 ;
      LAYER Metal1 ;
        RECT 80.030 23.470 80.320 23.760 ;
        RECT 80.160 23.400 80.320 23.470 ;
      LAYER Metal2 ;
        RECT 80.030 23.470 80.320 26.190 ;
    END
  END ON[89]
  PIN ONB[89]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 79.410 23.380 79.710 23.680 ;
        RECT 79.580 23.310 79.710 23.380 ;
        RECT 79.580 22.830 79.710 23.010 ;
      LAYER Metal1 ;
        RECT 79.480 23.470 79.770 23.760 ;
        RECT 79.480 23.400 79.640 23.470 ;
      LAYER Metal2 ;
        RECT 79.480 23.470 79.770 26.190 ;
    END
  END ONB[89]
  PIN ON[90]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 78.090 23.380 78.390 23.680 ;
        RECT 78.090 23.310 78.220 23.380 ;
        RECT 78.090 22.830 78.220 23.010 ;
      LAYER Metal1 ;
        RECT 78.030 23.470 78.320 23.760 ;
        RECT 78.160 23.400 78.320 23.470 ;
      LAYER Metal2 ;
        RECT 78.030 23.470 78.320 26.190 ;
    END
  END ON[90]
  PIN ONB[90]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 77.410 23.380 77.710 23.680 ;
        RECT 77.580 23.310 77.710 23.380 ;
        RECT 77.580 22.830 77.710 23.010 ;
      LAYER Metal1 ;
        RECT 77.480 23.470 77.770 23.760 ;
        RECT 77.480 23.400 77.640 23.470 ;
      LAYER Metal2 ;
        RECT 77.480 23.470 77.770 26.190 ;
    END
  END ONB[90]
  PIN ON[91]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 76.090 23.380 76.390 23.680 ;
        RECT 76.090 23.310 76.220 23.380 ;
        RECT 76.090 22.830 76.220 23.010 ;
      LAYER Metal1 ;
        RECT 76.030 23.470 76.320 23.760 ;
        RECT 76.160 23.400 76.320 23.470 ;
      LAYER Metal2 ;
        RECT 76.030 23.470 76.320 26.190 ;
    END
  END ON[91]
  PIN ONB[91]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 75.410 23.380 75.710 23.680 ;
        RECT 75.580 23.310 75.710 23.380 ;
        RECT 75.580 22.830 75.710 23.010 ;
      LAYER Metal1 ;
        RECT 75.480 23.470 75.770 23.760 ;
        RECT 75.480 23.400 75.640 23.470 ;
      LAYER Metal2 ;
        RECT 75.480 23.470 75.770 26.190 ;
    END
  END ONB[91]
  PIN ON[92]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 74.090 23.380 74.390 23.680 ;
        RECT 74.090 23.310 74.220 23.380 ;
        RECT 74.090 22.830 74.220 23.010 ;
      LAYER Metal1 ;
        RECT 74.030 23.470 74.320 23.760 ;
        RECT 74.160 23.400 74.320 23.470 ;
      LAYER Metal2 ;
        RECT 74.030 23.470 74.320 26.190 ;
    END
  END ON[92]
  PIN ONB[92]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 73.410 23.380 73.710 23.680 ;
        RECT 73.580 23.310 73.710 23.380 ;
        RECT 73.580 22.830 73.710 23.010 ;
      LAYER Metal1 ;
        RECT 73.480 23.470 73.770 23.760 ;
        RECT 73.480 23.400 73.640 23.470 ;
      LAYER Metal2 ;
        RECT 73.480 23.470 73.770 26.190 ;
    END
  END ONB[92]
  PIN ON[93]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 72.090 23.380 72.390 23.680 ;
        RECT 72.090 23.310 72.220 23.380 ;
        RECT 72.090 22.830 72.220 23.010 ;
      LAYER Metal1 ;
        RECT 72.030 23.470 72.320 23.760 ;
        RECT 72.160 23.400 72.320 23.470 ;
      LAYER Metal2 ;
        RECT 72.030 23.470 72.320 26.190 ;
    END
  END ON[93]
  PIN ONB[93]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 71.410 23.380 71.710 23.680 ;
        RECT 71.580 23.310 71.710 23.380 ;
        RECT 71.580 22.830 71.710 23.010 ;
      LAYER Metal1 ;
        RECT 71.480 23.470 71.770 23.760 ;
        RECT 71.480 23.400 71.640 23.470 ;
      LAYER Metal2 ;
        RECT 71.480 23.470 71.770 26.190 ;
    END
  END ONB[93]
  PIN ON[94]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 70.090 23.380 70.390 23.680 ;
        RECT 70.090 23.310 70.220 23.380 ;
        RECT 70.090 22.830 70.220 23.010 ;
      LAYER Metal1 ;
        RECT 70.030 23.470 70.320 23.760 ;
        RECT 70.160 23.400 70.320 23.470 ;
      LAYER Metal2 ;
        RECT 70.030 23.470 70.320 26.190 ;
    END
  END ON[94]
  PIN ONB[94]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 69.410 23.380 69.710 23.680 ;
        RECT 69.580 23.310 69.710 23.380 ;
        RECT 69.580 22.830 69.710 23.010 ;
      LAYER Metal1 ;
        RECT 69.480 23.470 69.770 23.760 ;
        RECT 69.480 23.400 69.640 23.470 ;
      LAYER Metal2 ;
        RECT 69.480 23.470 69.770 26.190 ;
    END
  END ONB[94]
  PIN ON[95]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 68.090 23.380 68.390 23.680 ;
        RECT 68.090 23.310 68.220 23.380 ;
        RECT 68.090 22.830 68.220 23.010 ;
      LAYER Metal1 ;
        RECT 68.030 23.470 68.320 23.760 ;
        RECT 68.160 23.400 68.320 23.470 ;
      LAYER Metal2 ;
        RECT 68.030 23.470 68.320 26.190 ;
    END
  END ON[95]
  PIN ONB[95]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 67.410 23.380 67.710 23.680 ;
        RECT 67.580 23.310 67.710 23.380 ;
        RECT 67.580 22.830 67.710 23.010 ;
      LAYER Metal1 ;
        RECT 67.480 23.470 67.770 23.760 ;
        RECT 67.480 23.400 67.640 23.470 ;
      LAYER Metal2 ;
        RECT 67.480 23.470 67.770 26.190 ;
    END
  END ONB[95]
  PIN EN[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 132.090 23.380 132.390 23.680 ;
        RECT 132.090 23.310 132.220 23.380 ;
        RECT 132.090 22.830 132.220 23.010 ;
      LAYER Metal1 ;
        RECT 132.030 23.470 132.320 23.760 ;
        RECT 132.160 23.400 132.320 23.470 ;
      LAYER Metal2 ;
        RECT 132.030 23.470 132.320 26.190 ;
    END
  END EN[2]
  PIN ENB[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 131.410 23.380 131.710 23.680 ;
        RECT 131.580 23.310 131.710 23.380 ;
        RECT 131.580 22.830 131.710 23.010 ;
      LAYER Metal1 ;
        RECT 131.480 23.470 131.770 23.760 ;
        RECT 131.480 23.400 131.640 23.470 ;
      LAYER Metal2 ;
        RECT 131.480 23.470 131.770 26.190 ;
    END
  END ENB[2]
  PIN ON[97]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 64.090 23.380 64.390 23.680 ;
        RECT 64.090 23.310 64.220 23.380 ;
        RECT 64.090 22.830 64.220 23.010 ;
      LAYER Metal1 ;
        RECT 64.030 23.470 64.320 23.760 ;
        RECT 64.160 23.400 64.320 23.470 ;
      LAYER Metal2 ;
        RECT 64.030 23.470 64.320 26.190 ;
    END
  END ON[97]
  PIN ONB[97]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 63.410 23.380 63.710 23.680 ;
        RECT 63.580 23.310 63.710 23.380 ;
        RECT 63.580 22.830 63.710 23.010 ;
      LAYER Metal1 ;
        RECT 63.480 23.470 63.770 23.760 ;
        RECT 63.480 23.400 63.640 23.470 ;
      LAYER Metal2 ;
        RECT 63.480 23.470 63.770 26.190 ;
    END
  END ONB[97]
  PIN ON[98]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 62.090 23.380 62.390 23.680 ;
        RECT 62.090 23.310 62.220 23.380 ;
        RECT 62.090 22.830 62.220 23.010 ;
      LAYER Metal1 ;
        RECT 62.030 23.470 62.320 23.760 ;
        RECT 62.160 23.400 62.320 23.470 ;
      LAYER Metal2 ;
        RECT 62.030 23.470 62.320 26.190 ;
    END
  END ON[98]
  PIN ONB[98]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 61.410 23.380 61.710 23.680 ;
        RECT 61.580 23.310 61.710 23.380 ;
        RECT 61.580 22.830 61.710 23.010 ;
      LAYER Metal1 ;
        RECT 61.480 23.470 61.770 23.760 ;
        RECT 61.480 23.400 61.640 23.470 ;
      LAYER Metal2 ;
        RECT 61.480 23.470 61.770 26.190 ;
    END
  END ONB[98]
  PIN ON[99]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 60.090 23.380 60.390 23.680 ;
        RECT 60.090 23.310 60.220 23.380 ;
        RECT 60.090 22.830 60.220 23.010 ;
      LAYER Metal1 ;
        RECT 60.030 23.470 60.320 23.760 ;
        RECT 60.160 23.400 60.320 23.470 ;
      LAYER Metal2 ;
        RECT 60.030 23.470 60.320 26.190 ;
    END
  END ON[99]
  PIN ONB[99]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 59.410 23.380 59.710 23.680 ;
        RECT 59.580 23.310 59.710 23.380 ;
        RECT 59.580 22.830 59.710 23.010 ;
      LAYER Metal1 ;
        RECT 59.480 23.470 59.770 23.760 ;
        RECT 59.480 23.400 59.640 23.470 ;
      LAYER Metal2 ;
        RECT 59.480 23.470 59.770 26.190 ;
    END
  END ONB[99]
  PIN ON[100]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 58.090 23.380 58.390 23.680 ;
        RECT 58.090 23.310 58.220 23.380 ;
        RECT 58.090 22.830 58.220 23.010 ;
      LAYER Metal1 ;
        RECT 58.030 23.470 58.320 23.760 ;
        RECT 58.160 23.400 58.320 23.470 ;
      LAYER Metal2 ;
        RECT 58.030 23.470 58.320 26.190 ;
    END
  END ON[100]
  PIN ONB[100]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 57.410 23.380 57.710 23.680 ;
        RECT 57.580 23.310 57.710 23.380 ;
        RECT 57.580 22.830 57.710 23.010 ;
      LAYER Metal1 ;
        RECT 57.480 23.470 57.770 23.760 ;
        RECT 57.480 23.400 57.640 23.470 ;
      LAYER Metal2 ;
        RECT 57.480 23.470 57.770 26.190 ;
    END
  END ONB[100]
  PIN ON[101]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 56.090 23.380 56.390 23.680 ;
        RECT 56.090 23.310 56.220 23.380 ;
        RECT 56.090 22.830 56.220 23.010 ;
      LAYER Metal1 ;
        RECT 56.030 23.470 56.320 23.760 ;
        RECT 56.160 23.400 56.320 23.470 ;
      LAYER Metal2 ;
        RECT 56.030 23.470 56.320 26.190 ;
    END
  END ON[101]
  PIN ONB[101]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 55.410 23.380 55.710 23.680 ;
        RECT 55.580 23.310 55.710 23.380 ;
        RECT 55.580 22.830 55.710 23.010 ;
      LAYER Metal1 ;
        RECT 55.480 23.470 55.770 23.760 ;
        RECT 55.480 23.400 55.640 23.470 ;
      LAYER Metal2 ;
        RECT 55.480 23.470 55.770 26.190 ;
    END
  END ONB[101]
  PIN ON[102]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 54.090 23.380 54.390 23.680 ;
        RECT 54.090 23.310 54.220 23.380 ;
        RECT 54.090 22.830 54.220 23.010 ;
      LAYER Metal1 ;
        RECT 54.030 23.470 54.320 23.760 ;
        RECT 54.160 23.400 54.320 23.470 ;
      LAYER Metal2 ;
        RECT 54.030 23.470 54.320 26.190 ;
    END
  END ON[102]
  PIN ONB[102]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 53.410 23.380 53.710 23.680 ;
        RECT 53.580 23.310 53.710 23.380 ;
        RECT 53.580 22.830 53.710 23.010 ;
      LAYER Metal1 ;
        RECT 53.480 23.470 53.770 23.760 ;
        RECT 53.480 23.400 53.640 23.470 ;
      LAYER Metal2 ;
        RECT 53.480 23.470 53.770 26.190 ;
    END
  END ONB[102]
  PIN ON[103]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 52.090 23.380 52.390 23.680 ;
        RECT 52.090 23.310 52.220 23.380 ;
        RECT 52.090 22.830 52.220 23.010 ;
      LAYER Metal1 ;
        RECT 52.030 23.470 52.320 23.760 ;
        RECT 52.160 23.400 52.320 23.470 ;
      LAYER Metal2 ;
        RECT 52.030 23.470 52.320 26.190 ;
    END
  END ON[103]
  PIN ONB[103]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 51.410 23.380 51.710 23.680 ;
        RECT 51.580 23.310 51.710 23.380 ;
        RECT 51.580 22.830 51.710 23.010 ;
      LAYER Metal1 ;
        RECT 51.480 23.470 51.770 23.760 ;
        RECT 51.480 23.400 51.640 23.470 ;
      LAYER Metal2 ;
        RECT 51.480 23.470 51.770 26.190 ;
    END
  END ONB[103]
  PIN ON[104]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 50.090 23.380 50.390 23.680 ;
        RECT 50.090 23.310 50.220 23.380 ;
        RECT 50.090 22.830 50.220 23.010 ;
      LAYER Metal1 ;
        RECT 50.030 23.470 50.320 23.760 ;
        RECT 50.160 23.400 50.320 23.470 ;
      LAYER Metal2 ;
        RECT 50.030 23.470 50.320 26.190 ;
    END
  END ON[104]
  PIN ONB[104]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 49.410 23.380 49.710 23.680 ;
        RECT 49.580 23.310 49.710 23.380 ;
        RECT 49.580 22.830 49.710 23.010 ;
      LAYER Metal1 ;
        RECT 49.480 23.470 49.770 23.760 ;
        RECT 49.480 23.400 49.640 23.470 ;
      LAYER Metal2 ;
        RECT 49.480 23.470 49.770 26.190 ;
    END
  END ONB[104]
  PIN ON[105]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 48.090 23.380 48.390 23.680 ;
        RECT 48.090 23.310 48.220 23.380 ;
        RECT 48.090 22.830 48.220 23.010 ;
      LAYER Metal1 ;
        RECT 48.030 23.470 48.320 23.760 ;
        RECT 48.160 23.400 48.320 23.470 ;
      LAYER Metal2 ;
        RECT 48.030 23.470 48.320 26.190 ;
    END
  END ON[105]
  PIN ONB[105]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 47.410 23.380 47.710 23.680 ;
        RECT 47.580 23.310 47.710 23.380 ;
        RECT 47.580 22.830 47.710 23.010 ;
      LAYER Metal1 ;
        RECT 47.480 23.470 47.770 23.760 ;
        RECT 47.480 23.400 47.640 23.470 ;
      LAYER Metal2 ;
        RECT 47.480 23.470 47.770 26.190 ;
    END
  END ONB[105]
  PIN ON[106]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 46.090 23.380 46.390 23.680 ;
        RECT 46.090 23.310 46.220 23.380 ;
        RECT 46.090 22.830 46.220 23.010 ;
      LAYER Metal1 ;
        RECT 46.030 23.470 46.320 23.760 ;
        RECT 46.160 23.400 46.320 23.470 ;
      LAYER Metal2 ;
        RECT 46.030 23.470 46.320 26.190 ;
    END
  END ON[106]
  PIN ONB[106]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 45.410 23.380 45.710 23.680 ;
        RECT 45.580 23.310 45.710 23.380 ;
        RECT 45.580 22.830 45.710 23.010 ;
      LAYER Metal1 ;
        RECT 45.480 23.470 45.770 23.760 ;
        RECT 45.480 23.400 45.640 23.470 ;
      LAYER Metal2 ;
        RECT 45.480 23.470 45.770 26.190 ;
    END
  END ONB[106]
  PIN ON[107]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 44.090 23.380 44.390 23.680 ;
        RECT 44.090 23.310 44.220 23.380 ;
        RECT 44.090 22.830 44.220 23.010 ;
      LAYER Metal1 ;
        RECT 44.030 23.470 44.320 23.760 ;
        RECT 44.160 23.400 44.320 23.470 ;
      LAYER Metal2 ;
        RECT 44.030 23.470 44.320 26.190 ;
    END
  END ON[107]
  PIN ONB[107]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 43.410 23.380 43.710 23.680 ;
        RECT 43.580 23.310 43.710 23.380 ;
        RECT 43.580 22.830 43.710 23.010 ;
      LAYER Metal1 ;
        RECT 43.480 23.470 43.770 23.760 ;
        RECT 43.480 23.400 43.640 23.470 ;
      LAYER Metal2 ;
        RECT 43.480 23.470 43.770 26.190 ;
    END
  END ONB[107]
  PIN ON[108]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 42.090 23.380 42.390 23.680 ;
        RECT 42.090 23.310 42.220 23.380 ;
        RECT 42.090 22.830 42.220 23.010 ;
      LAYER Metal1 ;
        RECT 42.030 23.470 42.320 23.760 ;
        RECT 42.160 23.400 42.320 23.470 ;
      LAYER Metal2 ;
        RECT 42.030 23.470 42.320 26.190 ;
    END
  END ON[108]
  PIN ONB[108]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 41.410 23.380 41.710 23.680 ;
        RECT 41.580 23.310 41.710 23.380 ;
        RECT 41.580 22.830 41.710 23.010 ;
      LAYER Metal1 ;
        RECT 41.480 23.470 41.770 23.760 ;
        RECT 41.480 23.400 41.640 23.470 ;
      LAYER Metal2 ;
        RECT 41.480 23.470 41.770 26.190 ;
    END
  END ONB[108]
  PIN ON[109]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 40.090 23.380 40.390 23.680 ;
        RECT 40.090 23.310 40.220 23.380 ;
        RECT 40.090 22.830 40.220 23.010 ;
      LAYER Metal1 ;
        RECT 40.030 23.470 40.320 23.760 ;
        RECT 40.160 23.400 40.320 23.470 ;
      LAYER Metal2 ;
        RECT 40.030 23.470 40.320 26.190 ;
    END
  END ON[109]
  PIN ONB[109]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 39.410 23.380 39.710 23.680 ;
        RECT 39.580 23.310 39.710 23.380 ;
        RECT 39.580 22.830 39.710 23.010 ;
      LAYER Metal1 ;
        RECT 39.480 23.470 39.770 23.760 ;
        RECT 39.480 23.400 39.640 23.470 ;
      LAYER Metal2 ;
        RECT 39.480 23.470 39.770 26.190 ;
    END
  END ONB[109]
  PIN ON[110]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 38.090 23.380 38.390 23.680 ;
        RECT 38.090 23.310 38.220 23.380 ;
        RECT 38.090 22.830 38.220 23.010 ;
      LAYER Metal1 ;
        RECT 38.030 23.470 38.320 23.760 ;
        RECT 38.160 23.400 38.320 23.470 ;
      LAYER Metal2 ;
        RECT 38.030 23.470 38.320 26.190 ;
    END
  END ON[110]
  PIN ONB[110]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 37.410 23.380 37.710 23.680 ;
        RECT 37.580 23.310 37.710 23.380 ;
        RECT 37.580 22.830 37.710 23.010 ;
      LAYER Metal1 ;
        RECT 37.480 23.470 37.770 23.760 ;
        RECT 37.480 23.400 37.640 23.470 ;
      LAYER Metal2 ;
        RECT 37.480 23.470 37.770 26.190 ;
    END
  END ONB[110]
  PIN ON[111]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 36.090 23.380 36.390 23.680 ;
        RECT 36.090 23.310 36.220 23.380 ;
        RECT 36.090 22.830 36.220 23.010 ;
      LAYER Metal1 ;
        RECT 36.030 23.470 36.320 23.760 ;
        RECT 36.160 23.400 36.320 23.470 ;
      LAYER Metal2 ;
        RECT 36.030 23.470 36.320 26.190 ;
    END
  END ON[111]
  PIN ONB[111]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 35.410 23.380 35.710 23.680 ;
        RECT 35.580 23.310 35.710 23.380 ;
        RECT 35.580 22.830 35.710 23.010 ;
      LAYER Metal1 ;
        RECT 35.480 23.470 35.770 23.760 ;
        RECT 35.480 23.400 35.640 23.470 ;
      LAYER Metal2 ;
        RECT 35.480 23.470 35.770 26.190 ;
    END
  END ONB[111]
  PIN ON[112]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 34.090 23.380 34.390 23.680 ;
        RECT 34.090 23.310 34.220 23.380 ;
        RECT 34.090 22.830 34.220 23.010 ;
      LAYER Metal1 ;
        RECT 34.030 23.470 34.320 23.760 ;
        RECT 34.160 23.400 34.320 23.470 ;
      LAYER Metal2 ;
        RECT 34.030 23.470 34.320 26.190 ;
    END
  END ON[112]
  PIN ONB[112]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 33.410 23.380 33.710 23.680 ;
        RECT 33.580 23.310 33.710 23.380 ;
        RECT 33.580 22.830 33.710 23.010 ;
      LAYER Metal1 ;
        RECT 33.480 23.470 33.770 23.760 ;
        RECT 33.480 23.400 33.640 23.470 ;
      LAYER Metal2 ;
        RECT 33.480 23.470 33.770 26.190 ;
    END
  END ONB[112]
  PIN ON[113]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 32.090 23.380 32.390 23.680 ;
        RECT 32.090 23.310 32.220 23.380 ;
        RECT 32.090 22.830 32.220 23.010 ;
      LAYER Metal1 ;
        RECT 32.030 23.470 32.320 23.760 ;
        RECT 32.160 23.400 32.320 23.470 ;
      LAYER Metal2 ;
        RECT 32.030 23.470 32.320 26.190 ;
    END
  END ON[113]
  PIN ONB[113]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 31.410 23.380 31.710 23.680 ;
        RECT 31.580 23.310 31.710 23.380 ;
        RECT 31.580 22.830 31.710 23.010 ;
      LAYER Metal1 ;
        RECT 31.480 23.470 31.770 23.760 ;
        RECT 31.480 23.400 31.640 23.470 ;
      LAYER Metal2 ;
        RECT 31.480 23.470 31.770 26.190 ;
    END
  END ONB[113]
  PIN ON[114]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 30.090 23.380 30.390 23.680 ;
        RECT 30.090 23.310 30.220 23.380 ;
        RECT 30.090 22.830 30.220 23.010 ;
      LAYER Metal1 ;
        RECT 30.030 23.470 30.320 23.760 ;
        RECT 30.160 23.400 30.320 23.470 ;
      LAYER Metal2 ;
        RECT 30.030 23.470 30.320 26.190 ;
    END
  END ON[114]
  PIN ONB[114]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 29.410 23.380 29.710 23.680 ;
        RECT 29.580 23.310 29.710 23.380 ;
        RECT 29.580 22.830 29.710 23.010 ;
      LAYER Metal1 ;
        RECT 29.480 23.470 29.770 23.760 ;
        RECT 29.480 23.400 29.640 23.470 ;
      LAYER Metal2 ;
        RECT 29.480 23.470 29.770 26.190 ;
    END
  END ONB[114]
  PIN ON[115]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 28.090 23.380 28.390 23.680 ;
        RECT 28.090 23.310 28.220 23.380 ;
        RECT 28.090 22.830 28.220 23.010 ;
      LAYER Metal1 ;
        RECT 28.030 23.470 28.320 23.760 ;
        RECT 28.160 23.400 28.320 23.470 ;
      LAYER Metal2 ;
        RECT 28.030 23.470 28.320 26.190 ;
    END
  END ON[115]
  PIN ONB[115]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 27.410 23.380 27.710 23.680 ;
        RECT 27.580 23.310 27.710 23.380 ;
        RECT 27.580 22.830 27.710 23.010 ;
      LAYER Metal1 ;
        RECT 27.480 23.470 27.770 23.760 ;
        RECT 27.480 23.400 27.640 23.470 ;
      LAYER Metal2 ;
        RECT 27.480 23.470 27.770 26.190 ;
    END
  END ONB[115]
  PIN ON[116]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 26.090 23.380 26.390 23.680 ;
        RECT 26.090 23.310 26.220 23.380 ;
        RECT 26.090 22.830 26.220 23.010 ;
      LAYER Metal1 ;
        RECT 26.030 23.470 26.320 23.760 ;
        RECT 26.160 23.400 26.320 23.470 ;
      LAYER Metal2 ;
        RECT 26.030 23.470 26.320 26.190 ;
    END
  END ON[116]
  PIN ONB[116]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 25.410 23.380 25.710 23.680 ;
        RECT 25.580 23.310 25.710 23.380 ;
        RECT 25.580 22.830 25.710 23.010 ;
      LAYER Metal1 ;
        RECT 25.480 23.470 25.770 23.760 ;
        RECT 25.480 23.400 25.640 23.470 ;
      LAYER Metal2 ;
        RECT 25.480 23.470 25.770 26.190 ;
    END
  END ONB[116]
  PIN ON[117]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 24.090 23.380 24.390 23.680 ;
        RECT 24.090 23.310 24.220 23.380 ;
        RECT 24.090 22.830 24.220 23.010 ;
      LAYER Metal1 ;
        RECT 24.030 23.470 24.320 23.760 ;
        RECT 24.160 23.400 24.320 23.470 ;
      LAYER Metal2 ;
        RECT 24.030 23.470 24.320 26.190 ;
    END
  END ON[117]
  PIN ONB[117]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 23.410 23.380 23.710 23.680 ;
        RECT 23.580 23.310 23.710 23.380 ;
        RECT 23.580 22.830 23.710 23.010 ;
      LAYER Metal1 ;
        RECT 23.480 23.470 23.770 23.760 ;
        RECT 23.480 23.400 23.640 23.470 ;
      LAYER Metal2 ;
        RECT 23.480 23.470 23.770 26.190 ;
    END
  END ONB[117]
  PIN ON[118]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 22.090 23.380 22.390 23.680 ;
        RECT 22.090 23.310 22.220 23.380 ;
        RECT 22.090 22.830 22.220 23.010 ;
      LAYER Metal1 ;
        RECT 22.030 23.470 22.320 23.760 ;
        RECT 22.160 23.400 22.320 23.470 ;
      LAYER Metal2 ;
        RECT 22.030 23.470 22.320 26.190 ;
    END
  END ON[118]
  PIN ONB[118]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 21.410 23.380 21.710 23.680 ;
        RECT 21.580 23.310 21.710 23.380 ;
        RECT 21.580 22.830 21.710 23.010 ;
      LAYER Metal1 ;
        RECT 21.480 23.470 21.770 23.760 ;
        RECT 21.480 23.400 21.640 23.470 ;
      LAYER Metal2 ;
        RECT 21.480 23.470 21.770 26.190 ;
    END
  END ONB[118]
  PIN ON[119]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 20.090 23.380 20.390 23.680 ;
        RECT 20.090 23.310 20.220 23.380 ;
        RECT 20.090 22.830 20.220 23.010 ;
      LAYER Metal1 ;
        RECT 20.030 23.470 20.320 23.760 ;
        RECT 20.160 23.400 20.320 23.470 ;
      LAYER Metal2 ;
        RECT 20.030 23.470 20.320 26.190 ;
    END
  END ON[119]
  PIN ONB[119]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 19.410 23.380 19.710 23.680 ;
        RECT 19.580 23.310 19.710 23.380 ;
        RECT 19.580 22.830 19.710 23.010 ;
      LAYER Metal1 ;
        RECT 19.480 23.470 19.770 23.760 ;
        RECT 19.480 23.400 19.640 23.470 ;
      LAYER Metal2 ;
        RECT 19.480 23.470 19.770 26.190 ;
    END
  END ONB[119]
  PIN ON[120]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 18.090 23.380 18.390 23.680 ;
        RECT 18.090 23.310 18.220 23.380 ;
        RECT 18.090 22.830 18.220 23.010 ;
      LAYER Metal1 ;
        RECT 18.030 23.470 18.320 23.760 ;
        RECT 18.160 23.400 18.320 23.470 ;
      LAYER Metal2 ;
        RECT 18.030 23.470 18.320 26.190 ;
    END
  END ON[120]
  PIN ONB[120]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 17.410 23.380 17.710 23.680 ;
        RECT 17.580 23.310 17.710 23.380 ;
        RECT 17.580 22.830 17.710 23.010 ;
      LAYER Metal1 ;
        RECT 17.480 23.470 17.770 23.760 ;
        RECT 17.480 23.400 17.640 23.470 ;
      LAYER Metal2 ;
        RECT 17.480 23.470 17.770 26.190 ;
    END
  END ONB[120]
  PIN ON[121]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 16.090 23.380 16.390 23.680 ;
        RECT 16.090 23.310 16.220 23.380 ;
        RECT 16.090 22.830 16.220 23.010 ;
      LAYER Metal1 ;
        RECT 16.030 23.470 16.320 23.760 ;
        RECT 16.160 23.400 16.320 23.470 ;
      LAYER Metal2 ;
        RECT 16.030 23.470 16.320 26.190 ;
    END
  END ON[121]
  PIN ONB[121]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 15.410 23.380 15.710 23.680 ;
        RECT 15.580 23.310 15.710 23.380 ;
        RECT 15.580 22.830 15.710 23.010 ;
      LAYER Metal1 ;
        RECT 15.480 23.470 15.770 23.760 ;
        RECT 15.480 23.400 15.640 23.470 ;
      LAYER Metal2 ;
        RECT 15.480 23.470 15.770 26.190 ;
    END
  END ONB[121]
  PIN ON[122]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 14.090 23.380 14.390 23.680 ;
        RECT 14.090 23.310 14.220 23.380 ;
        RECT 14.090 22.830 14.220 23.010 ;
      LAYER Metal1 ;
        RECT 14.030 23.470 14.320 23.760 ;
        RECT 14.160 23.400 14.320 23.470 ;
      LAYER Metal2 ;
        RECT 14.030 23.470 14.320 26.190 ;
    END
  END ON[122]
  PIN ONB[122]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 13.410 23.380 13.710 23.680 ;
        RECT 13.580 23.310 13.710 23.380 ;
        RECT 13.580 22.830 13.710 23.010 ;
      LAYER Metal1 ;
        RECT 13.480 23.470 13.770 23.760 ;
        RECT 13.480 23.400 13.640 23.470 ;
      LAYER Metal2 ;
        RECT 13.480 23.470 13.770 26.190 ;
    END
  END ONB[122]
  PIN ON[123]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 12.090 23.380 12.390 23.680 ;
        RECT 12.090 23.310 12.220 23.380 ;
        RECT 12.090 22.830 12.220 23.010 ;
      LAYER Metal1 ;
        RECT 12.030 23.470 12.320 23.760 ;
        RECT 12.160 23.400 12.320 23.470 ;
      LAYER Metal2 ;
        RECT 12.030 23.470 12.320 26.190 ;
    END
  END ON[123]
  PIN ONB[123]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 11.410 23.380 11.710 23.680 ;
        RECT 11.580 23.310 11.710 23.380 ;
        RECT 11.580 22.830 11.710 23.010 ;
      LAYER Metal1 ;
        RECT 11.480 23.470 11.770 23.760 ;
        RECT 11.480 23.400 11.640 23.470 ;
      LAYER Metal2 ;
        RECT 11.480 23.470 11.770 26.190 ;
    END
  END ONB[123]
  PIN ON[124]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 10.090 23.380 10.390 23.680 ;
        RECT 10.090 23.310 10.220 23.380 ;
        RECT 10.090 22.830 10.220 23.010 ;
      LAYER Metal1 ;
        RECT 10.030 23.470 10.320 23.760 ;
        RECT 10.160 23.400 10.320 23.470 ;
      LAYER Metal2 ;
        RECT 10.030 23.470 10.320 26.190 ;
    END
  END ON[124]
  PIN ONB[124]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 9.410 23.380 9.710 23.680 ;
        RECT 9.580 23.310 9.710 23.380 ;
        RECT 9.580 22.830 9.710 23.010 ;
      LAYER Metal1 ;
        RECT 9.480 23.470 9.770 23.760 ;
        RECT 9.480 23.400 9.640 23.470 ;
      LAYER Metal2 ;
        RECT 9.480 23.470 9.770 26.190 ;
    END
  END ONB[124]
  PIN ON[125]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 8.090 23.380 8.390 23.680 ;
        RECT 8.090 23.310 8.220 23.380 ;
        RECT 8.090 22.830 8.220 23.010 ;
      LAYER Metal1 ;
        RECT 8.030 23.470 8.320 23.760 ;
        RECT 8.160 23.400 8.320 23.470 ;
      LAYER Metal2 ;
        RECT 8.030 23.470 8.320 26.190 ;
    END
  END ON[125]
  PIN ONB[125]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 7.410 23.380 7.710 23.680 ;
        RECT 7.580 23.310 7.710 23.380 ;
        RECT 7.580 22.830 7.710 23.010 ;
      LAYER Metal1 ;
        RECT 7.480 23.470 7.770 23.760 ;
        RECT 7.480 23.400 7.640 23.470 ;
      LAYER Metal2 ;
        RECT 7.480 23.470 7.770 26.190 ;
    END
  END ONB[125]
  PIN ON[126]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 6.090 23.380 6.390 23.680 ;
        RECT 6.090 23.310 6.220 23.380 ;
        RECT 6.090 22.830 6.220 23.010 ;
      LAYER Metal1 ;
        RECT 6.030 23.470 6.320 23.760 ;
        RECT 6.160 23.400 6.320 23.470 ;
      LAYER Metal2 ;
        RECT 6.030 23.470 6.320 26.190 ;
    END
  END ON[126]
  PIN ONB[126]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 5.410 23.380 5.710 23.680 ;
        RECT 5.580 23.310 5.710 23.380 ;
        RECT 5.580 22.830 5.710 23.010 ;
      LAYER Metal1 ;
        RECT 5.480 23.470 5.770 23.760 ;
        RECT 5.480 23.400 5.640 23.470 ;
      LAYER Metal2 ;
        RECT 5.480 23.470 5.770 26.190 ;
    END
  END ONB[126]
  PIN ON[127]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 4.090 23.380 4.390 23.680 ;
        RECT 4.090 23.310 4.220 23.380 ;
        RECT 4.090 22.830 4.220 23.010 ;
      LAYER Metal1 ;
        RECT 4.030 23.470 4.320 23.760 ;
        RECT 4.160 23.400 4.320 23.470 ;
      LAYER Metal2 ;
        RECT 4.030 23.470 4.320 26.190 ;
    END
  END ON[127]
  PIN ONB[127]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.410 23.380 3.710 23.680 ;
        RECT 3.580 23.310 3.710 23.380 ;
        RECT 3.580 22.830 3.710 23.010 ;
      LAYER Metal1 ;
        RECT 3.480 23.470 3.770 23.760 ;
        RECT 3.480 23.400 3.640 23.470 ;
      LAYER Metal2 ;
        RECT 3.480 23.470 3.770 26.190 ;
    END
  END ONB[127]
  PIN ON[96]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 66.090 23.380 66.390 23.680 ;
        RECT 66.090 23.310 66.220 23.380 ;
        RECT 66.090 22.830 66.220 23.010 ;
      LAYER Metal1 ;
        RECT 66.030 23.470 66.320 23.760 ;
        RECT 66.160 23.400 66.320 23.470 ;
      LAYER Metal2 ;
        RECT 66.030 23.470 66.320 26.190 ;
    END
  END ON[96]
  PIN ONB[96]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 65.410 23.380 65.710 23.680 ;
        RECT 65.580 23.310 65.710 23.380 ;
        RECT 65.580 22.830 65.710 23.010 ;
      LAYER Metal1 ;
        RECT 65.480 23.470 65.770 23.760 ;
        RECT 65.480 23.400 65.640 23.470 ;
      LAYER Metal2 ;
        RECT 65.480 23.470 65.770 26.190 ;
    END
  END ONB[96]
  PIN EN[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.090 23.380 2.390 23.680 ;
        RECT 2.090 23.310 2.220 23.380 ;
        RECT 2.090 22.830 2.220 23.010 ;
      LAYER Metal1 ;
        RECT 2.030 23.470 2.320 23.760 ;
        RECT 2.160 23.400 2.320 23.470 ;
      LAYER Metal2 ;
        RECT 2.030 23.470 2.320 26.190 ;
    END
  END EN[3]
  PIN ENB[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.410 23.380 1.710 23.680 ;
        RECT 1.580 23.310 1.710 23.380 ;
        RECT 1.580 22.830 1.710 23.010 ;
      LAYER Metal1 ;
        RECT 1.480 23.470 1.770 23.760 ;
        RECT 1.480 23.400 1.640 23.470 ;
      LAYER Metal2 ;
        RECT 1.480 23.470 1.770 26.190 ;
    END
  END ENB[3]
  PIN ON[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 3.580 3.180 3.710 3.360 ;
        RECT 3.580 2.810 3.710 2.880 ;
        RECT 3.410 2.510 3.710 2.810 ;
      LAYER Metal1 ;
        RECT 3.480 2.720 3.640 2.790 ;
        RECT 3.480 2.430 3.770 2.720 ;
      LAYER Metal2 ;
        RECT 3.480 0.000 3.770 2.720 ;
    END
  END ON[0]
  PIN ONB[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 4.090 3.180 4.220 3.360 ;
        RECT 4.090 2.810 4.220 2.880 ;
        RECT 4.090 2.510 4.390 2.810 ;
      LAYER Metal1 ;
        RECT 4.160 2.720 4.320 2.790 ;
        RECT 4.030 2.430 4.320 2.720 ;
      LAYER Metal2 ;
        RECT 4.030 0.000 4.320 2.720 ;
    END
  END ONB[0]
  PIN ON[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 5.580 3.180 5.710 3.360 ;
        RECT 5.580 2.810 5.710 2.880 ;
        RECT 5.410 2.510 5.710 2.810 ;
      LAYER Metal1 ;
        RECT 5.480 2.720 5.640 2.790 ;
        RECT 5.480 2.430 5.770 2.720 ;
      LAYER Metal2 ;
        RECT 5.480 0.000 5.770 2.720 ;
    END
  END ON[1]
  PIN ONB[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 6.090 3.180 6.220 3.360 ;
        RECT 6.090 2.810 6.220 2.880 ;
        RECT 6.090 2.510 6.390 2.810 ;
      LAYER Metal1 ;
        RECT 6.160 2.720 6.320 2.790 ;
        RECT 6.030 2.430 6.320 2.720 ;
      LAYER Metal2 ;
        RECT 6.030 0.000 6.320 2.720 ;
    END
  END ONB[1]
  PIN ON[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 7.580 3.180 7.710 3.360 ;
        RECT 7.580 2.810 7.710 2.880 ;
        RECT 7.410 2.510 7.710 2.810 ;
      LAYER Metal1 ;
        RECT 7.480 2.720 7.640 2.790 ;
        RECT 7.480 2.430 7.770 2.720 ;
      LAYER Metal2 ;
        RECT 7.480 0.000 7.770 2.720 ;
    END
  END ON[2]
  PIN ONB[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 8.090 3.180 8.220 3.360 ;
        RECT 8.090 2.810 8.220 2.880 ;
        RECT 8.090 2.510 8.390 2.810 ;
      LAYER Metal1 ;
        RECT 8.160 2.720 8.320 2.790 ;
        RECT 8.030 2.430 8.320 2.720 ;
      LAYER Metal2 ;
        RECT 8.030 0.000 8.320 2.720 ;
    END
  END ONB[2]
  PIN ON[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 9.580 3.180 9.710 3.360 ;
        RECT 9.580 2.810 9.710 2.880 ;
        RECT 9.410 2.510 9.710 2.810 ;
      LAYER Metal1 ;
        RECT 9.480 2.720 9.640 2.790 ;
        RECT 9.480 2.430 9.770 2.720 ;
      LAYER Metal2 ;
        RECT 9.480 0.000 9.770 2.720 ;
    END
  END ON[3]
  PIN ONB[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 10.090 3.180 10.220 3.360 ;
        RECT 10.090 2.810 10.220 2.880 ;
        RECT 10.090 2.510 10.390 2.810 ;
      LAYER Metal1 ;
        RECT 10.160 2.720 10.320 2.790 ;
        RECT 10.030 2.430 10.320 2.720 ;
      LAYER Metal2 ;
        RECT 10.030 0.000 10.320 2.720 ;
    END
  END ONB[3]
  PIN ON[4]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 11.580 3.180 11.710 3.360 ;
        RECT 11.580 2.810 11.710 2.880 ;
        RECT 11.410 2.510 11.710 2.810 ;
      LAYER Metal1 ;
        RECT 11.480 2.720 11.640 2.790 ;
        RECT 11.480 2.430 11.770 2.720 ;
      LAYER Metal2 ;
        RECT 11.480 0.000 11.770 2.720 ;
    END
  END ON[4]
  PIN ONB[4]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 12.090 3.180 12.220 3.360 ;
        RECT 12.090 2.810 12.220 2.880 ;
        RECT 12.090 2.510 12.390 2.810 ;
      LAYER Metal1 ;
        RECT 12.160 2.720 12.320 2.790 ;
        RECT 12.030 2.430 12.320 2.720 ;
      LAYER Metal2 ;
        RECT 12.030 0.000 12.320 2.720 ;
    END
  END ONB[4]
  PIN ON[5]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 13.580 3.180 13.710 3.360 ;
        RECT 13.580 2.810 13.710 2.880 ;
        RECT 13.410 2.510 13.710 2.810 ;
      LAYER Metal1 ;
        RECT 13.480 2.720 13.640 2.790 ;
        RECT 13.480 2.430 13.770 2.720 ;
      LAYER Metal2 ;
        RECT 13.480 0.000 13.770 2.720 ;
    END
  END ON[5]
  PIN ONB[5]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 14.090 3.180 14.220 3.360 ;
        RECT 14.090 2.810 14.220 2.880 ;
        RECT 14.090 2.510 14.390 2.810 ;
      LAYER Metal1 ;
        RECT 14.160 2.720 14.320 2.790 ;
        RECT 14.030 2.430 14.320 2.720 ;
      LAYER Metal2 ;
        RECT 14.030 0.000 14.320 2.720 ;
    END
  END ONB[5]
  PIN ON[6]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 15.580 3.180 15.710 3.360 ;
        RECT 15.580 2.810 15.710 2.880 ;
        RECT 15.410 2.510 15.710 2.810 ;
      LAYER Metal1 ;
        RECT 15.480 2.720 15.640 2.790 ;
        RECT 15.480 2.430 15.770 2.720 ;
      LAYER Metal2 ;
        RECT 15.480 0.000 15.770 2.720 ;
    END
  END ON[6]
  PIN ONB[6]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 16.090 3.180 16.220 3.360 ;
        RECT 16.090 2.810 16.220 2.880 ;
        RECT 16.090 2.510 16.390 2.810 ;
      LAYER Metal1 ;
        RECT 16.160 2.720 16.320 2.790 ;
        RECT 16.030 2.430 16.320 2.720 ;
      LAYER Metal2 ;
        RECT 16.030 0.000 16.320 2.720 ;
    END
  END ONB[6]
  PIN ON[7]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 17.580 3.180 17.710 3.360 ;
        RECT 17.580 2.810 17.710 2.880 ;
        RECT 17.410 2.510 17.710 2.810 ;
      LAYER Metal1 ;
        RECT 17.480 2.720 17.640 2.790 ;
        RECT 17.480 2.430 17.770 2.720 ;
      LAYER Metal2 ;
        RECT 17.480 0.000 17.770 2.720 ;
    END
  END ON[7]
  PIN ONB[7]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 18.090 3.180 18.220 3.360 ;
        RECT 18.090 2.810 18.220 2.880 ;
        RECT 18.090 2.510 18.390 2.810 ;
      LAYER Metal1 ;
        RECT 18.160 2.720 18.320 2.790 ;
        RECT 18.030 2.430 18.320 2.720 ;
      LAYER Metal2 ;
        RECT 18.030 0.000 18.320 2.720 ;
    END
  END ONB[7]
  PIN ON[8]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 19.580 3.180 19.710 3.360 ;
        RECT 19.580 2.810 19.710 2.880 ;
        RECT 19.410 2.510 19.710 2.810 ;
      LAYER Metal1 ;
        RECT 19.480 2.720 19.640 2.790 ;
        RECT 19.480 2.430 19.770 2.720 ;
      LAYER Metal2 ;
        RECT 19.480 0.000 19.770 2.720 ;
    END
  END ON[8]
  PIN ONB[8]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 20.090 3.180 20.220 3.360 ;
        RECT 20.090 2.810 20.220 2.880 ;
        RECT 20.090 2.510 20.390 2.810 ;
      LAYER Metal1 ;
        RECT 20.160 2.720 20.320 2.790 ;
        RECT 20.030 2.430 20.320 2.720 ;
      LAYER Metal2 ;
        RECT 20.030 0.000 20.320 2.720 ;
    END
  END ONB[8]
  PIN ON[9]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 21.580 3.180 21.710 3.360 ;
        RECT 21.580 2.810 21.710 2.880 ;
        RECT 21.410 2.510 21.710 2.810 ;
      LAYER Metal1 ;
        RECT 21.480 2.720 21.640 2.790 ;
        RECT 21.480 2.430 21.770 2.720 ;
      LAYER Metal2 ;
        RECT 21.480 0.000 21.770 2.720 ;
    END
  END ON[9]
  PIN ONB[9]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 22.090 3.180 22.220 3.360 ;
        RECT 22.090 2.810 22.220 2.880 ;
        RECT 22.090 2.510 22.390 2.810 ;
      LAYER Metal1 ;
        RECT 22.160 2.720 22.320 2.790 ;
        RECT 22.030 2.430 22.320 2.720 ;
      LAYER Metal2 ;
        RECT 22.030 0.000 22.320 2.720 ;
    END
  END ONB[9]
  PIN ON[10]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 23.580 3.180 23.710 3.360 ;
        RECT 23.580 2.810 23.710 2.880 ;
        RECT 23.410 2.510 23.710 2.810 ;
      LAYER Metal1 ;
        RECT 23.480 2.720 23.640 2.790 ;
        RECT 23.480 2.430 23.770 2.720 ;
      LAYER Metal2 ;
        RECT 23.480 0.000 23.770 2.720 ;
    END
  END ON[10]
  PIN ONB[10]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 24.090 3.180 24.220 3.360 ;
        RECT 24.090 2.810 24.220 2.880 ;
        RECT 24.090 2.510 24.390 2.810 ;
      LAYER Metal1 ;
        RECT 24.160 2.720 24.320 2.790 ;
        RECT 24.030 2.430 24.320 2.720 ;
      LAYER Metal2 ;
        RECT 24.030 0.000 24.320 2.720 ;
    END
  END ONB[10]
  PIN ON[11]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 25.580 3.180 25.710 3.360 ;
        RECT 25.580 2.810 25.710 2.880 ;
        RECT 25.410 2.510 25.710 2.810 ;
      LAYER Metal1 ;
        RECT 25.480 2.720 25.640 2.790 ;
        RECT 25.480 2.430 25.770 2.720 ;
      LAYER Metal2 ;
        RECT 25.480 0.000 25.770 2.720 ;
    END
  END ON[11]
  PIN ONB[11]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 26.090 3.180 26.220 3.360 ;
        RECT 26.090 2.810 26.220 2.880 ;
        RECT 26.090 2.510 26.390 2.810 ;
      LAYER Metal1 ;
        RECT 26.160 2.720 26.320 2.790 ;
        RECT 26.030 2.430 26.320 2.720 ;
      LAYER Metal2 ;
        RECT 26.030 0.000 26.320 2.720 ;
    END
  END ONB[11]
  PIN ON[12]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 27.580 3.180 27.710 3.360 ;
        RECT 27.580 2.810 27.710 2.880 ;
        RECT 27.410 2.510 27.710 2.810 ;
      LAYER Metal1 ;
        RECT 27.480 2.720 27.640 2.790 ;
        RECT 27.480 2.430 27.770 2.720 ;
      LAYER Metal2 ;
        RECT 27.480 0.000 27.770 2.720 ;
    END
  END ON[12]
  PIN ONB[12]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 28.090 3.180 28.220 3.360 ;
        RECT 28.090 2.810 28.220 2.880 ;
        RECT 28.090 2.510 28.390 2.810 ;
      LAYER Metal1 ;
        RECT 28.160 2.720 28.320 2.790 ;
        RECT 28.030 2.430 28.320 2.720 ;
      LAYER Metal2 ;
        RECT 28.030 0.000 28.320 2.720 ;
    END
  END ONB[12]
  PIN ON[13]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 29.580 3.180 29.710 3.360 ;
        RECT 29.580 2.810 29.710 2.880 ;
        RECT 29.410 2.510 29.710 2.810 ;
      LAYER Metal1 ;
        RECT 29.480 2.720 29.640 2.790 ;
        RECT 29.480 2.430 29.770 2.720 ;
      LAYER Metal2 ;
        RECT 29.480 0.000 29.770 2.720 ;
    END
  END ON[13]
  PIN ONB[13]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 30.090 3.180 30.220 3.360 ;
        RECT 30.090 2.810 30.220 2.880 ;
        RECT 30.090 2.510 30.390 2.810 ;
      LAYER Metal1 ;
        RECT 30.160 2.720 30.320 2.790 ;
        RECT 30.030 2.430 30.320 2.720 ;
      LAYER Metal2 ;
        RECT 30.030 0.000 30.320 2.720 ;
    END
  END ONB[13]
  PIN ON[14]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 31.580 3.180 31.710 3.360 ;
        RECT 31.580 2.810 31.710 2.880 ;
        RECT 31.410 2.510 31.710 2.810 ;
      LAYER Metal1 ;
        RECT 31.480 2.720 31.640 2.790 ;
        RECT 31.480 2.430 31.770 2.720 ;
      LAYER Metal2 ;
        RECT 31.480 0.000 31.770 2.720 ;
    END
  END ON[14]
  PIN ONB[14]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 32.090 3.180 32.220 3.360 ;
        RECT 32.090 2.810 32.220 2.880 ;
        RECT 32.090 2.510 32.390 2.810 ;
      LAYER Metal1 ;
        RECT 32.160 2.720 32.320 2.790 ;
        RECT 32.030 2.430 32.320 2.720 ;
      LAYER Metal2 ;
        RECT 32.030 0.000 32.320 2.720 ;
    END
  END ONB[14]
  PIN ON[15]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 33.580 3.180 33.710 3.360 ;
        RECT 33.580 2.810 33.710 2.880 ;
        RECT 33.410 2.510 33.710 2.810 ;
      LAYER Metal1 ;
        RECT 33.480 2.720 33.640 2.790 ;
        RECT 33.480 2.430 33.770 2.720 ;
      LAYER Metal2 ;
        RECT 33.480 0.000 33.770 2.720 ;
    END
  END ON[15]
  PIN ONB[15]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 34.090 3.180 34.220 3.360 ;
        RECT 34.090 2.810 34.220 2.880 ;
        RECT 34.090 2.510 34.390 2.810 ;
      LAYER Metal1 ;
        RECT 34.160 2.720 34.320 2.790 ;
        RECT 34.030 2.430 34.320 2.720 ;
      LAYER Metal2 ;
        RECT 34.030 0.000 34.320 2.720 ;
    END
  END ONB[15]
  PIN ON[16]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 35.580 3.180 35.710 3.360 ;
        RECT 35.580 2.810 35.710 2.880 ;
        RECT 35.410 2.510 35.710 2.810 ;
      LAYER Metal1 ;
        RECT 35.480 2.720 35.640 2.790 ;
        RECT 35.480 2.430 35.770 2.720 ;
      LAYER Metal2 ;
        RECT 35.480 0.000 35.770 2.720 ;
    END
  END ON[16]
  PIN ONB[16]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 36.090 3.180 36.220 3.360 ;
        RECT 36.090 2.810 36.220 2.880 ;
        RECT 36.090 2.510 36.390 2.810 ;
      LAYER Metal1 ;
        RECT 36.160 2.720 36.320 2.790 ;
        RECT 36.030 2.430 36.320 2.720 ;
      LAYER Metal2 ;
        RECT 36.030 0.000 36.320 2.720 ;
    END
  END ONB[16]
  PIN ON[17]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 37.580 3.180 37.710 3.360 ;
        RECT 37.580 2.810 37.710 2.880 ;
        RECT 37.410 2.510 37.710 2.810 ;
      LAYER Metal1 ;
        RECT 37.480 2.720 37.640 2.790 ;
        RECT 37.480 2.430 37.770 2.720 ;
      LAYER Metal2 ;
        RECT 37.480 0.000 37.770 2.720 ;
    END
  END ON[17]
  PIN ONB[17]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 38.090 3.180 38.220 3.360 ;
        RECT 38.090 2.810 38.220 2.880 ;
        RECT 38.090 2.510 38.390 2.810 ;
      LAYER Metal1 ;
        RECT 38.160 2.720 38.320 2.790 ;
        RECT 38.030 2.430 38.320 2.720 ;
      LAYER Metal2 ;
        RECT 38.030 0.000 38.320 2.720 ;
    END
  END ONB[17]
  PIN ON[18]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 39.580 3.180 39.710 3.360 ;
        RECT 39.580 2.810 39.710 2.880 ;
        RECT 39.410 2.510 39.710 2.810 ;
      LAYER Metal1 ;
        RECT 39.480 2.720 39.640 2.790 ;
        RECT 39.480 2.430 39.770 2.720 ;
      LAYER Metal2 ;
        RECT 39.480 0.000 39.770 2.720 ;
    END
  END ON[18]
  PIN ONB[18]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 40.090 3.180 40.220 3.360 ;
        RECT 40.090 2.810 40.220 2.880 ;
        RECT 40.090 2.510 40.390 2.810 ;
      LAYER Metal1 ;
        RECT 40.160 2.720 40.320 2.790 ;
        RECT 40.030 2.430 40.320 2.720 ;
      LAYER Metal2 ;
        RECT 40.030 0.000 40.320 2.720 ;
    END
  END ONB[18]
  PIN ON[19]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 41.580 3.180 41.710 3.360 ;
        RECT 41.580 2.810 41.710 2.880 ;
        RECT 41.410 2.510 41.710 2.810 ;
      LAYER Metal1 ;
        RECT 41.480 2.720 41.640 2.790 ;
        RECT 41.480 2.430 41.770 2.720 ;
      LAYER Metal2 ;
        RECT 41.480 0.000 41.770 2.720 ;
    END
  END ON[19]
  PIN ONB[19]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 42.090 3.180 42.220 3.360 ;
        RECT 42.090 2.810 42.220 2.880 ;
        RECT 42.090 2.510 42.390 2.810 ;
      LAYER Metal1 ;
        RECT 42.160 2.720 42.320 2.790 ;
        RECT 42.030 2.430 42.320 2.720 ;
      LAYER Metal2 ;
        RECT 42.030 0.000 42.320 2.720 ;
    END
  END ONB[19]
  PIN ON[20]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 43.580 3.180 43.710 3.360 ;
        RECT 43.580 2.810 43.710 2.880 ;
        RECT 43.410 2.510 43.710 2.810 ;
      LAYER Metal1 ;
        RECT 43.480 2.720 43.640 2.790 ;
        RECT 43.480 2.430 43.770 2.720 ;
      LAYER Metal2 ;
        RECT 43.480 0.000 43.770 2.720 ;
    END
  END ON[20]
  PIN ONB[20]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 44.090 3.180 44.220 3.360 ;
        RECT 44.090 2.810 44.220 2.880 ;
        RECT 44.090 2.510 44.390 2.810 ;
      LAYER Metal1 ;
        RECT 44.160 2.720 44.320 2.790 ;
        RECT 44.030 2.430 44.320 2.720 ;
      LAYER Metal2 ;
        RECT 44.030 0.000 44.320 2.720 ;
    END
  END ONB[20]
  PIN ON[21]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 45.580 3.180 45.710 3.360 ;
        RECT 45.580 2.810 45.710 2.880 ;
        RECT 45.410 2.510 45.710 2.810 ;
      LAYER Metal1 ;
        RECT 45.480 2.720 45.640 2.790 ;
        RECT 45.480 2.430 45.770 2.720 ;
      LAYER Metal2 ;
        RECT 45.480 0.000 45.770 2.720 ;
    END
  END ON[21]
  PIN ONB[21]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 46.090 3.180 46.220 3.360 ;
        RECT 46.090 2.810 46.220 2.880 ;
        RECT 46.090 2.510 46.390 2.810 ;
      LAYER Metal1 ;
        RECT 46.160 2.720 46.320 2.790 ;
        RECT 46.030 2.430 46.320 2.720 ;
      LAYER Metal2 ;
        RECT 46.030 0.000 46.320 2.720 ;
    END
  END ONB[21]
  PIN ON[22]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 47.580 3.180 47.710 3.360 ;
        RECT 47.580 2.810 47.710 2.880 ;
        RECT 47.410 2.510 47.710 2.810 ;
      LAYER Metal1 ;
        RECT 47.480 2.720 47.640 2.790 ;
        RECT 47.480 2.430 47.770 2.720 ;
      LAYER Metal2 ;
        RECT 47.480 0.000 47.770 2.720 ;
    END
  END ON[22]
  PIN ONB[22]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 48.090 3.180 48.220 3.360 ;
        RECT 48.090 2.810 48.220 2.880 ;
        RECT 48.090 2.510 48.390 2.810 ;
      LAYER Metal1 ;
        RECT 48.160 2.720 48.320 2.790 ;
        RECT 48.030 2.430 48.320 2.720 ;
      LAYER Metal2 ;
        RECT 48.030 0.000 48.320 2.720 ;
    END
  END ONB[22]
  PIN ON[23]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 49.580 3.180 49.710 3.360 ;
        RECT 49.580 2.810 49.710 2.880 ;
        RECT 49.410 2.510 49.710 2.810 ;
      LAYER Metal1 ;
        RECT 49.480 2.720 49.640 2.790 ;
        RECT 49.480 2.430 49.770 2.720 ;
      LAYER Metal2 ;
        RECT 49.480 0.000 49.770 2.720 ;
    END
  END ON[23]
  PIN ONB[23]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 50.090 3.180 50.220 3.360 ;
        RECT 50.090 2.810 50.220 2.880 ;
        RECT 50.090 2.510 50.390 2.810 ;
      LAYER Metal1 ;
        RECT 50.160 2.720 50.320 2.790 ;
        RECT 50.030 2.430 50.320 2.720 ;
      LAYER Metal2 ;
        RECT 50.030 0.000 50.320 2.720 ;
    END
  END ONB[23]
  PIN ON[24]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 51.580 3.180 51.710 3.360 ;
        RECT 51.580 2.810 51.710 2.880 ;
        RECT 51.410 2.510 51.710 2.810 ;
      LAYER Metal1 ;
        RECT 51.480 2.720 51.640 2.790 ;
        RECT 51.480 2.430 51.770 2.720 ;
      LAYER Metal2 ;
        RECT 51.480 0.000 51.770 2.720 ;
    END
  END ON[24]
  PIN ONB[24]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 52.090 3.180 52.220 3.360 ;
        RECT 52.090 2.810 52.220 2.880 ;
        RECT 52.090 2.510 52.390 2.810 ;
      LAYER Metal1 ;
        RECT 52.160 2.720 52.320 2.790 ;
        RECT 52.030 2.430 52.320 2.720 ;
      LAYER Metal2 ;
        RECT 52.030 0.000 52.320 2.720 ;
    END
  END ONB[24]
  PIN ON[25]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 53.580 3.180 53.710 3.360 ;
        RECT 53.580 2.810 53.710 2.880 ;
        RECT 53.410 2.510 53.710 2.810 ;
      LAYER Metal1 ;
        RECT 53.480 2.720 53.640 2.790 ;
        RECT 53.480 2.430 53.770 2.720 ;
      LAYER Metal2 ;
        RECT 53.480 0.000 53.770 2.720 ;
    END
  END ON[25]
  PIN ONB[25]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 54.090 3.180 54.220 3.360 ;
        RECT 54.090 2.810 54.220 2.880 ;
        RECT 54.090 2.510 54.390 2.810 ;
      LAYER Metal1 ;
        RECT 54.160 2.720 54.320 2.790 ;
        RECT 54.030 2.430 54.320 2.720 ;
      LAYER Metal2 ;
        RECT 54.030 0.000 54.320 2.720 ;
    END
  END ONB[25]
  PIN ON[26]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 55.580 3.180 55.710 3.360 ;
        RECT 55.580 2.810 55.710 2.880 ;
        RECT 55.410 2.510 55.710 2.810 ;
      LAYER Metal1 ;
        RECT 55.480 2.720 55.640 2.790 ;
        RECT 55.480 2.430 55.770 2.720 ;
      LAYER Metal2 ;
        RECT 55.480 0.000 55.770 2.720 ;
    END
  END ON[26]
  PIN ONB[26]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 56.090 3.180 56.220 3.360 ;
        RECT 56.090 2.810 56.220 2.880 ;
        RECT 56.090 2.510 56.390 2.810 ;
      LAYER Metal1 ;
        RECT 56.160 2.720 56.320 2.790 ;
        RECT 56.030 2.430 56.320 2.720 ;
      LAYER Metal2 ;
        RECT 56.030 0.000 56.320 2.720 ;
    END
  END ONB[26]
  PIN ON[27]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 57.580 3.180 57.710 3.360 ;
        RECT 57.580 2.810 57.710 2.880 ;
        RECT 57.410 2.510 57.710 2.810 ;
      LAYER Metal1 ;
        RECT 57.480 2.720 57.640 2.790 ;
        RECT 57.480 2.430 57.770 2.720 ;
      LAYER Metal2 ;
        RECT 57.480 0.000 57.770 2.720 ;
    END
  END ON[27]
  PIN ONB[27]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 58.090 3.180 58.220 3.360 ;
        RECT 58.090 2.810 58.220 2.880 ;
        RECT 58.090 2.510 58.390 2.810 ;
      LAYER Metal1 ;
        RECT 58.160 2.720 58.320 2.790 ;
        RECT 58.030 2.430 58.320 2.720 ;
      LAYER Metal2 ;
        RECT 58.030 0.000 58.320 2.720 ;
    END
  END ONB[27]
  PIN ON[28]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 59.580 3.180 59.710 3.360 ;
        RECT 59.580 2.810 59.710 2.880 ;
        RECT 59.410 2.510 59.710 2.810 ;
      LAYER Metal1 ;
        RECT 59.480 2.720 59.640 2.790 ;
        RECT 59.480 2.430 59.770 2.720 ;
      LAYER Metal2 ;
        RECT 59.480 0.000 59.770 2.720 ;
    END
  END ON[28]
  PIN ONB[28]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 60.090 3.180 60.220 3.360 ;
        RECT 60.090 2.810 60.220 2.880 ;
        RECT 60.090 2.510 60.390 2.810 ;
      LAYER Metal1 ;
        RECT 60.160 2.720 60.320 2.790 ;
        RECT 60.030 2.430 60.320 2.720 ;
      LAYER Metal2 ;
        RECT 60.030 0.000 60.320 2.720 ;
    END
  END ONB[28]
  PIN ON[29]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 61.580 3.180 61.710 3.360 ;
        RECT 61.580 2.810 61.710 2.880 ;
        RECT 61.410 2.510 61.710 2.810 ;
      LAYER Metal1 ;
        RECT 61.480 2.720 61.640 2.790 ;
        RECT 61.480 2.430 61.770 2.720 ;
      LAYER Metal2 ;
        RECT 61.480 0.000 61.770 2.720 ;
    END
  END ON[29]
  PIN ONB[29]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 62.090 3.180 62.220 3.360 ;
        RECT 62.090 2.810 62.220 2.880 ;
        RECT 62.090 2.510 62.390 2.810 ;
      LAYER Metal1 ;
        RECT 62.160 2.720 62.320 2.790 ;
        RECT 62.030 2.430 62.320 2.720 ;
      LAYER Metal2 ;
        RECT 62.030 0.000 62.320 2.720 ;
    END
  END ONB[29]
  PIN ON[30]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 63.580 3.180 63.710 3.360 ;
        RECT 63.580 2.810 63.710 2.880 ;
        RECT 63.410 2.510 63.710 2.810 ;
      LAYER Metal1 ;
        RECT 63.480 2.720 63.640 2.790 ;
        RECT 63.480 2.430 63.770 2.720 ;
      LAYER Metal2 ;
        RECT 63.480 0.000 63.770 2.720 ;
    END
  END ON[30]
  PIN ONB[30]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 64.090 3.180 64.220 3.360 ;
        RECT 64.090 2.810 64.220 2.880 ;
        RECT 64.090 2.510 64.390 2.810 ;
      LAYER Metal1 ;
        RECT 64.160 2.720 64.320 2.790 ;
        RECT 64.030 2.430 64.320 2.720 ;
      LAYER Metal2 ;
        RECT 64.030 0.000 64.320 2.720 ;
    END
  END ONB[30]
  PIN ON[31]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 65.580 3.180 65.710 3.360 ;
        RECT 65.580 2.810 65.710 2.880 ;
        RECT 65.410 2.510 65.710 2.810 ;
      LAYER Metal1 ;
        RECT 65.480 2.720 65.640 2.790 ;
        RECT 65.480 2.430 65.770 2.720 ;
      LAYER Metal2 ;
        RECT 65.480 0.000 65.770 2.720 ;
    END
  END ON[31]
  PIN ONB[31]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 66.090 3.180 66.220 3.360 ;
        RECT 66.090 2.810 66.220 2.880 ;
        RECT 66.090 2.510 66.390 2.810 ;
      LAYER Metal1 ;
        RECT 66.160 2.720 66.320 2.790 ;
        RECT 66.030 2.430 66.320 2.720 ;
      LAYER Metal2 ;
        RECT 66.030 0.000 66.320 2.720 ;
    END
  END ONB[31]
  PIN EN[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 1.580 3.180 1.710 3.360 ;
        RECT 1.580 2.810 1.710 2.880 ;
        RECT 1.410 2.510 1.710 2.810 ;
      LAYER Metal1 ;
        RECT 1.480 2.720 1.640 2.790 ;
        RECT 1.480 2.430 1.770 2.720 ;
      LAYER Metal2 ;
        RECT 1.480 0.000 1.770 2.720 ;
    END
  END EN[0]
  PIN ENB[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 2.090 3.180 2.220 3.360 ;
        RECT 2.090 2.810 2.220 2.880 ;
        RECT 2.090 2.510 2.390 2.810 ;
      LAYER Metal1 ;
        RECT 2.160 2.720 2.320 2.790 ;
        RECT 2.030 2.430 2.320 2.720 ;
      LAYER Metal2 ;
        RECT 2.030 0.000 2.320 2.720 ;
    END
  END ENB[0]
  PIN ON[33]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 69.580 3.180 69.710 3.360 ;
        RECT 69.580 2.810 69.710 2.880 ;
        RECT 69.410 2.510 69.710 2.810 ;
      LAYER Metal1 ;
        RECT 69.480 2.720 69.640 2.790 ;
        RECT 69.480 2.430 69.770 2.720 ;
      LAYER Metal2 ;
        RECT 69.480 0.000 69.770 2.720 ;
    END
  END ON[33]
  PIN ONB[33]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 70.090 3.180 70.220 3.360 ;
        RECT 70.090 2.810 70.220 2.880 ;
        RECT 70.090 2.510 70.390 2.810 ;
      LAYER Metal1 ;
        RECT 70.160 2.720 70.320 2.790 ;
        RECT 70.030 2.430 70.320 2.720 ;
      LAYER Metal2 ;
        RECT 70.030 0.000 70.320 2.720 ;
    END
  END ONB[33]
  PIN ON[34]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 71.580 3.180 71.710 3.360 ;
        RECT 71.580 2.810 71.710 2.880 ;
        RECT 71.410 2.510 71.710 2.810 ;
      LAYER Metal1 ;
        RECT 71.480 2.720 71.640 2.790 ;
        RECT 71.480 2.430 71.770 2.720 ;
      LAYER Metal2 ;
        RECT 71.480 0.000 71.770 2.720 ;
    END
  END ON[34]
  PIN ONB[34]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 72.090 3.180 72.220 3.360 ;
        RECT 72.090 2.810 72.220 2.880 ;
        RECT 72.090 2.510 72.390 2.810 ;
      LAYER Metal1 ;
        RECT 72.160 2.720 72.320 2.790 ;
        RECT 72.030 2.430 72.320 2.720 ;
      LAYER Metal2 ;
        RECT 72.030 0.000 72.320 2.720 ;
    END
  END ONB[34]
  PIN ON[35]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 73.580 3.180 73.710 3.360 ;
        RECT 73.580 2.810 73.710 2.880 ;
        RECT 73.410 2.510 73.710 2.810 ;
      LAYER Metal1 ;
        RECT 73.480 2.720 73.640 2.790 ;
        RECT 73.480 2.430 73.770 2.720 ;
      LAYER Metal2 ;
        RECT 73.480 0.000 73.770 2.720 ;
    END
  END ON[35]
  PIN ONB[35]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 74.090 3.180 74.220 3.360 ;
        RECT 74.090 2.810 74.220 2.880 ;
        RECT 74.090 2.510 74.390 2.810 ;
      LAYER Metal1 ;
        RECT 74.160 2.720 74.320 2.790 ;
        RECT 74.030 2.430 74.320 2.720 ;
      LAYER Metal2 ;
        RECT 74.030 0.000 74.320 2.720 ;
    END
  END ONB[35]
  PIN ON[36]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 75.580 3.180 75.710 3.360 ;
        RECT 75.580 2.810 75.710 2.880 ;
        RECT 75.410 2.510 75.710 2.810 ;
      LAYER Metal1 ;
        RECT 75.480 2.720 75.640 2.790 ;
        RECT 75.480 2.430 75.770 2.720 ;
      LAYER Metal2 ;
        RECT 75.480 0.000 75.770 2.720 ;
    END
  END ON[36]
  PIN ONB[36]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 76.090 3.180 76.220 3.360 ;
        RECT 76.090 2.810 76.220 2.880 ;
        RECT 76.090 2.510 76.390 2.810 ;
      LAYER Metal1 ;
        RECT 76.160 2.720 76.320 2.790 ;
        RECT 76.030 2.430 76.320 2.720 ;
      LAYER Metal2 ;
        RECT 76.030 0.000 76.320 2.720 ;
    END
  END ONB[36]
  PIN ON[37]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 77.580 3.180 77.710 3.360 ;
        RECT 77.580 2.810 77.710 2.880 ;
        RECT 77.410 2.510 77.710 2.810 ;
      LAYER Metal1 ;
        RECT 77.480 2.720 77.640 2.790 ;
        RECT 77.480 2.430 77.770 2.720 ;
      LAYER Metal2 ;
        RECT 77.480 0.000 77.770 2.720 ;
    END
  END ON[37]
  PIN ONB[37]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 78.090 3.180 78.220 3.360 ;
        RECT 78.090 2.810 78.220 2.880 ;
        RECT 78.090 2.510 78.390 2.810 ;
      LAYER Metal1 ;
        RECT 78.160 2.720 78.320 2.790 ;
        RECT 78.030 2.430 78.320 2.720 ;
      LAYER Metal2 ;
        RECT 78.030 0.000 78.320 2.720 ;
    END
  END ONB[37]
  PIN ON[38]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 79.580 3.180 79.710 3.360 ;
        RECT 79.580 2.810 79.710 2.880 ;
        RECT 79.410 2.510 79.710 2.810 ;
      LAYER Metal1 ;
        RECT 79.480 2.720 79.640 2.790 ;
        RECT 79.480 2.430 79.770 2.720 ;
      LAYER Metal2 ;
        RECT 79.480 0.000 79.770 2.720 ;
    END
  END ON[38]
  PIN ONB[38]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 80.090 3.180 80.220 3.360 ;
        RECT 80.090 2.810 80.220 2.880 ;
        RECT 80.090 2.510 80.390 2.810 ;
      LAYER Metal1 ;
        RECT 80.160 2.720 80.320 2.790 ;
        RECT 80.030 2.430 80.320 2.720 ;
      LAYER Metal2 ;
        RECT 80.030 0.000 80.320 2.720 ;
    END
  END ONB[38]
  PIN ON[39]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 81.580 3.180 81.710 3.360 ;
        RECT 81.580 2.810 81.710 2.880 ;
        RECT 81.410 2.510 81.710 2.810 ;
      LAYER Metal1 ;
        RECT 81.480 2.720 81.640 2.790 ;
        RECT 81.480 2.430 81.770 2.720 ;
      LAYER Metal2 ;
        RECT 81.480 0.000 81.770 2.720 ;
    END
  END ON[39]
  PIN ONB[39]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 82.090 3.180 82.220 3.360 ;
        RECT 82.090 2.810 82.220 2.880 ;
        RECT 82.090 2.510 82.390 2.810 ;
      LAYER Metal1 ;
        RECT 82.160 2.720 82.320 2.790 ;
        RECT 82.030 2.430 82.320 2.720 ;
      LAYER Metal2 ;
        RECT 82.030 0.000 82.320 2.720 ;
    END
  END ONB[39]
  PIN ON[40]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 83.580 3.180 83.710 3.360 ;
        RECT 83.580 2.810 83.710 2.880 ;
        RECT 83.410 2.510 83.710 2.810 ;
      LAYER Metal1 ;
        RECT 83.480 2.720 83.640 2.790 ;
        RECT 83.480 2.430 83.770 2.720 ;
      LAYER Metal2 ;
        RECT 83.480 0.000 83.770 2.720 ;
    END
  END ON[40]
  PIN ONB[40]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 84.090 3.180 84.220 3.360 ;
        RECT 84.090 2.810 84.220 2.880 ;
        RECT 84.090 2.510 84.390 2.810 ;
      LAYER Metal1 ;
        RECT 84.160 2.720 84.320 2.790 ;
        RECT 84.030 2.430 84.320 2.720 ;
      LAYER Metal2 ;
        RECT 84.030 0.000 84.320 2.720 ;
    END
  END ONB[40]
  PIN ON[41]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 85.580 3.180 85.710 3.360 ;
        RECT 85.580 2.810 85.710 2.880 ;
        RECT 85.410 2.510 85.710 2.810 ;
      LAYER Metal1 ;
        RECT 85.480 2.720 85.640 2.790 ;
        RECT 85.480 2.430 85.770 2.720 ;
      LAYER Metal2 ;
        RECT 85.480 0.000 85.770 2.720 ;
    END
  END ON[41]
  PIN ONB[41]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 86.090 3.180 86.220 3.360 ;
        RECT 86.090 2.810 86.220 2.880 ;
        RECT 86.090 2.510 86.390 2.810 ;
      LAYER Metal1 ;
        RECT 86.160 2.720 86.320 2.790 ;
        RECT 86.030 2.430 86.320 2.720 ;
      LAYER Metal2 ;
        RECT 86.030 0.000 86.320 2.720 ;
    END
  END ONB[41]
  PIN ON[42]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 87.580 3.180 87.710 3.360 ;
        RECT 87.580 2.810 87.710 2.880 ;
        RECT 87.410 2.510 87.710 2.810 ;
      LAYER Metal1 ;
        RECT 87.480 2.720 87.640 2.790 ;
        RECT 87.480 2.430 87.770 2.720 ;
      LAYER Metal2 ;
        RECT 87.480 0.000 87.770 2.720 ;
    END
  END ON[42]
  PIN ONB[42]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 88.090 3.180 88.220 3.360 ;
        RECT 88.090 2.810 88.220 2.880 ;
        RECT 88.090 2.510 88.390 2.810 ;
      LAYER Metal1 ;
        RECT 88.160 2.720 88.320 2.790 ;
        RECT 88.030 2.430 88.320 2.720 ;
      LAYER Metal2 ;
        RECT 88.030 0.000 88.320 2.720 ;
    END
  END ONB[42]
  PIN ON[43]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 89.580 3.180 89.710 3.360 ;
        RECT 89.580 2.810 89.710 2.880 ;
        RECT 89.410 2.510 89.710 2.810 ;
      LAYER Metal1 ;
        RECT 89.480 2.720 89.640 2.790 ;
        RECT 89.480 2.430 89.770 2.720 ;
      LAYER Metal2 ;
        RECT 89.480 0.000 89.770 2.720 ;
    END
  END ON[43]
  PIN ONB[43]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 90.090 3.180 90.220 3.360 ;
        RECT 90.090 2.810 90.220 2.880 ;
        RECT 90.090 2.510 90.390 2.810 ;
      LAYER Metal1 ;
        RECT 90.160 2.720 90.320 2.790 ;
        RECT 90.030 2.430 90.320 2.720 ;
      LAYER Metal2 ;
        RECT 90.030 0.000 90.320 2.720 ;
    END
  END ONB[43]
  PIN ON[44]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 91.580 3.180 91.710 3.360 ;
        RECT 91.580 2.810 91.710 2.880 ;
        RECT 91.410 2.510 91.710 2.810 ;
      LAYER Metal1 ;
        RECT 91.480 2.720 91.640 2.790 ;
        RECT 91.480 2.430 91.770 2.720 ;
      LAYER Metal2 ;
        RECT 91.480 0.000 91.770 2.720 ;
    END
  END ON[44]
  PIN ONB[44]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 92.090 3.180 92.220 3.360 ;
        RECT 92.090 2.810 92.220 2.880 ;
        RECT 92.090 2.510 92.390 2.810 ;
      LAYER Metal1 ;
        RECT 92.160 2.720 92.320 2.790 ;
        RECT 92.030 2.430 92.320 2.720 ;
      LAYER Metal2 ;
        RECT 92.030 0.000 92.320 2.720 ;
    END
  END ONB[44]
  PIN ON[45]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 93.580 3.180 93.710 3.360 ;
        RECT 93.580 2.810 93.710 2.880 ;
        RECT 93.410 2.510 93.710 2.810 ;
      LAYER Metal1 ;
        RECT 93.480 2.720 93.640 2.790 ;
        RECT 93.480 2.430 93.770 2.720 ;
      LAYER Metal2 ;
        RECT 93.480 0.000 93.770 2.720 ;
    END
  END ON[45]
  PIN ONB[45]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 94.090 3.180 94.220 3.360 ;
        RECT 94.090 2.810 94.220 2.880 ;
        RECT 94.090 2.510 94.390 2.810 ;
      LAYER Metal1 ;
        RECT 94.160 2.720 94.320 2.790 ;
        RECT 94.030 2.430 94.320 2.720 ;
      LAYER Metal2 ;
        RECT 94.030 0.000 94.320 2.720 ;
    END
  END ONB[45]
  PIN ON[46]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 95.580 3.180 95.710 3.360 ;
        RECT 95.580 2.810 95.710 2.880 ;
        RECT 95.410 2.510 95.710 2.810 ;
      LAYER Metal1 ;
        RECT 95.480 2.720 95.640 2.790 ;
        RECT 95.480 2.430 95.770 2.720 ;
      LAYER Metal2 ;
        RECT 95.480 0.000 95.770 2.720 ;
    END
  END ON[46]
  PIN ONB[46]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 96.090 3.180 96.220 3.360 ;
        RECT 96.090 2.810 96.220 2.880 ;
        RECT 96.090 2.510 96.390 2.810 ;
      LAYER Metal1 ;
        RECT 96.160 2.720 96.320 2.790 ;
        RECT 96.030 2.430 96.320 2.720 ;
      LAYER Metal2 ;
        RECT 96.030 0.000 96.320 2.720 ;
    END
  END ONB[46]
  PIN ON[47]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 97.580 3.180 97.710 3.360 ;
        RECT 97.580 2.810 97.710 2.880 ;
        RECT 97.410 2.510 97.710 2.810 ;
      LAYER Metal1 ;
        RECT 97.480 2.720 97.640 2.790 ;
        RECT 97.480 2.430 97.770 2.720 ;
      LAYER Metal2 ;
        RECT 97.480 0.000 97.770 2.720 ;
    END
  END ON[47]
  PIN ONB[47]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 98.090 3.180 98.220 3.360 ;
        RECT 98.090 2.810 98.220 2.880 ;
        RECT 98.090 2.510 98.390 2.810 ;
      LAYER Metal1 ;
        RECT 98.160 2.720 98.320 2.790 ;
        RECT 98.030 2.430 98.320 2.720 ;
      LAYER Metal2 ;
        RECT 98.030 0.000 98.320 2.720 ;
    END
  END ONB[47]
  PIN ON[48]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 99.580 3.180 99.710 3.360 ;
        RECT 99.580 2.810 99.710 2.880 ;
        RECT 99.410 2.510 99.710 2.810 ;
      LAYER Metal1 ;
        RECT 99.480 2.720 99.640 2.790 ;
        RECT 99.480 2.430 99.770 2.720 ;
      LAYER Metal2 ;
        RECT 99.480 0.000 99.770 2.720 ;
    END
  END ON[48]
  PIN ONB[48]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 100.090 3.180 100.220 3.360 ;
        RECT 100.090 2.810 100.220 2.880 ;
        RECT 100.090 2.510 100.390 2.810 ;
      LAYER Metal1 ;
        RECT 100.160 2.720 100.320 2.790 ;
        RECT 100.030 2.430 100.320 2.720 ;
      LAYER Metal2 ;
        RECT 100.030 0.000 100.320 2.720 ;
    END
  END ONB[48]
  PIN ON[49]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 101.580 3.180 101.710 3.360 ;
        RECT 101.580 2.810 101.710 2.880 ;
        RECT 101.410 2.510 101.710 2.810 ;
      LAYER Metal1 ;
        RECT 101.480 2.720 101.640 2.790 ;
        RECT 101.480 2.430 101.770 2.720 ;
      LAYER Metal2 ;
        RECT 101.480 0.000 101.770 2.720 ;
    END
  END ON[49]
  PIN ONB[49]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 102.090 3.180 102.220 3.360 ;
        RECT 102.090 2.810 102.220 2.880 ;
        RECT 102.090 2.510 102.390 2.810 ;
      LAYER Metal1 ;
        RECT 102.160 2.720 102.320 2.790 ;
        RECT 102.030 2.430 102.320 2.720 ;
      LAYER Metal2 ;
        RECT 102.030 0.000 102.320 2.720 ;
    END
  END ONB[49]
  PIN ON[50]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 103.580 3.180 103.710 3.360 ;
        RECT 103.580 2.810 103.710 2.880 ;
        RECT 103.410 2.510 103.710 2.810 ;
      LAYER Metal1 ;
        RECT 103.480 2.720 103.640 2.790 ;
        RECT 103.480 2.430 103.770 2.720 ;
      LAYER Metal2 ;
        RECT 103.480 0.000 103.770 2.720 ;
    END
  END ON[50]
  PIN ONB[50]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 104.090 3.180 104.220 3.360 ;
        RECT 104.090 2.810 104.220 2.880 ;
        RECT 104.090 2.510 104.390 2.810 ;
      LAYER Metal1 ;
        RECT 104.160 2.720 104.320 2.790 ;
        RECT 104.030 2.430 104.320 2.720 ;
      LAYER Metal2 ;
        RECT 104.030 0.000 104.320 2.720 ;
    END
  END ONB[50]
  PIN ON[51]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 105.580 3.180 105.710 3.360 ;
        RECT 105.580 2.810 105.710 2.880 ;
        RECT 105.410 2.510 105.710 2.810 ;
      LAYER Metal1 ;
        RECT 105.480 2.720 105.640 2.790 ;
        RECT 105.480 2.430 105.770 2.720 ;
      LAYER Metal2 ;
        RECT 105.480 0.000 105.770 2.720 ;
    END
  END ON[51]
  PIN ONB[51]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 106.090 3.180 106.220 3.360 ;
        RECT 106.090 2.810 106.220 2.880 ;
        RECT 106.090 2.510 106.390 2.810 ;
      LAYER Metal1 ;
        RECT 106.160 2.720 106.320 2.790 ;
        RECT 106.030 2.430 106.320 2.720 ;
      LAYER Metal2 ;
        RECT 106.030 0.000 106.320 2.720 ;
    END
  END ONB[51]
  PIN ON[52]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 107.580 3.180 107.710 3.360 ;
        RECT 107.580 2.810 107.710 2.880 ;
        RECT 107.410 2.510 107.710 2.810 ;
      LAYER Metal1 ;
        RECT 107.480 2.720 107.640 2.790 ;
        RECT 107.480 2.430 107.770 2.720 ;
      LAYER Metal2 ;
        RECT 107.480 0.000 107.770 2.720 ;
    END
  END ON[52]
  PIN ONB[52]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 108.090 3.180 108.220 3.360 ;
        RECT 108.090 2.810 108.220 2.880 ;
        RECT 108.090 2.510 108.390 2.810 ;
      LAYER Metal1 ;
        RECT 108.160 2.720 108.320 2.790 ;
        RECT 108.030 2.430 108.320 2.720 ;
      LAYER Metal2 ;
        RECT 108.030 0.000 108.320 2.720 ;
    END
  END ONB[52]
  PIN ON[53]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 109.580 3.180 109.710 3.360 ;
        RECT 109.580 2.810 109.710 2.880 ;
        RECT 109.410 2.510 109.710 2.810 ;
      LAYER Metal1 ;
        RECT 109.480 2.720 109.640 2.790 ;
        RECT 109.480 2.430 109.770 2.720 ;
      LAYER Metal2 ;
        RECT 109.480 0.000 109.770 2.720 ;
    END
  END ON[53]
  PIN ONB[53]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 110.090 3.180 110.220 3.360 ;
        RECT 110.090 2.810 110.220 2.880 ;
        RECT 110.090 2.510 110.390 2.810 ;
      LAYER Metal1 ;
        RECT 110.160 2.720 110.320 2.790 ;
        RECT 110.030 2.430 110.320 2.720 ;
      LAYER Metal2 ;
        RECT 110.030 0.000 110.320 2.720 ;
    END
  END ONB[53]
  PIN ON[54]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 111.580 3.180 111.710 3.360 ;
        RECT 111.580 2.810 111.710 2.880 ;
        RECT 111.410 2.510 111.710 2.810 ;
      LAYER Metal1 ;
        RECT 111.480 2.720 111.640 2.790 ;
        RECT 111.480 2.430 111.770 2.720 ;
      LAYER Metal2 ;
        RECT 111.480 0.000 111.770 2.720 ;
    END
  END ON[54]
  PIN ONB[54]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 112.090 3.180 112.220 3.360 ;
        RECT 112.090 2.810 112.220 2.880 ;
        RECT 112.090 2.510 112.390 2.810 ;
      LAYER Metal1 ;
        RECT 112.160 2.720 112.320 2.790 ;
        RECT 112.030 2.430 112.320 2.720 ;
      LAYER Metal2 ;
        RECT 112.030 0.000 112.320 2.720 ;
    END
  END ONB[54]
  PIN ON[55]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 113.580 3.180 113.710 3.360 ;
        RECT 113.580 2.810 113.710 2.880 ;
        RECT 113.410 2.510 113.710 2.810 ;
      LAYER Metal1 ;
        RECT 113.480 2.720 113.640 2.790 ;
        RECT 113.480 2.430 113.770 2.720 ;
      LAYER Metal2 ;
        RECT 113.480 0.000 113.770 2.720 ;
    END
  END ON[55]
  PIN ONB[55]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 114.090 3.180 114.220 3.360 ;
        RECT 114.090 2.810 114.220 2.880 ;
        RECT 114.090 2.510 114.390 2.810 ;
      LAYER Metal1 ;
        RECT 114.160 2.720 114.320 2.790 ;
        RECT 114.030 2.430 114.320 2.720 ;
      LAYER Metal2 ;
        RECT 114.030 0.000 114.320 2.720 ;
    END
  END ONB[55]
  PIN ON[56]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 115.580 3.180 115.710 3.360 ;
        RECT 115.580 2.810 115.710 2.880 ;
        RECT 115.410 2.510 115.710 2.810 ;
      LAYER Metal1 ;
        RECT 115.480 2.720 115.640 2.790 ;
        RECT 115.480 2.430 115.770 2.720 ;
      LAYER Metal2 ;
        RECT 115.480 0.000 115.770 2.720 ;
    END
  END ON[56]
  PIN ONB[56]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 116.090 3.180 116.220 3.360 ;
        RECT 116.090 2.810 116.220 2.880 ;
        RECT 116.090 2.510 116.390 2.810 ;
      LAYER Metal1 ;
        RECT 116.160 2.720 116.320 2.790 ;
        RECT 116.030 2.430 116.320 2.720 ;
      LAYER Metal2 ;
        RECT 116.030 0.000 116.320 2.720 ;
    END
  END ONB[56]
  PIN ON[57]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 117.580 3.180 117.710 3.360 ;
        RECT 117.580 2.810 117.710 2.880 ;
        RECT 117.410 2.510 117.710 2.810 ;
      LAYER Metal1 ;
        RECT 117.480 2.720 117.640 2.790 ;
        RECT 117.480 2.430 117.770 2.720 ;
      LAYER Metal2 ;
        RECT 117.480 0.000 117.770 2.720 ;
    END
  END ON[57]
  PIN ONB[57]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 118.090 3.180 118.220 3.360 ;
        RECT 118.090 2.810 118.220 2.880 ;
        RECT 118.090 2.510 118.390 2.810 ;
      LAYER Metal1 ;
        RECT 118.160 2.720 118.320 2.790 ;
        RECT 118.030 2.430 118.320 2.720 ;
      LAYER Metal2 ;
        RECT 118.030 0.000 118.320 2.720 ;
    END
  END ONB[57]
  PIN ON[58]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 119.580 3.180 119.710 3.360 ;
        RECT 119.580 2.810 119.710 2.880 ;
        RECT 119.410 2.510 119.710 2.810 ;
      LAYER Metal1 ;
        RECT 119.480 2.720 119.640 2.790 ;
        RECT 119.480 2.430 119.770 2.720 ;
      LAYER Metal2 ;
        RECT 119.480 0.000 119.770 2.720 ;
    END
  END ON[58]
  PIN ONB[58]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 120.090 3.180 120.220 3.360 ;
        RECT 120.090 2.810 120.220 2.880 ;
        RECT 120.090 2.510 120.390 2.810 ;
      LAYER Metal1 ;
        RECT 120.160 2.720 120.320 2.790 ;
        RECT 120.030 2.430 120.320 2.720 ;
      LAYER Metal2 ;
        RECT 120.030 0.000 120.320 2.720 ;
    END
  END ONB[58]
  PIN ON[59]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 121.580 3.180 121.710 3.360 ;
        RECT 121.580 2.810 121.710 2.880 ;
        RECT 121.410 2.510 121.710 2.810 ;
      LAYER Metal1 ;
        RECT 121.480 2.720 121.640 2.790 ;
        RECT 121.480 2.430 121.770 2.720 ;
      LAYER Metal2 ;
        RECT 121.480 0.000 121.770 2.720 ;
    END
  END ON[59]
  PIN ONB[59]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 122.090 3.180 122.220 3.360 ;
        RECT 122.090 2.810 122.220 2.880 ;
        RECT 122.090 2.510 122.390 2.810 ;
      LAYER Metal1 ;
        RECT 122.160 2.720 122.320 2.790 ;
        RECT 122.030 2.430 122.320 2.720 ;
      LAYER Metal2 ;
        RECT 122.030 0.000 122.320 2.720 ;
    END
  END ONB[59]
  PIN ON[60]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 123.580 3.180 123.710 3.360 ;
        RECT 123.580 2.810 123.710 2.880 ;
        RECT 123.410 2.510 123.710 2.810 ;
      LAYER Metal1 ;
        RECT 123.480 2.720 123.640 2.790 ;
        RECT 123.480 2.430 123.770 2.720 ;
      LAYER Metal2 ;
        RECT 123.480 0.000 123.770 2.720 ;
    END
  END ON[60]
  PIN ONB[60]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 124.090 3.180 124.220 3.360 ;
        RECT 124.090 2.810 124.220 2.880 ;
        RECT 124.090 2.510 124.390 2.810 ;
      LAYER Metal1 ;
        RECT 124.160 2.720 124.320 2.790 ;
        RECT 124.030 2.430 124.320 2.720 ;
      LAYER Metal2 ;
        RECT 124.030 0.000 124.320 2.720 ;
    END
  END ONB[60]
  PIN ON[61]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 125.580 3.180 125.710 3.360 ;
        RECT 125.580 2.810 125.710 2.880 ;
        RECT 125.410 2.510 125.710 2.810 ;
      LAYER Metal1 ;
        RECT 125.480 2.720 125.640 2.790 ;
        RECT 125.480 2.430 125.770 2.720 ;
      LAYER Metal2 ;
        RECT 125.480 0.000 125.770 2.720 ;
    END
  END ON[61]
  PIN ONB[61]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 126.090 3.180 126.220 3.360 ;
        RECT 126.090 2.810 126.220 2.880 ;
        RECT 126.090 2.510 126.390 2.810 ;
      LAYER Metal1 ;
        RECT 126.160 2.720 126.320 2.790 ;
        RECT 126.030 2.430 126.320 2.720 ;
      LAYER Metal2 ;
        RECT 126.030 0.000 126.320 2.720 ;
    END
  END ONB[61]
  PIN ON[62]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 127.580 3.180 127.710 3.360 ;
        RECT 127.580 2.810 127.710 2.880 ;
        RECT 127.410 2.510 127.710 2.810 ;
      LAYER Metal1 ;
        RECT 127.480 2.720 127.640 2.790 ;
        RECT 127.480 2.430 127.770 2.720 ;
      LAYER Metal2 ;
        RECT 127.480 0.000 127.770 2.720 ;
    END
  END ON[62]
  PIN ONB[62]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 128.090 3.180 128.220 3.360 ;
        RECT 128.090 2.810 128.220 2.880 ;
        RECT 128.090 2.510 128.390 2.810 ;
      LAYER Metal1 ;
        RECT 128.160 2.720 128.320 2.790 ;
        RECT 128.030 2.430 128.320 2.720 ;
      LAYER Metal2 ;
        RECT 128.030 0.000 128.320 2.720 ;
    END
  END ONB[62]
  PIN ON[63]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 129.580 3.180 129.710 3.360 ;
        RECT 129.580 2.810 129.710 2.880 ;
        RECT 129.410 2.510 129.710 2.810 ;
      LAYER Metal1 ;
        RECT 129.480 2.720 129.640 2.790 ;
        RECT 129.480 2.430 129.770 2.720 ;
      LAYER Metal2 ;
        RECT 129.480 0.000 129.770 2.720 ;
    END
  END ON[63]
  PIN ONB[63]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 130.090 3.180 130.220 3.360 ;
        RECT 130.090 2.810 130.220 2.880 ;
        RECT 130.090 2.510 130.390 2.810 ;
      LAYER Metal1 ;
        RECT 130.160 2.720 130.320 2.790 ;
        RECT 130.030 2.430 130.320 2.720 ;
      LAYER Metal2 ;
        RECT 130.030 0.000 130.320 2.720 ;
    END
  END ONB[63]
  PIN ON[32]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 67.580 3.180 67.710 3.360 ;
        RECT 67.580 2.810 67.710 2.880 ;
        RECT 67.410 2.510 67.710 2.810 ;
      LAYER Metal1 ;
        RECT 67.480 2.720 67.640 2.790 ;
        RECT 67.480 2.430 67.770 2.720 ;
      LAYER Metal2 ;
        RECT 67.480 0.000 67.770 2.720 ;
    END
  END ON[32]
  PIN ONB[32]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 68.090 3.180 68.220 3.360 ;
        RECT 68.090 2.810 68.220 2.880 ;
        RECT 68.090 2.510 68.390 2.810 ;
      LAYER Metal1 ;
        RECT 68.160 2.720 68.320 2.790 ;
        RECT 68.030 2.430 68.320 2.720 ;
      LAYER Metal2 ;
        RECT 68.030 0.000 68.320 2.720 ;
    END
  END ONB[32]
  PIN EN[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 131.580 3.180 131.710 3.360 ;
        RECT 131.580 2.810 131.710 2.880 ;
        RECT 131.410 2.510 131.710 2.810 ;
      LAYER Metal1 ;
        RECT 131.480 2.720 131.640 2.790 ;
        RECT 131.480 2.430 131.770 2.720 ;
      LAYER Metal2 ;
        RECT 131.480 0.000 131.770 2.720 ;
    END
  END EN[1]
  PIN ENB[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER GatPoly ;
        RECT 132.090 3.180 132.220 3.360 ;
        RECT 132.090 2.810 132.220 2.880 ;
        RECT 132.090 2.510 132.390 2.810 ;
      LAYER Metal1 ;
        RECT 132.160 2.720 132.320 2.790 ;
        RECT 132.030 2.430 132.320 2.720 ;
      LAYER Metal2 ;
        RECT 132.030 0.000 132.320 2.720 ;
    END
  END ENB[1]
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 1.820 0.500 1.980 1.060 ;
        RECT 3.820 0.500 3.980 1.060 ;
        RECT 5.820 0.500 5.980 1.060 ;
        RECT 7.820 0.500 7.980 1.060 ;
        RECT 9.820 0.500 9.980 1.060 ;
        RECT 11.820 0.500 11.980 1.060 ;
        RECT 13.820 0.500 13.980 1.060 ;
        RECT 15.820 0.500 15.980 1.060 ;
        RECT 17.820 0.500 17.980 1.060 ;
        RECT 19.820 0.500 19.980 1.060 ;
        RECT 21.820 0.500 21.980 1.060 ;
        RECT 23.820 0.500 23.980 1.060 ;
        RECT 25.820 0.500 25.980 1.060 ;
        RECT 27.820 0.500 27.980 1.060 ;
        RECT 29.820 0.500 29.980 1.060 ;
        RECT 31.820 0.500 31.980 1.060 ;
        RECT 33.820 0.500 33.980 1.060 ;
        RECT 35.820 0.500 35.980 1.060 ;
        RECT 37.820 0.500 37.980 1.060 ;
        RECT 39.820 0.500 39.980 1.060 ;
        RECT 41.820 0.500 41.980 1.060 ;
        RECT 43.820 0.500 43.980 1.060 ;
        RECT 45.820 0.500 45.980 1.060 ;
        RECT 47.820 0.500 47.980 1.060 ;
        RECT 49.820 0.500 49.980 1.060 ;
        RECT 51.820 0.500 51.980 1.060 ;
        RECT 53.820 0.500 53.980 1.060 ;
        RECT 55.820 0.500 55.980 1.060 ;
        RECT 57.820 0.500 57.980 1.060 ;
        RECT 59.820 0.500 59.980 1.060 ;
        RECT 61.820 0.500 61.980 1.060 ;
        RECT 63.820 0.500 63.980 1.060 ;
        RECT 65.820 0.500 65.980 1.060 ;
        RECT 67.820 0.500 67.980 1.060 ;
        RECT 69.820 0.500 69.980 1.060 ;
        RECT 71.820 0.500 71.980 1.060 ;
        RECT 73.820 0.500 73.980 1.060 ;
        RECT 75.820 0.500 75.980 1.060 ;
        RECT 77.820 0.500 77.980 1.060 ;
        RECT 79.820 0.500 79.980 1.060 ;
        RECT 81.820 0.500 81.980 1.060 ;
        RECT 83.820 0.500 83.980 1.060 ;
        RECT 85.820 0.500 85.980 1.060 ;
        RECT 87.820 0.500 87.980 1.060 ;
        RECT 89.820 0.500 89.980 1.060 ;
        RECT 91.820 0.500 91.980 1.060 ;
        RECT 93.820 0.500 93.980 1.060 ;
        RECT 95.820 0.500 95.980 1.060 ;
        RECT 97.820 0.500 97.980 1.060 ;
        RECT 99.820 0.500 99.980 1.060 ;
        RECT 101.820 0.500 101.980 1.060 ;
        RECT 103.820 0.500 103.980 1.060 ;
        RECT 105.820 0.500 105.980 1.060 ;
        RECT 107.820 0.500 107.980 1.060 ;
        RECT 109.820 0.500 109.980 1.060 ;
        RECT 111.820 0.500 111.980 1.060 ;
        RECT 113.820 0.500 113.980 1.060 ;
        RECT 115.820 0.500 115.980 1.060 ;
        RECT 117.820 0.500 117.980 1.060 ;
        RECT 119.820 0.500 119.980 1.060 ;
        RECT 121.820 0.500 121.980 1.060 ;
        RECT 123.820 0.500 123.980 1.060 ;
        RECT 125.820 0.500 125.980 1.060 ;
        RECT 127.820 0.500 127.980 1.060 ;
        RECT 129.820 0.500 129.980 1.060 ;
        RECT 131.820 0.500 131.980 1.060 ;
        RECT 0.000 0.000 133.800 0.500 ;
      LAYER Metal2 ;
        RECT 0.980 0.000 1.270 0.500 ;
        RECT 2.980 0.000 3.270 0.500 ;
        RECT 4.980 0.000 5.270 0.500 ;
        RECT 6.980 0.000 7.270 0.500 ;
        RECT 8.980 0.000 9.270 0.500 ;
        RECT 10.980 0.000 11.270 0.500 ;
        RECT 12.980 0.000 13.270 0.500 ;
        RECT 14.980 0.000 15.270 0.500 ;
        RECT 16.980 0.000 17.270 0.500 ;
        RECT 18.980 0.000 19.270 0.500 ;
        RECT 20.980 0.000 21.270 0.500 ;
        RECT 22.980 0.000 23.270 0.500 ;
        RECT 24.980 0.000 25.270 0.500 ;
        RECT 26.980 0.000 27.270 0.500 ;
        RECT 28.980 0.000 29.270 0.500 ;
        RECT 30.980 0.000 31.270 0.500 ;
        RECT 32.980 0.000 33.270 0.500 ;
        RECT 34.980 0.000 35.270 0.500 ;
        RECT 36.980 0.000 37.270 0.500 ;
        RECT 38.980 0.000 39.270 0.500 ;
        RECT 40.980 0.000 41.270 0.500 ;
        RECT 42.980 0.000 43.270 0.500 ;
        RECT 44.980 0.000 45.270 0.500 ;
        RECT 46.980 0.000 47.270 0.500 ;
        RECT 48.980 0.000 49.270 0.500 ;
        RECT 50.980 0.000 51.270 0.500 ;
        RECT 52.980 0.000 53.270 0.500 ;
        RECT 54.980 0.000 55.270 0.500 ;
        RECT 56.980 0.000 57.270 0.500 ;
        RECT 58.980 0.000 59.270 0.500 ;
        RECT 60.980 0.000 61.270 0.500 ;
        RECT 62.980 0.000 63.270 0.500 ;
        RECT 64.980 0.000 65.270 0.500 ;
        RECT 66.980 0.000 67.270 0.500 ;
        RECT 68.980 0.000 69.270 0.500 ;
        RECT 70.980 0.000 71.270 0.500 ;
        RECT 72.980 0.000 73.270 0.500 ;
        RECT 74.980 0.000 75.270 0.500 ;
        RECT 76.980 0.000 77.270 0.500 ;
        RECT 78.980 0.000 79.270 0.500 ;
        RECT 80.980 0.000 81.270 0.500 ;
        RECT 82.980 0.000 83.270 0.500 ;
        RECT 84.980 0.000 85.270 0.500 ;
        RECT 86.980 0.000 87.270 0.500 ;
        RECT 88.980 0.000 89.270 0.500 ;
        RECT 90.980 0.000 91.270 0.500 ;
        RECT 92.980 0.000 93.270 0.500 ;
        RECT 94.980 0.000 95.270 0.500 ;
        RECT 96.980 0.000 97.270 0.500 ;
        RECT 98.980 0.000 99.270 0.500 ;
        RECT 100.980 0.000 101.270 0.500 ;
        RECT 102.980 0.000 103.270 0.500 ;
        RECT 104.980 0.000 105.270 0.500 ;
        RECT 106.980 0.000 107.270 0.500 ;
        RECT 108.980 0.000 109.270 0.500 ;
        RECT 110.980 0.000 111.270 0.500 ;
        RECT 112.980 0.000 113.270 0.500 ;
        RECT 114.980 0.000 115.270 0.500 ;
        RECT 116.980 0.000 117.270 0.500 ;
        RECT 118.980 0.000 119.270 0.500 ;
        RECT 120.980 0.000 121.270 0.500 ;
        RECT 122.980 0.000 123.270 0.500 ;
        RECT 124.980 0.000 125.270 0.500 ;
        RECT 126.980 0.000 127.270 0.500 ;
        RECT 128.980 0.000 129.270 0.500 ;
        RECT 130.980 0.000 131.270 0.500 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 133.800 1.730 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0.000 25.690 133.800 26.190 ;
        RECT 1.820 25.130 1.980 25.690 ;
        RECT 3.820 25.130 3.980 25.690 ;
        RECT 5.820 25.130 5.980 25.690 ;
        RECT 7.820 25.130 7.980 25.690 ;
        RECT 9.820 25.130 9.980 25.690 ;
        RECT 11.820 25.130 11.980 25.690 ;
        RECT 13.820 25.130 13.980 25.690 ;
        RECT 15.820 25.130 15.980 25.690 ;
        RECT 17.820 25.130 17.980 25.690 ;
        RECT 19.820 25.130 19.980 25.690 ;
        RECT 21.820 25.130 21.980 25.690 ;
        RECT 23.820 25.130 23.980 25.690 ;
        RECT 25.820 25.130 25.980 25.690 ;
        RECT 27.820 25.130 27.980 25.690 ;
        RECT 29.820 25.130 29.980 25.690 ;
        RECT 31.820 25.130 31.980 25.690 ;
        RECT 33.820 25.130 33.980 25.690 ;
        RECT 35.820 25.130 35.980 25.690 ;
        RECT 37.820 25.130 37.980 25.690 ;
        RECT 39.820 25.130 39.980 25.690 ;
        RECT 41.820 25.130 41.980 25.690 ;
        RECT 43.820 25.130 43.980 25.690 ;
        RECT 45.820 25.130 45.980 25.690 ;
        RECT 47.820 25.130 47.980 25.690 ;
        RECT 49.820 25.130 49.980 25.690 ;
        RECT 51.820 25.130 51.980 25.690 ;
        RECT 53.820 25.130 53.980 25.690 ;
        RECT 55.820 25.130 55.980 25.690 ;
        RECT 57.820 25.130 57.980 25.690 ;
        RECT 59.820 25.130 59.980 25.690 ;
        RECT 61.820 25.130 61.980 25.690 ;
        RECT 63.820 25.130 63.980 25.690 ;
        RECT 65.820 25.130 65.980 25.690 ;
        RECT 67.820 25.130 67.980 25.690 ;
        RECT 69.820 25.130 69.980 25.690 ;
        RECT 71.820 25.130 71.980 25.690 ;
        RECT 73.820 25.130 73.980 25.690 ;
        RECT 75.820 25.130 75.980 25.690 ;
        RECT 77.820 25.130 77.980 25.690 ;
        RECT 79.820 25.130 79.980 25.690 ;
        RECT 81.820 25.130 81.980 25.690 ;
        RECT 83.820 25.130 83.980 25.690 ;
        RECT 85.820 25.130 85.980 25.690 ;
        RECT 87.820 25.130 87.980 25.690 ;
        RECT 89.820 25.130 89.980 25.690 ;
        RECT 91.820 25.130 91.980 25.690 ;
        RECT 93.820 25.130 93.980 25.690 ;
        RECT 95.820 25.130 95.980 25.690 ;
        RECT 97.820 25.130 97.980 25.690 ;
        RECT 99.820 25.130 99.980 25.690 ;
        RECT 101.820 25.130 101.980 25.690 ;
        RECT 103.820 25.130 103.980 25.690 ;
        RECT 105.820 25.130 105.980 25.690 ;
        RECT 107.820 25.130 107.980 25.690 ;
        RECT 109.820 25.130 109.980 25.690 ;
        RECT 111.820 25.130 111.980 25.690 ;
        RECT 113.820 25.130 113.980 25.690 ;
        RECT 115.820 25.130 115.980 25.690 ;
        RECT 117.820 25.130 117.980 25.690 ;
        RECT 119.820 25.130 119.980 25.690 ;
        RECT 121.820 25.130 121.980 25.690 ;
        RECT 123.820 25.130 123.980 25.690 ;
        RECT 125.820 25.130 125.980 25.690 ;
        RECT 127.820 25.130 127.980 25.690 ;
        RECT 129.820 25.130 129.980 25.690 ;
        RECT 131.820 25.130 131.980 25.690 ;
      LAYER Metal2 ;
        RECT 2.530 25.690 2.820 26.190 ;
        RECT 4.530 25.690 4.820 26.190 ;
        RECT 6.530 25.690 6.820 26.190 ;
        RECT 8.530 25.690 8.820 26.190 ;
        RECT 10.530 25.690 10.820 26.190 ;
        RECT 12.530 25.690 12.820 26.190 ;
        RECT 14.530 25.690 14.820 26.190 ;
        RECT 16.530 25.690 16.820 26.190 ;
        RECT 18.530 25.690 18.820 26.190 ;
        RECT 20.530 25.690 20.820 26.190 ;
        RECT 22.530 25.690 22.820 26.190 ;
        RECT 24.530 25.690 24.820 26.190 ;
        RECT 26.530 25.690 26.820 26.190 ;
        RECT 28.530 25.690 28.820 26.190 ;
        RECT 30.530 25.690 30.820 26.190 ;
        RECT 32.530 25.690 32.820 26.190 ;
        RECT 34.530 25.690 34.820 26.190 ;
        RECT 36.530 25.690 36.820 26.190 ;
        RECT 38.530 25.690 38.820 26.190 ;
        RECT 40.530 25.690 40.820 26.190 ;
        RECT 42.530 25.690 42.820 26.190 ;
        RECT 44.530 25.690 44.820 26.190 ;
        RECT 46.530 25.690 46.820 26.190 ;
        RECT 48.530 25.690 48.820 26.190 ;
        RECT 50.530 25.690 50.820 26.190 ;
        RECT 52.530 25.690 52.820 26.190 ;
        RECT 54.530 25.690 54.820 26.190 ;
        RECT 56.530 25.690 56.820 26.190 ;
        RECT 58.530 25.690 58.820 26.190 ;
        RECT 60.530 25.690 60.820 26.190 ;
        RECT 62.530 25.690 62.820 26.190 ;
        RECT 64.530 25.690 64.820 26.190 ;
        RECT 66.530 25.690 66.820 26.190 ;
        RECT 68.530 25.690 68.820 26.190 ;
        RECT 70.530 25.690 70.820 26.190 ;
        RECT 72.530 25.690 72.820 26.190 ;
        RECT 74.530 25.690 74.820 26.190 ;
        RECT 76.530 25.690 76.820 26.190 ;
        RECT 78.530 25.690 78.820 26.190 ;
        RECT 80.530 25.690 80.820 26.190 ;
        RECT 82.530 25.690 82.820 26.190 ;
        RECT 84.530 25.690 84.820 26.190 ;
        RECT 86.530 25.690 86.820 26.190 ;
        RECT 88.530 25.690 88.820 26.190 ;
        RECT 90.530 25.690 90.820 26.190 ;
        RECT 92.530 25.690 92.820 26.190 ;
        RECT 94.530 25.690 94.820 26.190 ;
        RECT 96.530 25.690 96.820 26.190 ;
        RECT 98.530 25.690 98.820 26.190 ;
        RECT 100.530 25.690 100.820 26.190 ;
        RECT 102.530 25.690 102.820 26.190 ;
        RECT 104.530 25.690 104.820 26.190 ;
        RECT 106.530 25.690 106.820 26.190 ;
        RECT 108.530 25.690 108.820 26.190 ;
        RECT 110.530 25.690 110.820 26.190 ;
        RECT 112.530 25.690 112.820 26.190 ;
        RECT 114.530 25.690 114.820 26.190 ;
        RECT 116.530 25.690 116.820 26.190 ;
        RECT 118.530 25.690 118.820 26.190 ;
        RECT 120.530 25.690 120.820 26.190 ;
        RECT 122.530 25.690 122.820 26.190 ;
        RECT 124.530 25.690 124.820 26.190 ;
        RECT 126.530 25.690 126.820 26.190 ;
        RECT 128.530 25.690 128.820 26.190 ;
        RECT 130.530 25.690 130.820 26.190 ;
        RECT 132.530 25.690 132.820 26.190 ;
      LAYER Metal3 ;
        RECT 0.000 24.460 133.800 26.190 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 1.820 22.610 1.980 23.290 ;
        RECT 3.820 22.610 3.980 23.290 ;
        RECT 5.820 22.610 5.980 23.290 ;
        RECT 7.820 22.610 7.980 23.290 ;
        RECT 9.820 22.610 9.980 23.290 ;
        RECT 11.820 22.610 11.980 23.290 ;
        RECT 13.820 22.610 13.980 23.290 ;
        RECT 15.820 22.610 15.980 23.290 ;
        RECT 17.820 22.610 17.980 23.290 ;
        RECT 19.820 22.610 19.980 23.290 ;
        RECT 21.820 22.610 21.980 23.290 ;
        RECT 23.820 22.610 23.980 23.290 ;
        RECT 25.820 22.610 25.980 23.290 ;
        RECT 27.820 22.610 27.980 23.290 ;
        RECT 29.820 22.610 29.980 23.290 ;
        RECT 31.820 22.610 31.980 23.290 ;
        RECT 33.820 22.610 33.980 23.290 ;
        RECT 35.820 22.610 35.980 23.290 ;
        RECT 37.820 22.610 37.980 23.290 ;
        RECT 39.820 22.610 39.980 23.290 ;
        RECT 41.820 22.610 41.980 23.290 ;
        RECT 43.820 22.610 43.980 23.290 ;
        RECT 45.820 22.610 45.980 23.290 ;
        RECT 47.820 22.610 47.980 23.290 ;
        RECT 49.820 22.610 49.980 23.290 ;
        RECT 51.820 22.610 51.980 23.290 ;
        RECT 53.820 22.610 53.980 23.290 ;
        RECT 55.820 22.610 55.980 23.290 ;
        RECT 57.820 22.610 57.980 23.290 ;
        RECT 59.820 22.610 59.980 23.290 ;
        RECT 61.820 22.610 61.980 23.290 ;
        RECT 63.820 22.610 63.980 23.290 ;
        RECT 65.820 22.610 65.980 23.290 ;
        RECT 67.820 22.610 67.980 23.290 ;
        RECT 69.820 22.610 69.980 23.290 ;
        RECT 71.820 22.610 71.980 23.290 ;
        RECT 73.820 22.610 73.980 23.290 ;
        RECT 75.820 22.610 75.980 23.290 ;
        RECT 77.820 22.610 77.980 23.290 ;
        RECT 79.820 22.610 79.980 23.290 ;
        RECT 81.820 22.610 81.980 23.290 ;
        RECT 83.820 22.610 83.980 23.290 ;
        RECT 85.820 22.610 85.980 23.290 ;
        RECT 87.820 22.610 87.980 23.290 ;
        RECT 89.820 22.610 89.980 23.290 ;
        RECT 91.820 22.610 91.980 23.290 ;
        RECT 93.820 22.610 93.980 23.290 ;
        RECT 95.820 22.610 95.980 23.290 ;
        RECT 97.820 22.610 97.980 23.290 ;
        RECT 99.820 22.610 99.980 23.290 ;
        RECT 101.820 22.610 101.980 23.290 ;
        RECT 103.820 22.610 103.980 23.290 ;
        RECT 105.820 22.610 105.980 23.290 ;
        RECT 107.820 22.610 107.980 23.290 ;
        RECT 109.820 22.610 109.980 23.290 ;
        RECT 111.820 22.610 111.980 23.290 ;
        RECT 113.820 22.610 113.980 23.290 ;
        RECT 115.820 22.610 115.980 23.290 ;
        RECT 117.820 22.610 117.980 23.290 ;
        RECT 119.820 22.610 119.980 23.290 ;
        RECT 121.820 22.610 121.980 23.290 ;
        RECT 123.820 22.610 123.980 23.290 ;
        RECT 125.820 22.610 125.980 23.290 ;
        RECT 127.820 22.610 127.980 23.290 ;
        RECT 129.820 22.610 129.980 23.290 ;
        RECT 131.820 22.610 131.980 23.290 ;
        RECT 0.900 22.110 132.900 22.610 ;
        RECT 0.970 21.410 1.230 22.110 ;
        RECT 2.970 21.410 3.230 22.110 ;
        RECT 4.970 21.410 5.230 22.110 ;
        RECT 6.970 21.410 7.230 22.110 ;
        RECT 8.970 21.410 9.230 22.110 ;
        RECT 10.970 21.410 11.230 22.110 ;
        RECT 12.970 21.410 13.230 22.110 ;
        RECT 14.970 21.410 15.230 22.110 ;
        RECT 16.970 21.410 17.230 22.110 ;
        RECT 18.970 21.410 19.230 22.110 ;
        RECT 20.970 21.410 21.230 22.110 ;
        RECT 22.970 21.410 23.230 22.110 ;
        RECT 24.970 21.410 25.230 22.110 ;
        RECT 26.970 21.410 27.230 22.110 ;
        RECT 28.970 21.410 29.230 22.110 ;
        RECT 30.970 21.410 31.230 22.110 ;
        RECT 32.970 21.410 33.230 22.110 ;
        RECT 34.970 21.410 35.230 22.110 ;
        RECT 36.970 21.410 37.230 22.110 ;
        RECT 38.970 21.410 39.230 22.110 ;
        RECT 40.970 21.410 41.230 22.110 ;
        RECT 42.970 21.410 43.230 22.110 ;
        RECT 44.970 21.410 45.230 22.110 ;
        RECT 46.970 21.410 47.230 22.110 ;
        RECT 48.970 21.410 49.230 22.110 ;
        RECT 50.970 21.410 51.230 22.110 ;
        RECT 52.970 21.410 53.230 22.110 ;
        RECT 54.970 21.410 55.230 22.110 ;
        RECT 56.970 21.410 57.230 22.110 ;
        RECT 58.970 21.410 59.230 22.110 ;
        RECT 60.970 21.410 61.230 22.110 ;
        RECT 62.970 21.410 63.230 22.110 ;
        RECT 64.970 21.410 65.230 22.110 ;
        RECT 66.970 21.410 67.230 22.110 ;
        RECT 68.970 21.410 69.230 22.110 ;
        RECT 70.970 21.410 71.230 22.110 ;
        RECT 72.970 21.410 73.230 22.110 ;
        RECT 74.970 21.410 75.230 22.110 ;
        RECT 76.970 21.410 77.230 22.110 ;
        RECT 78.970 21.410 79.230 22.110 ;
        RECT 80.970 21.410 81.230 22.110 ;
        RECT 82.970 21.410 83.230 22.110 ;
        RECT 84.970 21.410 85.230 22.110 ;
        RECT 86.970 21.410 87.230 22.110 ;
        RECT 88.970 21.410 89.230 22.110 ;
        RECT 90.970 21.410 91.230 22.110 ;
        RECT 92.970 21.410 93.230 22.110 ;
        RECT 94.970 21.410 95.230 22.110 ;
        RECT 96.970 21.410 97.230 22.110 ;
        RECT 98.970 21.410 99.230 22.110 ;
        RECT 100.970 21.410 101.230 22.110 ;
        RECT 102.970 21.410 103.230 22.110 ;
        RECT 104.970 21.410 105.230 22.110 ;
        RECT 106.970 21.410 107.230 22.110 ;
        RECT 108.970 21.410 109.230 22.110 ;
        RECT 110.970 21.410 111.230 22.110 ;
        RECT 112.970 21.410 113.230 22.110 ;
        RECT 114.970 21.410 115.230 22.110 ;
        RECT 116.970 21.410 117.230 22.110 ;
        RECT 118.970 21.410 119.230 22.110 ;
        RECT 120.970 21.410 121.230 22.110 ;
        RECT 122.970 21.410 123.230 22.110 ;
        RECT 124.970 21.410 125.230 22.110 ;
        RECT 126.970 21.410 127.230 22.110 ;
        RECT 128.970 21.410 129.230 22.110 ;
        RECT 130.970 21.410 131.230 22.110 ;
        RECT 0.970 20.730 1.470 21.410 ;
        RECT 2.970 20.730 3.470 21.410 ;
        RECT 4.970 20.730 5.470 21.410 ;
        RECT 6.970 20.730 7.470 21.410 ;
        RECT 8.970 20.730 9.470 21.410 ;
        RECT 10.970 20.730 11.470 21.410 ;
        RECT 12.970 20.730 13.470 21.410 ;
        RECT 14.970 20.730 15.470 21.410 ;
        RECT 16.970 20.730 17.470 21.410 ;
        RECT 18.970 20.730 19.470 21.410 ;
        RECT 20.970 20.730 21.470 21.410 ;
        RECT 22.970 20.730 23.470 21.410 ;
        RECT 24.970 20.730 25.470 21.410 ;
        RECT 26.970 20.730 27.470 21.410 ;
        RECT 28.970 20.730 29.470 21.410 ;
        RECT 30.970 20.730 31.470 21.410 ;
        RECT 32.970 20.730 33.470 21.410 ;
        RECT 34.970 20.730 35.470 21.410 ;
        RECT 36.970 20.730 37.470 21.410 ;
        RECT 38.970 20.730 39.470 21.410 ;
        RECT 40.970 20.730 41.470 21.410 ;
        RECT 42.970 20.730 43.470 21.410 ;
        RECT 44.970 20.730 45.470 21.410 ;
        RECT 46.970 20.730 47.470 21.410 ;
        RECT 48.970 20.730 49.470 21.410 ;
        RECT 50.970 20.730 51.470 21.410 ;
        RECT 52.970 20.730 53.470 21.410 ;
        RECT 54.970 20.730 55.470 21.410 ;
        RECT 56.970 20.730 57.470 21.410 ;
        RECT 58.970 20.730 59.470 21.410 ;
        RECT 60.970 20.730 61.470 21.410 ;
        RECT 62.970 20.730 63.470 21.410 ;
        RECT 64.970 20.730 65.470 21.410 ;
        RECT 66.970 20.730 67.470 21.410 ;
        RECT 68.970 20.730 69.470 21.410 ;
        RECT 70.970 20.730 71.470 21.410 ;
        RECT 72.970 20.730 73.470 21.410 ;
        RECT 74.970 20.730 75.470 21.410 ;
        RECT 76.970 20.730 77.470 21.410 ;
        RECT 78.970 20.730 79.470 21.410 ;
        RECT 80.970 20.730 81.470 21.410 ;
        RECT 82.970 20.730 83.470 21.410 ;
        RECT 84.970 20.730 85.470 21.410 ;
        RECT 86.970 20.730 87.470 21.410 ;
        RECT 88.970 20.730 89.470 21.410 ;
        RECT 90.970 20.730 91.470 21.410 ;
        RECT 92.970 20.730 93.470 21.410 ;
        RECT 94.970 20.730 95.470 21.410 ;
        RECT 96.970 20.730 97.470 21.410 ;
        RECT 98.970 20.730 99.470 21.410 ;
        RECT 100.970 20.730 101.470 21.410 ;
        RECT 102.970 20.730 103.470 21.410 ;
        RECT 104.970 20.730 105.470 21.410 ;
        RECT 106.970 20.730 107.470 21.410 ;
        RECT 108.970 20.730 109.470 21.410 ;
        RECT 110.970 20.730 111.470 21.410 ;
        RECT 112.970 20.730 113.470 21.410 ;
        RECT 114.970 20.730 115.470 21.410 ;
        RECT 116.970 20.730 117.470 21.410 ;
        RECT 118.970 20.730 119.470 21.410 ;
        RECT 120.970 20.730 121.470 21.410 ;
        RECT 122.970 20.730 123.470 21.410 ;
        RECT 124.970 20.730 125.470 21.410 ;
        RECT 126.970 20.730 127.470 21.410 ;
        RECT 128.970 20.730 129.470 21.410 ;
        RECT 130.970 20.730 131.470 21.410 ;
        RECT 0.900 20.060 132.900 20.730 ;
        RECT 0.900 5.460 132.900 6.130 ;
        RECT 2.330 4.780 2.830 5.460 ;
        RECT 4.330 4.780 4.830 5.460 ;
        RECT 6.330 4.780 6.830 5.460 ;
        RECT 8.330 4.780 8.830 5.460 ;
        RECT 10.330 4.780 10.830 5.460 ;
        RECT 12.330 4.780 12.830 5.460 ;
        RECT 14.330 4.780 14.830 5.460 ;
        RECT 16.330 4.780 16.830 5.460 ;
        RECT 18.330 4.780 18.830 5.460 ;
        RECT 20.330 4.780 20.830 5.460 ;
        RECT 22.330 4.780 22.830 5.460 ;
        RECT 24.330 4.780 24.830 5.460 ;
        RECT 26.330 4.780 26.830 5.460 ;
        RECT 28.330 4.780 28.830 5.460 ;
        RECT 30.330 4.780 30.830 5.460 ;
        RECT 32.330 4.780 32.830 5.460 ;
        RECT 34.330 4.780 34.830 5.460 ;
        RECT 36.330 4.780 36.830 5.460 ;
        RECT 38.330 4.780 38.830 5.460 ;
        RECT 40.330 4.780 40.830 5.460 ;
        RECT 42.330 4.780 42.830 5.460 ;
        RECT 44.330 4.780 44.830 5.460 ;
        RECT 46.330 4.780 46.830 5.460 ;
        RECT 48.330 4.780 48.830 5.460 ;
        RECT 50.330 4.780 50.830 5.460 ;
        RECT 52.330 4.780 52.830 5.460 ;
        RECT 54.330 4.780 54.830 5.460 ;
        RECT 56.330 4.780 56.830 5.460 ;
        RECT 58.330 4.780 58.830 5.460 ;
        RECT 60.330 4.780 60.830 5.460 ;
        RECT 62.330 4.780 62.830 5.460 ;
        RECT 64.330 4.780 64.830 5.460 ;
        RECT 66.330 4.780 66.830 5.460 ;
        RECT 68.330 4.780 68.830 5.460 ;
        RECT 70.330 4.780 70.830 5.460 ;
        RECT 72.330 4.780 72.830 5.460 ;
        RECT 74.330 4.780 74.830 5.460 ;
        RECT 76.330 4.780 76.830 5.460 ;
        RECT 78.330 4.780 78.830 5.460 ;
        RECT 80.330 4.780 80.830 5.460 ;
        RECT 82.330 4.780 82.830 5.460 ;
        RECT 84.330 4.780 84.830 5.460 ;
        RECT 86.330 4.780 86.830 5.460 ;
        RECT 88.330 4.780 88.830 5.460 ;
        RECT 90.330 4.780 90.830 5.460 ;
        RECT 92.330 4.780 92.830 5.460 ;
        RECT 94.330 4.780 94.830 5.460 ;
        RECT 96.330 4.780 96.830 5.460 ;
        RECT 98.330 4.780 98.830 5.460 ;
        RECT 100.330 4.780 100.830 5.460 ;
        RECT 102.330 4.780 102.830 5.460 ;
        RECT 104.330 4.780 104.830 5.460 ;
        RECT 106.330 4.780 106.830 5.460 ;
        RECT 108.330 4.780 108.830 5.460 ;
        RECT 110.330 4.780 110.830 5.460 ;
        RECT 112.330 4.780 112.830 5.460 ;
        RECT 114.330 4.780 114.830 5.460 ;
        RECT 116.330 4.780 116.830 5.460 ;
        RECT 118.330 4.780 118.830 5.460 ;
        RECT 120.330 4.780 120.830 5.460 ;
        RECT 122.330 4.780 122.830 5.460 ;
        RECT 124.330 4.780 124.830 5.460 ;
        RECT 126.330 4.780 126.830 5.460 ;
        RECT 128.330 4.780 128.830 5.460 ;
        RECT 130.330 4.780 130.830 5.460 ;
        RECT 132.330 4.780 132.830 5.460 ;
        RECT 2.570 4.080 2.830 4.780 ;
        RECT 4.570 4.080 4.830 4.780 ;
        RECT 6.570 4.080 6.830 4.780 ;
        RECT 8.570 4.080 8.830 4.780 ;
        RECT 10.570 4.080 10.830 4.780 ;
        RECT 12.570 4.080 12.830 4.780 ;
        RECT 14.570 4.080 14.830 4.780 ;
        RECT 16.570 4.080 16.830 4.780 ;
        RECT 18.570 4.080 18.830 4.780 ;
        RECT 20.570 4.080 20.830 4.780 ;
        RECT 22.570 4.080 22.830 4.780 ;
        RECT 24.570 4.080 24.830 4.780 ;
        RECT 26.570 4.080 26.830 4.780 ;
        RECT 28.570 4.080 28.830 4.780 ;
        RECT 30.570 4.080 30.830 4.780 ;
        RECT 32.570 4.080 32.830 4.780 ;
        RECT 34.570 4.080 34.830 4.780 ;
        RECT 36.570 4.080 36.830 4.780 ;
        RECT 38.570 4.080 38.830 4.780 ;
        RECT 40.570 4.080 40.830 4.780 ;
        RECT 42.570 4.080 42.830 4.780 ;
        RECT 44.570 4.080 44.830 4.780 ;
        RECT 46.570 4.080 46.830 4.780 ;
        RECT 48.570 4.080 48.830 4.780 ;
        RECT 50.570 4.080 50.830 4.780 ;
        RECT 52.570 4.080 52.830 4.780 ;
        RECT 54.570 4.080 54.830 4.780 ;
        RECT 56.570 4.080 56.830 4.780 ;
        RECT 58.570 4.080 58.830 4.780 ;
        RECT 60.570 4.080 60.830 4.780 ;
        RECT 62.570 4.080 62.830 4.780 ;
        RECT 64.570 4.080 64.830 4.780 ;
        RECT 66.570 4.080 66.830 4.780 ;
        RECT 68.570 4.080 68.830 4.780 ;
        RECT 70.570 4.080 70.830 4.780 ;
        RECT 72.570 4.080 72.830 4.780 ;
        RECT 74.570 4.080 74.830 4.780 ;
        RECT 76.570 4.080 76.830 4.780 ;
        RECT 78.570 4.080 78.830 4.780 ;
        RECT 80.570 4.080 80.830 4.780 ;
        RECT 82.570 4.080 82.830 4.780 ;
        RECT 84.570 4.080 84.830 4.780 ;
        RECT 86.570 4.080 86.830 4.780 ;
        RECT 88.570 4.080 88.830 4.780 ;
        RECT 90.570 4.080 90.830 4.780 ;
        RECT 92.570 4.080 92.830 4.780 ;
        RECT 94.570 4.080 94.830 4.780 ;
        RECT 96.570 4.080 96.830 4.780 ;
        RECT 98.570 4.080 98.830 4.780 ;
        RECT 100.570 4.080 100.830 4.780 ;
        RECT 102.570 4.080 102.830 4.780 ;
        RECT 104.570 4.080 104.830 4.780 ;
        RECT 106.570 4.080 106.830 4.780 ;
        RECT 108.570 4.080 108.830 4.780 ;
        RECT 110.570 4.080 110.830 4.780 ;
        RECT 112.570 4.080 112.830 4.780 ;
        RECT 114.570 4.080 114.830 4.780 ;
        RECT 116.570 4.080 116.830 4.780 ;
        RECT 118.570 4.080 118.830 4.780 ;
        RECT 120.570 4.080 120.830 4.780 ;
        RECT 122.570 4.080 122.830 4.780 ;
        RECT 124.570 4.080 124.830 4.780 ;
        RECT 126.570 4.080 126.830 4.780 ;
        RECT 128.570 4.080 128.830 4.780 ;
        RECT 130.570 4.080 130.830 4.780 ;
        RECT 132.570 4.080 132.830 4.780 ;
        RECT 0.900 3.580 132.900 4.080 ;
        RECT 1.820 2.900 1.980 3.580 ;
        RECT 3.820 2.900 3.980 3.580 ;
        RECT 5.820 2.900 5.980 3.580 ;
        RECT 7.820 2.900 7.980 3.580 ;
        RECT 9.820 2.900 9.980 3.580 ;
        RECT 11.820 2.900 11.980 3.580 ;
        RECT 13.820 2.900 13.980 3.580 ;
        RECT 15.820 2.900 15.980 3.580 ;
        RECT 17.820 2.900 17.980 3.580 ;
        RECT 19.820 2.900 19.980 3.580 ;
        RECT 21.820 2.900 21.980 3.580 ;
        RECT 23.820 2.900 23.980 3.580 ;
        RECT 25.820 2.900 25.980 3.580 ;
        RECT 27.820 2.900 27.980 3.580 ;
        RECT 29.820 2.900 29.980 3.580 ;
        RECT 31.820 2.900 31.980 3.580 ;
        RECT 33.820 2.900 33.980 3.580 ;
        RECT 35.820 2.900 35.980 3.580 ;
        RECT 37.820 2.900 37.980 3.580 ;
        RECT 39.820 2.900 39.980 3.580 ;
        RECT 41.820 2.900 41.980 3.580 ;
        RECT 43.820 2.900 43.980 3.580 ;
        RECT 45.820 2.900 45.980 3.580 ;
        RECT 47.820 2.900 47.980 3.580 ;
        RECT 49.820 2.900 49.980 3.580 ;
        RECT 51.820 2.900 51.980 3.580 ;
        RECT 53.820 2.900 53.980 3.580 ;
        RECT 55.820 2.900 55.980 3.580 ;
        RECT 57.820 2.900 57.980 3.580 ;
        RECT 59.820 2.900 59.980 3.580 ;
        RECT 61.820 2.900 61.980 3.580 ;
        RECT 63.820 2.900 63.980 3.580 ;
        RECT 65.820 2.900 65.980 3.580 ;
        RECT 67.820 2.900 67.980 3.580 ;
        RECT 69.820 2.900 69.980 3.580 ;
        RECT 71.820 2.900 71.980 3.580 ;
        RECT 73.820 2.900 73.980 3.580 ;
        RECT 75.820 2.900 75.980 3.580 ;
        RECT 77.820 2.900 77.980 3.580 ;
        RECT 79.820 2.900 79.980 3.580 ;
        RECT 81.820 2.900 81.980 3.580 ;
        RECT 83.820 2.900 83.980 3.580 ;
        RECT 85.820 2.900 85.980 3.580 ;
        RECT 87.820 2.900 87.980 3.580 ;
        RECT 89.820 2.900 89.980 3.580 ;
        RECT 91.820 2.900 91.980 3.580 ;
        RECT 93.820 2.900 93.980 3.580 ;
        RECT 95.820 2.900 95.980 3.580 ;
        RECT 97.820 2.900 97.980 3.580 ;
        RECT 99.820 2.900 99.980 3.580 ;
        RECT 101.820 2.900 101.980 3.580 ;
        RECT 103.820 2.900 103.980 3.580 ;
        RECT 105.820 2.900 105.980 3.580 ;
        RECT 107.820 2.900 107.980 3.580 ;
        RECT 109.820 2.900 109.980 3.580 ;
        RECT 111.820 2.900 111.980 3.580 ;
        RECT 113.820 2.900 113.980 3.580 ;
        RECT 115.820 2.900 115.980 3.580 ;
        RECT 117.820 2.900 117.980 3.580 ;
        RECT 119.820 2.900 119.980 3.580 ;
        RECT 121.820 2.900 121.980 3.580 ;
        RECT 123.820 2.900 123.980 3.580 ;
        RECT 125.820 2.900 125.980 3.580 ;
        RECT 127.820 2.900 127.980 3.580 ;
        RECT 129.820 2.900 129.980 3.580 ;
        RECT 131.820 2.900 131.980 3.580 ;
      LAYER Metal2 ;
        RECT 1.550 22.215 2.250 22.505 ;
        RECT 3.550 22.215 4.250 22.505 ;
        RECT 5.550 22.215 6.250 22.505 ;
        RECT 7.550 22.215 8.250 22.505 ;
        RECT 9.550 22.215 10.250 22.505 ;
        RECT 11.550 22.215 12.250 22.505 ;
        RECT 13.550 22.215 14.250 22.505 ;
        RECT 15.550 22.215 16.250 22.505 ;
        RECT 17.550 22.215 18.250 22.505 ;
        RECT 19.550 22.215 20.250 22.505 ;
        RECT 21.550 22.215 22.250 22.505 ;
        RECT 23.550 22.215 24.250 22.505 ;
        RECT 25.550 22.215 26.250 22.505 ;
        RECT 27.550 22.215 28.250 22.505 ;
        RECT 29.550 22.215 30.250 22.505 ;
        RECT 31.550 22.215 32.250 22.505 ;
        RECT 33.550 22.215 34.250 22.505 ;
        RECT 35.550 22.215 36.250 22.505 ;
        RECT 37.550 22.215 38.250 22.505 ;
        RECT 39.550 22.215 40.250 22.505 ;
        RECT 41.550 22.215 42.250 22.505 ;
        RECT 43.550 22.215 44.250 22.505 ;
        RECT 45.550 22.215 46.250 22.505 ;
        RECT 47.550 22.215 48.250 22.505 ;
        RECT 49.550 22.215 50.250 22.505 ;
        RECT 51.550 22.215 52.250 22.505 ;
        RECT 53.550 22.215 54.250 22.505 ;
        RECT 55.550 22.215 56.250 22.505 ;
        RECT 57.550 22.215 58.250 22.505 ;
        RECT 59.550 22.215 60.250 22.505 ;
        RECT 61.550 22.215 62.250 22.505 ;
        RECT 63.550 22.215 64.250 22.505 ;
        RECT 65.550 22.215 66.250 22.505 ;
        RECT 67.550 22.215 68.250 22.505 ;
        RECT 69.550 22.215 70.250 22.505 ;
        RECT 71.550 22.215 72.250 22.505 ;
        RECT 73.550 22.215 74.250 22.505 ;
        RECT 75.550 22.215 76.250 22.505 ;
        RECT 77.550 22.215 78.250 22.505 ;
        RECT 79.550 22.215 80.250 22.505 ;
        RECT 81.550 22.215 82.250 22.505 ;
        RECT 83.550 22.215 84.250 22.505 ;
        RECT 85.550 22.215 86.250 22.505 ;
        RECT 87.550 22.215 88.250 22.505 ;
        RECT 89.550 22.215 90.250 22.505 ;
        RECT 91.550 22.215 92.250 22.505 ;
        RECT 93.550 22.215 94.250 22.505 ;
        RECT 95.550 22.215 96.250 22.505 ;
        RECT 97.550 22.215 98.250 22.505 ;
        RECT 99.550 22.215 100.250 22.505 ;
        RECT 101.550 22.215 102.250 22.505 ;
        RECT 103.550 22.215 104.250 22.505 ;
        RECT 105.550 22.215 106.250 22.505 ;
        RECT 107.550 22.215 108.250 22.505 ;
        RECT 109.550 22.215 110.250 22.505 ;
        RECT 111.550 22.215 112.250 22.505 ;
        RECT 113.550 22.215 114.250 22.505 ;
        RECT 115.550 22.215 116.250 22.505 ;
        RECT 117.550 22.215 118.250 22.505 ;
        RECT 119.550 22.215 120.250 22.505 ;
        RECT 121.550 22.215 122.250 22.505 ;
        RECT 123.550 22.215 124.250 22.505 ;
        RECT 125.550 22.215 126.250 22.505 ;
        RECT 127.550 22.215 128.250 22.505 ;
        RECT 129.550 22.215 130.250 22.505 ;
        RECT 131.550 22.215 132.250 22.505 ;
        RECT 1.105 20.060 1.395 20.760 ;
        RECT 3.105 20.060 3.395 20.760 ;
        RECT 5.105 20.060 5.395 20.760 ;
        RECT 7.105 20.060 7.395 20.760 ;
        RECT 9.105 20.060 9.395 20.760 ;
        RECT 11.105 20.060 11.395 20.760 ;
        RECT 13.105 20.060 13.395 20.760 ;
        RECT 15.105 20.060 15.395 20.760 ;
        RECT 17.105 20.060 17.395 20.760 ;
        RECT 19.105 20.060 19.395 20.760 ;
        RECT 21.105 20.060 21.395 20.760 ;
        RECT 23.105 20.060 23.395 20.760 ;
        RECT 25.105 20.060 25.395 20.760 ;
        RECT 27.105 20.060 27.395 20.760 ;
        RECT 29.105 20.060 29.395 20.760 ;
        RECT 31.105 20.060 31.395 20.760 ;
        RECT 33.105 20.060 33.395 20.760 ;
        RECT 35.105 20.060 35.395 20.760 ;
        RECT 37.105 20.060 37.395 20.760 ;
        RECT 39.105 20.060 39.395 20.760 ;
        RECT 41.105 20.060 41.395 20.760 ;
        RECT 43.105 20.060 43.395 20.760 ;
        RECT 45.105 20.060 45.395 20.760 ;
        RECT 47.105 20.060 47.395 20.760 ;
        RECT 49.105 20.060 49.395 20.760 ;
        RECT 51.105 20.060 51.395 20.760 ;
        RECT 53.105 20.060 53.395 20.760 ;
        RECT 55.105 20.060 55.395 20.760 ;
        RECT 57.105 20.060 57.395 20.760 ;
        RECT 59.105 20.060 59.395 20.760 ;
        RECT 61.105 20.060 61.395 20.760 ;
        RECT 63.105 20.060 63.395 20.760 ;
        RECT 65.105 20.060 65.395 20.760 ;
        RECT 67.105 20.060 67.395 20.760 ;
        RECT 69.105 20.060 69.395 20.760 ;
        RECT 71.105 20.060 71.395 20.760 ;
        RECT 73.105 20.060 73.395 20.760 ;
        RECT 75.105 20.060 75.395 20.760 ;
        RECT 77.105 20.060 77.395 20.760 ;
        RECT 79.105 20.060 79.395 20.760 ;
        RECT 81.105 20.060 81.395 20.760 ;
        RECT 83.105 20.060 83.395 20.760 ;
        RECT 85.105 20.060 85.395 20.760 ;
        RECT 87.105 20.060 87.395 20.760 ;
        RECT 89.105 20.060 89.395 20.760 ;
        RECT 91.105 20.060 91.395 20.760 ;
        RECT 93.105 20.060 93.395 20.760 ;
        RECT 95.105 20.060 95.395 20.760 ;
        RECT 97.105 20.060 97.395 20.760 ;
        RECT 99.105 20.060 99.395 20.760 ;
        RECT 101.105 20.060 101.395 20.760 ;
        RECT 103.105 20.060 103.395 20.760 ;
        RECT 105.105 20.060 105.395 20.760 ;
        RECT 107.105 20.060 107.395 20.760 ;
        RECT 109.105 20.060 109.395 20.760 ;
        RECT 111.105 20.060 111.395 20.760 ;
        RECT 113.105 20.060 113.395 20.760 ;
        RECT 115.105 20.060 115.395 20.760 ;
        RECT 117.105 20.060 117.395 20.760 ;
        RECT 119.105 20.060 119.395 20.760 ;
        RECT 121.105 20.060 121.395 20.760 ;
        RECT 123.105 20.060 123.395 20.760 ;
        RECT 125.105 20.060 125.395 20.760 ;
        RECT 127.105 20.060 127.395 20.760 ;
        RECT 129.105 20.060 129.395 20.760 ;
        RECT 131.105 20.060 131.395 20.760 ;
        RECT 2.405 5.430 2.695 6.130 ;
        RECT 4.405 5.430 4.695 6.130 ;
        RECT 6.405 5.430 6.695 6.130 ;
        RECT 8.405 5.430 8.695 6.130 ;
        RECT 10.405 5.430 10.695 6.130 ;
        RECT 12.405 5.430 12.695 6.130 ;
        RECT 14.405 5.430 14.695 6.130 ;
        RECT 16.405 5.430 16.695 6.130 ;
        RECT 18.405 5.430 18.695 6.130 ;
        RECT 20.405 5.430 20.695 6.130 ;
        RECT 22.405 5.430 22.695 6.130 ;
        RECT 24.405 5.430 24.695 6.130 ;
        RECT 26.405 5.430 26.695 6.130 ;
        RECT 28.405 5.430 28.695 6.130 ;
        RECT 30.405 5.430 30.695 6.130 ;
        RECT 32.405 5.430 32.695 6.130 ;
        RECT 34.405 5.430 34.695 6.130 ;
        RECT 36.405 5.430 36.695 6.130 ;
        RECT 38.405 5.430 38.695 6.130 ;
        RECT 40.405 5.430 40.695 6.130 ;
        RECT 42.405 5.430 42.695 6.130 ;
        RECT 44.405 5.430 44.695 6.130 ;
        RECT 46.405 5.430 46.695 6.130 ;
        RECT 48.405 5.430 48.695 6.130 ;
        RECT 50.405 5.430 50.695 6.130 ;
        RECT 52.405 5.430 52.695 6.130 ;
        RECT 54.405 5.430 54.695 6.130 ;
        RECT 56.405 5.430 56.695 6.130 ;
        RECT 58.405 5.430 58.695 6.130 ;
        RECT 60.405 5.430 60.695 6.130 ;
        RECT 62.405 5.430 62.695 6.130 ;
        RECT 64.405 5.430 64.695 6.130 ;
        RECT 66.405 5.430 66.695 6.130 ;
        RECT 68.405 5.430 68.695 6.130 ;
        RECT 70.405 5.430 70.695 6.130 ;
        RECT 72.405 5.430 72.695 6.130 ;
        RECT 74.405 5.430 74.695 6.130 ;
        RECT 76.405 5.430 76.695 6.130 ;
        RECT 78.405 5.430 78.695 6.130 ;
        RECT 80.405 5.430 80.695 6.130 ;
        RECT 82.405 5.430 82.695 6.130 ;
        RECT 84.405 5.430 84.695 6.130 ;
        RECT 86.405 5.430 86.695 6.130 ;
        RECT 88.405 5.430 88.695 6.130 ;
        RECT 90.405 5.430 90.695 6.130 ;
        RECT 92.405 5.430 92.695 6.130 ;
        RECT 94.405 5.430 94.695 6.130 ;
        RECT 96.405 5.430 96.695 6.130 ;
        RECT 98.405 5.430 98.695 6.130 ;
        RECT 100.405 5.430 100.695 6.130 ;
        RECT 102.405 5.430 102.695 6.130 ;
        RECT 104.405 5.430 104.695 6.130 ;
        RECT 106.405 5.430 106.695 6.130 ;
        RECT 108.405 5.430 108.695 6.130 ;
        RECT 110.405 5.430 110.695 6.130 ;
        RECT 112.405 5.430 112.695 6.130 ;
        RECT 114.405 5.430 114.695 6.130 ;
        RECT 116.405 5.430 116.695 6.130 ;
        RECT 118.405 5.430 118.695 6.130 ;
        RECT 120.405 5.430 120.695 6.130 ;
        RECT 122.405 5.430 122.695 6.130 ;
        RECT 124.405 5.430 124.695 6.130 ;
        RECT 126.405 5.430 126.695 6.130 ;
        RECT 128.405 5.430 128.695 6.130 ;
        RECT 130.405 5.430 130.695 6.130 ;
        RECT 132.405 5.430 132.695 6.130 ;
        RECT 1.550 3.685 2.250 3.975 ;
        RECT 3.550 3.685 4.250 3.975 ;
        RECT 5.550 3.685 6.250 3.975 ;
        RECT 7.550 3.685 8.250 3.975 ;
        RECT 9.550 3.685 10.250 3.975 ;
        RECT 11.550 3.685 12.250 3.975 ;
        RECT 13.550 3.685 14.250 3.975 ;
        RECT 15.550 3.685 16.250 3.975 ;
        RECT 17.550 3.685 18.250 3.975 ;
        RECT 19.550 3.685 20.250 3.975 ;
        RECT 21.550 3.685 22.250 3.975 ;
        RECT 23.550 3.685 24.250 3.975 ;
        RECT 25.550 3.685 26.250 3.975 ;
        RECT 27.550 3.685 28.250 3.975 ;
        RECT 29.550 3.685 30.250 3.975 ;
        RECT 31.550 3.685 32.250 3.975 ;
        RECT 33.550 3.685 34.250 3.975 ;
        RECT 35.550 3.685 36.250 3.975 ;
        RECT 37.550 3.685 38.250 3.975 ;
        RECT 39.550 3.685 40.250 3.975 ;
        RECT 41.550 3.685 42.250 3.975 ;
        RECT 43.550 3.685 44.250 3.975 ;
        RECT 45.550 3.685 46.250 3.975 ;
        RECT 47.550 3.685 48.250 3.975 ;
        RECT 49.550 3.685 50.250 3.975 ;
        RECT 51.550 3.685 52.250 3.975 ;
        RECT 53.550 3.685 54.250 3.975 ;
        RECT 55.550 3.685 56.250 3.975 ;
        RECT 57.550 3.685 58.250 3.975 ;
        RECT 59.550 3.685 60.250 3.975 ;
        RECT 61.550 3.685 62.250 3.975 ;
        RECT 63.550 3.685 64.250 3.975 ;
        RECT 65.550 3.685 66.250 3.975 ;
        RECT 67.550 3.685 68.250 3.975 ;
        RECT 69.550 3.685 70.250 3.975 ;
        RECT 71.550 3.685 72.250 3.975 ;
        RECT 73.550 3.685 74.250 3.975 ;
        RECT 75.550 3.685 76.250 3.975 ;
        RECT 77.550 3.685 78.250 3.975 ;
        RECT 79.550 3.685 80.250 3.975 ;
        RECT 81.550 3.685 82.250 3.975 ;
        RECT 83.550 3.685 84.250 3.975 ;
        RECT 85.550 3.685 86.250 3.975 ;
        RECT 87.550 3.685 88.250 3.975 ;
        RECT 89.550 3.685 90.250 3.975 ;
        RECT 91.550 3.685 92.250 3.975 ;
        RECT 93.550 3.685 94.250 3.975 ;
        RECT 95.550 3.685 96.250 3.975 ;
        RECT 97.550 3.685 98.250 3.975 ;
        RECT 99.550 3.685 100.250 3.975 ;
        RECT 101.550 3.685 102.250 3.975 ;
        RECT 103.550 3.685 104.250 3.975 ;
        RECT 105.550 3.685 106.250 3.975 ;
        RECT 107.550 3.685 108.250 3.975 ;
        RECT 109.550 3.685 110.250 3.975 ;
        RECT 111.550 3.685 112.250 3.975 ;
        RECT 113.550 3.685 114.250 3.975 ;
        RECT 115.550 3.685 116.250 3.975 ;
        RECT 117.550 3.685 118.250 3.975 ;
        RECT 119.550 3.685 120.250 3.975 ;
        RECT 121.550 3.685 122.250 3.975 ;
        RECT 123.550 3.685 124.250 3.975 ;
        RECT 125.550 3.685 126.250 3.975 ;
        RECT 127.550 3.685 128.250 3.975 ;
        RECT 129.550 3.685 130.250 3.975 ;
        RECT 131.550 3.685 132.250 3.975 ;
      LAYER Metal3 ;
        RECT 0.000 22.030 133.800 23.760 ;
        RECT 0.000 18.800 133.800 20.530 ;
        RECT 0.000 5.660 133.800 7.390 ;
        RECT 0.000 2.430 133.800 4.160 ;
    END
  END VDD
  PIN VcascP[1]
    ANTENNAGATEAREA 1.755000 ;
    ANTENNADIFFAREA 10.710000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.000 19.600 0.490 19.900 ;
        RECT 0.340 19.520 0.490 19.600 ;
        RECT 133.310 19.600 133.800 19.900 ;
        RECT 133.310 19.520 133.460 19.600 ;
        RECT 0.340 13.490 0.490 13.670 ;
        RECT 133.310 13.490 133.460 13.670 ;
      LAYER Metal1 ;
        RECT 2.260 21.130 2.560 21.430 ;
        RECT 4.260 21.130 4.560 21.430 ;
        RECT 6.260 21.130 6.560 21.430 ;
        RECT 8.260 21.130 8.560 21.430 ;
        RECT 10.260 21.130 10.560 21.430 ;
        RECT 12.260 21.130 12.560 21.430 ;
        RECT 14.260 21.130 14.560 21.430 ;
        RECT 16.260 21.130 16.560 21.430 ;
        RECT 18.260 21.130 18.560 21.430 ;
        RECT 20.260 21.130 20.560 21.430 ;
        RECT 22.260 21.130 22.560 21.430 ;
        RECT 24.260 21.130 24.560 21.430 ;
        RECT 26.260 21.130 26.560 21.430 ;
        RECT 28.260 21.130 28.560 21.430 ;
        RECT 30.260 21.130 30.560 21.430 ;
        RECT 32.260 21.130 32.560 21.430 ;
        RECT 34.260 21.130 34.560 21.430 ;
        RECT 36.260 21.130 36.560 21.430 ;
        RECT 38.260 21.130 38.560 21.430 ;
        RECT 40.260 21.130 40.560 21.430 ;
        RECT 42.260 21.130 42.560 21.430 ;
        RECT 44.260 21.130 44.560 21.430 ;
        RECT 46.260 21.130 46.560 21.430 ;
        RECT 48.260 21.130 48.560 21.430 ;
        RECT 50.260 21.130 50.560 21.430 ;
        RECT 52.260 21.130 52.560 21.430 ;
        RECT 54.260 21.130 54.560 21.430 ;
        RECT 56.260 21.130 56.560 21.430 ;
        RECT 58.260 21.130 58.560 21.430 ;
        RECT 60.260 21.130 60.560 21.430 ;
        RECT 62.260 21.130 62.560 21.430 ;
        RECT 64.260 21.130 64.560 21.430 ;
        RECT 66.260 21.130 66.560 21.430 ;
        RECT 68.260 21.130 68.560 21.430 ;
        RECT 70.260 21.130 70.560 21.430 ;
        RECT 72.260 21.130 72.560 21.430 ;
        RECT 74.260 21.130 74.560 21.430 ;
        RECT 76.260 21.130 76.560 21.430 ;
        RECT 78.260 21.130 78.560 21.430 ;
        RECT 80.260 21.130 80.560 21.430 ;
        RECT 82.260 21.130 82.560 21.430 ;
        RECT 84.260 21.130 84.560 21.430 ;
        RECT 86.260 21.130 86.560 21.430 ;
        RECT 88.260 21.130 88.560 21.430 ;
        RECT 90.260 21.130 90.560 21.430 ;
        RECT 92.260 21.130 92.560 21.430 ;
        RECT 94.260 21.130 94.560 21.430 ;
        RECT 96.260 21.130 96.560 21.430 ;
        RECT 98.260 21.130 98.560 21.430 ;
        RECT 100.260 21.130 100.560 21.430 ;
        RECT 102.260 21.130 102.560 21.430 ;
        RECT 104.260 21.130 104.560 21.430 ;
        RECT 106.260 21.130 106.560 21.430 ;
        RECT 108.260 21.130 108.560 21.430 ;
        RECT 110.260 21.130 110.560 21.430 ;
        RECT 112.260 21.130 112.560 21.430 ;
        RECT 114.260 21.130 114.560 21.430 ;
        RECT 116.260 21.130 116.560 21.430 ;
        RECT 118.260 21.130 118.560 21.430 ;
        RECT 120.260 21.130 120.560 21.430 ;
        RECT 122.260 21.130 122.560 21.430 ;
        RECT 124.260 21.130 124.560 21.430 ;
        RECT 126.260 21.130 126.560 21.430 ;
        RECT 128.260 21.130 128.560 21.430 ;
        RECT 130.260 21.130 130.560 21.430 ;
        RECT 132.260 21.130 132.560 21.430 ;
        RECT 0.005 13.670 0.295 19.880 ;
        RECT 133.505 13.670 133.795 19.880 ;
      LAYER Metal2 ;
        RECT 0.005 13.830 0.295 21.630 ;
        RECT 2.265 21.075 2.745 21.425 ;
        RECT 4.265 21.075 4.745 21.425 ;
        RECT 6.265 21.075 6.745 21.425 ;
        RECT 8.265 21.075 8.745 21.425 ;
        RECT 10.265 21.075 10.745 21.425 ;
        RECT 12.265 21.075 12.745 21.425 ;
        RECT 14.265 21.075 14.745 21.425 ;
        RECT 16.265 21.075 16.745 21.425 ;
        RECT 18.265 21.075 18.745 21.425 ;
        RECT 20.265 21.075 20.745 21.425 ;
        RECT 22.265 21.075 22.745 21.425 ;
        RECT 24.265 21.075 24.745 21.425 ;
        RECT 26.265 21.075 26.745 21.425 ;
        RECT 28.265 21.075 28.745 21.425 ;
        RECT 30.265 21.075 30.745 21.425 ;
        RECT 32.265 21.075 32.745 21.425 ;
        RECT 34.265 21.075 34.745 21.425 ;
        RECT 36.265 21.075 36.745 21.425 ;
        RECT 38.265 21.075 38.745 21.425 ;
        RECT 40.265 21.075 40.745 21.425 ;
        RECT 42.265 21.075 42.745 21.425 ;
        RECT 44.265 21.075 44.745 21.425 ;
        RECT 46.265 21.075 46.745 21.425 ;
        RECT 48.265 21.075 48.745 21.425 ;
        RECT 50.265 21.075 50.745 21.425 ;
        RECT 52.265 21.075 52.745 21.425 ;
        RECT 54.265 21.075 54.745 21.425 ;
        RECT 56.265 21.075 56.745 21.425 ;
        RECT 58.265 21.075 58.745 21.425 ;
        RECT 60.265 21.075 60.745 21.425 ;
        RECT 62.265 21.075 62.745 21.425 ;
        RECT 64.265 21.075 64.745 21.425 ;
        RECT 66.265 21.075 66.745 21.425 ;
        RECT 68.265 21.075 68.745 21.425 ;
        RECT 70.265 21.075 70.745 21.425 ;
        RECT 72.265 21.075 72.745 21.425 ;
        RECT 74.265 21.075 74.745 21.425 ;
        RECT 76.265 21.075 76.745 21.425 ;
        RECT 78.265 21.075 78.745 21.425 ;
        RECT 80.265 21.075 80.745 21.425 ;
        RECT 82.265 21.075 82.745 21.425 ;
        RECT 84.265 21.075 84.745 21.425 ;
        RECT 86.265 21.075 86.745 21.425 ;
        RECT 88.265 21.075 88.745 21.425 ;
        RECT 90.265 21.075 90.745 21.425 ;
        RECT 92.265 21.075 92.745 21.425 ;
        RECT 94.265 21.075 94.745 21.425 ;
        RECT 96.265 21.075 96.745 21.425 ;
        RECT 98.265 21.075 98.745 21.425 ;
        RECT 100.265 21.075 100.745 21.425 ;
        RECT 102.265 21.075 102.745 21.425 ;
        RECT 104.265 21.075 104.745 21.425 ;
        RECT 106.265 21.075 106.745 21.425 ;
        RECT 108.265 21.075 108.745 21.425 ;
        RECT 110.265 21.075 110.745 21.425 ;
        RECT 112.265 21.075 112.745 21.425 ;
        RECT 114.265 21.075 114.745 21.425 ;
        RECT 116.265 21.075 116.745 21.425 ;
        RECT 118.265 21.075 118.745 21.425 ;
        RECT 120.265 21.075 120.745 21.425 ;
        RECT 122.265 21.075 122.745 21.425 ;
        RECT 124.265 21.075 124.745 21.425 ;
        RECT 126.265 21.075 126.745 21.425 ;
        RECT 128.265 21.075 128.745 21.425 ;
        RECT 130.265 21.075 130.745 21.425 ;
        RECT 132.265 21.075 132.745 21.425 ;
        RECT 133.505 13.830 133.795 21.630 ;
      LAYER Metal3 ;
        RECT 0.000 20.930 133.800 21.630 ;
    END
  END VcascP[1]
  PIN VcascP[0]
    ANTENNAGATEAREA 1.755000 ;
    ANTENNADIFFAREA 10.710000 ;
    PORT
      LAYER GatPoly ;
        RECT 0.340 12.520 0.490 12.700 ;
        RECT 133.310 12.520 133.460 12.700 ;
        RECT 0.340 6.590 0.490 6.670 ;
        RECT 0.000 6.290 0.490 6.590 ;
        RECT 133.310 6.590 133.460 6.670 ;
        RECT 133.310 6.290 133.800 6.590 ;
      LAYER Metal1 ;
        RECT 0.005 6.310 0.295 12.520 ;
        RECT 133.505 6.310 133.795 12.520 ;
        RECT 1.240 4.760 1.540 5.060 ;
        RECT 3.240 4.760 3.540 5.060 ;
        RECT 5.240 4.760 5.540 5.060 ;
        RECT 7.240 4.760 7.540 5.060 ;
        RECT 9.240 4.760 9.540 5.060 ;
        RECT 11.240 4.760 11.540 5.060 ;
        RECT 13.240 4.760 13.540 5.060 ;
        RECT 15.240 4.760 15.540 5.060 ;
        RECT 17.240 4.760 17.540 5.060 ;
        RECT 19.240 4.760 19.540 5.060 ;
        RECT 21.240 4.760 21.540 5.060 ;
        RECT 23.240 4.760 23.540 5.060 ;
        RECT 25.240 4.760 25.540 5.060 ;
        RECT 27.240 4.760 27.540 5.060 ;
        RECT 29.240 4.760 29.540 5.060 ;
        RECT 31.240 4.760 31.540 5.060 ;
        RECT 33.240 4.760 33.540 5.060 ;
        RECT 35.240 4.760 35.540 5.060 ;
        RECT 37.240 4.760 37.540 5.060 ;
        RECT 39.240 4.760 39.540 5.060 ;
        RECT 41.240 4.760 41.540 5.060 ;
        RECT 43.240 4.760 43.540 5.060 ;
        RECT 45.240 4.760 45.540 5.060 ;
        RECT 47.240 4.760 47.540 5.060 ;
        RECT 49.240 4.760 49.540 5.060 ;
        RECT 51.240 4.760 51.540 5.060 ;
        RECT 53.240 4.760 53.540 5.060 ;
        RECT 55.240 4.760 55.540 5.060 ;
        RECT 57.240 4.760 57.540 5.060 ;
        RECT 59.240 4.760 59.540 5.060 ;
        RECT 61.240 4.760 61.540 5.060 ;
        RECT 63.240 4.760 63.540 5.060 ;
        RECT 65.240 4.760 65.540 5.060 ;
        RECT 67.240 4.760 67.540 5.060 ;
        RECT 69.240 4.760 69.540 5.060 ;
        RECT 71.240 4.760 71.540 5.060 ;
        RECT 73.240 4.760 73.540 5.060 ;
        RECT 75.240 4.760 75.540 5.060 ;
        RECT 77.240 4.760 77.540 5.060 ;
        RECT 79.240 4.760 79.540 5.060 ;
        RECT 81.240 4.760 81.540 5.060 ;
        RECT 83.240 4.760 83.540 5.060 ;
        RECT 85.240 4.760 85.540 5.060 ;
        RECT 87.240 4.760 87.540 5.060 ;
        RECT 89.240 4.760 89.540 5.060 ;
        RECT 91.240 4.760 91.540 5.060 ;
        RECT 93.240 4.760 93.540 5.060 ;
        RECT 95.240 4.760 95.540 5.060 ;
        RECT 97.240 4.760 97.540 5.060 ;
        RECT 99.240 4.760 99.540 5.060 ;
        RECT 101.240 4.760 101.540 5.060 ;
        RECT 103.240 4.760 103.540 5.060 ;
        RECT 105.240 4.760 105.540 5.060 ;
        RECT 107.240 4.760 107.540 5.060 ;
        RECT 109.240 4.760 109.540 5.060 ;
        RECT 111.240 4.760 111.540 5.060 ;
        RECT 113.240 4.760 113.540 5.060 ;
        RECT 115.240 4.760 115.540 5.060 ;
        RECT 117.240 4.760 117.540 5.060 ;
        RECT 119.240 4.760 119.540 5.060 ;
        RECT 121.240 4.760 121.540 5.060 ;
        RECT 123.240 4.760 123.540 5.060 ;
        RECT 125.240 4.760 125.540 5.060 ;
        RECT 127.240 4.760 127.540 5.060 ;
        RECT 129.240 4.760 129.540 5.060 ;
        RECT 131.240 4.760 131.540 5.060 ;
      LAYER Metal2 ;
        RECT 0.005 4.560 0.295 12.360 ;
        RECT 1.055 4.765 1.535 5.115 ;
        RECT 3.055 4.765 3.535 5.115 ;
        RECT 5.055 4.765 5.535 5.115 ;
        RECT 7.055 4.765 7.535 5.115 ;
        RECT 9.055 4.765 9.535 5.115 ;
        RECT 11.055 4.765 11.535 5.115 ;
        RECT 13.055 4.765 13.535 5.115 ;
        RECT 15.055 4.765 15.535 5.115 ;
        RECT 17.055 4.765 17.535 5.115 ;
        RECT 19.055 4.765 19.535 5.115 ;
        RECT 21.055 4.765 21.535 5.115 ;
        RECT 23.055 4.765 23.535 5.115 ;
        RECT 25.055 4.765 25.535 5.115 ;
        RECT 27.055 4.765 27.535 5.115 ;
        RECT 29.055 4.765 29.535 5.115 ;
        RECT 31.055 4.765 31.535 5.115 ;
        RECT 33.055 4.765 33.535 5.115 ;
        RECT 35.055 4.765 35.535 5.115 ;
        RECT 37.055 4.765 37.535 5.115 ;
        RECT 39.055 4.765 39.535 5.115 ;
        RECT 41.055 4.765 41.535 5.115 ;
        RECT 43.055 4.765 43.535 5.115 ;
        RECT 45.055 4.765 45.535 5.115 ;
        RECT 47.055 4.765 47.535 5.115 ;
        RECT 49.055 4.765 49.535 5.115 ;
        RECT 51.055 4.765 51.535 5.115 ;
        RECT 53.055 4.765 53.535 5.115 ;
        RECT 55.055 4.765 55.535 5.115 ;
        RECT 57.055 4.765 57.535 5.115 ;
        RECT 59.055 4.765 59.535 5.115 ;
        RECT 61.055 4.765 61.535 5.115 ;
        RECT 63.055 4.765 63.535 5.115 ;
        RECT 65.055 4.765 65.535 5.115 ;
        RECT 67.055 4.765 67.535 5.115 ;
        RECT 69.055 4.765 69.535 5.115 ;
        RECT 71.055 4.765 71.535 5.115 ;
        RECT 73.055 4.765 73.535 5.115 ;
        RECT 75.055 4.765 75.535 5.115 ;
        RECT 77.055 4.765 77.535 5.115 ;
        RECT 79.055 4.765 79.535 5.115 ;
        RECT 81.055 4.765 81.535 5.115 ;
        RECT 83.055 4.765 83.535 5.115 ;
        RECT 85.055 4.765 85.535 5.115 ;
        RECT 87.055 4.765 87.535 5.115 ;
        RECT 89.055 4.765 89.535 5.115 ;
        RECT 91.055 4.765 91.535 5.115 ;
        RECT 93.055 4.765 93.535 5.115 ;
        RECT 95.055 4.765 95.535 5.115 ;
        RECT 97.055 4.765 97.535 5.115 ;
        RECT 99.055 4.765 99.535 5.115 ;
        RECT 101.055 4.765 101.535 5.115 ;
        RECT 103.055 4.765 103.535 5.115 ;
        RECT 105.055 4.765 105.535 5.115 ;
        RECT 107.055 4.765 107.535 5.115 ;
        RECT 109.055 4.765 109.535 5.115 ;
        RECT 111.055 4.765 111.535 5.115 ;
        RECT 113.055 4.765 113.535 5.115 ;
        RECT 115.055 4.765 115.535 5.115 ;
        RECT 117.055 4.765 117.535 5.115 ;
        RECT 119.055 4.765 119.535 5.115 ;
        RECT 121.055 4.765 121.535 5.115 ;
        RECT 123.055 4.765 123.535 5.115 ;
        RECT 125.055 4.765 125.535 5.115 ;
        RECT 127.055 4.765 127.535 5.115 ;
        RECT 129.055 4.765 129.535 5.115 ;
        RECT 131.055 4.765 131.535 5.115 ;
        RECT 133.505 4.560 133.795 12.360 ;
      LAYER Metal3 ;
        RECT 0.000 4.560 133.800 5.260 ;
    END
  END VcascP[0]
  OBS
      LAYER GatPoly ;
        RECT 1.235 24.860 1.755 25.040 ;
        RECT 2.045 24.860 2.565 25.040 ;
        RECT 3.235 24.860 3.755 25.040 ;
        RECT 4.045 24.860 4.565 25.040 ;
        RECT 5.235 24.860 5.755 25.040 ;
        RECT 6.045 24.860 6.565 25.040 ;
        RECT 7.235 24.860 7.755 25.040 ;
        RECT 8.045 24.860 8.565 25.040 ;
        RECT 9.235 24.860 9.755 25.040 ;
        RECT 10.045 24.860 10.565 25.040 ;
        RECT 11.235 24.860 11.755 25.040 ;
        RECT 12.045 24.860 12.565 25.040 ;
        RECT 13.235 24.860 13.755 25.040 ;
        RECT 14.045 24.860 14.565 25.040 ;
        RECT 15.235 24.860 15.755 25.040 ;
        RECT 16.045 24.860 16.565 25.040 ;
        RECT 17.235 24.860 17.755 25.040 ;
        RECT 18.045 24.860 18.565 25.040 ;
        RECT 19.235 24.860 19.755 25.040 ;
        RECT 20.045 24.860 20.565 25.040 ;
        RECT 21.235 24.860 21.755 25.040 ;
        RECT 22.045 24.860 22.565 25.040 ;
        RECT 23.235 24.860 23.755 25.040 ;
        RECT 24.045 24.860 24.565 25.040 ;
        RECT 25.235 24.860 25.755 25.040 ;
        RECT 26.045 24.860 26.565 25.040 ;
        RECT 27.235 24.860 27.755 25.040 ;
        RECT 28.045 24.860 28.565 25.040 ;
        RECT 29.235 24.860 29.755 25.040 ;
        RECT 30.045 24.860 30.565 25.040 ;
        RECT 31.235 24.860 31.755 25.040 ;
        RECT 32.045 24.860 32.565 25.040 ;
        RECT 33.235 24.860 33.755 25.040 ;
        RECT 34.045 24.860 34.565 25.040 ;
        RECT 35.235 24.860 35.755 25.040 ;
        RECT 36.045 24.860 36.565 25.040 ;
        RECT 37.235 24.860 37.755 25.040 ;
        RECT 38.045 24.860 38.565 25.040 ;
        RECT 39.235 24.860 39.755 25.040 ;
        RECT 40.045 24.860 40.565 25.040 ;
        RECT 41.235 24.860 41.755 25.040 ;
        RECT 42.045 24.860 42.565 25.040 ;
        RECT 43.235 24.860 43.755 25.040 ;
        RECT 44.045 24.860 44.565 25.040 ;
        RECT 45.235 24.860 45.755 25.040 ;
        RECT 46.045 24.860 46.565 25.040 ;
        RECT 47.235 24.860 47.755 25.040 ;
        RECT 48.045 24.860 48.565 25.040 ;
        RECT 49.235 24.860 49.755 25.040 ;
        RECT 50.045 24.860 50.565 25.040 ;
        RECT 51.235 24.860 51.755 25.040 ;
        RECT 52.045 24.860 52.565 25.040 ;
        RECT 53.235 24.860 53.755 25.040 ;
        RECT 54.045 24.860 54.565 25.040 ;
        RECT 55.235 24.860 55.755 25.040 ;
        RECT 56.045 24.860 56.565 25.040 ;
        RECT 57.235 24.860 57.755 25.040 ;
        RECT 58.045 24.860 58.565 25.040 ;
        RECT 59.235 24.860 59.755 25.040 ;
        RECT 60.045 24.860 60.565 25.040 ;
        RECT 61.235 24.860 61.755 25.040 ;
        RECT 62.045 24.860 62.565 25.040 ;
        RECT 63.235 24.860 63.755 25.040 ;
        RECT 64.045 24.860 64.565 25.040 ;
        RECT 65.235 24.860 65.755 25.040 ;
        RECT 66.045 24.860 66.565 25.040 ;
        RECT 67.235 24.860 67.755 25.040 ;
        RECT 68.045 24.860 68.565 25.040 ;
        RECT 69.235 24.860 69.755 25.040 ;
        RECT 70.045 24.860 70.565 25.040 ;
        RECT 71.235 24.860 71.755 25.040 ;
        RECT 72.045 24.860 72.565 25.040 ;
        RECT 73.235 24.860 73.755 25.040 ;
        RECT 74.045 24.860 74.565 25.040 ;
        RECT 75.235 24.860 75.755 25.040 ;
        RECT 76.045 24.860 76.565 25.040 ;
        RECT 77.235 24.860 77.755 25.040 ;
        RECT 78.045 24.860 78.565 25.040 ;
        RECT 79.235 24.860 79.755 25.040 ;
        RECT 80.045 24.860 80.565 25.040 ;
        RECT 81.235 24.860 81.755 25.040 ;
        RECT 82.045 24.860 82.565 25.040 ;
        RECT 83.235 24.860 83.755 25.040 ;
        RECT 84.045 24.860 84.565 25.040 ;
        RECT 85.235 24.860 85.755 25.040 ;
        RECT 86.045 24.860 86.565 25.040 ;
        RECT 87.235 24.860 87.755 25.040 ;
        RECT 88.045 24.860 88.565 25.040 ;
        RECT 89.235 24.860 89.755 25.040 ;
        RECT 90.045 24.860 90.565 25.040 ;
        RECT 91.235 24.860 91.755 25.040 ;
        RECT 92.045 24.860 92.565 25.040 ;
        RECT 93.235 24.860 93.755 25.040 ;
        RECT 94.045 24.860 94.565 25.040 ;
        RECT 95.235 24.860 95.755 25.040 ;
        RECT 96.045 24.860 96.565 25.040 ;
        RECT 97.235 24.860 97.755 25.040 ;
        RECT 98.045 24.860 98.565 25.040 ;
        RECT 99.235 24.860 99.755 25.040 ;
        RECT 100.045 24.860 100.565 25.040 ;
        RECT 101.235 24.860 101.755 25.040 ;
        RECT 102.045 24.860 102.565 25.040 ;
        RECT 103.235 24.860 103.755 25.040 ;
        RECT 104.045 24.860 104.565 25.040 ;
        RECT 105.235 24.860 105.755 25.040 ;
        RECT 106.045 24.860 106.565 25.040 ;
        RECT 107.235 24.860 107.755 25.040 ;
        RECT 108.045 24.860 108.565 25.040 ;
        RECT 109.235 24.860 109.755 25.040 ;
        RECT 110.045 24.860 110.565 25.040 ;
        RECT 111.235 24.860 111.755 25.040 ;
        RECT 112.045 24.860 112.565 25.040 ;
        RECT 113.235 24.860 113.755 25.040 ;
        RECT 114.045 24.860 114.565 25.040 ;
        RECT 115.235 24.860 115.755 25.040 ;
        RECT 116.045 24.860 116.565 25.040 ;
        RECT 117.235 24.860 117.755 25.040 ;
        RECT 118.045 24.860 118.565 25.040 ;
        RECT 119.235 24.860 119.755 25.040 ;
        RECT 120.045 24.860 120.565 25.040 ;
        RECT 121.235 24.860 121.755 25.040 ;
        RECT 122.045 24.860 122.565 25.040 ;
        RECT 123.235 24.860 123.755 25.040 ;
        RECT 124.045 24.860 124.565 25.040 ;
        RECT 125.235 24.860 125.755 25.040 ;
        RECT 126.045 24.860 126.565 25.040 ;
        RECT 127.235 24.860 127.755 25.040 ;
        RECT 128.045 24.860 128.565 25.040 ;
        RECT 129.235 24.860 129.755 25.040 ;
        RECT 130.045 24.860 130.565 25.040 ;
        RECT 131.235 24.860 131.755 25.040 ;
        RECT 132.045 24.860 132.565 25.040 ;
        RECT 1.235 24.530 1.755 24.710 ;
        RECT 1.455 24.340 1.755 24.530 ;
        RECT 2.045 24.530 2.565 24.710 ;
        RECT 3.235 24.530 3.755 24.710 ;
        RECT 2.045 24.160 2.345 24.530 ;
        RECT 3.455 24.340 3.755 24.530 ;
        RECT 4.045 24.530 4.565 24.710 ;
        RECT 5.235 24.530 5.755 24.710 ;
        RECT 4.045 24.160 4.345 24.530 ;
        RECT 5.455 24.340 5.755 24.530 ;
        RECT 6.045 24.530 6.565 24.710 ;
        RECT 7.235 24.530 7.755 24.710 ;
        RECT 6.045 24.160 6.345 24.530 ;
        RECT 7.455 24.340 7.755 24.530 ;
        RECT 8.045 24.530 8.565 24.710 ;
        RECT 9.235 24.530 9.755 24.710 ;
        RECT 8.045 24.160 8.345 24.530 ;
        RECT 9.455 24.340 9.755 24.530 ;
        RECT 10.045 24.530 10.565 24.710 ;
        RECT 11.235 24.530 11.755 24.710 ;
        RECT 10.045 24.160 10.345 24.530 ;
        RECT 11.455 24.340 11.755 24.530 ;
        RECT 12.045 24.530 12.565 24.710 ;
        RECT 13.235 24.530 13.755 24.710 ;
        RECT 12.045 24.160 12.345 24.530 ;
        RECT 13.455 24.340 13.755 24.530 ;
        RECT 14.045 24.530 14.565 24.710 ;
        RECT 15.235 24.530 15.755 24.710 ;
        RECT 14.045 24.160 14.345 24.530 ;
        RECT 15.455 24.340 15.755 24.530 ;
        RECT 16.045 24.530 16.565 24.710 ;
        RECT 17.235 24.530 17.755 24.710 ;
        RECT 16.045 24.160 16.345 24.530 ;
        RECT 17.455 24.340 17.755 24.530 ;
        RECT 18.045 24.530 18.565 24.710 ;
        RECT 19.235 24.530 19.755 24.710 ;
        RECT 18.045 24.160 18.345 24.530 ;
        RECT 19.455 24.340 19.755 24.530 ;
        RECT 20.045 24.530 20.565 24.710 ;
        RECT 21.235 24.530 21.755 24.710 ;
        RECT 20.045 24.160 20.345 24.530 ;
        RECT 21.455 24.340 21.755 24.530 ;
        RECT 22.045 24.530 22.565 24.710 ;
        RECT 23.235 24.530 23.755 24.710 ;
        RECT 22.045 24.160 22.345 24.530 ;
        RECT 23.455 24.340 23.755 24.530 ;
        RECT 24.045 24.530 24.565 24.710 ;
        RECT 25.235 24.530 25.755 24.710 ;
        RECT 24.045 24.160 24.345 24.530 ;
        RECT 25.455 24.340 25.755 24.530 ;
        RECT 26.045 24.530 26.565 24.710 ;
        RECT 27.235 24.530 27.755 24.710 ;
        RECT 26.045 24.160 26.345 24.530 ;
        RECT 27.455 24.340 27.755 24.530 ;
        RECT 28.045 24.530 28.565 24.710 ;
        RECT 29.235 24.530 29.755 24.710 ;
        RECT 28.045 24.160 28.345 24.530 ;
        RECT 29.455 24.340 29.755 24.530 ;
        RECT 30.045 24.530 30.565 24.710 ;
        RECT 31.235 24.530 31.755 24.710 ;
        RECT 30.045 24.160 30.345 24.530 ;
        RECT 31.455 24.340 31.755 24.530 ;
        RECT 32.045 24.530 32.565 24.710 ;
        RECT 33.235 24.530 33.755 24.710 ;
        RECT 32.045 24.160 32.345 24.530 ;
        RECT 33.455 24.340 33.755 24.530 ;
        RECT 34.045 24.530 34.565 24.710 ;
        RECT 35.235 24.530 35.755 24.710 ;
        RECT 34.045 24.160 34.345 24.530 ;
        RECT 35.455 24.340 35.755 24.530 ;
        RECT 36.045 24.530 36.565 24.710 ;
        RECT 37.235 24.530 37.755 24.710 ;
        RECT 36.045 24.160 36.345 24.530 ;
        RECT 37.455 24.340 37.755 24.530 ;
        RECT 38.045 24.530 38.565 24.710 ;
        RECT 39.235 24.530 39.755 24.710 ;
        RECT 38.045 24.160 38.345 24.530 ;
        RECT 39.455 24.340 39.755 24.530 ;
        RECT 40.045 24.530 40.565 24.710 ;
        RECT 41.235 24.530 41.755 24.710 ;
        RECT 40.045 24.160 40.345 24.530 ;
        RECT 41.455 24.340 41.755 24.530 ;
        RECT 42.045 24.530 42.565 24.710 ;
        RECT 43.235 24.530 43.755 24.710 ;
        RECT 42.045 24.160 42.345 24.530 ;
        RECT 43.455 24.340 43.755 24.530 ;
        RECT 44.045 24.530 44.565 24.710 ;
        RECT 45.235 24.530 45.755 24.710 ;
        RECT 44.045 24.160 44.345 24.530 ;
        RECT 45.455 24.340 45.755 24.530 ;
        RECT 46.045 24.530 46.565 24.710 ;
        RECT 47.235 24.530 47.755 24.710 ;
        RECT 46.045 24.160 46.345 24.530 ;
        RECT 47.455 24.340 47.755 24.530 ;
        RECT 48.045 24.530 48.565 24.710 ;
        RECT 49.235 24.530 49.755 24.710 ;
        RECT 48.045 24.160 48.345 24.530 ;
        RECT 49.455 24.340 49.755 24.530 ;
        RECT 50.045 24.530 50.565 24.710 ;
        RECT 51.235 24.530 51.755 24.710 ;
        RECT 50.045 24.160 50.345 24.530 ;
        RECT 51.455 24.340 51.755 24.530 ;
        RECT 52.045 24.530 52.565 24.710 ;
        RECT 53.235 24.530 53.755 24.710 ;
        RECT 52.045 24.160 52.345 24.530 ;
        RECT 53.455 24.340 53.755 24.530 ;
        RECT 54.045 24.530 54.565 24.710 ;
        RECT 55.235 24.530 55.755 24.710 ;
        RECT 54.045 24.160 54.345 24.530 ;
        RECT 55.455 24.340 55.755 24.530 ;
        RECT 56.045 24.530 56.565 24.710 ;
        RECT 57.235 24.530 57.755 24.710 ;
        RECT 56.045 24.160 56.345 24.530 ;
        RECT 57.455 24.340 57.755 24.530 ;
        RECT 58.045 24.530 58.565 24.710 ;
        RECT 59.235 24.530 59.755 24.710 ;
        RECT 58.045 24.160 58.345 24.530 ;
        RECT 59.455 24.340 59.755 24.530 ;
        RECT 60.045 24.530 60.565 24.710 ;
        RECT 61.235 24.530 61.755 24.710 ;
        RECT 60.045 24.160 60.345 24.530 ;
        RECT 61.455 24.340 61.755 24.530 ;
        RECT 62.045 24.530 62.565 24.710 ;
        RECT 63.235 24.530 63.755 24.710 ;
        RECT 62.045 24.160 62.345 24.530 ;
        RECT 63.455 24.340 63.755 24.530 ;
        RECT 64.045 24.530 64.565 24.710 ;
        RECT 65.235 24.530 65.755 24.710 ;
        RECT 64.045 24.160 64.345 24.530 ;
        RECT 65.455 24.340 65.755 24.530 ;
        RECT 66.045 24.530 66.565 24.710 ;
        RECT 67.235 24.530 67.755 24.710 ;
        RECT 66.045 24.160 66.345 24.530 ;
        RECT 67.455 24.340 67.755 24.530 ;
        RECT 68.045 24.530 68.565 24.710 ;
        RECT 69.235 24.530 69.755 24.710 ;
        RECT 68.045 24.160 68.345 24.530 ;
        RECT 69.455 24.340 69.755 24.530 ;
        RECT 70.045 24.530 70.565 24.710 ;
        RECT 71.235 24.530 71.755 24.710 ;
        RECT 70.045 24.160 70.345 24.530 ;
        RECT 71.455 24.340 71.755 24.530 ;
        RECT 72.045 24.530 72.565 24.710 ;
        RECT 73.235 24.530 73.755 24.710 ;
        RECT 72.045 24.160 72.345 24.530 ;
        RECT 73.455 24.340 73.755 24.530 ;
        RECT 74.045 24.530 74.565 24.710 ;
        RECT 75.235 24.530 75.755 24.710 ;
        RECT 74.045 24.160 74.345 24.530 ;
        RECT 75.455 24.340 75.755 24.530 ;
        RECT 76.045 24.530 76.565 24.710 ;
        RECT 77.235 24.530 77.755 24.710 ;
        RECT 76.045 24.160 76.345 24.530 ;
        RECT 77.455 24.340 77.755 24.530 ;
        RECT 78.045 24.530 78.565 24.710 ;
        RECT 79.235 24.530 79.755 24.710 ;
        RECT 78.045 24.160 78.345 24.530 ;
        RECT 79.455 24.340 79.755 24.530 ;
        RECT 80.045 24.530 80.565 24.710 ;
        RECT 81.235 24.530 81.755 24.710 ;
        RECT 80.045 24.160 80.345 24.530 ;
        RECT 81.455 24.340 81.755 24.530 ;
        RECT 82.045 24.530 82.565 24.710 ;
        RECT 83.235 24.530 83.755 24.710 ;
        RECT 82.045 24.160 82.345 24.530 ;
        RECT 83.455 24.340 83.755 24.530 ;
        RECT 84.045 24.530 84.565 24.710 ;
        RECT 85.235 24.530 85.755 24.710 ;
        RECT 84.045 24.160 84.345 24.530 ;
        RECT 85.455 24.340 85.755 24.530 ;
        RECT 86.045 24.530 86.565 24.710 ;
        RECT 87.235 24.530 87.755 24.710 ;
        RECT 86.045 24.160 86.345 24.530 ;
        RECT 87.455 24.340 87.755 24.530 ;
        RECT 88.045 24.530 88.565 24.710 ;
        RECT 89.235 24.530 89.755 24.710 ;
        RECT 88.045 24.160 88.345 24.530 ;
        RECT 89.455 24.340 89.755 24.530 ;
        RECT 90.045 24.530 90.565 24.710 ;
        RECT 91.235 24.530 91.755 24.710 ;
        RECT 90.045 24.160 90.345 24.530 ;
        RECT 91.455 24.340 91.755 24.530 ;
        RECT 92.045 24.530 92.565 24.710 ;
        RECT 93.235 24.530 93.755 24.710 ;
        RECT 92.045 24.160 92.345 24.530 ;
        RECT 93.455 24.340 93.755 24.530 ;
        RECT 94.045 24.530 94.565 24.710 ;
        RECT 95.235 24.530 95.755 24.710 ;
        RECT 94.045 24.160 94.345 24.530 ;
        RECT 95.455 24.340 95.755 24.530 ;
        RECT 96.045 24.530 96.565 24.710 ;
        RECT 97.235 24.530 97.755 24.710 ;
        RECT 96.045 24.160 96.345 24.530 ;
        RECT 97.455 24.340 97.755 24.530 ;
        RECT 98.045 24.530 98.565 24.710 ;
        RECT 99.235 24.530 99.755 24.710 ;
        RECT 98.045 24.160 98.345 24.530 ;
        RECT 99.455 24.340 99.755 24.530 ;
        RECT 100.045 24.530 100.565 24.710 ;
        RECT 101.235 24.530 101.755 24.710 ;
        RECT 100.045 24.160 100.345 24.530 ;
        RECT 101.455 24.340 101.755 24.530 ;
        RECT 102.045 24.530 102.565 24.710 ;
        RECT 103.235 24.530 103.755 24.710 ;
        RECT 102.045 24.160 102.345 24.530 ;
        RECT 103.455 24.340 103.755 24.530 ;
        RECT 104.045 24.530 104.565 24.710 ;
        RECT 105.235 24.530 105.755 24.710 ;
        RECT 104.045 24.160 104.345 24.530 ;
        RECT 105.455 24.340 105.755 24.530 ;
        RECT 106.045 24.530 106.565 24.710 ;
        RECT 107.235 24.530 107.755 24.710 ;
        RECT 106.045 24.160 106.345 24.530 ;
        RECT 107.455 24.340 107.755 24.530 ;
        RECT 108.045 24.530 108.565 24.710 ;
        RECT 109.235 24.530 109.755 24.710 ;
        RECT 108.045 24.160 108.345 24.530 ;
        RECT 109.455 24.340 109.755 24.530 ;
        RECT 110.045 24.530 110.565 24.710 ;
        RECT 111.235 24.530 111.755 24.710 ;
        RECT 110.045 24.160 110.345 24.530 ;
        RECT 111.455 24.340 111.755 24.530 ;
        RECT 112.045 24.530 112.565 24.710 ;
        RECT 113.235 24.530 113.755 24.710 ;
        RECT 112.045 24.160 112.345 24.530 ;
        RECT 113.455 24.340 113.755 24.530 ;
        RECT 114.045 24.530 114.565 24.710 ;
        RECT 115.235 24.530 115.755 24.710 ;
        RECT 114.045 24.160 114.345 24.530 ;
        RECT 115.455 24.340 115.755 24.530 ;
        RECT 116.045 24.530 116.565 24.710 ;
        RECT 117.235 24.530 117.755 24.710 ;
        RECT 116.045 24.160 116.345 24.530 ;
        RECT 117.455 24.340 117.755 24.530 ;
        RECT 118.045 24.530 118.565 24.710 ;
        RECT 119.235 24.530 119.755 24.710 ;
        RECT 118.045 24.160 118.345 24.530 ;
        RECT 119.455 24.340 119.755 24.530 ;
        RECT 120.045 24.530 120.565 24.710 ;
        RECT 121.235 24.530 121.755 24.710 ;
        RECT 120.045 24.160 120.345 24.530 ;
        RECT 121.455 24.340 121.755 24.530 ;
        RECT 122.045 24.530 122.565 24.710 ;
        RECT 123.235 24.530 123.755 24.710 ;
        RECT 122.045 24.160 122.345 24.530 ;
        RECT 123.455 24.340 123.755 24.530 ;
        RECT 124.045 24.530 124.565 24.710 ;
        RECT 125.235 24.530 125.755 24.710 ;
        RECT 124.045 24.160 124.345 24.530 ;
        RECT 125.455 24.340 125.755 24.530 ;
        RECT 126.045 24.530 126.565 24.710 ;
        RECT 127.235 24.530 127.755 24.710 ;
        RECT 126.045 24.160 126.345 24.530 ;
        RECT 127.455 24.340 127.755 24.530 ;
        RECT 128.045 24.530 128.565 24.710 ;
        RECT 129.235 24.530 129.755 24.710 ;
        RECT 128.045 24.160 128.345 24.530 ;
        RECT 129.455 24.340 129.755 24.530 ;
        RECT 130.045 24.530 130.565 24.710 ;
        RECT 131.235 24.530 131.755 24.710 ;
        RECT 130.045 24.160 130.345 24.530 ;
        RECT 131.455 24.340 131.755 24.530 ;
        RECT 132.045 24.530 132.565 24.710 ;
        RECT 132.045 24.160 132.345 24.530 ;
        RECT 1.005 23.860 2.345 24.160 ;
        RECT 3.005 23.860 4.345 24.160 ;
        RECT 5.005 23.860 6.345 24.160 ;
        RECT 7.005 23.860 8.345 24.160 ;
        RECT 9.005 23.860 10.345 24.160 ;
        RECT 11.005 23.860 12.345 24.160 ;
        RECT 13.005 23.860 14.345 24.160 ;
        RECT 15.005 23.860 16.345 24.160 ;
        RECT 17.005 23.860 18.345 24.160 ;
        RECT 19.005 23.860 20.345 24.160 ;
        RECT 21.005 23.860 22.345 24.160 ;
        RECT 23.005 23.860 24.345 24.160 ;
        RECT 25.005 23.860 26.345 24.160 ;
        RECT 27.005 23.860 28.345 24.160 ;
        RECT 29.005 23.860 30.345 24.160 ;
        RECT 31.005 23.860 32.345 24.160 ;
        RECT 33.005 23.860 34.345 24.160 ;
        RECT 35.005 23.860 36.345 24.160 ;
        RECT 37.005 23.860 38.345 24.160 ;
        RECT 39.005 23.860 40.345 24.160 ;
        RECT 41.005 23.860 42.345 24.160 ;
        RECT 43.005 23.860 44.345 24.160 ;
        RECT 45.005 23.860 46.345 24.160 ;
        RECT 47.005 23.860 48.345 24.160 ;
        RECT 49.005 23.860 50.345 24.160 ;
        RECT 51.005 23.860 52.345 24.160 ;
        RECT 53.005 23.860 54.345 24.160 ;
        RECT 55.005 23.860 56.345 24.160 ;
        RECT 57.005 23.860 58.345 24.160 ;
        RECT 59.005 23.860 60.345 24.160 ;
        RECT 61.005 23.860 62.345 24.160 ;
        RECT 63.005 23.860 64.345 24.160 ;
        RECT 65.005 23.860 66.345 24.160 ;
        RECT 67.005 23.860 68.345 24.160 ;
        RECT 69.005 23.860 70.345 24.160 ;
        RECT 71.005 23.860 72.345 24.160 ;
        RECT 73.005 23.860 74.345 24.160 ;
        RECT 75.005 23.860 76.345 24.160 ;
        RECT 77.005 23.860 78.345 24.160 ;
        RECT 79.005 23.860 80.345 24.160 ;
        RECT 81.005 23.860 82.345 24.160 ;
        RECT 83.005 23.860 84.345 24.160 ;
        RECT 85.005 23.860 86.345 24.160 ;
        RECT 87.005 23.860 88.345 24.160 ;
        RECT 89.005 23.860 90.345 24.160 ;
        RECT 91.005 23.860 92.345 24.160 ;
        RECT 93.005 23.860 94.345 24.160 ;
        RECT 95.005 23.860 96.345 24.160 ;
        RECT 97.005 23.860 98.345 24.160 ;
        RECT 99.005 23.860 100.345 24.160 ;
        RECT 101.005 23.860 102.345 24.160 ;
        RECT 103.005 23.860 104.345 24.160 ;
        RECT 105.005 23.860 106.345 24.160 ;
        RECT 107.005 23.860 108.345 24.160 ;
        RECT 109.005 23.860 110.345 24.160 ;
        RECT 111.005 23.860 112.345 24.160 ;
        RECT 113.005 23.860 114.345 24.160 ;
        RECT 115.005 23.860 116.345 24.160 ;
        RECT 117.005 23.860 118.345 24.160 ;
        RECT 119.005 23.860 120.345 24.160 ;
        RECT 121.005 23.860 122.345 24.160 ;
        RECT 123.005 23.860 124.345 24.160 ;
        RECT 125.005 23.860 126.345 24.160 ;
        RECT 127.005 23.860 128.345 24.160 ;
        RECT 129.005 23.860 130.345 24.160 ;
        RECT 131.005 23.860 132.345 24.160 ;
        RECT 1.410 21.630 1.710 21.930 ;
        RECT 1.580 21.430 1.710 21.630 ;
        RECT 2.090 21.630 2.390 21.930 ;
        RECT 3.410 21.630 3.710 21.930 ;
        RECT 2.090 21.430 2.220 21.630 ;
        RECT 3.580 21.430 3.710 21.630 ;
        RECT 4.090 21.630 4.390 21.930 ;
        RECT 5.410 21.630 5.710 21.930 ;
        RECT 4.090 21.430 4.220 21.630 ;
        RECT 5.580 21.430 5.710 21.630 ;
        RECT 6.090 21.630 6.390 21.930 ;
        RECT 7.410 21.630 7.710 21.930 ;
        RECT 6.090 21.430 6.220 21.630 ;
        RECT 7.580 21.430 7.710 21.630 ;
        RECT 8.090 21.630 8.390 21.930 ;
        RECT 9.410 21.630 9.710 21.930 ;
        RECT 8.090 21.430 8.220 21.630 ;
        RECT 9.580 21.430 9.710 21.630 ;
        RECT 10.090 21.630 10.390 21.930 ;
        RECT 11.410 21.630 11.710 21.930 ;
        RECT 10.090 21.430 10.220 21.630 ;
        RECT 11.580 21.430 11.710 21.630 ;
        RECT 12.090 21.630 12.390 21.930 ;
        RECT 13.410 21.630 13.710 21.930 ;
        RECT 12.090 21.430 12.220 21.630 ;
        RECT 13.580 21.430 13.710 21.630 ;
        RECT 14.090 21.630 14.390 21.930 ;
        RECT 15.410 21.630 15.710 21.930 ;
        RECT 14.090 21.430 14.220 21.630 ;
        RECT 15.580 21.430 15.710 21.630 ;
        RECT 16.090 21.630 16.390 21.930 ;
        RECT 17.410 21.630 17.710 21.930 ;
        RECT 16.090 21.430 16.220 21.630 ;
        RECT 17.580 21.430 17.710 21.630 ;
        RECT 18.090 21.630 18.390 21.930 ;
        RECT 19.410 21.630 19.710 21.930 ;
        RECT 18.090 21.430 18.220 21.630 ;
        RECT 19.580 21.430 19.710 21.630 ;
        RECT 20.090 21.630 20.390 21.930 ;
        RECT 21.410 21.630 21.710 21.930 ;
        RECT 20.090 21.430 20.220 21.630 ;
        RECT 21.580 21.430 21.710 21.630 ;
        RECT 22.090 21.630 22.390 21.930 ;
        RECT 23.410 21.630 23.710 21.930 ;
        RECT 22.090 21.430 22.220 21.630 ;
        RECT 23.580 21.430 23.710 21.630 ;
        RECT 24.090 21.630 24.390 21.930 ;
        RECT 25.410 21.630 25.710 21.930 ;
        RECT 24.090 21.430 24.220 21.630 ;
        RECT 25.580 21.430 25.710 21.630 ;
        RECT 26.090 21.630 26.390 21.930 ;
        RECT 27.410 21.630 27.710 21.930 ;
        RECT 26.090 21.430 26.220 21.630 ;
        RECT 27.580 21.430 27.710 21.630 ;
        RECT 28.090 21.630 28.390 21.930 ;
        RECT 29.410 21.630 29.710 21.930 ;
        RECT 28.090 21.430 28.220 21.630 ;
        RECT 29.580 21.430 29.710 21.630 ;
        RECT 30.090 21.630 30.390 21.930 ;
        RECT 31.410 21.630 31.710 21.930 ;
        RECT 30.090 21.430 30.220 21.630 ;
        RECT 31.580 21.430 31.710 21.630 ;
        RECT 32.090 21.630 32.390 21.930 ;
        RECT 33.410 21.630 33.710 21.930 ;
        RECT 32.090 21.430 32.220 21.630 ;
        RECT 33.580 21.430 33.710 21.630 ;
        RECT 34.090 21.630 34.390 21.930 ;
        RECT 35.410 21.630 35.710 21.930 ;
        RECT 34.090 21.430 34.220 21.630 ;
        RECT 35.580 21.430 35.710 21.630 ;
        RECT 36.090 21.630 36.390 21.930 ;
        RECT 37.410 21.630 37.710 21.930 ;
        RECT 36.090 21.430 36.220 21.630 ;
        RECT 37.580 21.430 37.710 21.630 ;
        RECT 38.090 21.630 38.390 21.930 ;
        RECT 39.410 21.630 39.710 21.930 ;
        RECT 38.090 21.430 38.220 21.630 ;
        RECT 39.580 21.430 39.710 21.630 ;
        RECT 40.090 21.630 40.390 21.930 ;
        RECT 41.410 21.630 41.710 21.930 ;
        RECT 40.090 21.430 40.220 21.630 ;
        RECT 41.580 21.430 41.710 21.630 ;
        RECT 42.090 21.630 42.390 21.930 ;
        RECT 43.410 21.630 43.710 21.930 ;
        RECT 42.090 21.430 42.220 21.630 ;
        RECT 43.580 21.430 43.710 21.630 ;
        RECT 44.090 21.630 44.390 21.930 ;
        RECT 45.410 21.630 45.710 21.930 ;
        RECT 44.090 21.430 44.220 21.630 ;
        RECT 45.580 21.430 45.710 21.630 ;
        RECT 46.090 21.630 46.390 21.930 ;
        RECT 47.410 21.630 47.710 21.930 ;
        RECT 46.090 21.430 46.220 21.630 ;
        RECT 47.580 21.430 47.710 21.630 ;
        RECT 48.090 21.630 48.390 21.930 ;
        RECT 49.410 21.630 49.710 21.930 ;
        RECT 48.090 21.430 48.220 21.630 ;
        RECT 49.580 21.430 49.710 21.630 ;
        RECT 50.090 21.630 50.390 21.930 ;
        RECT 51.410 21.630 51.710 21.930 ;
        RECT 50.090 21.430 50.220 21.630 ;
        RECT 51.580 21.430 51.710 21.630 ;
        RECT 52.090 21.630 52.390 21.930 ;
        RECT 53.410 21.630 53.710 21.930 ;
        RECT 52.090 21.430 52.220 21.630 ;
        RECT 53.580 21.430 53.710 21.630 ;
        RECT 54.090 21.630 54.390 21.930 ;
        RECT 55.410 21.630 55.710 21.930 ;
        RECT 54.090 21.430 54.220 21.630 ;
        RECT 55.580 21.430 55.710 21.630 ;
        RECT 56.090 21.630 56.390 21.930 ;
        RECT 57.410 21.630 57.710 21.930 ;
        RECT 56.090 21.430 56.220 21.630 ;
        RECT 57.580 21.430 57.710 21.630 ;
        RECT 58.090 21.630 58.390 21.930 ;
        RECT 59.410 21.630 59.710 21.930 ;
        RECT 58.090 21.430 58.220 21.630 ;
        RECT 59.580 21.430 59.710 21.630 ;
        RECT 60.090 21.630 60.390 21.930 ;
        RECT 61.410 21.630 61.710 21.930 ;
        RECT 60.090 21.430 60.220 21.630 ;
        RECT 61.580 21.430 61.710 21.630 ;
        RECT 62.090 21.630 62.390 21.930 ;
        RECT 63.410 21.630 63.710 21.930 ;
        RECT 62.090 21.430 62.220 21.630 ;
        RECT 63.580 21.430 63.710 21.630 ;
        RECT 64.090 21.630 64.390 21.930 ;
        RECT 65.410 21.630 65.710 21.930 ;
        RECT 64.090 21.430 64.220 21.630 ;
        RECT 65.580 21.430 65.710 21.630 ;
        RECT 66.090 21.630 66.390 21.930 ;
        RECT 67.410 21.630 67.710 21.930 ;
        RECT 66.090 21.430 66.220 21.630 ;
        RECT 67.580 21.430 67.710 21.630 ;
        RECT 68.090 21.630 68.390 21.930 ;
        RECT 69.410 21.630 69.710 21.930 ;
        RECT 68.090 21.430 68.220 21.630 ;
        RECT 69.580 21.430 69.710 21.630 ;
        RECT 70.090 21.630 70.390 21.930 ;
        RECT 71.410 21.630 71.710 21.930 ;
        RECT 70.090 21.430 70.220 21.630 ;
        RECT 71.580 21.430 71.710 21.630 ;
        RECT 72.090 21.630 72.390 21.930 ;
        RECT 73.410 21.630 73.710 21.930 ;
        RECT 72.090 21.430 72.220 21.630 ;
        RECT 73.580 21.430 73.710 21.630 ;
        RECT 74.090 21.630 74.390 21.930 ;
        RECT 75.410 21.630 75.710 21.930 ;
        RECT 74.090 21.430 74.220 21.630 ;
        RECT 75.580 21.430 75.710 21.630 ;
        RECT 76.090 21.630 76.390 21.930 ;
        RECT 77.410 21.630 77.710 21.930 ;
        RECT 76.090 21.430 76.220 21.630 ;
        RECT 77.580 21.430 77.710 21.630 ;
        RECT 78.090 21.630 78.390 21.930 ;
        RECT 79.410 21.630 79.710 21.930 ;
        RECT 78.090 21.430 78.220 21.630 ;
        RECT 79.580 21.430 79.710 21.630 ;
        RECT 80.090 21.630 80.390 21.930 ;
        RECT 81.410 21.630 81.710 21.930 ;
        RECT 80.090 21.430 80.220 21.630 ;
        RECT 81.580 21.430 81.710 21.630 ;
        RECT 82.090 21.630 82.390 21.930 ;
        RECT 83.410 21.630 83.710 21.930 ;
        RECT 82.090 21.430 82.220 21.630 ;
        RECT 83.580 21.430 83.710 21.630 ;
        RECT 84.090 21.630 84.390 21.930 ;
        RECT 85.410 21.630 85.710 21.930 ;
        RECT 84.090 21.430 84.220 21.630 ;
        RECT 85.580 21.430 85.710 21.630 ;
        RECT 86.090 21.630 86.390 21.930 ;
        RECT 87.410 21.630 87.710 21.930 ;
        RECT 86.090 21.430 86.220 21.630 ;
        RECT 87.580 21.430 87.710 21.630 ;
        RECT 88.090 21.630 88.390 21.930 ;
        RECT 89.410 21.630 89.710 21.930 ;
        RECT 88.090 21.430 88.220 21.630 ;
        RECT 89.580 21.430 89.710 21.630 ;
        RECT 90.090 21.630 90.390 21.930 ;
        RECT 91.410 21.630 91.710 21.930 ;
        RECT 90.090 21.430 90.220 21.630 ;
        RECT 91.580 21.430 91.710 21.630 ;
        RECT 92.090 21.630 92.390 21.930 ;
        RECT 93.410 21.630 93.710 21.930 ;
        RECT 92.090 21.430 92.220 21.630 ;
        RECT 93.580 21.430 93.710 21.630 ;
        RECT 94.090 21.630 94.390 21.930 ;
        RECT 95.410 21.630 95.710 21.930 ;
        RECT 94.090 21.430 94.220 21.630 ;
        RECT 95.580 21.430 95.710 21.630 ;
        RECT 96.090 21.630 96.390 21.930 ;
        RECT 97.410 21.630 97.710 21.930 ;
        RECT 96.090 21.430 96.220 21.630 ;
        RECT 97.580 21.430 97.710 21.630 ;
        RECT 98.090 21.630 98.390 21.930 ;
        RECT 99.410 21.630 99.710 21.930 ;
        RECT 98.090 21.430 98.220 21.630 ;
        RECT 99.580 21.430 99.710 21.630 ;
        RECT 100.090 21.630 100.390 21.930 ;
        RECT 101.410 21.630 101.710 21.930 ;
        RECT 100.090 21.430 100.220 21.630 ;
        RECT 101.580 21.430 101.710 21.630 ;
        RECT 102.090 21.630 102.390 21.930 ;
        RECT 103.410 21.630 103.710 21.930 ;
        RECT 102.090 21.430 102.220 21.630 ;
        RECT 103.580 21.430 103.710 21.630 ;
        RECT 104.090 21.630 104.390 21.930 ;
        RECT 105.410 21.630 105.710 21.930 ;
        RECT 104.090 21.430 104.220 21.630 ;
        RECT 105.580 21.430 105.710 21.630 ;
        RECT 106.090 21.630 106.390 21.930 ;
        RECT 107.410 21.630 107.710 21.930 ;
        RECT 106.090 21.430 106.220 21.630 ;
        RECT 107.580 21.430 107.710 21.630 ;
        RECT 108.090 21.630 108.390 21.930 ;
        RECT 109.410 21.630 109.710 21.930 ;
        RECT 108.090 21.430 108.220 21.630 ;
        RECT 109.580 21.430 109.710 21.630 ;
        RECT 110.090 21.630 110.390 21.930 ;
        RECT 111.410 21.630 111.710 21.930 ;
        RECT 110.090 21.430 110.220 21.630 ;
        RECT 111.580 21.430 111.710 21.630 ;
        RECT 112.090 21.630 112.390 21.930 ;
        RECT 113.410 21.630 113.710 21.930 ;
        RECT 112.090 21.430 112.220 21.630 ;
        RECT 113.580 21.430 113.710 21.630 ;
        RECT 114.090 21.630 114.390 21.930 ;
        RECT 115.410 21.630 115.710 21.930 ;
        RECT 114.090 21.430 114.220 21.630 ;
        RECT 115.580 21.430 115.710 21.630 ;
        RECT 116.090 21.630 116.390 21.930 ;
        RECT 117.410 21.630 117.710 21.930 ;
        RECT 116.090 21.430 116.220 21.630 ;
        RECT 117.580 21.430 117.710 21.630 ;
        RECT 118.090 21.630 118.390 21.930 ;
        RECT 119.410 21.630 119.710 21.930 ;
        RECT 118.090 21.430 118.220 21.630 ;
        RECT 119.580 21.430 119.710 21.630 ;
        RECT 120.090 21.630 120.390 21.930 ;
        RECT 121.410 21.630 121.710 21.930 ;
        RECT 120.090 21.430 120.220 21.630 ;
        RECT 121.580 21.430 121.710 21.630 ;
        RECT 122.090 21.630 122.390 21.930 ;
        RECT 123.410 21.630 123.710 21.930 ;
        RECT 122.090 21.430 122.220 21.630 ;
        RECT 123.580 21.430 123.710 21.630 ;
        RECT 124.090 21.630 124.390 21.930 ;
        RECT 125.410 21.630 125.710 21.930 ;
        RECT 124.090 21.430 124.220 21.630 ;
        RECT 125.580 21.430 125.710 21.630 ;
        RECT 126.090 21.630 126.390 21.930 ;
        RECT 127.410 21.630 127.710 21.930 ;
        RECT 126.090 21.430 126.220 21.630 ;
        RECT 127.580 21.430 127.710 21.630 ;
        RECT 128.090 21.630 128.390 21.930 ;
        RECT 129.410 21.630 129.710 21.930 ;
        RECT 128.090 21.430 128.220 21.630 ;
        RECT 129.580 21.430 129.710 21.630 ;
        RECT 130.090 21.630 130.390 21.930 ;
        RECT 131.410 21.630 131.710 21.930 ;
        RECT 130.090 21.430 130.220 21.630 ;
        RECT 131.580 21.430 131.710 21.630 ;
        RECT 132.090 21.630 132.390 21.930 ;
        RECT 132.090 21.430 132.220 21.630 ;
        RECT 1.580 20.950 1.710 21.130 ;
        RECT 2.090 20.950 2.220 21.130 ;
        RECT 3.580 20.950 3.710 21.130 ;
        RECT 4.090 20.950 4.220 21.130 ;
        RECT 5.580 20.950 5.710 21.130 ;
        RECT 6.090 20.950 6.220 21.130 ;
        RECT 7.580 20.950 7.710 21.130 ;
        RECT 8.090 20.950 8.220 21.130 ;
        RECT 9.580 20.950 9.710 21.130 ;
        RECT 10.090 20.950 10.220 21.130 ;
        RECT 11.580 20.950 11.710 21.130 ;
        RECT 12.090 20.950 12.220 21.130 ;
        RECT 13.580 20.950 13.710 21.130 ;
        RECT 14.090 20.950 14.220 21.130 ;
        RECT 15.580 20.950 15.710 21.130 ;
        RECT 16.090 20.950 16.220 21.130 ;
        RECT 17.580 20.950 17.710 21.130 ;
        RECT 18.090 20.950 18.220 21.130 ;
        RECT 19.580 20.950 19.710 21.130 ;
        RECT 20.090 20.950 20.220 21.130 ;
        RECT 21.580 20.950 21.710 21.130 ;
        RECT 22.090 20.950 22.220 21.130 ;
        RECT 23.580 20.950 23.710 21.130 ;
        RECT 24.090 20.950 24.220 21.130 ;
        RECT 25.580 20.950 25.710 21.130 ;
        RECT 26.090 20.950 26.220 21.130 ;
        RECT 27.580 20.950 27.710 21.130 ;
        RECT 28.090 20.950 28.220 21.130 ;
        RECT 29.580 20.950 29.710 21.130 ;
        RECT 30.090 20.950 30.220 21.130 ;
        RECT 31.580 20.950 31.710 21.130 ;
        RECT 32.090 20.950 32.220 21.130 ;
        RECT 33.580 20.950 33.710 21.130 ;
        RECT 34.090 20.950 34.220 21.130 ;
        RECT 35.580 20.950 35.710 21.130 ;
        RECT 36.090 20.950 36.220 21.130 ;
        RECT 37.580 20.950 37.710 21.130 ;
        RECT 38.090 20.950 38.220 21.130 ;
        RECT 39.580 20.950 39.710 21.130 ;
        RECT 40.090 20.950 40.220 21.130 ;
        RECT 41.580 20.950 41.710 21.130 ;
        RECT 42.090 20.950 42.220 21.130 ;
        RECT 43.580 20.950 43.710 21.130 ;
        RECT 44.090 20.950 44.220 21.130 ;
        RECT 45.580 20.950 45.710 21.130 ;
        RECT 46.090 20.950 46.220 21.130 ;
        RECT 47.580 20.950 47.710 21.130 ;
        RECT 48.090 20.950 48.220 21.130 ;
        RECT 49.580 20.950 49.710 21.130 ;
        RECT 50.090 20.950 50.220 21.130 ;
        RECT 51.580 20.950 51.710 21.130 ;
        RECT 52.090 20.950 52.220 21.130 ;
        RECT 53.580 20.950 53.710 21.130 ;
        RECT 54.090 20.950 54.220 21.130 ;
        RECT 55.580 20.950 55.710 21.130 ;
        RECT 56.090 20.950 56.220 21.130 ;
        RECT 57.580 20.950 57.710 21.130 ;
        RECT 58.090 20.950 58.220 21.130 ;
        RECT 59.580 20.950 59.710 21.130 ;
        RECT 60.090 20.950 60.220 21.130 ;
        RECT 61.580 20.950 61.710 21.130 ;
        RECT 62.090 20.950 62.220 21.130 ;
        RECT 63.580 20.950 63.710 21.130 ;
        RECT 64.090 20.950 64.220 21.130 ;
        RECT 65.580 20.950 65.710 21.130 ;
        RECT 66.090 20.950 66.220 21.130 ;
        RECT 67.580 20.950 67.710 21.130 ;
        RECT 68.090 20.950 68.220 21.130 ;
        RECT 69.580 20.950 69.710 21.130 ;
        RECT 70.090 20.950 70.220 21.130 ;
        RECT 71.580 20.950 71.710 21.130 ;
        RECT 72.090 20.950 72.220 21.130 ;
        RECT 73.580 20.950 73.710 21.130 ;
        RECT 74.090 20.950 74.220 21.130 ;
        RECT 75.580 20.950 75.710 21.130 ;
        RECT 76.090 20.950 76.220 21.130 ;
        RECT 77.580 20.950 77.710 21.130 ;
        RECT 78.090 20.950 78.220 21.130 ;
        RECT 79.580 20.950 79.710 21.130 ;
        RECT 80.090 20.950 80.220 21.130 ;
        RECT 81.580 20.950 81.710 21.130 ;
        RECT 82.090 20.950 82.220 21.130 ;
        RECT 83.580 20.950 83.710 21.130 ;
        RECT 84.090 20.950 84.220 21.130 ;
        RECT 85.580 20.950 85.710 21.130 ;
        RECT 86.090 20.950 86.220 21.130 ;
        RECT 87.580 20.950 87.710 21.130 ;
        RECT 88.090 20.950 88.220 21.130 ;
        RECT 89.580 20.950 89.710 21.130 ;
        RECT 90.090 20.950 90.220 21.130 ;
        RECT 91.580 20.950 91.710 21.130 ;
        RECT 92.090 20.950 92.220 21.130 ;
        RECT 93.580 20.950 93.710 21.130 ;
        RECT 94.090 20.950 94.220 21.130 ;
        RECT 95.580 20.950 95.710 21.130 ;
        RECT 96.090 20.950 96.220 21.130 ;
        RECT 97.580 20.950 97.710 21.130 ;
        RECT 98.090 20.950 98.220 21.130 ;
        RECT 99.580 20.950 99.710 21.130 ;
        RECT 100.090 20.950 100.220 21.130 ;
        RECT 101.580 20.950 101.710 21.130 ;
        RECT 102.090 20.950 102.220 21.130 ;
        RECT 103.580 20.950 103.710 21.130 ;
        RECT 104.090 20.950 104.220 21.130 ;
        RECT 105.580 20.950 105.710 21.130 ;
        RECT 106.090 20.950 106.220 21.130 ;
        RECT 107.580 20.950 107.710 21.130 ;
        RECT 108.090 20.950 108.220 21.130 ;
        RECT 109.580 20.950 109.710 21.130 ;
        RECT 110.090 20.950 110.220 21.130 ;
        RECT 111.580 20.950 111.710 21.130 ;
        RECT 112.090 20.950 112.220 21.130 ;
        RECT 113.580 20.950 113.710 21.130 ;
        RECT 114.090 20.950 114.220 21.130 ;
        RECT 115.580 20.950 115.710 21.130 ;
        RECT 116.090 20.950 116.220 21.130 ;
        RECT 117.580 20.950 117.710 21.130 ;
        RECT 118.090 20.950 118.220 21.130 ;
        RECT 119.580 20.950 119.710 21.130 ;
        RECT 120.090 20.950 120.220 21.130 ;
        RECT 121.580 20.950 121.710 21.130 ;
        RECT 122.090 20.950 122.220 21.130 ;
        RECT 123.580 20.950 123.710 21.130 ;
        RECT 124.090 20.950 124.220 21.130 ;
        RECT 125.580 20.950 125.710 21.130 ;
        RECT 126.090 20.950 126.220 21.130 ;
        RECT 127.580 20.950 127.710 21.130 ;
        RECT 128.090 20.950 128.220 21.130 ;
        RECT 129.580 20.950 129.710 21.130 ;
        RECT 130.090 20.950 130.220 21.130 ;
        RECT 131.580 20.950 131.710 21.130 ;
        RECT 132.090 20.950 132.220 21.130 ;
        RECT 0.900 14.050 1.080 14.650 ;
        RECT 2.280 14.050 2.720 14.650 ;
        RECT 2.900 14.050 3.080 14.650 ;
        RECT 4.280 14.050 4.720 14.650 ;
        RECT 4.900 14.050 5.080 14.650 ;
        RECT 6.280 14.050 6.720 14.650 ;
        RECT 6.900 14.050 7.080 14.650 ;
        RECT 8.280 14.050 8.720 14.650 ;
        RECT 8.900 14.050 9.080 14.650 ;
        RECT 10.280 14.050 10.720 14.650 ;
        RECT 10.900 14.050 11.080 14.650 ;
        RECT 12.280 14.050 12.720 14.650 ;
        RECT 12.900 14.050 13.080 14.650 ;
        RECT 14.280 14.050 14.720 14.650 ;
        RECT 14.900 14.050 15.080 14.650 ;
        RECT 16.280 14.050 16.720 14.650 ;
        RECT 16.900 14.050 17.080 14.650 ;
        RECT 18.280 14.050 18.720 14.650 ;
        RECT 18.900 14.050 19.080 14.650 ;
        RECT 20.280 14.050 20.720 14.650 ;
        RECT 20.900 14.050 21.080 14.650 ;
        RECT 22.280 14.050 22.720 14.650 ;
        RECT 22.900 14.050 23.080 14.650 ;
        RECT 24.280 14.050 24.720 14.650 ;
        RECT 24.900 14.050 25.080 14.650 ;
        RECT 26.280 14.050 26.720 14.650 ;
        RECT 26.900 14.050 27.080 14.650 ;
        RECT 28.280 14.050 28.720 14.650 ;
        RECT 28.900 14.050 29.080 14.650 ;
        RECT 30.280 14.050 30.720 14.650 ;
        RECT 30.900 14.050 31.080 14.650 ;
        RECT 32.280 14.050 32.720 14.650 ;
        RECT 32.900 14.050 33.080 14.650 ;
        RECT 34.280 14.050 34.720 14.650 ;
        RECT 34.900 14.050 35.080 14.650 ;
        RECT 36.280 14.050 36.720 14.650 ;
        RECT 36.900 14.050 37.080 14.650 ;
        RECT 38.280 14.050 38.720 14.650 ;
        RECT 38.900 14.050 39.080 14.650 ;
        RECT 40.280 14.050 40.720 14.650 ;
        RECT 40.900 14.050 41.080 14.650 ;
        RECT 42.280 14.050 42.720 14.650 ;
        RECT 42.900 14.050 43.080 14.650 ;
        RECT 44.280 14.050 44.720 14.650 ;
        RECT 44.900 14.050 45.080 14.650 ;
        RECT 46.280 14.050 46.720 14.650 ;
        RECT 46.900 14.050 47.080 14.650 ;
        RECT 48.280 14.050 48.720 14.650 ;
        RECT 48.900 14.050 49.080 14.650 ;
        RECT 50.280 14.050 50.720 14.650 ;
        RECT 50.900 14.050 51.080 14.650 ;
        RECT 52.280 14.050 52.720 14.650 ;
        RECT 52.900 14.050 53.080 14.650 ;
        RECT 54.280 14.050 54.720 14.650 ;
        RECT 54.900 14.050 55.080 14.650 ;
        RECT 56.280 14.050 56.720 14.650 ;
        RECT 56.900 14.050 57.080 14.650 ;
        RECT 58.280 14.050 58.720 14.650 ;
        RECT 58.900 14.050 59.080 14.650 ;
        RECT 60.280 14.050 60.720 14.650 ;
        RECT 60.900 14.050 61.080 14.650 ;
        RECT 62.280 14.050 62.720 14.650 ;
        RECT 62.900 14.050 63.080 14.650 ;
        RECT 64.280 14.050 64.720 14.650 ;
        RECT 64.900 14.050 65.080 14.650 ;
        RECT 66.280 14.050 66.720 14.650 ;
        RECT 66.900 14.050 67.080 14.650 ;
        RECT 68.280 14.050 68.720 14.650 ;
        RECT 68.900 14.050 69.080 14.650 ;
        RECT 70.280 14.050 70.720 14.650 ;
        RECT 70.900 14.050 71.080 14.650 ;
        RECT 72.280 14.050 72.720 14.650 ;
        RECT 72.900 14.050 73.080 14.650 ;
        RECT 74.280 14.050 74.720 14.650 ;
        RECT 74.900 14.050 75.080 14.650 ;
        RECT 76.280 14.050 76.720 14.650 ;
        RECT 76.900 14.050 77.080 14.650 ;
        RECT 78.280 14.050 78.720 14.650 ;
        RECT 78.900 14.050 79.080 14.650 ;
        RECT 80.280 14.050 80.720 14.650 ;
        RECT 80.900 14.050 81.080 14.650 ;
        RECT 82.280 14.050 82.720 14.650 ;
        RECT 82.900 14.050 83.080 14.650 ;
        RECT 84.280 14.050 84.720 14.650 ;
        RECT 84.900 14.050 85.080 14.650 ;
        RECT 86.280 14.050 86.720 14.650 ;
        RECT 86.900 14.050 87.080 14.650 ;
        RECT 88.280 14.050 88.720 14.650 ;
        RECT 88.900 14.050 89.080 14.650 ;
        RECT 90.280 14.050 90.720 14.650 ;
        RECT 90.900 14.050 91.080 14.650 ;
        RECT 92.280 14.050 92.720 14.650 ;
        RECT 92.900 14.050 93.080 14.650 ;
        RECT 94.280 14.050 94.720 14.650 ;
        RECT 94.900 14.050 95.080 14.650 ;
        RECT 96.280 14.050 96.720 14.650 ;
        RECT 96.900 14.050 97.080 14.650 ;
        RECT 98.280 14.050 98.720 14.650 ;
        RECT 98.900 14.050 99.080 14.650 ;
        RECT 100.280 14.050 100.720 14.650 ;
        RECT 100.900 14.050 101.080 14.650 ;
        RECT 102.280 14.050 102.720 14.650 ;
        RECT 102.900 14.050 103.080 14.650 ;
        RECT 104.280 14.050 104.720 14.650 ;
        RECT 104.900 14.050 105.080 14.650 ;
        RECT 106.280 14.050 106.720 14.650 ;
        RECT 106.900 14.050 107.080 14.650 ;
        RECT 108.280 14.050 108.720 14.650 ;
        RECT 108.900 14.050 109.080 14.650 ;
        RECT 110.280 14.050 110.720 14.650 ;
        RECT 110.900 14.050 111.080 14.650 ;
        RECT 112.280 14.050 112.720 14.650 ;
        RECT 112.900 14.050 113.080 14.650 ;
        RECT 114.280 14.050 114.720 14.650 ;
        RECT 114.900 14.050 115.080 14.650 ;
        RECT 116.280 14.050 116.720 14.650 ;
        RECT 116.900 14.050 117.080 14.650 ;
        RECT 118.280 14.050 118.720 14.650 ;
        RECT 118.900 14.050 119.080 14.650 ;
        RECT 120.280 14.050 120.720 14.650 ;
        RECT 120.900 14.050 121.080 14.650 ;
        RECT 122.280 14.050 122.720 14.650 ;
        RECT 122.900 14.050 123.080 14.650 ;
        RECT 124.280 14.050 124.720 14.650 ;
        RECT 124.900 14.050 125.080 14.650 ;
        RECT 126.280 14.050 126.720 14.650 ;
        RECT 126.900 14.050 127.080 14.650 ;
        RECT 128.280 14.050 128.720 14.650 ;
        RECT 128.900 14.050 129.080 14.650 ;
        RECT 130.280 14.050 130.720 14.650 ;
        RECT 130.900 14.050 131.080 14.650 ;
        RECT 132.280 14.050 132.720 14.650 ;
        RECT 1.080 11.540 1.520 12.140 ;
        RECT 2.720 11.540 2.900 12.140 ;
        RECT 3.080 11.540 3.520 12.140 ;
        RECT 4.720 11.540 4.900 12.140 ;
        RECT 5.080 11.540 5.520 12.140 ;
        RECT 6.720 11.540 6.900 12.140 ;
        RECT 7.080 11.540 7.520 12.140 ;
        RECT 8.720 11.540 8.900 12.140 ;
        RECT 9.080 11.540 9.520 12.140 ;
        RECT 10.720 11.540 10.900 12.140 ;
        RECT 11.080 11.540 11.520 12.140 ;
        RECT 12.720 11.540 12.900 12.140 ;
        RECT 13.080 11.540 13.520 12.140 ;
        RECT 14.720 11.540 14.900 12.140 ;
        RECT 15.080 11.540 15.520 12.140 ;
        RECT 16.720 11.540 16.900 12.140 ;
        RECT 17.080 11.540 17.520 12.140 ;
        RECT 18.720 11.540 18.900 12.140 ;
        RECT 19.080 11.540 19.520 12.140 ;
        RECT 20.720 11.540 20.900 12.140 ;
        RECT 21.080 11.540 21.520 12.140 ;
        RECT 22.720 11.540 22.900 12.140 ;
        RECT 23.080 11.540 23.520 12.140 ;
        RECT 24.720 11.540 24.900 12.140 ;
        RECT 25.080 11.540 25.520 12.140 ;
        RECT 26.720 11.540 26.900 12.140 ;
        RECT 27.080 11.540 27.520 12.140 ;
        RECT 28.720 11.540 28.900 12.140 ;
        RECT 29.080 11.540 29.520 12.140 ;
        RECT 30.720 11.540 30.900 12.140 ;
        RECT 31.080 11.540 31.520 12.140 ;
        RECT 32.720 11.540 32.900 12.140 ;
        RECT 33.080 11.540 33.520 12.140 ;
        RECT 34.720 11.540 34.900 12.140 ;
        RECT 35.080 11.540 35.520 12.140 ;
        RECT 36.720 11.540 36.900 12.140 ;
        RECT 37.080 11.540 37.520 12.140 ;
        RECT 38.720 11.540 38.900 12.140 ;
        RECT 39.080 11.540 39.520 12.140 ;
        RECT 40.720 11.540 40.900 12.140 ;
        RECT 41.080 11.540 41.520 12.140 ;
        RECT 42.720 11.540 42.900 12.140 ;
        RECT 43.080 11.540 43.520 12.140 ;
        RECT 44.720 11.540 44.900 12.140 ;
        RECT 45.080 11.540 45.520 12.140 ;
        RECT 46.720 11.540 46.900 12.140 ;
        RECT 47.080 11.540 47.520 12.140 ;
        RECT 48.720 11.540 48.900 12.140 ;
        RECT 49.080 11.540 49.520 12.140 ;
        RECT 50.720 11.540 50.900 12.140 ;
        RECT 51.080 11.540 51.520 12.140 ;
        RECT 52.720 11.540 52.900 12.140 ;
        RECT 53.080 11.540 53.520 12.140 ;
        RECT 54.720 11.540 54.900 12.140 ;
        RECT 55.080 11.540 55.520 12.140 ;
        RECT 56.720 11.540 56.900 12.140 ;
        RECT 57.080 11.540 57.520 12.140 ;
        RECT 58.720 11.540 58.900 12.140 ;
        RECT 59.080 11.540 59.520 12.140 ;
        RECT 60.720 11.540 60.900 12.140 ;
        RECT 61.080 11.540 61.520 12.140 ;
        RECT 62.720 11.540 62.900 12.140 ;
        RECT 63.080 11.540 63.520 12.140 ;
        RECT 64.720 11.540 64.900 12.140 ;
        RECT 65.080 11.540 65.520 12.140 ;
        RECT 66.720 11.540 66.900 12.140 ;
        RECT 67.080 11.540 67.520 12.140 ;
        RECT 68.720 11.540 68.900 12.140 ;
        RECT 69.080 11.540 69.520 12.140 ;
        RECT 70.720 11.540 70.900 12.140 ;
        RECT 71.080 11.540 71.520 12.140 ;
        RECT 72.720 11.540 72.900 12.140 ;
        RECT 73.080 11.540 73.520 12.140 ;
        RECT 74.720 11.540 74.900 12.140 ;
        RECT 75.080 11.540 75.520 12.140 ;
        RECT 76.720 11.540 76.900 12.140 ;
        RECT 77.080 11.540 77.520 12.140 ;
        RECT 78.720 11.540 78.900 12.140 ;
        RECT 79.080 11.540 79.520 12.140 ;
        RECT 80.720 11.540 80.900 12.140 ;
        RECT 81.080 11.540 81.520 12.140 ;
        RECT 82.720 11.540 82.900 12.140 ;
        RECT 83.080 11.540 83.520 12.140 ;
        RECT 84.720 11.540 84.900 12.140 ;
        RECT 85.080 11.540 85.520 12.140 ;
        RECT 86.720 11.540 86.900 12.140 ;
        RECT 87.080 11.540 87.520 12.140 ;
        RECT 88.720 11.540 88.900 12.140 ;
        RECT 89.080 11.540 89.520 12.140 ;
        RECT 90.720 11.540 90.900 12.140 ;
        RECT 91.080 11.540 91.520 12.140 ;
        RECT 92.720 11.540 92.900 12.140 ;
        RECT 93.080 11.540 93.520 12.140 ;
        RECT 94.720 11.540 94.900 12.140 ;
        RECT 95.080 11.540 95.520 12.140 ;
        RECT 96.720 11.540 96.900 12.140 ;
        RECT 97.080 11.540 97.520 12.140 ;
        RECT 98.720 11.540 98.900 12.140 ;
        RECT 99.080 11.540 99.520 12.140 ;
        RECT 100.720 11.540 100.900 12.140 ;
        RECT 101.080 11.540 101.520 12.140 ;
        RECT 102.720 11.540 102.900 12.140 ;
        RECT 103.080 11.540 103.520 12.140 ;
        RECT 104.720 11.540 104.900 12.140 ;
        RECT 105.080 11.540 105.520 12.140 ;
        RECT 106.720 11.540 106.900 12.140 ;
        RECT 107.080 11.540 107.520 12.140 ;
        RECT 108.720 11.540 108.900 12.140 ;
        RECT 109.080 11.540 109.520 12.140 ;
        RECT 110.720 11.540 110.900 12.140 ;
        RECT 111.080 11.540 111.520 12.140 ;
        RECT 112.720 11.540 112.900 12.140 ;
        RECT 113.080 11.540 113.520 12.140 ;
        RECT 114.720 11.540 114.900 12.140 ;
        RECT 115.080 11.540 115.520 12.140 ;
        RECT 116.720 11.540 116.900 12.140 ;
        RECT 117.080 11.540 117.520 12.140 ;
        RECT 118.720 11.540 118.900 12.140 ;
        RECT 119.080 11.540 119.520 12.140 ;
        RECT 120.720 11.540 120.900 12.140 ;
        RECT 121.080 11.540 121.520 12.140 ;
        RECT 122.720 11.540 122.900 12.140 ;
        RECT 123.080 11.540 123.520 12.140 ;
        RECT 124.720 11.540 124.900 12.140 ;
        RECT 125.080 11.540 125.520 12.140 ;
        RECT 126.720 11.540 126.900 12.140 ;
        RECT 127.080 11.540 127.520 12.140 ;
        RECT 128.720 11.540 128.900 12.140 ;
        RECT 129.080 11.540 129.520 12.140 ;
        RECT 130.720 11.540 130.900 12.140 ;
        RECT 131.080 11.540 131.520 12.140 ;
        RECT 132.720 11.540 132.900 12.140 ;
        RECT 1.580 5.060 1.710 5.240 ;
        RECT 2.090 5.060 2.220 5.240 ;
        RECT 3.580 5.060 3.710 5.240 ;
        RECT 4.090 5.060 4.220 5.240 ;
        RECT 5.580 5.060 5.710 5.240 ;
        RECT 6.090 5.060 6.220 5.240 ;
        RECT 7.580 5.060 7.710 5.240 ;
        RECT 8.090 5.060 8.220 5.240 ;
        RECT 9.580 5.060 9.710 5.240 ;
        RECT 10.090 5.060 10.220 5.240 ;
        RECT 11.580 5.060 11.710 5.240 ;
        RECT 12.090 5.060 12.220 5.240 ;
        RECT 13.580 5.060 13.710 5.240 ;
        RECT 14.090 5.060 14.220 5.240 ;
        RECT 15.580 5.060 15.710 5.240 ;
        RECT 16.090 5.060 16.220 5.240 ;
        RECT 17.580 5.060 17.710 5.240 ;
        RECT 18.090 5.060 18.220 5.240 ;
        RECT 19.580 5.060 19.710 5.240 ;
        RECT 20.090 5.060 20.220 5.240 ;
        RECT 21.580 5.060 21.710 5.240 ;
        RECT 22.090 5.060 22.220 5.240 ;
        RECT 23.580 5.060 23.710 5.240 ;
        RECT 24.090 5.060 24.220 5.240 ;
        RECT 25.580 5.060 25.710 5.240 ;
        RECT 26.090 5.060 26.220 5.240 ;
        RECT 27.580 5.060 27.710 5.240 ;
        RECT 28.090 5.060 28.220 5.240 ;
        RECT 29.580 5.060 29.710 5.240 ;
        RECT 30.090 5.060 30.220 5.240 ;
        RECT 31.580 5.060 31.710 5.240 ;
        RECT 32.090 5.060 32.220 5.240 ;
        RECT 33.580 5.060 33.710 5.240 ;
        RECT 34.090 5.060 34.220 5.240 ;
        RECT 35.580 5.060 35.710 5.240 ;
        RECT 36.090 5.060 36.220 5.240 ;
        RECT 37.580 5.060 37.710 5.240 ;
        RECT 38.090 5.060 38.220 5.240 ;
        RECT 39.580 5.060 39.710 5.240 ;
        RECT 40.090 5.060 40.220 5.240 ;
        RECT 41.580 5.060 41.710 5.240 ;
        RECT 42.090 5.060 42.220 5.240 ;
        RECT 43.580 5.060 43.710 5.240 ;
        RECT 44.090 5.060 44.220 5.240 ;
        RECT 45.580 5.060 45.710 5.240 ;
        RECT 46.090 5.060 46.220 5.240 ;
        RECT 47.580 5.060 47.710 5.240 ;
        RECT 48.090 5.060 48.220 5.240 ;
        RECT 49.580 5.060 49.710 5.240 ;
        RECT 50.090 5.060 50.220 5.240 ;
        RECT 51.580 5.060 51.710 5.240 ;
        RECT 52.090 5.060 52.220 5.240 ;
        RECT 53.580 5.060 53.710 5.240 ;
        RECT 54.090 5.060 54.220 5.240 ;
        RECT 55.580 5.060 55.710 5.240 ;
        RECT 56.090 5.060 56.220 5.240 ;
        RECT 57.580 5.060 57.710 5.240 ;
        RECT 58.090 5.060 58.220 5.240 ;
        RECT 59.580 5.060 59.710 5.240 ;
        RECT 60.090 5.060 60.220 5.240 ;
        RECT 61.580 5.060 61.710 5.240 ;
        RECT 62.090 5.060 62.220 5.240 ;
        RECT 63.580 5.060 63.710 5.240 ;
        RECT 64.090 5.060 64.220 5.240 ;
        RECT 65.580 5.060 65.710 5.240 ;
        RECT 66.090 5.060 66.220 5.240 ;
        RECT 67.580 5.060 67.710 5.240 ;
        RECT 68.090 5.060 68.220 5.240 ;
        RECT 69.580 5.060 69.710 5.240 ;
        RECT 70.090 5.060 70.220 5.240 ;
        RECT 71.580 5.060 71.710 5.240 ;
        RECT 72.090 5.060 72.220 5.240 ;
        RECT 73.580 5.060 73.710 5.240 ;
        RECT 74.090 5.060 74.220 5.240 ;
        RECT 75.580 5.060 75.710 5.240 ;
        RECT 76.090 5.060 76.220 5.240 ;
        RECT 77.580 5.060 77.710 5.240 ;
        RECT 78.090 5.060 78.220 5.240 ;
        RECT 79.580 5.060 79.710 5.240 ;
        RECT 80.090 5.060 80.220 5.240 ;
        RECT 81.580 5.060 81.710 5.240 ;
        RECT 82.090 5.060 82.220 5.240 ;
        RECT 83.580 5.060 83.710 5.240 ;
        RECT 84.090 5.060 84.220 5.240 ;
        RECT 85.580 5.060 85.710 5.240 ;
        RECT 86.090 5.060 86.220 5.240 ;
        RECT 87.580 5.060 87.710 5.240 ;
        RECT 88.090 5.060 88.220 5.240 ;
        RECT 89.580 5.060 89.710 5.240 ;
        RECT 90.090 5.060 90.220 5.240 ;
        RECT 91.580 5.060 91.710 5.240 ;
        RECT 92.090 5.060 92.220 5.240 ;
        RECT 93.580 5.060 93.710 5.240 ;
        RECT 94.090 5.060 94.220 5.240 ;
        RECT 95.580 5.060 95.710 5.240 ;
        RECT 96.090 5.060 96.220 5.240 ;
        RECT 97.580 5.060 97.710 5.240 ;
        RECT 98.090 5.060 98.220 5.240 ;
        RECT 99.580 5.060 99.710 5.240 ;
        RECT 100.090 5.060 100.220 5.240 ;
        RECT 101.580 5.060 101.710 5.240 ;
        RECT 102.090 5.060 102.220 5.240 ;
        RECT 103.580 5.060 103.710 5.240 ;
        RECT 104.090 5.060 104.220 5.240 ;
        RECT 105.580 5.060 105.710 5.240 ;
        RECT 106.090 5.060 106.220 5.240 ;
        RECT 107.580 5.060 107.710 5.240 ;
        RECT 108.090 5.060 108.220 5.240 ;
        RECT 109.580 5.060 109.710 5.240 ;
        RECT 110.090 5.060 110.220 5.240 ;
        RECT 111.580 5.060 111.710 5.240 ;
        RECT 112.090 5.060 112.220 5.240 ;
        RECT 113.580 5.060 113.710 5.240 ;
        RECT 114.090 5.060 114.220 5.240 ;
        RECT 115.580 5.060 115.710 5.240 ;
        RECT 116.090 5.060 116.220 5.240 ;
        RECT 117.580 5.060 117.710 5.240 ;
        RECT 118.090 5.060 118.220 5.240 ;
        RECT 119.580 5.060 119.710 5.240 ;
        RECT 120.090 5.060 120.220 5.240 ;
        RECT 121.580 5.060 121.710 5.240 ;
        RECT 122.090 5.060 122.220 5.240 ;
        RECT 123.580 5.060 123.710 5.240 ;
        RECT 124.090 5.060 124.220 5.240 ;
        RECT 125.580 5.060 125.710 5.240 ;
        RECT 126.090 5.060 126.220 5.240 ;
        RECT 127.580 5.060 127.710 5.240 ;
        RECT 128.090 5.060 128.220 5.240 ;
        RECT 129.580 5.060 129.710 5.240 ;
        RECT 130.090 5.060 130.220 5.240 ;
        RECT 131.580 5.060 131.710 5.240 ;
        RECT 132.090 5.060 132.220 5.240 ;
        RECT 1.580 4.560 1.710 4.760 ;
        RECT 1.410 4.260 1.710 4.560 ;
        RECT 2.090 4.560 2.220 4.760 ;
        RECT 3.580 4.560 3.710 4.760 ;
        RECT 2.090 4.260 2.390 4.560 ;
        RECT 3.410 4.260 3.710 4.560 ;
        RECT 4.090 4.560 4.220 4.760 ;
        RECT 5.580 4.560 5.710 4.760 ;
        RECT 4.090 4.260 4.390 4.560 ;
        RECT 5.410 4.260 5.710 4.560 ;
        RECT 6.090 4.560 6.220 4.760 ;
        RECT 7.580 4.560 7.710 4.760 ;
        RECT 6.090 4.260 6.390 4.560 ;
        RECT 7.410 4.260 7.710 4.560 ;
        RECT 8.090 4.560 8.220 4.760 ;
        RECT 9.580 4.560 9.710 4.760 ;
        RECT 8.090 4.260 8.390 4.560 ;
        RECT 9.410 4.260 9.710 4.560 ;
        RECT 10.090 4.560 10.220 4.760 ;
        RECT 11.580 4.560 11.710 4.760 ;
        RECT 10.090 4.260 10.390 4.560 ;
        RECT 11.410 4.260 11.710 4.560 ;
        RECT 12.090 4.560 12.220 4.760 ;
        RECT 13.580 4.560 13.710 4.760 ;
        RECT 12.090 4.260 12.390 4.560 ;
        RECT 13.410 4.260 13.710 4.560 ;
        RECT 14.090 4.560 14.220 4.760 ;
        RECT 15.580 4.560 15.710 4.760 ;
        RECT 14.090 4.260 14.390 4.560 ;
        RECT 15.410 4.260 15.710 4.560 ;
        RECT 16.090 4.560 16.220 4.760 ;
        RECT 17.580 4.560 17.710 4.760 ;
        RECT 16.090 4.260 16.390 4.560 ;
        RECT 17.410 4.260 17.710 4.560 ;
        RECT 18.090 4.560 18.220 4.760 ;
        RECT 19.580 4.560 19.710 4.760 ;
        RECT 18.090 4.260 18.390 4.560 ;
        RECT 19.410 4.260 19.710 4.560 ;
        RECT 20.090 4.560 20.220 4.760 ;
        RECT 21.580 4.560 21.710 4.760 ;
        RECT 20.090 4.260 20.390 4.560 ;
        RECT 21.410 4.260 21.710 4.560 ;
        RECT 22.090 4.560 22.220 4.760 ;
        RECT 23.580 4.560 23.710 4.760 ;
        RECT 22.090 4.260 22.390 4.560 ;
        RECT 23.410 4.260 23.710 4.560 ;
        RECT 24.090 4.560 24.220 4.760 ;
        RECT 25.580 4.560 25.710 4.760 ;
        RECT 24.090 4.260 24.390 4.560 ;
        RECT 25.410 4.260 25.710 4.560 ;
        RECT 26.090 4.560 26.220 4.760 ;
        RECT 27.580 4.560 27.710 4.760 ;
        RECT 26.090 4.260 26.390 4.560 ;
        RECT 27.410 4.260 27.710 4.560 ;
        RECT 28.090 4.560 28.220 4.760 ;
        RECT 29.580 4.560 29.710 4.760 ;
        RECT 28.090 4.260 28.390 4.560 ;
        RECT 29.410 4.260 29.710 4.560 ;
        RECT 30.090 4.560 30.220 4.760 ;
        RECT 31.580 4.560 31.710 4.760 ;
        RECT 30.090 4.260 30.390 4.560 ;
        RECT 31.410 4.260 31.710 4.560 ;
        RECT 32.090 4.560 32.220 4.760 ;
        RECT 33.580 4.560 33.710 4.760 ;
        RECT 32.090 4.260 32.390 4.560 ;
        RECT 33.410 4.260 33.710 4.560 ;
        RECT 34.090 4.560 34.220 4.760 ;
        RECT 35.580 4.560 35.710 4.760 ;
        RECT 34.090 4.260 34.390 4.560 ;
        RECT 35.410 4.260 35.710 4.560 ;
        RECT 36.090 4.560 36.220 4.760 ;
        RECT 37.580 4.560 37.710 4.760 ;
        RECT 36.090 4.260 36.390 4.560 ;
        RECT 37.410 4.260 37.710 4.560 ;
        RECT 38.090 4.560 38.220 4.760 ;
        RECT 39.580 4.560 39.710 4.760 ;
        RECT 38.090 4.260 38.390 4.560 ;
        RECT 39.410 4.260 39.710 4.560 ;
        RECT 40.090 4.560 40.220 4.760 ;
        RECT 41.580 4.560 41.710 4.760 ;
        RECT 40.090 4.260 40.390 4.560 ;
        RECT 41.410 4.260 41.710 4.560 ;
        RECT 42.090 4.560 42.220 4.760 ;
        RECT 43.580 4.560 43.710 4.760 ;
        RECT 42.090 4.260 42.390 4.560 ;
        RECT 43.410 4.260 43.710 4.560 ;
        RECT 44.090 4.560 44.220 4.760 ;
        RECT 45.580 4.560 45.710 4.760 ;
        RECT 44.090 4.260 44.390 4.560 ;
        RECT 45.410 4.260 45.710 4.560 ;
        RECT 46.090 4.560 46.220 4.760 ;
        RECT 47.580 4.560 47.710 4.760 ;
        RECT 46.090 4.260 46.390 4.560 ;
        RECT 47.410 4.260 47.710 4.560 ;
        RECT 48.090 4.560 48.220 4.760 ;
        RECT 49.580 4.560 49.710 4.760 ;
        RECT 48.090 4.260 48.390 4.560 ;
        RECT 49.410 4.260 49.710 4.560 ;
        RECT 50.090 4.560 50.220 4.760 ;
        RECT 51.580 4.560 51.710 4.760 ;
        RECT 50.090 4.260 50.390 4.560 ;
        RECT 51.410 4.260 51.710 4.560 ;
        RECT 52.090 4.560 52.220 4.760 ;
        RECT 53.580 4.560 53.710 4.760 ;
        RECT 52.090 4.260 52.390 4.560 ;
        RECT 53.410 4.260 53.710 4.560 ;
        RECT 54.090 4.560 54.220 4.760 ;
        RECT 55.580 4.560 55.710 4.760 ;
        RECT 54.090 4.260 54.390 4.560 ;
        RECT 55.410 4.260 55.710 4.560 ;
        RECT 56.090 4.560 56.220 4.760 ;
        RECT 57.580 4.560 57.710 4.760 ;
        RECT 56.090 4.260 56.390 4.560 ;
        RECT 57.410 4.260 57.710 4.560 ;
        RECT 58.090 4.560 58.220 4.760 ;
        RECT 59.580 4.560 59.710 4.760 ;
        RECT 58.090 4.260 58.390 4.560 ;
        RECT 59.410 4.260 59.710 4.560 ;
        RECT 60.090 4.560 60.220 4.760 ;
        RECT 61.580 4.560 61.710 4.760 ;
        RECT 60.090 4.260 60.390 4.560 ;
        RECT 61.410 4.260 61.710 4.560 ;
        RECT 62.090 4.560 62.220 4.760 ;
        RECT 63.580 4.560 63.710 4.760 ;
        RECT 62.090 4.260 62.390 4.560 ;
        RECT 63.410 4.260 63.710 4.560 ;
        RECT 64.090 4.560 64.220 4.760 ;
        RECT 65.580 4.560 65.710 4.760 ;
        RECT 64.090 4.260 64.390 4.560 ;
        RECT 65.410 4.260 65.710 4.560 ;
        RECT 66.090 4.560 66.220 4.760 ;
        RECT 67.580 4.560 67.710 4.760 ;
        RECT 66.090 4.260 66.390 4.560 ;
        RECT 67.410 4.260 67.710 4.560 ;
        RECT 68.090 4.560 68.220 4.760 ;
        RECT 69.580 4.560 69.710 4.760 ;
        RECT 68.090 4.260 68.390 4.560 ;
        RECT 69.410 4.260 69.710 4.560 ;
        RECT 70.090 4.560 70.220 4.760 ;
        RECT 71.580 4.560 71.710 4.760 ;
        RECT 70.090 4.260 70.390 4.560 ;
        RECT 71.410 4.260 71.710 4.560 ;
        RECT 72.090 4.560 72.220 4.760 ;
        RECT 73.580 4.560 73.710 4.760 ;
        RECT 72.090 4.260 72.390 4.560 ;
        RECT 73.410 4.260 73.710 4.560 ;
        RECT 74.090 4.560 74.220 4.760 ;
        RECT 75.580 4.560 75.710 4.760 ;
        RECT 74.090 4.260 74.390 4.560 ;
        RECT 75.410 4.260 75.710 4.560 ;
        RECT 76.090 4.560 76.220 4.760 ;
        RECT 77.580 4.560 77.710 4.760 ;
        RECT 76.090 4.260 76.390 4.560 ;
        RECT 77.410 4.260 77.710 4.560 ;
        RECT 78.090 4.560 78.220 4.760 ;
        RECT 79.580 4.560 79.710 4.760 ;
        RECT 78.090 4.260 78.390 4.560 ;
        RECT 79.410 4.260 79.710 4.560 ;
        RECT 80.090 4.560 80.220 4.760 ;
        RECT 81.580 4.560 81.710 4.760 ;
        RECT 80.090 4.260 80.390 4.560 ;
        RECT 81.410 4.260 81.710 4.560 ;
        RECT 82.090 4.560 82.220 4.760 ;
        RECT 83.580 4.560 83.710 4.760 ;
        RECT 82.090 4.260 82.390 4.560 ;
        RECT 83.410 4.260 83.710 4.560 ;
        RECT 84.090 4.560 84.220 4.760 ;
        RECT 85.580 4.560 85.710 4.760 ;
        RECT 84.090 4.260 84.390 4.560 ;
        RECT 85.410 4.260 85.710 4.560 ;
        RECT 86.090 4.560 86.220 4.760 ;
        RECT 87.580 4.560 87.710 4.760 ;
        RECT 86.090 4.260 86.390 4.560 ;
        RECT 87.410 4.260 87.710 4.560 ;
        RECT 88.090 4.560 88.220 4.760 ;
        RECT 89.580 4.560 89.710 4.760 ;
        RECT 88.090 4.260 88.390 4.560 ;
        RECT 89.410 4.260 89.710 4.560 ;
        RECT 90.090 4.560 90.220 4.760 ;
        RECT 91.580 4.560 91.710 4.760 ;
        RECT 90.090 4.260 90.390 4.560 ;
        RECT 91.410 4.260 91.710 4.560 ;
        RECT 92.090 4.560 92.220 4.760 ;
        RECT 93.580 4.560 93.710 4.760 ;
        RECT 92.090 4.260 92.390 4.560 ;
        RECT 93.410 4.260 93.710 4.560 ;
        RECT 94.090 4.560 94.220 4.760 ;
        RECT 95.580 4.560 95.710 4.760 ;
        RECT 94.090 4.260 94.390 4.560 ;
        RECT 95.410 4.260 95.710 4.560 ;
        RECT 96.090 4.560 96.220 4.760 ;
        RECT 97.580 4.560 97.710 4.760 ;
        RECT 96.090 4.260 96.390 4.560 ;
        RECT 97.410 4.260 97.710 4.560 ;
        RECT 98.090 4.560 98.220 4.760 ;
        RECT 99.580 4.560 99.710 4.760 ;
        RECT 98.090 4.260 98.390 4.560 ;
        RECT 99.410 4.260 99.710 4.560 ;
        RECT 100.090 4.560 100.220 4.760 ;
        RECT 101.580 4.560 101.710 4.760 ;
        RECT 100.090 4.260 100.390 4.560 ;
        RECT 101.410 4.260 101.710 4.560 ;
        RECT 102.090 4.560 102.220 4.760 ;
        RECT 103.580 4.560 103.710 4.760 ;
        RECT 102.090 4.260 102.390 4.560 ;
        RECT 103.410 4.260 103.710 4.560 ;
        RECT 104.090 4.560 104.220 4.760 ;
        RECT 105.580 4.560 105.710 4.760 ;
        RECT 104.090 4.260 104.390 4.560 ;
        RECT 105.410 4.260 105.710 4.560 ;
        RECT 106.090 4.560 106.220 4.760 ;
        RECT 107.580 4.560 107.710 4.760 ;
        RECT 106.090 4.260 106.390 4.560 ;
        RECT 107.410 4.260 107.710 4.560 ;
        RECT 108.090 4.560 108.220 4.760 ;
        RECT 109.580 4.560 109.710 4.760 ;
        RECT 108.090 4.260 108.390 4.560 ;
        RECT 109.410 4.260 109.710 4.560 ;
        RECT 110.090 4.560 110.220 4.760 ;
        RECT 111.580 4.560 111.710 4.760 ;
        RECT 110.090 4.260 110.390 4.560 ;
        RECT 111.410 4.260 111.710 4.560 ;
        RECT 112.090 4.560 112.220 4.760 ;
        RECT 113.580 4.560 113.710 4.760 ;
        RECT 112.090 4.260 112.390 4.560 ;
        RECT 113.410 4.260 113.710 4.560 ;
        RECT 114.090 4.560 114.220 4.760 ;
        RECT 115.580 4.560 115.710 4.760 ;
        RECT 114.090 4.260 114.390 4.560 ;
        RECT 115.410 4.260 115.710 4.560 ;
        RECT 116.090 4.560 116.220 4.760 ;
        RECT 117.580 4.560 117.710 4.760 ;
        RECT 116.090 4.260 116.390 4.560 ;
        RECT 117.410 4.260 117.710 4.560 ;
        RECT 118.090 4.560 118.220 4.760 ;
        RECT 119.580 4.560 119.710 4.760 ;
        RECT 118.090 4.260 118.390 4.560 ;
        RECT 119.410 4.260 119.710 4.560 ;
        RECT 120.090 4.560 120.220 4.760 ;
        RECT 121.580 4.560 121.710 4.760 ;
        RECT 120.090 4.260 120.390 4.560 ;
        RECT 121.410 4.260 121.710 4.560 ;
        RECT 122.090 4.560 122.220 4.760 ;
        RECT 123.580 4.560 123.710 4.760 ;
        RECT 122.090 4.260 122.390 4.560 ;
        RECT 123.410 4.260 123.710 4.560 ;
        RECT 124.090 4.560 124.220 4.760 ;
        RECT 125.580 4.560 125.710 4.760 ;
        RECT 124.090 4.260 124.390 4.560 ;
        RECT 125.410 4.260 125.710 4.560 ;
        RECT 126.090 4.560 126.220 4.760 ;
        RECT 127.580 4.560 127.710 4.760 ;
        RECT 126.090 4.260 126.390 4.560 ;
        RECT 127.410 4.260 127.710 4.560 ;
        RECT 128.090 4.560 128.220 4.760 ;
        RECT 129.580 4.560 129.710 4.760 ;
        RECT 128.090 4.260 128.390 4.560 ;
        RECT 129.410 4.260 129.710 4.560 ;
        RECT 130.090 4.560 130.220 4.760 ;
        RECT 131.580 4.560 131.710 4.760 ;
        RECT 130.090 4.260 130.390 4.560 ;
        RECT 131.410 4.260 131.710 4.560 ;
        RECT 132.090 4.560 132.220 4.760 ;
        RECT 132.090 4.260 132.390 4.560 ;
        RECT 1.455 2.030 2.795 2.330 ;
        RECT 3.455 2.030 4.795 2.330 ;
        RECT 5.455 2.030 6.795 2.330 ;
        RECT 7.455 2.030 8.795 2.330 ;
        RECT 9.455 2.030 10.795 2.330 ;
        RECT 11.455 2.030 12.795 2.330 ;
        RECT 13.455 2.030 14.795 2.330 ;
        RECT 15.455 2.030 16.795 2.330 ;
        RECT 17.455 2.030 18.795 2.330 ;
        RECT 19.455 2.030 20.795 2.330 ;
        RECT 21.455 2.030 22.795 2.330 ;
        RECT 23.455 2.030 24.795 2.330 ;
        RECT 25.455 2.030 26.795 2.330 ;
        RECT 27.455 2.030 28.795 2.330 ;
        RECT 29.455 2.030 30.795 2.330 ;
        RECT 31.455 2.030 32.795 2.330 ;
        RECT 33.455 2.030 34.795 2.330 ;
        RECT 35.455 2.030 36.795 2.330 ;
        RECT 37.455 2.030 38.795 2.330 ;
        RECT 39.455 2.030 40.795 2.330 ;
        RECT 41.455 2.030 42.795 2.330 ;
        RECT 43.455 2.030 44.795 2.330 ;
        RECT 45.455 2.030 46.795 2.330 ;
        RECT 47.455 2.030 48.795 2.330 ;
        RECT 49.455 2.030 50.795 2.330 ;
        RECT 51.455 2.030 52.795 2.330 ;
        RECT 53.455 2.030 54.795 2.330 ;
        RECT 55.455 2.030 56.795 2.330 ;
        RECT 57.455 2.030 58.795 2.330 ;
        RECT 59.455 2.030 60.795 2.330 ;
        RECT 61.455 2.030 62.795 2.330 ;
        RECT 63.455 2.030 64.795 2.330 ;
        RECT 65.455 2.030 66.795 2.330 ;
        RECT 67.455 2.030 68.795 2.330 ;
        RECT 69.455 2.030 70.795 2.330 ;
        RECT 71.455 2.030 72.795 2.330 ;
        RECT 73.455 2.030 74.795 2.330 ;
        RECT 75.455 2.030 76.795 2.330 ;
        RECT 77.455 2.030 78.795 2.330 ;
        RECT 79.455 2.030 80.795 2.330 ;
        RECT 81.455 2.030 82.795 2.330 ;
        RECT 83.455 2.030 84.795 2.330 ;
        RECT 85.455 2.030 86.795 2.330 ;
        RECT 87.455 2.030 88.795 2.330 ;
        RECT 89.455 2.030 90.795 2.330 ;
        RECT 91.455 2.030 92.795 2.330 ;
        RECT 93.455 2.030 94.795 2.330 ;
        RECT 95.455 2.030 96.795 2.330 ;
        RECT 97.455 2.030 98.795 2.330 ;
        RECT 99.455 2.030 100.795 2.330 ;
        RECT 101.455 2.030 102.795 2.330 ;
        RECT 103.455 2.030 104.795 2.330 ;
        RECT 105.455 2.030 106.795 2.330 ;
        RECT 107.455 2.030 108.795 2.330 ;
        RECT 109.455 2.030 110.795 2.330 ;
        RECT 111.455 2.030 112.795 2.330 ;
        RECT 113.455 2.030 114.795 2.330 ;
        RECT 115.455 2.030 116.795 2.330 ;
        RECT 117.455 2.030 118.795 2.330 ;
        RECT 119.455 2.030 120.795 2.330 ;
        RECT 121.455 2.030 122.795 2.330 ;
        RECT 123.455 2.030 124.795 2.330 ;
        RECT 125.455 2.030 126.795 2.330 ;
        RECT 127.455 2.030 128.795 2.330 ;
        RECT 129.455 2.030 130.795 2.330 ;
        RECT 131.455 2.030 132.795 2.330 ;
        RECT 1.455 1.660 1.755 2.030 ;
        RECT 1.235 1.480 1.755 1.660 ;
        RECT 2.045 1.660 2.345 1.850 ;
        RECT 3.455 1.660 3.755 2.030 ;
        RECT 2.045 1.480 2.565 1.660 ;
        RECT 3.235 1.480 3.755 1.660 ;
        RECT 4.045 1.660 4.345 1.850 ;
        RECT 5.455 1.660 5.755 2.030 ;
        RECT 4.045 1.480 4.565 1.660 ;
        RECT 5.235 1.480 5.755 1.660 ;
        RECT 6.045 1.660 6.345 1.850 ;
        RECT 7.455 1.660 7.755 2.030 ;
        RECT 6.045 1.480 6.565 1.660 ;
        RECT 7.235 1.480 7.755 1.660 ;
        RECT 8.045 1.660 8.345 1.850 ;
        RECT 9.455 1.660 9.755 2.030 ;
        RECT 8.045 1.480 8.565 1.660 ;
        RECT 9.235 1.480 9.755 1.660 ;
        RECT 10.045 1.660 10.345 1.850 ;
        RECT 11.455 1.660 11.755 2.030 ;
        RECT 10.045 1.480 10.565 1.660 ;
        RECT 11.235 1.480 11.755 1.660 ;
        RECT 12.045 1.660 12.345 1.850 ;
        RECT 13.455 1.660 13.755 2.030 ;
        RECT 12.045 1.480 12.565 1.660 ;
        RECT 13.235 1.480 13.755 1.660 ;
        RECT 14.045 1.660 14.345 1.850 ;
        RECT 15.455 1.660 15.755 2.030 ;
        RECT 14.045 1.480 14.565 1.660 ;
        RECT 15.235 1.480 15.755 1.660 ;
        RECT 16.045 1.660 16.345 1.850 ;
        RECT 17.455 1.660 17.755 2.030 ;
        RECT 16.045 1.480 16.565 1.660 ;
        RECT 17.235 1.480 17.755 1.660 ;
        RECT 18.045 1.660 18.345 1.850 ;
        RECT 19.455 1.660 19.755 2.030 ;
        RECT 18.045 1.480 18.565 1.660 ;
        RECT 19.235 1.480 19.755 1.660 ;
        RECT 20.045 1.660 20.345 1.850 ;
        RECT 21.455 1.660 21.755 2.030 ;
        RECT 20.045 1.480 20.565 1.660 ;
        RECT 21.235 1.480 21.755 1.660 ;
        RECT 22.045 1.660 22.345 1.850 ;
        RECT 23.455 1.660 23.755 2.030 ;
        RECT 22.045 1.480 22.565 1.660 ;
        RECT 23.235 1.480 23.755 1.660 ;
        RECT 24.045 1.660 24.345 1.850 ;
        RECT 25.455 1.660 25.755 2.030 ;
        RECT 24.045 1.480 24.565 1.660 ;
        RECT 25.235 1.480 25.755 1.660 ;
        RECT 26.045 1.660 26.345 1.850 ;
        RECT 27.455 1.660 27.755 2.030 ;
        RECT 26.045 1.480 26.565 1.660 ;
        RECT 27.235 1.480 27.755 1.660 ;
        RECT 28.045 1.660 28.345 1.850 ;
        RECT 29.455 1.660 29.755 2.030 ;
        RECT 28.045 1.480 28.565 1.660 ;
        RECT 29.235 1.480 29.755 1.660 ;
        RECT 30.045 1.660 30.345 1.850 ;
        RECT 31.455 1.660 31.755 2.030 ;
        RECT 30.045 1.480 30.565 1.660 ;
        RECT 31.235 1.480 31.755 1.660 ;
        RECT 32.045 1.660 32.345 1.850 ;
        RECT 33.455 1.660 33.755 2.030 ;
        RECT 32.045 1.480 32.565 1.660 ;
        RECT 33.235 1.480 33.755 1.660 ;
        RECT 34.045 1.660 34.345 1.850 ;
        RECT 35.455 1.660 35.755 2.030 ;
        RECT 34.045 1.480 34.565 1.660 ;
        RECT 35.235 1.480 35.755 1.660 ;
        RECT 36.045 1.660 36.345 1.850 ;
        RECT 37.455 1.660 37.755 2.030 ;
        RECT 36.045 1.480 36.565 1.660 ;
        RECT 37.235 1.480 37.755 1.660 ;
        RECT 38.045 1.660 38.345 1.850 ;
        RECT 39.455 1.660 39.755 2.030 ;
        RECT 38.045 1.480 38.565 1.660 ;
        RECT 39.235 1.480 39.755 1.660 ;
        RECT 40.045 1.660 40.345 1.850 ;
        RECT 41.455 1.660 41.755 2.030 ;
        RECT 40.045 1.480 40.565 1.660 ;
        RECT 41.235 1.480 41.755 1.660 ;
        RECT 42.045 1.660 42.345 1.850 ;
        RECT 43.455 1.660 43.755 2.030 ;
        RECT 42.045 1.480 42.565 1.660 ;
        RECT 43.235 1.480 43.755 1.660 ;
        RECT 44.045 1.660 44.345 1.850 ;
        RECT 45.455 1.660 45.755 2.030 ;
        RECT 44.045 1.480 44.565 1.660 ;
        RECT 45.235 1.480 45.755 1.660 ;
        RECT 46.045 1.660 46.345 1.850 ;
        RECT 47.455 1.660 47.755 2.030 ;
        RECT 46.045 1.480 46.565 1.660 ;
        RECT 47.235 1.480 47.755 1.660 ;
        RECT 48.045 1.660 48.345 1.850 ;
        RECT 49.455 1.660 49.755 2.030 ;
        RECT 48.045 1.480 48.565 1.660 ;
        RECT 49.235 1.480 49.755 1.660 ;
        RECT 50.045 1.660 50.345 1.850 ;
        RECT 51.455 1.660 51.755 2.030 ;
        RECT 50.045 1.480 50.565 1.660 ;
        RECT 51.235 1.480 51.755 1.660 ;
        RECT 52.045 1.660 52.345 1.850 ;
        RECT 53.455 1.660 53.755 2.030 ;
        RECT 52.045 1.480 52.565 1.660 ;
        RECT 53.235 1.480 53.755 1.660 ;
        RECT 54.045 1.660 54.345 1.850 ;
        RECT 55.455 1.660 55.755 2.030 ;
        RECT 54.045 1.480 54.565 1.660 ;
        RECT 55.235 1.480 55.755 1.660 ;
        RECT 56.045 1.660 56.345 1.850 ;
        RECT 57.455 1.660 57.755 2.030 ;
        RECT 56.045 1.480 56.565 1.660 ;
        RECT 57.235 1.480 57.755 1.660 ;
        RECT 58.045 1.660 58.345 1.850 ;
        RECT 59.455 1.660 59.755 2.030 ;
        RECT 58.045 1.480 58.565 1.660 ;
        RECT 59.235 1.480 59.755 1.660 ;
        RECT 60.045 1.660 60.345 1.850 ;
        RECT 61.455 1.660 61.755 2.030 ;
        RECT 60.045 1.480 60.565 1.660 ;
        RECT 61.235 1.480 61.755 1.660 ;
        RECT 62.045 1.660 62.345 1.850 ;
        RECT 63.455 1.660 63.755 2.030 ;
        RECT 62.045 1.480 62.565 1.660 ;
        RECT 63.235 1.480 63.755 1.660 ;
        RECT 64.045 1.660 64.345 1.850 ;
        RECT 65.455 1.660 65.755 2.030 ;
        RECT 64.045 1.480 64.565 1.660 ;
        RECT 65.235 1.480 65.755 1.660 ;
        RECT 66.045 1.660 66.345 1.850 ;
        RECT 67.455 1.660 67.755 2.030 ;
        RECT 66.045 1.480 66.565 1.660 ;
        RECT 67.235 1.480 67.755 1.660 ;
        RECT 68.045 1.660 68.345 1.850 ;
        RECT 69.455 1.660 69.755 2.030 ;
        RECT 68.045 1.480 68.565 1.660 ;
        RECT 69.235 1.480 69.755 1.660 ;
        RECT 70.045 1.660 70.345 1.850 ;
        RECT 71.455 1.660 71.755 2.030 ;
        RECT 70.045 1.480 70.565 1.660 ;
        RECT 71.235 1.480 71.755 1.660 ;
        RECT 72.045 1.660 72.345 1.850 ;
        RECT 73.455 1.660 73.755 2.030 ;
        RECT 72.045 1.480 72.565 1.660 ;
        RECT 73.235 1.480 73.755 1.660 ;
        RECT 74.045 1.660 74.345 1.850 ;
        RECT 75.455 1.660 75.755 2.030 ;
        RECT 74.045 1.480 74.565 1.660 ;
        RECT 75.235 1.480 75.755 1.660 ;
        RECT 76.045 1.660 76.345 1.850 ;
        RECT 77.455 1.660 77.755 2.030 ;
        RECT 76.045 1.480 76.565 1.660 ;
        RECT 77.235 1.480 77.755 1.660 ;
        RECT 78.045 1.660 78.345 1.850 ;
        RECT 79.455 1.660 79.755 2.030 ;
        RECT 78.045 1.480 78.565 1.660 ;
        RECT 79.235 1.480 79.755 1.660 ;
        RECT 80.045 1.660 80.345 1.850 ;
        RECT 81.455 1.660 81.755 2.030 ;
        RECT 80.045 1.480 80.565 1.660 ;
        RECT 81.235 1.480 81.755 1.660 ;
        RECT 82.045 1.660 82.345 1.850 ;
        RECT 83.455 1.660 83.755 2.030 ;
        RECT 82.045 1.480 82.565 1.660 ;
        RECT 83.235 1.480 83.755 1.660 ;
        RECT 84.045 1.660 84.345 1.850 ;
        RECT 85.455 1.660 85.755 2.030 ;
        RECT 84.045 1.480 84.565 1.660 ;
        RECT 85.235 1.480 85.755 1.660 ;
        RECT 86.045 1.660 86.345 1.850 ;
        RECT 87.455 1.660 87.755 2.030 ;
        RECT 86.045 1.480 86.565 1.660 ;
        RECT 87.235 1.480 87.755 1.660 ;
        RECT 88.045 1.660 88.345 1.850 ;
        RECT 89.455 1.660 89.755 2.030 ;
        RECT 88.045 1.480 88.565 1.660 ;
        RECT 89.235 1.480 89.755 1.660 ;
        RECT 90.045 1.660 90.345 1.850 ;
        RECT 91.455 1.660 91.755 2.030 ;
        RECT 90.045 1.480 90.565 1.660 ;
        RECT 91.235 1.480 91.755 1.660 ;
        RECT 92.045 1.660 92.345 1.850 ;
        RECT 93.455 1.660 93.755 2.030 ;
        RECT 92.045 1.480 92.565 1.660 ;
        RECT 93.235 1.480 93.755 1.660 ;
        RECT 94.045 1.660 94.345 1.850 ;
        RECT 95.455 1.660 95.755 2.030 ;
        RECT 94.045 1.480 94.565 1.660 ;
        RECT 95.235 1.480 95.755 1.660 ;
        RECT 96.045 1.660 96.345 1.850 ;
        RECT 97.455 1.660 97.755 2.030 ;
        RECT 96.045 1.480 96.565 1.660 ;
        RECT 97.235 1.480 97.755 1.660 ;
        RECT 98.045 1.660 98.345 1.850 ;
        RECT 99.455 1.660 99.755 2.030 ;
        RECT 98.045 1.480 98.565 1.660 ;
        RECT 99.235 1.480 99.755 1.660 ;
        RECT 100.045 1.660 100.345 1.850 ;
        RECT 101.455 1.660 101.755 2.030 ;
        RECT 100.045 1.480 100.565 1.660 ;
        RECT 101.235 1.480 101.755 1.660 ;
        RECT 102.045 1.660 102.345 1.850 ;
        RECT 103.455 1.660 103.755 2.030 ;
        RECT 102.045 1.480 102.565 1.660 ;
        RECT 103.235 1.480 103.755 1.660 ;
        RECT 104.045 1.660 104.345 1.850 ;
        RECT 105.455 1.660 105.755 2.030 ;
        RECT 104.045 1.480 104.565 1.660 ;
        RECT 105.235 1.480 105.755 1.660 ;
        RECT 106.045 1.660 106.345 1.850 ;
        RECT 107.455 1.660 107.755 2.030 ;
        RECT 106.045 1.480 106.565 1.660 ;
        RECT 107.235 1.480 107.755 1.660 ;
        RECT 108.045 1.660 108.345 1.850 ;
        RECT 109.455 1.660 109.755 2.030 ;
        RECT 108.045 1.480 108.565 1.660 ;
        RECT 109.235 1.480 109.755 1.660 ;
        RECT 110.045 1.660 110.345 1.850 ;
        RECT 111.455 1.660 111.755 2.030 ;
        RECT 110.045 1.480 110.565 1.660 ;
        RECT 111.235 1.480 111.755 1.660 ;
        RECT 112.045 1.660 112.345 1.850 ;
        RECT 113.455 1.660 113.755 2.030 ;
        RECT 112.045 1.480 112.565 1.660 ;
        RECT 113.235 1.480 113.755 1.660 ;
        RECT 114.045 1.660 114.345 1.850 ;
        RECT 115.455 1.660 115.755 2.030 ;
        RECT 114.045 1.480 114.565 1.660 ;
        RECT 115.235 1.480 115.755 1.660 ;
        RECT 116.045 1.660 116.345 1.850 ;
        RECT 117.455 1.660 117.755 2.030 ;
        RECT 116.045 1.480 116.565 1.660 ;
        RECT 117.235 1.480 117.755 1.660 ;
        RECT 118.045 1.660 118.345 1.850 ;
        RECT 119.455 1.660 119.755 2.030 ;
        RECT 118.045 1.480 118.565 1.660 ;
        RECT 119.235 1.480 119.755 1.660 ;
        RECT 120.045 1.660 120.345 1.850 ;
        RECT 121.455 1.660 121.755 2.030 ;
        RECT 120.045 1.480 120.565 1.660 ;
        RECT 121.235 1.480 121.755 1.660 ;
        RECT 122.045 1.660 122.345 1.850 ;
        RECT 123.455 1.660 123.755 2.030 ;
        RECT 122.045 1.480 122.565 1.660 ;
        RECT 123.235 1.480 123.755 1.660 ;
        RECT 124.045 1.660 124.345 1.850 ;
        RECT 125.455 1.660 125.755 2.030 ;
        RECT 124.045 1.480 124.565 1.660 ;
        RECT 125.235 1.480 125.755 1.660 ;
        RECT 126.045 1.660 126.345 1.850 ;
        RECT 127.455 1.660 127.755 2.030 ;
        RECT 126.045 1.480 126.565 1.660 ;
        RECT 127.235 1.480 127.755 1.660 ;
        RECT 128.045 1.660 128.345 1.850 ;
        RECT 129.455 1.660 129.755 2.030 ;
        RECT 128.045 1.480 128.565 1.660 ;
        RECT 129.235 1.480 129.755 1.660 ;
        RECT 130.045 1.660 130.345 1.850 ;
        RECT 131.455 1.660 131.755 2.030 ;
        RECT 130.045 1.480 130.565 1.660 ;
        RECT 131.235 1.480 131.755 1.660 ;
        RECT 132.045 1.660 132.345 1.850 ;
        RECT 132.045 1.480 132.565 1.660 ;
        RECT 1.235 1.150 1.755 1.330 ;
        RECT 2.045 1.150 2.565 1.330 ;
        RECT 3.235 1.150 3.755 1.330 ;
        RECT 4.045 1.150 4.565 1.330 ;
        RECT 5.235 1.150 5.755 1.330 ;
        RECT 6.045 1.150 6.565 1.330 ;
        RECT 7.235 1.150 7.755 1.330 ;
        RECT 8.045 1.150 8.565 1.330 ;
        RECT 9.235 1.150 9.755 1.330 ;
        RECT 10.045 1.150 10.565 1.330 ;
        RECT 11.235 1.150 11.755 1.330 ;
        RECT 12.045 1.150 12.565 1.330 ;
        RECT 13.235 1.150 13.755 1.330 ;
        RECT 14.045 1.150 14.565 1.330 ;
        RECT 15.235 1.150 15.755 1.330 ;
        RECT 16.045 1.150 16.565 1.330 ;
        RECT 17.235 1.150 17.755 1.330 ;
        RECT 18.045 1.150 18.565 1.330 ;
        RECT 19.235 1.150 19.755 1.330 ;
        RECT 20.045 1.150 20.565 1.330 ;
        RECT 21.235 1.150 21.755 1.330 ;
        RECT 22.045 1.150 22.565 1.330 ;
        RECT 23.235 1.150 23.755 1.330 ;
        RECT 24.045 1.150 24.565 1.330 ;
        RECT 25.235 1.150 25.755 1.330 ;
        RECT 26.045 1.150 26.565 1.330 ;
        RECT 27.235 1.150 27.755 1.330 ;
        RECT 28.045 1.150 28.565 1.330 ;
        RECT 29.235 1.150 29.755 1.330 ;
        RECT 30.045 1.150 30.565 1.330 ;
        RECT 31.235 1.150 31.755 1.330 ;
        RECT 32.045 1.150 32.565 1.330 ;
        RECT 33.235 1.150 33.755 1.330 ;
        RECT 34.045 1.150 34.565 1.330 ;
        RECT 35.235 1.150 35.755 1.330 ;
        RECT 36.045 1.150 36.565 1.330 ;
        RECT 37.235 1.150 37.755 1.330 ;
        RECT 38.045 1.150 38.565 1.330 ;
        RECT 39.235 1.150 39.755 1.330 ;
        RECT 40.045 1.150 40.565 1.330 ;
        RECT 41.235 1.150 41.755 1.330 ;
        RECT 42.045 1.150 42.565 1.330 ;
        RECT 43.235 1.150 43.755 1.330 ;
        RECT 44.045 1.150 44.565 1.330 ;
        RECT 45.235 1.150 45.755 1.330 ;
        RECT 46.045 1.150 46.565 1.330 ;
        RECT 47.235 1.150 47.755 1.330 ;
        RECT 48.045 1.150 48.565 1.330 ;
        RECT 49.235 1.150 49.755 1.330 ;
        RECT 50.045 1.150 50.565 1.330 ;
        RECT 51.235 1.150 51.755 1.330 ;
        RECT 52.045 1.150 52.565 1.330 ;
        RECT 53.235 1.150 53.755 1.330 ;
        RECT 54.045 1.150 54.565 1.330 ;
        RECT 55.235 1.150 55.755 1.330 ;
        RECT 56.045 1.150 56.565 1.330 ;
        RECT 57.235 1.150 57.755 1.330 ;
        RECT 58.045 1.150 58.565 1.330 ;
        RECT 59.235 1.150 59.755 1.330 ;
        RECT 60.045 1.150 60.565 1.330 ;
        RECT 61.235 1.150 61.755 1.330 ;
        RECT 62.045 1.150 62.565 1.330 ;
        RECT 63.235 1.150 63.755 1.330 ;
        RECT 64.045 1.150 64.565 1.330 ;
        RECT 65.235 1.150 65.755 1.330 ;
        RECT 66.045 1.150 66.565 1.330 ;
        RECT 67.235 1.150 67.755 1.330 ;
        RECT 68.045 1.150 68.565 1.330 ;
        RECT 69.235 1.150 69.755 1.330 ;
        RECT 70.045 1.150 70.565 1.330 ;
        RECT 71.235 1.150 71.755 1.330 ;
        RECT 72.045 1.150 72.565 1.330 ;
        RECT 73.235 1.150 73.755 1.330 ;
        RECT 74.045 1.150 74.565 1.330 ;
        RECT 75.235 1.150 75.755 1.330 ;
        RECT 76.045 1.150 76.565 1.330 ;
        RECT 77.235 1.150 77.755 1.330 ;
        RECT 78.045 1.150 78.565 1.330 ;
        RECT 79.235 1.150 79.755 1.330 ;
        RECT 80.045 1.150 80.565 1.330 ;
        RECT 81.235 1.150 81.755 1.330 ;
        RECT 82.045 1.150 82.565 1.330 ;
        RECT 83.235 1.150 83.755 1.330 ;
        RECT 84.045 1.150 84.565 1.330 ;
        RECT 85.235 1.150 85.755 1.330 ;
        RECT 86.045 1.150 86.565 1.330 ;
        RECT 87.235 1.150 87.755 1.330 ;
        RECT 88.045 1.150 88.565 1.330 ;
        RECT 89.235 1.150 89.755 1.330 ;
        RECT 90.045 1.150 90.565 1.330 ;
        RECT 91.235 1.150 91.755 1.330 ;
        RECT 92.045 1.150 92.565 1.330 ;
        RECT 93.235 1.150 93.755 1.330 ;
        RECT 94.045 1.150 94.565 1.330 ;
        RECT 95.235 1.150 95.755 1.330 ;
        RECT 96.045 1.150 96.565 1.330 ;
        RECT 97.235 1.150 97.755 1.330 ;
        RECT 98.045 1.150 98.565 1.330 ;
        RECT 99.235 1.150 99.755 1.330 ;
        RECT 100.045 1.150 100.565 1.330 ;
        RECT 101.235 1.150 101.755 1.330 ;
        RECT 102.045 1.150 102.565 1.330 ;
        RECT 103.235 1.150 103.755 1.330 ;
        RECT 104.045 1.150 104.565 1.330 ;
        RECT 105.235 1.150 105.755 1.330 ;
        RECT 106.045 1.150 106.565 1.330 ;
        RECT 107.235 1.150 107.755 1.330 ;
        RECT 108.045 1.150 108.565 1.330 ;
        RECT 109.235 1.150 109.755 1.330 ;
        RECT 110.045 1.150 110.565 1.330 ;
        RECT 111.235 1.150 111.755 1.330 ;
        RECT 112.045 1.150 112.565 1.330 ;
        RECT 113.235 1.150 113.755 1.330 ;
        RECT 114.045 1.150 114.565 1.330 ;
        RECT 115.235 1.150 115.755 1.330 ;
        RECT 116.045 1.150 116.565 1.330 ;
        RECT 117.235 1.150 117.755 1.330 ;
        RECT 118.045 1.150 118.565 1.330 ;
        RECT 119.235 1.150 119.755 1.330 ;
        RECT 120.045 1.150 120.565 1.330 ;
        RECT 121.235 1.150 121.755 1.330 ;
        RECT 122.045 1.150 122.565 1.330 ;
        RECT 123.235 1.150 123.755 1.330 ;
        RECT 124.045 1.150 124.565 1.330 ;
        RECT 125.235 1.150 125.755 1.330 ;
        RECT 126.045 1.150 126.565 1.330 ;
        RECT 127.235 1.150 127.755 1.330 ;
        RECT 128.045 1.150 128.565 1.330 ;
        RECT 129.235 1.150 129.755 1.330 ;
        RECT 130.045 1.150 130.565 1.330 ;
        RECT 131.235 1.150 131.755 1.330 ;
        RECT 132.045 1.150 132.565 1.330 ;
      LAYER Metal1 ;
        RECT 1.075 23.280 1.235 25.390 ;
        RECT 2.565 24.570 2.725 25.390 ;
        RECT 1.475 24.410 2.725 24.570 ;
        RECT 2.565 23.280 2.725 24.410 ;
        RECT 3.075 23.280 3.235 25.390 ;
        RECT 4.565 24.570 4.725 25.390 ;
        RECT 3.475 24.410 4.725 24.570 ;
        RECT 4.565 23.280 4.725 24.410 ;
        RECT 5.075 23.280 5.235 25.390 ;
        RECT 6.565 24.570 6.725 25.390 ;
        RECT 5.475 24.410 6.725 24.570 ;
        RECT 6.565 23.280 6.725 24.410 ;
        RECT 7.075 23.280 7.235 25.390 ;
        RECT 8.565 24.570 8.725 25.390 ;
        RECT 7.475 24.410 8.725 24.570 ;
        RECT 8.565 23.280 8.725 24.410 ;
        RECT 9.075 23.280 9.235 25.390 ;
        RECT 10.565 24.570 10.725 25.390 ;
        RECT 9.475 24.410 10.725 24.570 ;
        RECT 10.565 23.280 10.725 24.410 ;
        RECT 11.075 23.280 11.235 25.390 ;
        RECT 12.565 24.570 12.725 25.390 ;
        RECT 11.475 24.410 12.725 24.570 ;
        RECT 12.565 23.280 12.725 24.410 ;
        RECT 13.075 23.280 13.235 25.390 ;
        RECT 14.565 24.570 14.725 25.390 ;
        RECT 13.475 24.410 14.725 24.570 ;
        RECT 14.565 23.280 14.725 24.410 ;
        RECT 15.075 23.280 15.235 25.390 ;
        RECT 16.565 24.570 16.725 25.390 ;
        RECT 15.475 24.410 16.725 24.570 ;
        RECT 16.565 23.280 16.725 24.410 ;
        RECT 17.075 23.280 17.235 25.390 ;
        RECT 18.565 24.570 18.725 25.390 ;
        RECT 17.475 24.410 18.725 24.570 ;
        RECT 18.565 23.280 18.725 24.410 ;
        RECT 19.075 23.280 19.235 25.390 ;
        RECT 20.565 24.570 20.725 25.390 ;
        RECT 19.475 24.410 20.725 24.570 ;
        RECT 20.565 23.280 20.725 24.410 ;
        RECT 21.075 23.280 21.235 25.390 ;
        RECT 22.565 24.570 22.725 25.390 ;
        RECT 21.475 24.410 22.725 24.570 ;
        RECT 22.565 23.280 22.725 24.410 ;
        RECT 23.075 23.280 23.235 25.390 ;
        RECT 24.565 24.570 24.725 25.390 ;
        RECT 23.475 24.410 24.725 24.570 ;
        RECT 24.565 23.280 24.725 24.410 ;
        RECT 25.075 23.280 25.235 25.390 ;
        RECT 26.565 24.570 26.725 25.390 ;
        RECT 25.475 24.410 26.725 24.570 ;
        RECT 26.565 23.280 26.725 24.410 ;
        RECT 27.075 23.280 27.235 25.390 ;
        RECT 28.565 24.570 28.725 25.390 ;
        RECT 27.475 24.410 28.725 24.570 ;
        RECT 28.565 23.280 28.725 24.410 ;
        RECT 29.075 23.280 29.235 25.390 ;
        RECT 30.565 24.570 30.725 25.390 ;
        RECT 29.475 24.410 30.725 24.570 ;
        RECT 30.565 23.280 30.725 24.410 ;
        RECT 31.075 23.280 31.235 25.390 ;
        RECT 32.565 24.570 32.725 25.390 ;
        RECT 31.475 24.410 32.725 24.570 ;
        RECT 32.565 23.280 32.725 24.410 ;
        RECT 33.075 23.280 33.235 25.390 ;
        RECT 34.565 24.570 34.725 25.390 ;
        RECT 33.475 24.410 34.725 24.570 ;
        RECT 34.565 23.280 34.725 24.410 ;
        RECT 35.075 23.280 35.235 25.390 ;
        RECT 36.565 24.570 36.725 25.390 ;
        RECT 35.475 24.410 36.725 24.570 ;
        RECT 36.565 23.280 36.725 24.410 ;
        RECT 37.075 23.280 37.235 25.390 ;
        RECT 38.565 24.570 38.725 25.390 ;
        RECT 37.475 24.410 38.725 24.570 ;
        RECT 38.565 23.280 38.725 24.410 ;
        RECT 39.075 23.280 39.235 25.390 ;
        RECT 40.565 24.570 40.725 25.390 ;
        RECT 39.475 24.410 40.725 24.570 ;
        RECT 40.565 23.280 40.725 24.410 ;
        RECT 41.075 23.280 41.235 25.390 ;
        RECT 42.565 24.570 42.725 25.390 ;
        RECT 41.475 24.410 42.725 24.570 ;
        RECT 42.565 23.280 42.725 24.410 ;
        RECT 43.075 23.280 43.235 25.390 ;
        RECT 44.565 24.570 44.725 25.390 ;
        RECT 43.475 24.410 44.725 24.570 ;
        RECT 44.565 23.280 44.725 24.410 ;
        RECT 45.075 23.280 45.235 25.390 ;
        RECT 46.565 24.570 46.725 25.390 ;
        RECT 45.475 24.410 46.725 24.570 ;
        RECT 46.565 23.280 46.725 24.410 ;
        RECT 47.075 23.280 47.235 25.390 ;
        RECT 48.565 24.570 48.725 25.390 ;
        RECT 47.475 24.410 48.725 24.570 ;
        RECT 48.565 23.280 48.725 24.410 ;
        RECT 49.075 23.280 49.235 25.390 ;
        RECT 50.565 24.570 50.725 25.390 ;
        RECT 49.475 24.410 50.725 24.570 ;
        RECT 50.565 23.280 50.725 24.410 ;
        RECT 51.075 23.280 51.235 25.390 ;
        RECT 52.565 24.570 52.725 25.390 ;
        RECT 51.475 24.410 52.725 24.570 ;
        RECT 52.565 23.280 52.725 24.410 ;
        RECT 53.075 23.280 53.235 25.390 ;
        RECT 54.565 24.570 54.725 25.390 ;
        RECT 53.475 24.410 54.725 24.570 ;
        RECT 54.565 23.280 54.725 24.410 ;
        RECT 55.075 23.280 55.235 25.390 ;
        RECT 56.565 24.570 56.725 25.390 ;
        RECT 55.475 24.410 56.725 24.570 ;
        RECT 56.565 23.280 56.725 24.410 ;
        RECT 57.075 23.280 57.235 25.390 ;
        RECT 58.565 24.570 58.725 25.390 ;
        RECT 57.475 24.410 58.725 24.570 ;
        RECT 58.565 23.280 58.725 24.410 ;
        RECT 59.075 23.280 59.235 25.390 ;
        RECT 60.565 24.570 60.725 25.390 ;
        RECT 59.475 24.410 60.725 24.570 ;
        RECT 60.565 23.280 60.725 24.410 ;
        RECT 61.075 23.280 61.235 25.390 ;
        RECT 62.565 24.570 62.725 25.390 ;
        RECT 61.475 24.410 62.725 24.570 ;
        RECT 62.565 23.280 62.725 24.410 ;
        RECT 63.075 23.280 63.235 25.390 ;
        RECT 64.565 24.570 64.725 25.390 ;
        RECT 63.475 24.410 64.725 24.570 ;
        RECT 64.565 23.280 64.725 24.410 ;
        RECT 65.075 23.280 65.235 25.390 ;
        RECT 66.565 24.570 66.725 25.390 ;
        RECT 65.475 24.410 66.725 24.570 ;
        RECT 66.565 23.280 66.725 24.410 ;
        RECT 67.075 23.280 67.235 25.390 ;
        RECT 68.565 24.570 68.725 25.390 ;
        RECT 67.475 24.410 68.725 24.570 ;
        RECT 68.565 23.280 68.725 24.410 ;
        RECT 69.075 23.280 69.235 25.390 ;
        RECT 70.565 24.570 70.725 25.390 ;
        RECT 69.475 24.410 70.725 24.570 ;
        RECT 70.565 23.280 70.725 24.410 ;
        RECT 71.075 23.280 71.235 25.390 ;
        RECT 72.565 24.570 72.725 25.390 ;
        RECT 71.475 24.410 72.725 24.570 ;
        RECT 72.565 23.280 72.725 24.410 ;
        RECT 73.075 23.280 73.235 25.390 ;
        RECT 74.565 24.570 74.725 25.390 ;
        RECT 73.475 24.410 74.725 24.570 ;
        RECT 74.565 23.280 74.725 24.410 ;
        RECT 75.075 23.280 75.235 25.390 ;
        RECT 76.565 24.570 76.725 25.390 ;
        RECT 75.475 24.410 76.725 24.570 ;
        RECT 76.565 23.280 76.725 24.410 ;
        RECT 77.075 23.280 77.235 25.390 ;
        RECT 78.565 24.570 78.725 25.390 ;
        RECT 77.475 24.410 78.725 24.570 ;
        RECT 78.565 23.280 78.725 24.410 ;
        RECT 79.075 23.280 79.235 25.390 ;
        RECT 80.565 24.570 80.725 25.390 ;
        RECT 79.475 24.410 80.725 24.570 ;
        RECT 80.565 23.280 80.725 24.410 ;
        RECT 81.075 23.280 81.235 25.390 ;
        RECT 82.565 24.570 82.725 25.390 ;
        RECT 81.475 24.410 82.725 24.570 ;
        RECT 82.565 23.280 82.725 24.410 ;
        RECT 83.075 23.280 83.235 25.390 ;
        RECT 84.565 24.570 84.725 25.390 ;
        RECT 83.475 24.410 84.725 24.570 ;
        RECT 84.565 23.280 84.725 24.410 ;
        RECT 85.075 23.280 85.235 25.390 ;
        RECT 86.565 24.570 86.725 25.390 ;
        RECT 85.475 24.410 86.725 24.570 ;
        RECT 86.565 23.280 86.725 24.410 ;
        RECT 87.075 23.280 87.235 25.390 ;
        RECT 88.565 24.570 88.725 25.390 ;
        RECT 87.475 24.410 88.725 24.570 ;
        RECT 88.565 23.280 88.725 24.410 ;
        RECT 89.075 23.280 89.235 25.390 ;
        RECT 90.565 24.570 90.725 25.390 ;
        RECT 89.475 24.410 90.725 24.570 ;
        RECT 90.565 23.280 90.725 24.410 ;
        RECT 91.075 23.280 91.235 25.390 ;
        RECT 92.565 24.570 92.725 25.390 ;
        RECT 91.475 24.410 92.725 24.570 ;
        RECT 92.565 23.280 92.725 24.410 ;
        RECT 93.075 23.280 93.235 25.390 ;
        RECT 94.565 24.570 94.725 25.390 ;
        RECT 93.475 24.410 94.725 24.570 ;
        RECT 94.565 23.280 94.725 24.410 ;
        RECT 95.075 23.280 95.235 25.390 ;
        RECT 96.565 24.570 96.725 25.390 ;
        RECT 95.475 24.410 96.725 24.570 ;
        RECT 96.565 23.280 96.725 24.410 ;
        RECT 97.075 23.280 97.235 25.390 ;
        RECT 98.565 24.570 98.725 25.390 ;
        RECT 97.475 24.410 98.725 24.570 ;
        RECT 98.565 23.280 98.725 24.410 ;
        RECT 99.075 23.280 99.235 25.390 ;
        RECT 100.565 24.570 100.725 25.390 ;
        RECT 99.475 24.410 100.725 24.570 ;
        RECT 100.565 23.280 100.725 24.410 ;
        RECT 101.075 23.280 101.235 25.390 ;
        RECT 102.565 24.570 102.725 25.390 ;
        RECT 101.475 24.410 102.725 24.570 ;
        RECT 102.565 23.280 102.725 24.410 ;
        RECT 103.075 23.280 103.235 25.390 ;
        RECT 104.565 24.570 104.725 25.390 ;
        RECT 103.475 24.410 104.725 24.570 ;
        RECT 104.565 23.280 104.725 24.410 ;
        RECT 105.075 23.280 105.235 25.390 ;
        RECT 106.565 24.570 106.725 25.390 ;
        RECT 105.475 24.410 106.725 24.570 ;
        RECT 106.565 23.280 106.725 24.410 ;
        RECT 107.075 23.280 107.235 25.390 ;
        RECT 108.565 24.570 108.725 25.390 ;
        RECT 107.475 24.410 108.725 24.570 ;
        RECT 108.565 23.280 108.725 24.410 ;
        RECT 109.075 23.280 109.235 25.390 ;
        RECT 110.565 24.570 110.725 25.390 ;
        RECT 109.475 24.410 110.725 24.570 ;
        RECT 110.565 23.280 110.725 24.410 ;
        RECT 111.075 23.280 111.235 25.390 ;
        RECT 112.565 24.570 112.725 25.390 ;
        RECT 111.475 24.410 112.725 24.570 ;
        RECT 112.565 23.280 112.725 24.410 ;
        RECT 113.075 23.280 113.235 25.390 ;
        RECT 114.565 24.570 114.725 25.390 ;
        RECT 113.475 24.410 114.725 24.570 ;
        RECT 114.565 23.280 114.725 24.410 ;
        RECT 115.075 23.280 115.235 25.390 ;
        RECT 116.565 24.570 116.725 25.390 ;
        RECT 115.475 24.410 116.725 24.570 ;
        RECT 116.565 23.280 116.725 24.410 ;
        RECT 117.075 23.280 117.235 25.390 ;
        RECT 118.565 24.570 118.725 25.390 ;
        RECT 117.475 24.410 118.725 24.570 ;
        RECT 118.565 23.280 118.725 24.410 ;
        RECT 119.075 23.280 119.235 25.390 ;
        RECT 120.565 24.570 120.725 25.390 ;
        RECT 119.475 24.410 120.725 24.570 ;
        RECT 120.565 23.280 120.725 24.410 ;
        RECT 121.075 23.280 121.235 25.390 ;
        RECT 122.565 24.570 122.725 25.390 ;
        RECT 121.475 24.410 122.725 24.570 ;
        RECT 122.565 23.280 122.725 24.410 ;
        RECT 123.075 23.280 123.235 25.390 ;
        RECT 124.565 24.570 124.725 25.390 ;
        RECT 123.475 24.410 124.725 24.570 ;
        RECT 124.565 23.280 124.725 24.410 ;
        RECT 125.075 23.280 125.235 25.390 ;
        RECT 126.565 24.570 126.725 25.390 ;
        RECT 125.475 24.410 126.725 24.570 ;
        RECT 126.565 23.280 126.725 24.410 ;
        RECT 127.075 23.280 127.235 25.390 ;
        RECT 128.565 24.570 128.725 25.390 ;
        RECT 127.475 24.410 128.725 24.570 ;
        RECT 128.565 23.280 128.725 24.410 ;
        RECT 129.075 23.280 129.235 25.390 ;
        RECT 130.565 24.570 130.725 25.390 ;
        RECT 129.475 24.410 130.725 24.570 ;
        RECT 130.565 23.280 130.725 24.410 ;
        RECT 131.075 23.280 131.235 25.390 ;
        RECT 132.565 24.570 132.725 25.390 ;
        RECT 131.475 24.410 132.725 24.570 ;
        RECT 132.565 23.280 132.725 24.410 ;
        RECT 1.010 22.990 1.300 23.280 ;
        RECT 2.500 22.990 2.790 23.280 ;
        RECT 3.010 22.990 3.300 23.280 ;
        RECT 4.500 22.990 4.790 23.280 ;
        RECT 5.010 22.990 5.300 23.280 ;
        RECT 6.500 22.990 6.790 23.280 ;
        RECT 7.010 22.990 7.300 23.280 ;
        RECT 8.500 22.990 8.790 23.280 ;
        RECT 9.010 22.990 9.300 23.280 ;
        RECT 10.500 22.990 10.790 23.280 ;
        RECT 11.010 22.990 11.300 23.280 ;
        RECT 12.500 22.990 12.790 23.280 ;
        RECT 13.010 22.990 13.300 23.280 ;
        RECT 14.500 22.990 14.790 23.280 ;
        RECT 15.010 22.990 15.300 23.280 ;
        RECT 16.500 22.990 16.790 23.280 ;
        RECT 17.010 22.990 17.300 23.280 ;
        RECT 18.500 22.990 18.790 23.280 ;
        RECT 19.010 22.990 19.300 23.280 ;
        RECT 20.500 22.990 20.790 23.280 ;
        RECT 21.010 22.990 21.300 23.280 ;
        RECT 22.500 22.990 22.790 23.280 ;
        RECT 23.010 22.990 23.300 23.280 ;
        RECT 24.500 22.990 24.790 23.280 ;
        RECT 25.010 22.990 25.300 23.280 ;
        RECT 26.500 22.990 26.790 23.280 ;
        RECT 27.010 22.990 27.300 23.280 ;
        RECT 28.500 22.990 28.790 23.280 ;
        RECT 29.010 22.990 29.300 23.280 ;
        RECT 30.500 22.990 30.790 23.280 ;
        RECT 31.010 22.990 31.300 23.280 ;
        RECT 32.500 22.990 32.790 23.280 ;
        RECT 33.010 22.990 33.300 23.280 ;
        RECT 34.500 22.990 34.790 23.280 ;
        RECT 35.010 22.990 35.300 23.280 ;
        RECT 36.500 22.990 36.790 23.280 ;
        RECT 37.010 22.990 37.300 23.280 ;
        RECT 38.500 22.990 38.790 23.280 ;
        RECT 39.010 22.990 39.300 23.280 ;
        RECT 40.500 22.990 40.790 23.280 ;
        RECT 41.010 22.990 41.300 23.280 ;
        RECT 42.500 22.990 42.790 23.280 ;
        RECT 43.010 22.990 43.300 23.280 ;
        RECT 44.500 22.990 44.790 23.280 ;
        RECT 45.010 22.990 45.300 23.280 ;
        RECT 46.500 22.990 46.790 23.280 ;
        RECT 47.010 22.990 47.300 23.280 ;
        RECT 48.500 22.990 48.790 23.280 ;
        RECT 49.010 22.990 49.300 23.280 ;
        RECT 50.500 22.990 50.790 23.280 ;
        RECT 51.010 22.990 51.300 23.280 ;
        RECT 52.500 22.990 52.790 23.280 ;
        RECT 53.010 22.990 53.300 23.280 ;
        RECT 54.500 22.990 54.790 23.280 ;
        RECT 55.010 22.990 55.300 23.280 ;
        RECT 56.500 22.990 56.790 23.280 ;
        RECT 57.010 22.990 57.300 23.280 ;
        RECT 58.500 22.990 58.790 23.280 ;
        RECT 59.010 22.990 59.300 23.280 ;
        RECT 60.500 22.990 60.790 23.280 ;
        RECT 61.010 22.990 61.300 23.280 ;
        RECT 62.500 22.990 62.790 23.280 ;
        RECT 63.010 22.990 63.300 23.280 ;
        RECT 64.500 22.990 64.790 23.280 ;
        RECT 65.010 22.990 65.300 23.280 ;
        RECT 66.500 22.990 66.790 23.280 ;
        RECT 67.010 22.990 67.300 23.280 ;
        RECT 68.500 22.990 68.790 23.280 ;
        RECT 69.010 22.990 69.300 23.280 ;
        RECT 70.500 22.990 70.790 23.280 ;
        RECT 71.010 22.990 71.300 23.280 ;
        RECT 72.500 22.990 72.790 23.280 ;
        RECT 73.010 22.990 73.300 23.280 ;
        RECT 74.500 22.990 74.790 23.280 ;
        RECT 75.010 22.990 75.300 23.280 ;
        RECT 76.500 22.990 76.790 23.280 ;
        RECT 77.010 22.990 77.300 23.280 ;
        RECT 78.500 22.990 78.790 23.280 ;
        RECT 79.010 22.990 79.300 23.280 ;
        RECT 80.500 22.990 80.790 23.280 ;
        RECT 81.010 22.990 81.300 23.280 ;
        RECT 82.500 22.990 82.790 23.280 ;
        RECT 83.010 22.990 83.300 23.280 ;
        RECT 84.500 22.990 84.790 23.280 ;
        RECT 85.010 22.990 85.300 23.280 ;
        RECT 86.500 22.990 86.790 23.280 ;
        RECT 87.010 22.990 87.300 23.280 ;
        RECT 88.500 22.990 88.790 23.280 ;
        RECT 89.010 22.990 89.300 23.280 ;
        RECT 90.500 22.990 90.790 23.280 ;
        RECT 91.010 22.990 91.300 23.280 ;
        RECT 92.500 22.990 92.790 23.280 ;
        RECT 93.010 22.990 93.300 23.280 ;
        RECT 94.500 22.990 94.790 23.280 ;
        RECT 95.010 22.990 95.300 23.280 ;
        RECT 96.500 22.990 96.790 23.280 ;
        RECT 97.010 22.990 97.300 23.280 ;
        RECT 98.500 22.990 98.790 23.280 ;
        RECT 99.010 22.990 99.300 23.280 ;
        RECT 100.500 22.990 100.790 23.280 ;
        RECT 101.010 22.990 101.300 23.280 ;
        RECT 102.500 22.990 102.790 23.280 ;
        RECT 103.010 22.990 103.300 23.280 ;
        RECT 104.500 22.990 104.790 23.280 ;
        RECT 105.010 22.990 105.300 23.280 ;
        RECT 106.500 22.990 106.790 23.280 ;
        RECT 107.010 22.990 107.300 23.280 ;
        RECT 108.500 22.990 108.790 23.280 ;
        RECT 109.010 22.990 109.300 23.280 ;
        RECT 110.500 22.990 110.790 23.280 ;
        RECT 111.010 22.990 111.300 23.280 ;
        RECT 112.500 22.990 112.790 23.280 ;
        RECT 113.010 22.990 113.300 23.280 ;
        RECT 114.500 22.990 114.790 23.280 ;
        RECT 115.010 22.990 115.300 23.280 ;
        RECT 116.500 22.990 116.790 23.280 ;
        RECT 117.010 22.990 117.300 23.280 ;
        RECT 118.500 22.990 118.790 23.280 ;
        RECT 119.010 22.990 119.300 23.280 ;
        RECT 120.500 22.990 120.790 23.280 ;
        RECT 121.010 22.990 121.300 23.280 ;
        RECT 122.500 22.990 122.790 23.280 ;
        RECT 123.010 22.990 123.300 23.280 ;
        RECT 124.500 22.990 124.790 23.280 ;
        RECT 125.010 22.990 125.300 23.280 ;
        RECT 126.500 22.990 126.790 23.280 ;
        RECT 127.010 22.990 127.300 23.280 ;
        RECT 128.500 22.990 128.790 23.280 ;
        RECT 129.010 22.990 129.300 23.280 ;
        RECT 130.500 22.990 130.790 23.280 ;
        RECT 131.010 22.990 131.300 23.280 ;
        RECT 132.500 22.990 132.790 23.280 ;
        RECT 1.410 21.630 1.710 21.930 ;
        RECT 2.090 21.630 2.390 21.930 ;
        RECT 3.410 21.630 3.710 21.930 ;
        RECT 4.090 21.630 4.390 21.930 ;
        RECT 5.410 21.630 5.710 21.930 ;
        RECT 6.090 21.630 6.390 21.930 ;
        RECT 7.410 21.630 7.710 21.930 ;
        RECT 8.090 21.630 8.390 21.930 ;
        RECT 9.410 21.630 9.710 21.930 ;
        RECT 10.090 21.630 10.390 21.930 ;
        RECT 11.410 21.630 11.710 21.930 ;
        RECT 12.090 21.630 12.390 21.930 ;
        RECT 13.410 21.630 13.710 21.930 ;
        RECT 14.090 21.630 14.390 21.930 ;
        RECT 15.410 21.630 15.710 21.930 ;
        RECT 16.090 21.630 16.390 21.930 ;
        RECT 17.410 21.630 17.710 21.930 ;
        RECT 18.090 21.630 18.390 21.930 ;
        RECT 19.410 21.630 19.710 21.930 ;
        RECT 20.090 21.630 20.390 21.930 ;
        RECT 21.410 21.630 21.710 21.930 ;
        RECT 22.090 21.630 22.390 21.930 ;
        RECT 23.410 21.630 23.710 21.930 ;
        RECT 24.090 21.630 24.390 21.930 ;
        RECT 25.410 21.630 25.710 21.930 ;
        RECT 26.090 21.630 26.390 21.930 ;
        RECT 27.410 21.630 27.710 21.930 ;
        RECT 28.090 21.630 28.390 21.930 ;
        RECT 29.410 21.630 29.710 21.930 ;
        RECT 30.090 21.630 30.390 21.930 ;
        RECT 31.410 21.630 31.710 21.930 ;
        RECT 32.090 21.630 32.390 21.930 ;
        RECT 33.410 21.630 33.710 21.930 ;
        RECT 34.090 21.630 34.390 21.930 ;
        RECT 35.410 21.630 35.710 21.930 ;
        RECT 36.090 21.630 36.390 21.930 ;
        RECT 37.410 21.630 37.710 21.930 ;
        RECT 38.090 21.630 38.390 21.930 ;
        RECT 39.410 21.630 39.710 21.930 ;
        RECT 40.090 21.630 40.390 21.930 ;
        RECT 41.410 21.630 41.710 21.930 ;
        RECT 42.090 21.630 42.390 21.930 ;
        RECT 43.410 21.630 43.710 21.930 ;
        RECT 44.090 21.630 44.390 21.930 ;
        RECT 45.410 21.630 45.710 21.930 ;
        RECT 46.090 21.630 46.390 21.930 ;
        RECT 47.410 21.630 47.710 21.930 ;
        RECT 48.090 21.630 48.390 21.930 ;
        RECT 49.410 21.630 49.710 21.930 ;
        RECT 50.090 21.630 50.390 21.930 ;
        RECT 51.410 21.630 51.710 21.930 ;
        RECT 52.090 21.630 52.390 21.930 ;
        RECT 53.410 21.630 53.710 21.930 ;
        RECT 54.090 21.630 54.390 21.930 ;
        RECT 55.410 21.630 55.710 21.930 ;
        RECT 56.090 21.630 56.390 21.930 ;
        RECT 57.410 21.630 57.710 21.930 ;
        RECT 58.090 21.630 58.390 21.930 ;
        RECT 59.410 21.630 59.710 21.930 ;
        RECT 60.090 21.630 60.390 21.930 ;
        RECT 61.410 21.630 61.710 21.930 ;
        RECT 62.090 21.630 62.390 21.930 ;
        RECT 63.410 21.630 63.710 21.930 ;
        RECT 64.090 21.630 64.390 21.930 ;
        RECT 65.410 21.630 65.710 21.930 ;
        RECT 66.090 21.630 66.390 21.930 ;
        RECT 67.410 21.630 67.710 21.930 ;
        RECT 68.090 21.630 68.390 21.930 ;
        RECT 69.410 21.630 69.710 21.930 ;
        RECT 70.090 21.630 70.390 21.930 ;
        RECT 71.410 21.630 71.710 21.930 ;
        RECT 72.090 21.630 72.390 21.930 ;
        RECT 73.410 21.630 73.710 21.930 ;
        RECT 74.090 21.630 74.390 21.930 ;
        RECT 75.410 21.630 75.710 21.930 ;
        RECT 76.090 21.630 76.390 21.930 ;
        RECT 77.410 21.630 77.710 21.930 ;
        RECT 78.090 21.630 78.390 21.930 ;
        RECT 79.410 21.630 79.710 21.930 ;
        RECT 80.090 21.630 80.390 21.930 ;
        RECT 81.410 21.630 81.710 21.930 ;
        RECT 82.090 21.630 82.390 21.930 ;
        RECT 83.410 21.630 83.710 21.930 ;
        RECT 84.090 21.630 84.390 21.930 ;
        RECT 85.410 21.630 85.710 21.930 ;
        RECT 86.090 21.630 86.390 21.930 ;
        RECT 87.410 21.630 87.710 21.930 ;
        RECT 88.090 21.630 88.390 21.930 ;
        RECT 89.410 21.630 89.710 21.930 ;
        RECT 90.090 21.630 90.390 21.930 ;
        RECT 91.410 21.630 91.710 21.930 ;
        RECT 92.090 21.630 92.390 21.930 ;
        RECT 93.410 21.630 93.710 21.930 ;
        RECT 94.090 21.630 94.390 21.930 ;
        RECT 95.410 21.630 95.710 21.930 ;
        RECT 96.090 21.630 96.390 21.930 ;
        RECT 97.410 21.630 97.710 21.930 ;
        RECT 98.090 21.630 98.390 21.930 ;
        RECT 99.410 21.630 99.710 21.930 ;
        RECT 100.090 21.630 100.390 21.930 ;
        RECT 101.410 21.630 101.710 21.930 ;
        RECT 102.090 21.630 102.390 21.930 ;
        RECT 103.410 21.630 103.710 21.930 ;
        RECT 104.090 21.630 104.390 21.930 ;
        RECT 105.410 21.630 105.710 21.930 ;
        RECT 106.090 21.630 106.390 21.930 ;
        RECT 107.410 21.630 107.710 21.930 ;
        RECT 108.090 21.630 108.390 21.930 ;
        RECT 109.410 21.630 109.710 21.930 ;
        RECT 110.090 21.630 110.390 21.930 ;
        RECT 111.410 21.630 111.710 21.930 ;
        RECT 112.090 21.630 112.390 21.930 ;
        RECT 113.410 21.630 113.710 21.930 ;
        RECT 114.090 21.630 114.390 21.930 ;
        RECT 115.410 21.630 115.710 21.930 ;
        RECT 116.090 21.630 116.390 21.930 ;
        RECT 117.410 21.630 117.710 21.930 ;
        RECT 118.090 21.630 118.390 21.930 ;
        RECT 119.410 21.630 119.710 21.930 ;
        RECT 120.090 21.630 120.390 21.930 ;
        RECT 121.410 21.630 121.710 21.930 ;
        RECT 122.090 21.630 122.390 21.930 ;
        RECT 123.410 21.630 123.710 21.930 ;
        RECT 124.090 21.630 124.390 21.930 ;
        RECT 125.410 21.630 125.710 21.930 ;
        RECT 126.090 21.630 126.390 21.930 ;
        RECT 127.410 21.630 127.710 21.930 ;
        RECT 128.090 21.630 128.390 21.930 ;
        RECT 129.410 21.630 129.710 21.930 ;
        RECT 130.090 21.630 130.390 21.930 ;
        RECT 131.410 21.630 131.710 21.930 ;
        RECT 132.090 21.630 132.390 21.930 ;
        RECT 1.750 21.130 2.050 21.430 ;
        RECT 3.750 21.130 4.050 21.430 ;
        RECT 5.750 21.130 6.050 21.430 ;
        RECT 7.750 21.130 8.050 21.430 ;
        RECT 9.750 21.130 10.050 21.430 ;
        RECT 11.750 21.130 12.050 21.430 ;
        RECT 13.750 21.130 14.050 21.430 ;
        RECT 15.750 21.130 16.050 21.430 ;
        RECT 17.750 21.130 18.050 21.430 ;
        RECT 19.750 21.130 20.050 21.430 ;
        RECT 21.750 21.130 22.050 21.430 ;
        RECT 23.750 21.130 24.050 21.430 ;
        RECT 25.750 21.130 26.050 21.430 ;
        RECT 27.750 21.130 28.050 21.430 ;
        RECT 29.750 21.130 30.050 21.430 ;
        RECT 31.750 21.130 32.050 21.430 ;
        RECT 33.750 21.130 34.050 21.430 ;
        RECT 35.750 21.130 36.050 21.430 ;
        RECT 37.750 21.130 38.050 21.430 ;
        RECT 39.750 21.130 40.050 21.430 ;
        RECT 41.750 21.130 42.050 21.430 ;
        RECT 43.750 21.130 44.050 21.430 ;
        RECT 45.750 21.130 46.050 21.430 ;
        RECT 47.750 21.130 48.050 21.430 ;
        RECT 49.750 21.130 50.050 21.430 ;
        RECT 51.750 21.130 52.050 21.430 ;
        RECT 53.750 21.130 54.050 21.430 ;
        RECT 55.750 21.130 56.050 21.430 ;
        RECT 57.750 21.130 58.050 21.430 ;
        RECT 59.750 21.130 60.050 21.430 ;
        RECT 61.750 21.130 62.050 21.430 ;
        RECT 63.750 21.130 64.050 21.430 ;
        RECT 65.750 21.130 66.050 21.430 ;
        RECT 67.750 21.130 68.050 21.430 ;
        RECT 69.750 21.130 70.050 21.430 ;
        RECT 71.750 21.130 72.050 21.430 ;
        RECT 73.750 21.130 74.050 21.430 ;
        RECT 75.750 21.130 76.050 21.430 ;
        RECT 77.750 21.130 78.050 21.430 ;
        RECT 79.750 21.130 80.050 21.430 ;
        RECT 81.750 21.130 82.050 21.430 ;
        RECT 83.750 21.130 84.050 21.430 ;
        RECT 85.750 21.130 86.050 21.430 ;
        RECT 87.750 21.130 88.050 21.430 ;
        RECT 89.750 21.130 90.050 21.430 ;
        RECT 91.750 21.130 92.050 21.430 ;
        RECT 93.750 21.130 94.050 21.430 ;
        RECT 95.750 21.130 96.050 21.430 ;
        RECT 97.750 21.130 98.050 21.430 ;
        RECT 99.750 21.130 100.050 21.430 ;
        RECT 101.750 21.130 102.050 21.430 ;
        RECT 103.750 21.130 104.050 21.430 ;
        RECT 105.750 21.130 106.050 21.430 ;
        RECT 107.750 21.130 108.050 21.430 ;
        RECT 109.750 21.130 110.050 21.430 ;
        RECT 111.750 21.130 112.050 21.430 ;
        RECT 113.750 21.130 114.050 21.430 ;
        RECT 115.750 21.130 116.050 21.430 ;
        RECT 117.750 21.130 118.050 21.430 ;
        RECT 119.750 21.130 120.050 21.430 ;
        RECT 121.750 21.130 122.050 21.430 ;
        RECT 123.750 21.130 124.050 21.430 ;
        RECT 125.750 21.130 126.050 21.430 ;
        RECT 127.750 21.130 128.050 21.430 ;
        RECT 129.750 21.130 130.050 21.430 ;
        RECT 131.750 21.130 132.050 21.430 ;
        RECT 2.460 14.055 2.680 14.765 ;
        RECT 4.460 14.055 4.680 14.765 ;
        RECT 6.460 14.055 6.680 14.765 ;
        RECT 8.460 14.055 8.680 14.765 ;
        RECT 10.460 14.055 10.680 14.765 ;
        RECT 12.460 14.055 12.680 14.765 ;
        RECT 14.460 14.055 14.680 14.765 ;
        RECT 16.460 14.055 16.680 14.765 ;
        RECT 18.460 14.055 18.680 14.765 ;
        RECT 20.460 14.055 20.680 14.765 ;
        RECT 22.460 14.055 22.680 14.765 ;
        RECT 24.460 14.055 24.680 14.765 ;
        RECT 26.460 14.055 26.680 14.765 ;
        RECT 28.460 14.055 28.680 14.765 ;
        RECT 30.460 14.055 30.680 14.765 ;
        RECT 32.460 14.055 32.680 14.765 ;
        RECT 34.460 14.055 34.680 14.765 ;
        RECT 36.460 14.055 36.680 14.765 ;
        RECT 38.460 14.055 38.680 14.765 ;
        RECT 40.460 14.055 40.680 14.765 ;
        RECT 42.460 14.055 42.680 14.765 ;
        RECT 44.460 14.055 44.680 14.765 ;
        RECT 46.460 14.055 46.680 14.765 ;
        RECT 48.460 14.055 48.680 14.765 ;
        RECT 50.460 14.055 50.680 14.765 ;
        RECT 52.460 14.055 52.680 14.765 ;
        RECT 54.460 14.055 54.680 14.765 ;
        RECT 56.460 14.055 56.680 14.765 ;
        RECT 58.460 14.055 58.680 14.765 ;
        RECT 60.460 14.055 60.680 14.765 ;
        RECT 62.460 14.055 62.680 14.765 ;
        RECT 64.460 14.055 64.680 14.765 ;
        RECT 66.460 14.055 66.680 14.765 ;
        RECT 68.460 14.055 68.680 14.765 ;
        RECT 70.460 14.055 70.680 14.765 ;
        RECT 72.460 14.055 72.680 14.765 ;
        RECT 74.460 14.055 74.680 14.765 ;
        RECT 76.460 14.055 76.680 14.765 ;
        RECT 78.460 14.055 78.680 14.765 ;
        RECT 80.460 14.055 80.680 14.765 ;
        RECT 82.460 14.055 82.680 14.765 ;
        RECT 84.460 14.055 84.680 14.765 ;
        RECT 86.460 14.055 86.680 14.765 ;
        RECT 88.460 14.055 88.680 14.765 ;
        RECT 90.460 14.055 90.680 14.765 ;
        RECT 92.460 14.055 92.680 14.765 ;
        RECT 94.460 14.055 94.680 14.765 ;
        RECT 96.460 14.055 96.680 14.765 ;
        RECT 98.460 14.055 98.680 14.765 ;
        RECT 100.460 14.055 100.680 14.765 ;
        RECT 102.460 14.055 102.680 14.765 ;
        RECT 104.460 14.055 104.680 14.765 ;
        RECT 106.460 14.055 106.680 14.765 ;
        RECT 108.460 14.055 108.680 14.765 ;
        RECT 110.460 14.055 110.680 14.765 ;
        RECT 112.460 14.055 112.680 14.765 ;
        RECT 114.460 14.055 114.680 14.765 ;
        RECT 116.460 14.055 116.680 14.765 ;
        RECT 118.460 14.055 118.680 14.765 ;
        RECT 120.460 14.055 120.680 14.765 ;
        RECT 122.460 14.055 122.680 14.765 ;
        RECT 124.460 14.055 124.680 14.765 ;
        RECT 126.460 14.055 126.680 14.765 ;
        RECT 128.460 14.055 128.680 14.765 ;
        RECT 130.460 14.055 130.680 14.765 ;
        RECT 132.460 14.055 132.680 14.765 ;
        RECT 1.120 11.425 1.340 12.135 ;
        RECT 3.120 11.425 3.340 12.135 ;
        RECT 5.120 11.425 5.340 12.135 ;
        RECT 7.120 11.425 7.340 12.135 ;
        RECT 9.120 11.425 9.340 12.135 ;
        RECT 11.120 11.425 11.340 12.135 ;
        RECT 13.120 11.425 13.340 12.135 ;
        RECT 15.120 11.425 15.340 12.135 ;
        RECT 17.120 11.425 17.340 12.135 ;
        RECT 19.120 11.425 19.340 12.135 ;
        RECT 21.120 11.425 21.340 12.135 ;
        RECT 23.120 11.425 23.340 12.135 ;
        RECT 25.120 11.425 25.340 12.135 ;
        RECT 27.120 11.425 27.340 12.135 ;
        RECT 29.120 11.425 29.340 12.135 ;
        RECT 31.120 11.425 31.340 12.135 ;
        RECT 33.120 11.425 33.340 12.135 ;
        RECT 35.120 11.425 35.340 12.135 ;
        RECT 37.120 11.425 37.340 12.135 ;
        RECT 39.120 11.425 39.340 12.135 ;
        RECT 41.120 11.425 41.340 12.135 ;
        RECT 43.120 11.425 43.340 12.135 ;
        RECT 45.120 11.425 45.340 12.135 ;
        RECT 47.120 11.425 47.340 12.135 ;
        RECT 49.120 11.425 49.340 12.135 ;
        RECT 51.120 11.425 51.340 12.135 ;
        RECT 53.120 11.425 53.340 12.135 ;
        RECT 55.120 11.425 55.340 12.135 ;
        RECT 57.120 11.425 57.340 12.135 ;
        RECT 59.120 11.425 59.340 12.135 ;
        RECT 61.120 11.425 61.340 12.135 ;
        RECT 63.120 11.425 63.340 12.135 ;
        RECT 65.120 11.425 65.340 12.135 ;
        RECT 67.120 11.425 67.340 12.135 ;
        RECT 69.120 11.425 69.340 12.135 ;
        RECT 71.120 11.425 71.340 12.135 ;
        RECT 73.120 11.425 73.340 12.135 ;
        RECT 75.120 11.425 75.340 12.135 ;
        RECT 77.120 11.425 77.340 12.135 ;
        RECT 79.120 11.425 79.340 12.135 ;
        RECT 81.120 11.425 81.340 12.135 ;
        RECT 83.120 11.425 83.340 12.135 ;
        RECT 85.120 11.425 85.340 12.135 ;
        RECT 87.120 11.425 87.340 12.135 ;
        RECT 89.120 11.425 89.340 12.135 ;
        RECT 91.120 11.425 91.340 12.135 ;
        RECT 93.120 11.425 93.340 12.135 ;
        RECT 95.120 11.425 95.340 12.135 ;
        RECT 97.120 11.425 97.340 12.135 ;
        RECT 99.120 11.425 99.340 12.135 ;
        RECT 101.120 11.425 101.340 12.135 ;
        RECT 103.120 11.425 103.340 12.135 ;
        RECT 105.120 11.425 105.340 12.135 ;
        RECT 107.120 11.425 107.340 12.135 ;
        RECT 109.120 11.425 109.340 12.135 ;
        RECT 111.120 11.425 111.340 12.135 ;
        RECT 113.120 11.425 113.340 12.135 ;
        RECT 115.120 11.425 115.340 12.135 ;
        RECT 117.120 11.425 117.340 12.135 ;
        RECT 119.120 11.425 119.340 12.135 ;
        RECT 121.120 11.425 121.340 12.135 ;
        RECT 123.120 11.425 123.340 12.135 ;
        RECT 125.120 11.425 125.340 12.135 ;
        RECT 127.120 11.425 127.340 12.135 ;
        RECT 129.120 11.425 129.340 12.135 ;
        RECT 131.120 11.425 131.340 12.135 ;
        RECT 1.750 4.760 2.050 5.060 ;
        RECT 3.750 4.760 4.050 5.060 ;
        RECT 5.750 4.760 6.050 5.060 ;
        RECT 7.750 4.760 8.050 5.060 ;
        RECT 9.750 4.760 10.050 5.060 ;
        RECT 11.750 4.760 12.050 5.060 ;
        RECT 13.750 4.760 14.050 5.060 ;
        RECT 15.750 4.760 16.050 5.060 ;
        RECT 17.750 4.760 18.050 5.060 ;
        RECT 19.750 4.760 20.050 5.060 ;
        RECT 21.750 4.760 22.050 5.060 ;
        RECT 23.750 4.760 24.050 5.060 ;
        RECT 25.750 4.760 26.050 5.060 ;
        RECT 27.750 4.760 28.050 5.060 ;
        RECT 29.750 4.760 30.050 5.060 ;
        RECT 31.750 4.760 32.050 5.060 ;
        RECT 33.750 4.760 34.050 5.060 ;
        RECT 35.750 4.760 36.050 5.060 ;
        RECT 37.750 4.760 38.050 5.060 ;
        RECT 39.750 4.760 40.050 5.060 ;
        RECT 41.750 4.760 42.050 5.060 ;
        RECT 43.750 4.760 44.050 5.060 ;
        RECT 45.750 4.760 46.050 5.060 ;
        RECT 47.750 4.760 48.050 5.060 ;
        RECT 49.750 4.760 50.050 5.060 ;
        RECT 51.750 4.760 52.050 5.060 ;
        RECT 53.750 4.760 54.050 5.060 ;
        RECT 55.750 4.760 56.050 5.060 ;
        RECT 57.750 4.760 58.050 5.060 ;
        RECT 59.750 4.760 60.050 5.060 ;
        RECT 61.750 4.760 62.050 5.060 ;
        RECT 63.750 4.760 64.050 5.060 ;
        RECT 65.750 4.760 66.050 5.060 ;
        RECT 67.750 4.760 68.050 5.060 ;
        RECT 69.750 4.760 70.050 5.060 ;
        RECT 71.750 4.760 72.050 5.060 ;
        RECT 73.750 4.760 74.050 5.060 ;
        RECT 75.750 4.760 76.050 5.060 ;
        RECT 77.750 4.760 78.050 5.060 ;
        RECT 79.750 4.760 80.050 5.060 ;
        RECT 81.750 4.760 82.050 5.060 ;
        RECT 83.750 4.760 84.050 5.060 ;
        RECT 85.750 4.760 86.050 5.060 ;
        RECT 87.750 4.760 88.050 5.060 ;
        RECT 89.750 4.760 90.050 5.060 ;
        RECT 91.750 4.760 92.050 5.060 ;
        RECT 93.750 4.760 94.050 5.060 ;
        RECT 95.750 4.760 96.050 5.060 ;
        RECT 97.750 4.760 98.050 5.060 ;
        RECT 99.750 4.760 100.050 5.060 ;
        RECT 101.750 4.760 102.050 5.060 ;
        RECT 103.750 4.760 104.050 5.060 ;
        RECT 105.750 4.760 106.050 5.060 ;
        RECT 107.750 4.760 108.050 5.060 ;
        RECT 109.750 4.760 110.050 5.060 ;
        RECT 111.750 4.760 112.050 5.060 ;
        RECT 113.750 4.760 114.050 5.060 ;
        RECT 115.750 4.760 116.050 5.060 ;
        RECT 117.750 4.760 118.050 5.060 ;
        RECT 119.750 4.760 120.050 5.060 ;
        RECT 121.750 4.760 122.050 5.060 ;
        RECT 123.750 4.760 124.050 5.060 ;
        RECT 125.750 4.760 126.050 5.060 ;
        RECT 127.750 4.760 128.050 5.060 ;
        RECT 129.750 4.760 130.050 5.060 ;
        RECT 131.750 4.760 132.050 5.060 ;
        RECT 1.410 4.260 1.710 4.560 ;
        RECT 2.090 4.260 2.390 4.560 ;
        RECT 3.410 4.260 3.710 4.560 ;
        RECT 4.090 4.260 4.390 4.560 ;
        RECT 5.410 4.260 5.710 4.560 ;
        RECT 6.090 4.260 6.390 4.560 ;
        RECT 7.410 4.260 7.710 4.560 ;
        RECT 8.090 4.260 8.390 4.560 ;
        RECT 9.410 4.260 9.710 4.560 ;
        RECT 10.090 4.260 10.390 4.560 ;
        RECT 11.410 4.260 11.710 4.560 ;
        RECT 12.090 4.260 12.390 4.560 ;
        RECT 13.410 4.260 13.710 4.560 ;
        RECT 14.090 4.260 14.390 4.560 ;
        RECT 15.410 4.260 15.710 4.560 ;
        RECT 16.090 4.260 16.390 4.560 ;
        RECT 17.410 4.260 17.710 4.560 ;
        RECT 18.090 4.260 18.390 4.560 ;
        RECT 19.410 4.260 19.710 4.560 ;
        RECT 20.090 4.260 20.390 4.560 ;
        RECT 21.410 4.260 21.710 4.560 ;
        RECT 22.090 4.260 22.390 4.560 ;
        RECT 23.410 4.260 23.710 4.560 ;
        RECT 24.090 4.260 24.390 4.560 ;
        RECT 25.410 4.260 25.710 4.560 ;
        RECT 26.090 4.260 26.390 4.560 ;
        RECT 27.410 4.260 27.710 4.560 ;
        RECT 28.090 4.260 28.390 4.560 ;
        RECT 29.410 4.260 29.710 4.560 ;
        RECT 30.090 4.260 30.390 4.560 ;
        RECT 31.410 4.260 31.710 4.560 ;
        RECT 32.090 4.260 32.390 4.560 ;
        RECT 33.410 4.260 33.710 4.560 ;
        RECT 34.090 4.260 34.390 4.560 ;
        RECT 35.410 4.260 35.710 4.560 ;
        RECT 36.090 4.260 36.390 4.560 ;
        RECT 37.410 4.260 37.710 4.560 ;
        RECT 38.090 4.260 38.390 4.560 ;
        RECT 39.410 4.260 39.710 4.560 ;
        RECT 40.090 4.260 40.390 4.560 ;
        RECT 41.410 4.260 41.710 4.560 ;
        RECT 42.090 4.260 42.390 4.560 ;
        RECT 43.410 4.260 43.710 4.560 ;
        RECT 44.090 4.260 44.390 4.560 ;
        RECT 45.410 4.260 45.710 4.560 ;
        RECT 46.090 4.260 46.390 4.560 ;
        RECT 47.410 4.260 47.710 4.560 ;
        RECT 48.090 4.260 48.390 4.560 ;
        RECT 49.410 4.260 49.710 4.560 ;
        RECT 50.090 4.260 50.390 4.560 ;
        RECT 51.410 4.260 51.710 4.560 ;
        RECT 52.090 4.260 52.390 4.560 ;
        RECT 53.410 4.260 53.710 4.560 ;
        RECT 54.090 4.260 54.390 4.560 ;
        RECT 55.410 4.260 55.710 4.560 ;
        RECT 56.090 4.260 56.390 4.560 ;
        RECT 57.410 4.260 57.710 4.560 ;
        RECT 58.090 4.260 58.390 4.560 ;
        RECT 59.410 4.260 59.710 4.560 ;
        RECT 60.090 4.260 60.390 4.560 ;
        RECT 61.410 4.260 61.710 4.560 ;
        RECT 62.090 4.260 62.390 4.560 ;
        RECT 63.410 4.260 63.710 4.560 ;
        RECT 64.090 4.260 64.390 4.560 ;
        RECT 65.410 4.260 65.710 4.560 ;
        RECT 66.090 4.260 66.390 4.560 ;
        RECT 67.410 4.260 67.710 4.560 ;
        RECT 68.090 4.260 68.390 4.560 ;
        RECT 69.410 4.260 69.710 4.560 ;
        RECT 70.090 4.260 70.390 4.560 ;
        RECT 71.410 4.260 71.710 4.560 ;
        RECT 72.090 4.260 72.390 4.560 ;
        RECT 73.410 4.260 73.710 4.560 ;
        RECT 74.090 4.260 74.390 4.560 ;
        RECT 75.410 4.260 75.710 4.560 ;
        RECT 76.090 4.260 76.390 4.560 ;
        RECT 77.410 4.260 77.710 4.560 ;
        RECT 78.090 4.260 78.390 4.560 ;
        RECT 79.410 4.260 79.710 4.560 ;
        RECT 80.090 4.260 80.390 4.560 ;
        RECT 81.410 4.260 81.710 4.560 ;
        RECT 82.090 4.260 82.390 4.560 ;
        RECT 83.410 4.260 83.710 4.560 ;
        RECT 84.090 4.260 84.390 4.560 ;
        RECT 85.410 4.260 85.710 4.560 ;
        RECT 86.090 4.260 86.390 4.560 ;
        RECT 87.410 4.260 87.710 4.560 ;
        RECT 88.090 4.260 88.390 4.560 ;
        RECT 89.410 4.260 89.710 4.560 ;
        RECT 90.090 4.260 90.390 4.560 ;
        RECT 91.410 4.260 91.710 4.560 ;
        RECT 92.090 4.260 92.390 4.560 ;
        RECT 93.410 4.260 93.710 4.560 ;
        RECT 94.090 4.260 94.390 4.560 ;
        RECT 95.410 4.260 95.710 4.560 ;
        RECT 96.090 4.260 96.390 4.560 ;
        RECT 97.410 4.260 97.710 4.560 ;
        RECT 98.090 4.260 98.390 4.560 ;
        RECT 99.410 4.260 99.710 4.560 ;
        RECT 100.090 4.260 100.390 4.560 ;
        RECT 101.410 4.260 101.710 4.560 ;
        RECT 102.090 4.260 102.390 4.560 ;
        RECT 103.410 4.260 103.710 4.560 ;
        RECT 104.090 4.260 104.390 4.560 ;
        RECT 105.410 4.260 105.710 4.560 ;
        RECT 106.090 4.260 106.390 4.560 ;
        RECT 107.410 4.260 107.710 4.560 ;
        RECT 108.090 4.260 108.390 4.560 ;
        RECT 109.410 4.260 109.710 4.560 ;
        RECT 110.090 4.260 110.390 4.560 ;
        RECT 111.410 4.260 111.710 4.560 ;
        RECT 112.090 4.260 112.390 4.560 ;
        RECT 113.410 4.260 113.710 4.560 ;
        RECT 114.090 4.260 114.390 4.560 ;
        RECT 115.410 4.260 115.710 4.560 ;
        RECT 116.090 4.260 116.390 4.560 ;
        RECT 117.410 4.260 117.710 4.560 ;
        RECT 118.090 4.260 118.390 4.560 ;
        RECT 119.410 4.260 119.710 4.560 ;
        RECT 120.090 4.260 120.390 4.560 ;
        RECT 121.410 4.260 121.710 4.560 ;
        RECT 122.090 4.260 122.390 4.560 ;
        RECT 123.410 4.260 123.710 4.560 ;
        RECT 124.090 4.260 124.390 4.560 ;
        RECT 125.410 4.260 125.710 4.560 ;
        RECT 126.090 4.260 126.390 4.560 ;
        RECT 127.410 4.260 127.710 4.560 ;
        RECT 128.090 4.260 128.390 4.560 ;
        RECT 129.410 4.260 129.710 4.560 ;
        RECT 130.090 4.260 130.390 4.560 ;
        RECT 131.410 4.260 131.710 4.560 ;
        RECT 132.090 4.260 132.390 4.560 ;
        RECT 1.010 2.910 1.300 3.200 ;
        RECT 2.500 2.910 2.790 3.200 ;
        RECT 3.010 2.910 3.300 3.200 ;
        RECT 4.500 2.910 4.790 3.200 ;
        RECT 5.010 2.910 5.300 3.200 ;
        RECT 6.500 2.910 6.790 3.200 ;
        RECT 7.010 2.910 7.300 3.200 ;
        RECT 8.500 2.910 8.790 3.200 ;
        RECT 9.010 2.910 9.300 3.200 ;
        RECT 10.500 2.910 10.790 3.200 ;
        RECT 11.010 2.910 11.300 3.200 ;
        RECT 12.500 2.910 12.790 3.200 ;
        RECT 13.010 2.910 13.300 3.200 ;
        RECT 14.500 2.910 14.790 3.200 ;
        RECT 15.010 2.910 15.300 3.200 ;
        RECT 16.500 2.910 16.790 3.200 ;
        RECT 17.010 2.910 17.300 3.200 ;
        RECT 18.500 2.910 18.790 3.200 ;
        RECT 19.010 2.910 19.300 3.200 ;
        RECT 20.500 2.910 20.790 3.200 ;
        RECT 21.010 2.910 21.300 3.200 ;
        RECT 22.500 2.910 22.790 3.200 ;
        RECT 23.010 2.910 23.300 3.200 ;
        RECT 24.500 2.910 24.790 3.200 ;
        RECT 25.010 2.910 25.300 3.200 ;
        RECT 26.500 2.910 26.790 3.200 ;
        RECT 27.010 2.910 27.300 3.200 ;
        RECT 28.500 2.910 28.790 3.200 ;
        RECT 29.010 2.910 29.300 3.200 ;
        RECT 30.500 2.910 30.790 3.200 ;
        RECT 31.010 2.910 31.300 3.200 ;
        RECT 32.500 2.910 32.790 3.200 ;
        RECT 33.010 2.910 33.300 3.200 ;
        RECT 34.500 2.910 34.790 3.200 ;
        RECT 35.010 2.910 35.300 3.200 ;
        RECT 36.500 2.910 36.790 3.200 ;
        RECT 37.010 2.910 37.300 3.200 ;
        RECT 38.500 2.910 38.790 3.200 ;
        RECT 39.010 2.910 39.300 3.200 ;
        RECT 40.500 2.910 40.790 3.200 ;
        RECT 41.010 2.910 41.300 3.200 ;
        RECT 42.500 2.910 42.790 3.200 ;
        RECT 43.010 2.910 43.300 3.200 ;
        RECT 44.500 2.910 44.790 3.200 ;
        RECT 45.010 2.910 45.300 3.200 ;
        RECT 46.500 2.910 46.790 3.200 ;
        RECT 47.010 2.910 47.300 3.200 ;
        RECT 48.500 2.910 48.790 3.200 ;
        RECT 49.010 2.910 49.300 3.200 ;
        RECT 50.500 2.910 50.790 3.200 ;
        RECT 51.010 2.910 51.300 3.200 ;
        RECT 52.500 2.910 52.790 3.200 ;
        RECT 53.010 2.910 53.300 3.200 ;
        RECT 54.500 2.910 54.790 3.200 ;
        RECT 55.010 2.910 55.300 3.200 ;
        RECT 56.500 2.910 56.790 3.200 ;
        RECT 57.010 2.910 57.300 3.200 ;
        RECT 58.500 2.910 58.790 3.200 ;
        RECT 59.010 2.910 59.300 3.200 ;
        RECT 60.500 2.910 60.790 3.200 ;
        RECT 61.010 2.910 61.300 3.200 ;
        RECT 62.500 2.910 62.790 3.200 ;
        RECT 63.010 2.910 63.300 3.200 ;
        RECT 64.500 2.910 64.790 3.200 ;
        RECT 65.010 2.910 65.300 3.200 ;
        RECT 66.500 2.910 66.790 3.200 ;
        RECT 67.010 2.910 67.300 3.200 ;
        RECT 68.500 2.910 68.790 3.200 ;
        RECT 69.010 2.910 69.300 3.200 ;
        RECT 70.500 2.910 70.790 3.200 ;
        RECT 71.010 2.910 71.300 3.200 ;
        RECT 72.500 2.910 72.790 3.200 ;
        RECT 73.010 2.910 73.300 3.200 ;
        RECT 74.500 2.910 74.790 3.200 ;
        RECT 75.010 2.910 75.300 3.200 ;
        RECT 76.500 2.910 76.790 3.200 ;
        RECT 77.010 2.910 77.300 3.200 ;
        RECT 78.500 2.910 78.790 3.200 ;
        RECT 79.010 2.910 79.300 3.200 ;
        RECT 80.500 2.910 80.790 3.200 ;
        RECT 81.010 2.910 81.300 3.200 ;
        RECT 82.500 2.910 82.790 3.200 ;
        RECT 83.010 2.910 83.300 3.200 ;
        RECT 84.500 2.910 84.790 3.200 ;
        RECT 85.010 2.910 85.300 3.200 ;
        RECT 86.500 2.910 86.790 3.200 ;
        RECT 87.010 2.910 87.300 3.200 ;
        RECT 88.500 2.910 88.790 3.200 ;
        RECT 89.010 2.910 89.300 3.200 ;
        RECT 90.500 2.910 90.790 3.200 ;
        RECT 91.010 2.910 91.300 3.200 ;
        RECT 92.500 2.910 92.790 3.200 ;
        RECT 93.010 2.910 93.300 3.200 ;
        RECT 94.500 2.910 94.790 3.200 ;
        RECT 95.010 2.910 95.300 3.200 ;
        RECT 96.500 2.910 96.790 3.200 ;
        RECT 97.010 2.910 97.300 3.200 ;
        RECT 98.500 2.910 98.790 3.200 ;
        RECT 99.010 2.910 99.300 3.200 ;
        RECT 100.500 2.910 100.790 3.200 ;
        RECT 101.010 2.910 101.300 3.200 ;
        RECT 102.500 2.910 102.790 3.200 ;
        RECT 103.010 2.910 103.300 3.200 ;
        RECT 104.500 2.910 104.790 3.200 ;
        RECT 105.010 2.910 105.300 3.200 ;
        RECT 106.500 2.910 106.790 3.200 ;
        RECT 107.010 2.910 107.300 3.200 ;
        RECT 108.500 2.910 108.790 3.200 ;
        RECT 109.010 2.910 109.300 3.200 ;
        RECT 110.500 2.910 110.790 3.200 ;
        RECT 111.010 2.910 111.300 3.200 ;
        RECT 112.500 2.910 112.790 3.200 ;
        RECT 113.010 2.910 113.300 3.200 ;
        RECT 114.500 2.910 114.790 3.200 ;
        RECT 115.010 2.910 115.300 3.200 ;
        RECT 116.500 2.910 116.790 3.200 ;
        RECT 117.010 2.910 117.300 3.200 ;
        RECT 118.500 2.910 118.790 3.200 ;
        RECT 119.010 2.910 119.300 3.200 ;
        RECT 120.500 2.910 120.790 3.200 ;
        RECT 121.010 2.910 121.300 3.200 ;
        RECT 122.500 2.910 122.790 3.200 ;
        RECT 123.010 2.910 123.300 3.200 ;
        RECT 124.500 2.910 124.790 3.200 ;
        RECT 125.010 2.910 125.300 3.200 ;
        RECT 126.500 2.910 126.790 3.200 ;
        RECT 127.010 2.910 127.300 3.200 ;
        RECT 128.500 2.910 128.790 3.200 ;
        RECT 129.010 2.910 129.300 3.200 ;
        RECT 130.500 2.910 130.790 3.200 ;
        RECT 131.010 2.910 131.300 3.200 ;
        RECT 132.500 2.910 132.790 3.200 ;
        RECT 1.075 1.780 1.235 2.910 ;
        RECT 1.075 1.620 2.325 1.780 ;
        RECT 1.075 0.800 1.235 1.620 ;
        RECT 2.565 0.800 2.725 2.910 ;
        RECT 3.075 1.780 3.235 2.910 ;
        RECT 3.075 1.620 4.325 1.780 ;
        RECT 3.075 0.800 3.235 1.620 ;
        RECT 4.565 0.800 4.725 2.910 ;
        RECT 5.075 1.780 5.235 2.910 ;
        RECT 5.075 1.620 6.325 1.780 ;
        RECT 5.075 0.800 5.235 1.620 ;
        RECT 6.565 0.800 6.725 2.910 ;
        RECT 7.075 1.780 7.235 2.910 ;
        RECT 7.075 1.620 8.325 1.780 ;
        RECT 7.075 0.800 7.235 1.620 ;
        RECT 8.565 0.800 8.725 2.910 ;
        RECT 9.075 1.780 9.235 2.910 ;
        RECT 9.075 1.620 10.325 1.780 ;
        RECT 9.075 0.800 9.235 1.620 ;
        RECT 10.565 0.800 10.725 2.910 ;
        RECT 11.075 1.780 11.235 2.910 ;
        RECT 11.075 1.620 12.325 1.780 ;
        RECT 11.075 0.800 11.235 1.620 ;
        RECT 12.565 0.800 12.725 2.910 ;
        RECT 13.075 1.780 13.235 2.910 ;
        RECT 13.075 1.620 14.325 1.780 ;
        RECT 13.075 0.800 13.235 1.620 ;
        RECT 14.565 0.800 14.725 2.910 ;
        RECT 15.075 1.780 15.235 2.910 ;
        RECT 15.075 1.620 16.325 1.780 ;
        RECT 15.075 0.800 15.235 1.620 ;
        RECT 16.565 0.800 16.725 2.910 ;
        RECT 17.075 1.780 17.235 2.910 ;
        RECT 17.075 1.620 18.325 1.780 ;
        RECT 17.075 0.800 17.235 1.620 ;
        RECT 18.565 0.800 18.725 2.910 ;
        RECT 19.075 1.780 19.235 2.910 ;
        RECT 19.075 1.620 20.325 1.780 ;
        RECT 19.075 0.800 19.235 1.620 ;
        RECT 20.565 0.800 20.725 2.910 ;
        RECT 21.075 1.780 21.235 2.910 ;
        RECT 21.075 1.620 22.325 1.780 ;
        RECT 21.075 0.800 21.235 1.620 ;
        RECT 22.565 0.800 22.725 2.910 ;
        RECT 23.075 1.780 23.235 2.910 ;
        RECT 23.075 1.620 24.325 1.780 ;
        RECT 23.075 0.800 23.235 1.620 ;
        RECT 24.565 0.800 24.725 2.910 ;
        RECT 25.075 1.780 25.235 2.910 ;
        RECT 25.075 1.620 26.325 1.780 ;
        RECT 25.075 0.800 25.235 1.620 ;
        RECT 26.565 0.800 26.725 2.910 ;
        RECT 27.075 1.780 27.235 2.910 ;
        RECT 27.075 1.620 28.325 1.780 ;
        RECT 27.075 0.800 27.235 1.620 ;
        RECT 28.565 0.800 28.725 2.910 ;
        RECT 29.075 1.780 29.235 2.910 ;
        RECT 29.075 1.620 30.325 1.780 ;
        RECT 29.075 0.800 29.235 1.620 ;
        RECT 30.565 0.800 30.725 2.910 ;
        RECT 31.075 1.780 31.235 2.910 ;
        RECT 31.075 1.620 32.325 1.780 ;
        RECT 31.075 0.800 31.235 1.620 ;
        RECT 32.565 0.800 32.725 2.910 ;
        RECT 33.075 1.780 33.235 2.910 ;
        RECT 33.075 1.620 34.325 1.780 ;
        RECT 33.075 0.800 33.235 1.620 ;
        RECT 34.565 0.800 34.725 2.910 ;
        RECT 35.075 1.780 35.235 2.910 ;
        RECT 35.075 1.620 36.325 1.780 ;
        RECT 35.075 0.800 35.235 1.620 ;
        RECT 36.565 0.800 36.725 2.910 ;
        RECT 37.075 1.780 37.235 2.910 ;
        RECT 37.075 1.620 38.325 1.780 ;
        RECT 37.075 0.800 37.235 1.620 ;
        RECT 38.565 0.800 38.725 2.910 ;
        RECT 39.075 1.780 39.235 2.910 ;
        RECT 39.075 1.620 40.325 1.780 ;
        RECT 39.075 0.800 39.235 1.620 ;
        RECT 40.565 0.800 40.725 2.910 ;
        RECT 41.075 1.780 41.235 2.910 ;
        RECT 41.075 1.620 42.325 1.780 ;
        RECT 41.075 0.800 41.235 1.620 ;
        RECT 42.565 0.800 42.725 2.910 ;
        RECT 43.075 1.780 43.235 2.910 ;
        RECT 43.075 1.620 44.325 1.780 ;
        RECT 43.075 0.800 43.235 1.620 ;
        RECT 44.565 0.800 44.725 2.910 ;
        RECT 45.075 1.780 45.235 2.910 ;
        RECT 45.075 1.620 46.325 1.780 ;
        RECT 45.075 0.800 45.235 1.620 ;
        RECT 46.565 0.800 46.725 2.910 ;
        RECT 47.075 1.780 47.235 2.910 ;
        RECT 47.075 1.620 48.325 1.780 ;
        RECT 47.075 0.800 47.235 1.620 ;
        RECT 48.565 0.800 48.725 2.910 ;
        RECT 49.075 1.780 49.235 2.910 ;
        RECT 49.075 1.620 50.325 1.780 ;
        RECT 49.075 0.800 49.235 1.620 ;
        RECT 50.565 0.800 50.725 2.910 ;
        RECT 51.075 1.780 51.235 2.910 ;
        RECT 51.075 1.620 52.325 1.780 ;
        RECT 51.075 0.800 51.235 1.620 ;
        RECT 52.565 0.800 52.725 2.910 ;
        RECT 53.075 1.780 53.235 2.910 ;
        RECT 53.075 1.620 54.325 1.780 ;
        RECT 53.075 0.800 53.235 1.620 ;
        RECT 54.565 0.800 54.725 2.910 ;
        RECT 55.075 1.780 55.235 2.910 ;
        RECT 55.075 1.620 56.325 1.780 ;
        RECT 55.075 0.800 55.235 1.620 ;
        RECT 56.565 0.800 56.725 2.910 ;
        RECT 57.075 1.780 57.235 2.910 ;
        RECT 57.075 1.620 58.325 1.780 ;
        RECT 57.075 0.800 57.235 1.620 ;
        RECT 58.565 0.800 58.725 2.910 ;
        RECT 59.075 1.780 59.235 2.910 ;
        RECT 59.075 1.620 60.325 1.780 ;
        RECT 59.075 0.800 59.235 1.620 ;
        RECT 60.565 0.800 60.725 2.910 ;
        RECT 61.075 1.780 61.235 2.910 ;
        RECT 61.075 1.620 62.325 1.780 ;
        RECT 61.075 0.800 61.235 1.620 ;
        RECT 62.565 0.800 62.725 2.910 ;
        RECT 63.075 1.780 63.235 2.910 ;
        RECT 63.075 1.620 64.325 1.780 ;
        RECT 63.075 0.800 63.235 1.620 ;
        RECT 64.565 0.800 64.725 2.910 ;
        RECT 65.075 1.780 65.235 2.910 ;
        RECT 65.075 1.620 66.325 1.780 ;
        RECT 65.075 0.800 65.235 1.620 ;
        RECT 66.565 0.800 66.725 2.910 ;
        RECT 67.075 1.780 67.235 2.910 ;
        RECT 67.075 1.620 68.325 1.780 ;
        RECT 67.075 0.800 67.235 1.620 ;
        RECT 68.565 0.800 68.725 2.910 ;
        RECT 69.075 1.780 69.235 2.910 ;
        RECT 69.075 1.620 70.325 1.780 ;
        RECT 69.075 0.800 69.235 1.620 ;
        RECT 70.565 0.800 70.725 2.910 ;
        RECT 71.075 1.780 71.235 2.910 ;
        RECT 71.075 1.620 72.325 1.780 ;
        RECT 71.075 0.800 71.235 1.620 ;
        RECT 72.565 0.800 72.725 2.910 ;
        RECT 73.075 1.780 73.235 2.910 ;
        RECT 73.075 1.620 74.325 1.780 ;
        RECT 73.075 0.800 73.235 1.620 ;
        RECT 74.565 0.800 74.725 2.910 ;
        RECT 75.075 1.780 75.235 2.910 ;
        RECT 75.075 1.620 76.325 1.780 ;
        RECT 75.075 0.800 75.235 1.620 ;
        RECT 76.565 0.800 76.725 2.910 ;
        RECT 77.075 1.780 77.235 2.910 ;
        RECT 77.075 1.620 78.325 1.780 ;
        RECT 77.075 0.800 77.235 1.620 ;
        RECT 78.565 0.800 78.725 2.910 ;
        RECT 79.075 1.780 79.235 2.910 ;
        RECT 79.075 1.620 80.325 1.780 ;
        RECT 79.075 0.800 79.235 1.620 ;
        RECT 80.565 0.800 80.725 2.910 ;
        RECT 81.075 1.780 81.235 2.910 ;
        RECT 81.075 1.620 82.325 1.780 ;
        RECT 81.075 0.800 81.235 1.620 ;
        RECT 82.565 0.800 82.725 2.910 ;
        RECT 83.075 1.780 83.235 2.910 ;
        RECT 83.075 1.620 84.325 1.780 ;
        RECT 83.075 0.800 83.235 1.620 ;
        RECT 84.565 0.800 84.725 2.910 ;
        RECT 85.075 1.780 85.235 2.910 ;
        RECT 85.075 1.620 86.325 1.780 ;
        RECT 85.075 0.800 85.235 1.620 ;
        RECT 86.565 0.800 86.725 2.910 ;
        RECT 87.075 1.780 87.235 2.910 ;
        RECT 87.075 1.620 88.325 1.780 ;
        RECT 87.075 0.800 87.235 1.620 ;
        RECT 88.565 0.800 88.725 2.910 ;
        RECT 89.075 1.780 89.235 2.910 ;
        RECT 89.075 1.620 90.325 1.780 ;
        RECT 89.075 0.800 89.235 1.620 ;
        RECT 90.565 0.800 90.725 2.910 ;
        RECT 91.075 1.780 91.235 2.910 ;
        RECT 91.075 1.620 92.325 1.780 ;
        RECT 91.075 0.800 91.235 1.620 ;
        RECT 92.565 0.800 92.725 2.910 ;
        RECT 93.075 1.780 93.235 2.910 ;
        RECT 93.075 1.620 94.325 1.780 ;
        RECT 93.075 0.800 93.235 1.620 ;
        RECT 94.565 0.800 94.725 2.910 ;
        RECT 95.075 1.780 95.235 2.910 ;
        RECT 95.075 1.620 96.325 1.780 ;
        RECT 95.075 0.800 95.235 1.620 ;
        RECT 96.565 0.800 96.725 2.910 ;
        RECT 97.075 1.780 97.235 2.910 ;
        RECT 97.075 1.620 98.325 1.780 ;
        RECT 97.075 0.800 97.235 1.620 ;
        RECT 98.565 0.800 98.725 2.910 ;
        RECT 99.075 1.780 99.235 2.910 ;
        RECT 99.075 1.620 100.325 1.780 ;
        RECT 99.075 0.800 99.235 1.620 ;
        RECT 100.565 0.800 100.725 2.910 ;
        RECT 101.075 1.780 101.235 2.910 ;
        RECT 101.075 1.620 102.325 1.780 ;
        RECT 101.075 0.800 101.235 1.620 ;
        RECT 102.565 0.800 102.725 2.910 ;
        RECT 103.075 1.780 103.235 2.910 ;
        RECT 103.075 1.620 104.325 1.780 ;
        RECT 103.075 0.800 103.235 1.620 ;
        RECT 104.565 0.800 104.725 2.910 ;
        RECT 105.075 1.780 105.235 2.910 ;
        RECT 105.075 1.620 106.325 1.780 ;
        RECT 105.075 0.800 105.235 1.620 ;
        RECT 106.565 0.800 106.725 2.910 ;
        RECT 107.075 1.780 107.235 2.910 ;
        RECT 107.075 1.620 108.325 1.780 ;
        RECT 107.075 0.800 107.235 1.620 ;
        RECT 108.565 0.800 108.725 2.910 ;
        RECT 109.075 1.780 109.235 2.910 ;
        RECT 109.075 1.620 110.325 1.780 ;
        RECT 109.075 0.800 109.235 1.620 ;
        RECT 110.565 0.800 110.725 2.910 ;
        RECT 111.075 1.780 111.235 2.910 ;
        RECT 111.075 1.620 112.325 1.780 ;
        RECT 111.075 0.800 111.235 1.620 ;
        RECT 112.565 0.800 112.725 2.910 ;
        RECT 113.075 1.780 113.235 2.910 ;
        RECT 113.075 1.620 114.325 1.780 ;
        RECT 113.075 0.800 113.235 1.620 ;
        RECT 114.565 0.800 114.725 2.910 ;
        RECT 115.075 1.780 115.235 2.910 ;
        RECT 115.075 1.620 116.325 1.780 ;
        RECT 115.075 0.800 115.235 1.620 ;
        RECT 116.565 0.800 116.725 2.910 ;
        RECT 117.075 1.780 117.235 2.910 ;
        RECT 117.075 1.620 118.325 1.780 ;
        RECT 117.075 0.800 117.235 1.620 ;
        RECT 118.565 0.800 118.725 2.910 ;
        RECT 119.075 1.780 119.235 2.910 ;
        RECT 119.075 1.620 120.325 1.780 ;
        RECT 119.075 0.800 119.235 1.620 ;
        RECT 120.565 0.800 120.725 2.910 ;
        RECT 121.075 1.780 121.235 2.910 ;
        RECT 121.075 1.620 122.325 1.780 ;
        RECT 121.075 0.800 121.235 1.620 ;
        RECT 122.565 0.800 122.725 2.910 ;
        RECT 123.075 1.780 123.235 2.910 ;
        RECT 123.075 1.620 124.325 1.780 ;
        RECT 123.075 0.800 123.235 1.620 ;
        RECT 124.565 0.800 124.725 2.910 ;
        RECT 125.075 1.780 125.235 2.910 ;
        RECT 125.075 1.620 126.325 1.780 ;
        RECT 125.075 0.800 125.235 1.620 ;
        RECT 126.565 0.800 126.725 2.910 ;
        RECT 127.075 1.780 127.235 2.910 ;
        RECT 127.075 1.620 128.325 1.780 ;
        RECT 127.075 0.800 127.235 1.620 ;
        RECT 128.565 0.800 128.725 2.910 ;
        RECT 129.075 1.780 129.235 2.910 ;
        RECT 129.075 1.620 130.325 1.780 ;
        RECT 129.075 0.800 129.235 1.620 ;
        RECT 130.565 0.800 130.725 2.910 ;
        RECT 131.075 1.780 131.235 2.910 ;
        RECT 131.075 1.620 132.325 1.780 ;
        RECT 131.075 0.800 131.235 1.620 ;
        RECT 132.565 0.800 132.725 2.910 ;
      LAYER Metal2 ;
        RECT 1.010 22.990 1.300 23.280 ;
        RECT 2.500 22.990 2.790 23.280 ;
        RECT 3.010 22.990 3.300 23.280 ;
        RECT 4.500 22.990 4.790 23.280 ;
        RECT 5.010 22.990 5.300 23.280 ;
        RECT 6.500 22.990 6.790 23.280 ;
        RECT 7.010 22.990 7.300 23.280 ;
        RECT 8.500 22.990 8.790 23.280 ;
        RECT 9.010 22.990 9.300 23.280 ;
        RECT 10.500 22.990 10.790 23.280 ;
        RECT 11.010 22.990 11.300 23.280 ;
        RECT 12.500 22.990 12.790 23.280 ;
        RECT 13.010 22.990 13.300 23.280 ;
        RECT 14.500 22.990 14.790 23.280 ;
        RECT 15.010 22.990 15.300 23.280 ;
        RECT 16.500 22.990 16.790 23.280 ;
        RECT 17.010 22.990 17.300 23.280 ;
        RECT 18.500 22.990 18.790 23.280 ;
        RECT 19.010 22.990 19.300 23.280 ;
        RECT 20.500 22.990 20.790 23.280 ;
        RECT 21.010 22.990 21.300 23.280 ;
        RECT 22.500 22.990 22.790 23.280 ;
        RECT 23.010 22.990 23.300 23.280 ;
        RECT 24.500 22.990 24.790 23.280 ;
        RECT 25.010 22.990 25.300 23.280 ;
        RECT 26.500 22.990 26.790 23.280 ;
        RECT 27.010 22.990 27.300 23.280 ;
        RECT 28.500 22.990 28.790 23.280 ;
        RECT 29.010 22.990 29.300 23.280 ;
        RECT 30.500 22.990 30.790 23.280 ;
        RECT 31.010 22.990 31.300 23.280 ;
        RECT 32.500 22.990 32.790 23.280 ;
        RECT 33.010 22.990 33.300 23.280 ;
        RECT 34.500 22.990 34.790 23.280 ;
        RECT 35.010 22.990 35.300 23.280 ;
        RECT 36.500 22.990 36.790 23.280 ;
        RECT 37.010 22.990 37.300 23.280 ;
        RECT 38.500 22.990 38.790 23.280 ;
        RECT 39.010 22.990 39.300 23.280 ;
        RECT 40.500 22.990 40.790 23.280 ;
        RECT 41.010 22.990 41.300 23.280 ;
        RECT 42.500 22.990 42.790 23.280 ;
        RECT 43.010 22.990 43.300 23.280 ;
        RECT 44.500 22.990 44.790 23.280 ;
        RECT 45.010 22.990 45.300 23.280 ;
        RECT 46.500 22.990 46.790 23.280 ;
        RECT 47.010 22.990 47.300 23.280 ;
        RECT 48.500 22.990 48.790 23.280 ;
        RECT 49.010 22.990 49.300 23.280 ;
        RECT 50.500 22.990 50.790 23.280 ;
        RECT 51.010 22.990 51.300 23.280 ;
        RECT 52.500 22.990 52.790 23.280 ;
        RECT 53.010 22.990 53.300 23.280 ;
        RECT 54.500 22.990 54.790 23.280 ;
        RECT 55.010 22.990 55.300 23.280 ;
        RECT 56.500 22.990 56.790 23.280 ;
        RECT 57.010 22.990 57.300 23.280 ;
        RECT 58.500 22.990 58.790 23.280 ;
        RECT 59.010 22.990 59.300 23.280 ;
        RECT 60.500 22.990 60.790 23.280 ;
        RECT 61.010 22.990 61.300 23.280 ;
        RECT 62.500 22.990 62.790 23.280 ;
        RECT 63.010 22.990 63.300 23.280 ;
        RECT 64.500 22.990 64.790 23.280 ;
        RECT 65.010 22.990 65.300 23.280 ;
        RECT 66.500 22.990 66.790 23.280 ;
        RECT 67.010 22.990 67.300 23.280 ;
        RECT 68.500 22.990 68.790 23.280 ;
        RECT 69.010 22.990 69.300 23.280 ;
        RECT 70.500 22.990 70.790 23.280 ;
        RECT 71.010 22.990 71.300 23.280 ;
        RECT 72.500 22.990 72.790 23.280 ;
        RECT 73.010 22.990 73.300 23.280 ;
        RECT 74.500 22.990 74.790 23.280 ;
        RECT 75.010 22.990 75.300 23.280 ;
        RECT 76.500 22.990 76.790 23.280 ;
        RECT 77.010 22.990 77.300 23.280 ;
        RECT 78.500 22.990 78.790 23.280 ;
        RECT 79.010 22.990 79.300 23.280 ;
        RECT 80.500 22.990 80.790 23.280 ;
        RECT 81.010 22.990 81.300 23.280 ;
        RECT 82.500 22.990 82.790 23.280 ;
        RECT 83.010 22.990 83.300 23.280 ;
        RECT 84.500 22.990 84.790 23.280 ;
        RECT 85.010 22.990 85.300 23.280 ;
        RECT 86.500 22.990 86.790 23.280 ;
        RECT 87.010 22.990 87.300 23.280 ;
        RECT 88.500 22.990 88.790 23.280 ;
        RECT 89.010 22.990 89.300 23.280 ;
        RECT 90.500 22.990 90.790 23.280 ;
        RECT 91.010 22.990 91.300 23.280 ;
        RECT 92.500 22.990 92.790 23.280 ;
        RECT 93.010 22.990 93.300 23.280 ;
        RECT 94.500 22.990 94.790 23.280 ;
        RECT 95.010 22.990 95.300 23.280 ;
        RECT 96.500 22.990 96.790 23.280 ;
        RECT 97.010 22.990 97.300 23.280 ;
        RECT 98.500 22.990 98.790 23.280 ;
        RECT 99.010 22.990 99.300 23.280 ;
        RECT 100.500 22.990 100.790 23.280 ;
        RECT 101.010 22.990 101.300 23.280 ;
        RECT 102.500 22.990 102.790 23.280 ;
        RECT 103.010 22.990 103.300 23.280 ;
        RECT 104.500 22.990 104.790 23.280 ;
        RECT 105.010 22.990 105.300 23.280 ;
        RECT 106.500 22.990 106.790 23.280 ;
        RECT 107.010 22.990 107.300 23.280 ;
        RECT 108.500 22.990 108.790 23.280 ;
        RECT 109.010 22.990 109.300 23.280 ;
        RECT 110.500 22.990 110.790 23.280 ;
        RECT 111.010 22.990 111.300 23.280 ;
        RECT 112.500 22.990 112.790 23.280 ;
        RECT 113.010 22.990 113.300 23.280 ;
        RECT 114.500 22.990 114.790 23.280 ;
        RECT 115.010 22.990 115.300 23.280 ;
        RECT 116.500 22.990 116.790 23.280 ;
        RECT 117.010 22.990 117.300 23.280 ;
        RECT 118.500 22.990 118.790 23.280 ;
        RECT 119.010 22.990 119.300 23.280 ;
        RECT 120.500 22.990 120.790 23.280 ;
        RECT 121.010 22.990 121.300 23.280 ;
        RECT 122.500 22.990 122.790 23.280 ;
        RECT 123.010 22.990 123.300 23.280 ;
        RECT 124.500 22.990 124.790 23.280 ;
        RECT 125.010 22.990 125.300 23.280 ;
        RECT 126.500 22.990 126.790 23.280 ;
        RECT 127.010 22.990 127.300 23.280 ;
        RECT 128.500 22.990 128.790 23.280 ;
        RECT 129.010 22.990 129.300 23.280 ;
        RECT 130.500 22.990 130.790 23.280 ;
        RECT 131.010 22.990 131.300 23.280 ;
        RECT 132.500 22.990 132.790 23.280 ;
        RECT 1.060 21.925 1.260 22.990 ;
        RECT 2.545 21.925 2.745 22.990 ;
        RECT 1.060 21.725 1.705 21.925 ;
        RECT 1.415 21.635 1.705 21.725 ;
        RECT 2.095 21.725 2.745 21.925 ;
        RECT 3.060 21.925 3.260 22.990 ;
        RECT 4.545 21.925 4.745 22.990 ;
        RECT 3.060 21.725 3.705 21.925 ;
        RECT 2.095 21.635 2.385 21.725 ;
        RECT 3.415 21.635 3.705 21.725 ;
        RECT 4.095 21.725 4.745 21.925 ;
        RECT 5.060 21.925 5.260 22.990 ;
        RECT 6.545 21.925 6.745 22.990 ;
        RECT 5.060 21.725 5.705 21.925 ;
        RECT 4.095 21.635 4.385 21.725 ;
        RECT 5.415 21.635 5.705 21.725 ;
        RECT 6.095 21.725 6.745 21.925 ;
        RECT 7.060 21.925 7.260 22.990 ;
        RECT 8.545 21.925 8.745 22.990 ;
        RECT 7.060 21.725 7.705 21.925 ;
        RECT 6.095 21.635 6.385 21.725 ;
        RECT 7.415 21.635 7.705 21.725 ;
        RECT 8.095 21.725 8.745 21.925 ;
        RECT 9.060 21.925 9.260 22.990 ;
        RECT 10.545 21.925 10.745 22.990 ;
        RECT 9.060 21.725 9.705 21.925 ;
        RECT 8.095 21.635 8.385 21.725 ;
        RECT 9.415 21.635 9.705 21.725 ;
        RECT 10.095 21.725 10.745 21.925 ;
        RECT 11.060 21.925 11.260 22.990 ;
        RECT 12.545 21.925 12.745 22.990 ;
        RECT 11.060 21.725 11.705 21.925 ;
        RECT 10.095 21.635 10.385 21.725 ;
        RECT 11.415 21.635 11.705 21.725 ;
        RECT 12.095 21.725 12.745 21.925 ;
        RECT 13.060 21.925 13.260 22.990 ;
        RECT 14.545 21.925 14.745 22.990 ;
        RECT 13.060 21.725 13.705 21.925 ;
        RECT 12.095 21.635 12.385 21.725 ;
        RECT 13.415 21.635 13.705 21.725 ;
        RECT 14.095 21.725 14.745 21.925 ;
        RECT 15.060 21.925 15.260 22.990 ;
        RECT 16.545 21.925 16.745 22.990 ;
        RECT 15.060 21.725 15.705 21.925 ;
        RECT 14.095 21.635 14.385 21.725 ;
        RECT 15.415 21.635 15.705 21.725 ;
        RECT 16.095 21.725 16.745 21.925 ;
        RECT 17.060 21.925 17.260 22.990 ;
        RECT 18.545 21.925 18.745 22.990 ;
        RECT 17.060 21.725 17.705 21.925 ;
        RECT 16.095 21.635 16.385 21.725 ;
        RECT 17.415 21.635 17.705 21.725 ;
        RECT 18.095 21.725 18.745 21.925 ;
        RECT 19.060 21.925 19.260 22.990 ;
        RECT 20.545 21.925 20.745 22.990 ;
        RECT 19.060 21.725 19.705 21.925 ;
        RECT 18.095 21.635 18.385 21.725 ;
        RECT 19.415 21.635 19.705 21.725 ;
        RECT 20.095 21.725 20.745 21.925 ;
        RECT 21.060 21.925 21.260 22.990 ;
        RECT 22.545 21.925 22.745 22.990 ;
        RECT 21.060 21.725 21.705 21.925 ;
        RECT 20.095 21.635 20.385 21.725 ;
        RECT 21.415 21.635 21.705 21.725 ;
        RECT 22.095 21.725 22.745 21.925 ;
        RECT 23.060 21.925 23.260 22.990 ;
        RECT 24.545 21.925 24.745 22.990 ;
        RECT 23.060 21.725 23.705 21.925 ;
        RECT 22.095 21.635 22.385 21.725 ;
        RECT 23.415 21.635 23.705 21.725 ;
        RECT 24.095 21.725 24.745 21.925 ;
        RECT 25.060 21.925 25.260 22.990 ;
        RECT 26.545 21.925 26.745 22.990 ;
        RECT 25.060 21.725 25.705 21.925 ;
        RECT 24.095 21.635 24.385 21.725 ;
        RECT 25.415 21.635 25.705 21.725 ;
        RECT 26.095 21.725 26.745 21.925 ;
        RECT 27.060 21.925 27.260 22.990 ;
        RECT 28.545 21.925 28.745 22.990 ;
        RECT 27.060 21.725 27.705 21.925 ;
        RECT 26.095 21.635 26.385 21.725 ;
        RECT 27.415 21.635 27.705 21.725 ;
        RECT 28.095 21.725 28.745 21.925 ;
        RECT 29.060 21.925 29.260 22.990 ;
        RECT 30.545 21.925 30.745 22.990 ;
        RECT 29.060 21.725 29.705 21.925 ;
        RECT 28.095 21.635 28.385 21.725 ;
        RECT 29.415 21.635 29.705 21.725 ;
        RECT 30.095 21.725 30.745 21.925 ;
        RECT 31.060 21.925 31.260 22.990 ;
        RECT 32.545 21.925 32.745 22.990 ;
        RECT 31.060 21.725 31.705 21.925 ;
        RECT 30.095 21.635 30.385 21.725 ;
        RECT 31.415 21.635 31.705 21.725 ;
        RECT 32.095 21.725 32.745 21.925 ;
        RECT 33.060 21.925 33.260 22.990 ;
        RECT 34.545 21.925 34.745 22.990 ;
        RECT 33.060 21.725 33.705 21.925 ;
        RECT 32.095 21.635 32.385 21.725 ;
        RECT 33.415 21.635 33.705 21.725 ;
        RECT 34.095 21.725 34.745 21.925 ;
        RECT 35.060 21.925 35.260 22.990 ;
        RECT 36.545 21.925 36.745 22.990 ;
        RECT 35.060 21.725 35.705 21.925 ;
        RECT 34.095 21.635 34.385 21.725 ;
        RECT 35.415 21.635 35.705 21.725 ;
        RECT 36.095 21.725 36.745 21.925 ;
        RECT 37.060 21.925 37.260 22.990 ;
        RECT 38.545 21.925 38.745 22.990 ;
        RECT 37.060 21.725 37.705 21.925 ;
        RECT 36.095 21.635 36.385 21.725 ;
        RECT 37.415 21.635 37.705 21.725 ;
        RECT 38.095 21.725 38.745 21.925 ;
        RECT 39.060 21.925 39.260 22.990 ;
        RECT 40.545 21.925 40.745 22.990 ;
        RECT 39.060 21.725 39.705 21.925 ;
        RECT 38.095 21.635 38.385 21.725 ;
        RECT 39.415 21.635 39.705 21.725 ;
        RECT 40.095 21.725 40.745 21.925 ;
        RECT 41.060 21.925 41.260 22.990 ;
        RECT 42.545 21.925 42.745 22.990 ;
        RECT 41.060 21.725 41.705 21.925 ;
        RECT 40.095 21.635 40.385 21.725 ;
        RECT 41.415 21.635 41.705 21.725 ;
        RECT 42.095 21.725 42.745 21.925 ;
        RECT 43.060 21.925 43.260 22.990 ;
        RECT 44.545 21.925 44.745 22.990 ;
        RECT 43.060 21.725 43.705 21.925 ;
        RECT 42.095 21.635 42.385 21.725 ;
        RECT 43.415 21.635 43.705 21.725 ;
        RECT 44.095 21.725 44.745 21.925 ;
        RECT 45.060 21.925 45.260 22.990 ;
        RECT 46.545 21.925 46.745 22.990 ;
        RECT 45.060 21.725 45.705 21.925 ;
        RECT 44.095 21.635 44.385 21.725 ;
        RECT 45.415 21.635 45.705 21.725 ;
        RECT 46.095 21.725 46.745 21.925 ;
        RECT 47.060 21.925 47.260 22.990 ;
        RECT 48.545 21.925 48.745 22.990 ;
        RECT 47.060 21.725 47.705 21.925 ;
        RECT 46.095 21.635 46.385 21.725 ;
        RECT 47.415 21.635 47.705 21.725 ;
        RECT 48.095 21.725 48.745 21.925 ;
        RECT 49.060 21.925 49.260 22.990 ;
        RECT 50.545 21.925 50.745 22.990 ;
        RECT 49.060 21.725 49.705 21.925 ;
        RECT 48.095 21.635 48.385 21.725 ;
        RECT 49.415 21.635 49.705 21.725 ;
        RECT 50.095 21.725 50.745 21.925 ;
        RECT 51.060 21.925 51.260 22.990 ;
        RECT 52.545 21.925 52.745 22.990 ;
        RECT 51.060 21.725 51.705 21.925 ;
        RECT 50.095 21.635 50.385 21.725 ;
        RECT 51.415 21.635 51.705 21.725 ;
        RECT 52.095 21.725 52.745 21.925 ;
        RECT 53.060 21.925 53.260 22.990 ;
        RECT 54.545 21.925 54.745 22.990 ;
        RECT 53.060 21.725 53.705 21.925 ;
        RECT 52.095 21.635 52.385 21.725 ;
        RECT 53.415 21.635 53.705 21.725 ;
        RECT 54.095 21.725 54.745 21.925 ;
        RECT 55.060 21.925 55.260 22.990 ;
        RECT 56.545 21.925 56.745 22.990 ;
        RECT 55.060 21.725 55.705 21.925 ;
        RECT 54.095 21.635 54.385 21.725 ;
        RECT 55.415 21.635 55.705 21.725 ;
        RECT 56.095 21.725 56.745 21.925 ;
        RECT 57.060 21.925 57.260 22.990 ;
        RECT 58.545 21.925 58.745 22.990 ;
        RECT 57.060 21.725 57.705 21.925 ;
        RECT 56.095 21.635 56.385 21.725 ;
        RECT 57.415 21.635 57.705 21.725 ;
        RECT 58.095 21.725 58.745 21.925 ;
        RECT 59.060 21.925 59.260 22.990 ;
        RECT 60.545 21.925 60.745 22.990 ;
        RECT 59.060 21.725 59.705 21.925 ;
        RECT 58.095 21.635 58.385 21.725 ;
        RECT 59.415 21.635 59.705 21.725 ;
        RECT 60.095 21.725 60.745 21.925 ;
        RECT 61.060 21.925 61.260 22.990 ;
        RECT 62.545 21.925 62.745 22.990 ;
        RECT 61.060 21.725 61.705 21.925 ;
        RECT 60.095 21.635 60.385 21.725 ;
        RECT 61.415 21.635 61.705 21.725 ;
        RECT 62.095 21.725 62.745 21.925 ;
        RECT 63.060 21.925 63.260 22.990 ;
        RECT 64.545 21.925 64.745 22.990 ;
        RECT 63.060 21.725 63.705 21.925 ;
        RECT 62.095 21.635 62.385 21.725 ;
        RECT 63.415 21.635 63.705 21.725 ;
        RECT 64.095 21.725 64.745 21.925 ;
        RECT 65.060 21.925 65.260 22.990 ;
        RECT 66.545 21.925 66.745 22.990 ;
        RECT 65.060 21.725 65.705 21.925 ;
        RECT 64.095 21.635 64.385 21.725 ;
        RECT 65.415 21.635 65.705 21.725 ;
        RECT 66.095 21.725 66.745 21.925 ;
        RECT 67.060 21.925 67.260 22.990 ;
        RECT 68.545 21.925 68.745 22.990 ;
        RECT 67.060 21.725 67.705 21.925 ;
        RECT 66.095 21.635 66.385 21.725 ;
        RECT 67.415 21.635 67.705 21.725 ;
        RECT 68.095 21.725 68.745 21.925 ;
        RECT 69.060 21.925 69.260 22.990 ;
        RECT 70.545 21.925 70.745 22.990 ;
        RECT 69.060 21.725 69.705 21.925 ;
        RECT 68.095 21.635 68.385 21.725 ;
        RECT 69.415 21.635 69.705 21.725 ;
        RECT 70.095 21.725 70.745 21.925 ;
        RECT 71.060 21.925 71.260 22.990 ;
        RECT 72.545 21.925 72.745 22.990 ;
        RECT 71.060 21.725 71.705 21.925 ;
        RECT 70.095 21.635 70.385 21.725 ;
        RECT 71.415 21.635 71.705 21.725 ;
        RECT 72.095 21.725 72.745 21.925 ;
        RECT 73.060 21.925 73.260 22.990 ;
        RECT 74.545 21.925 74.745 22.990 ;
        RECT 73.060 21.725 73.705 21.925 ;
        RECT 72.095 21.635 72.385 21.725 ;
        RECT 73.415 21.635 73.705 21.725 ;
        RECT 74.095 21.725 74.745 21.925 ;
        RECT 75.060 21.925 75.260 22.990 ;
        RECT 76.545 21.925 76.745 22.990 ;
        RECT 75.060 21.725 75.705 21.925 ;
        RECT 74.095 21.635 74.385 21.725 ;
        RECT 75.415 21.635 75.705 21.725 ;
        RECT 76.095 21.725 76.745 21.925 ;
        RECT 77.060 21.925 77.260 22.990 ;
        RECT 78.545 21.925 78.745 22.990 ;
        RECT 77.060 21.725 77.705 21.925 ;
        RECT 76.095 21.635 76.385 21.725 ;
        RECT 77.415 21.635 77.705 21.725 ;
        RECT 78.095 21.725 78.745 21.925 ;
        RECT 79.060 21.925 79.260 22.990 ;
        RECT 80.545 21.925 80.745 22.990 ;
        RECT 79.060 21.725 79.705 21.925 ;
        RECT 78.095 21.635 78.385 21.725 ;
        RECT 79.415 21.635 79.705 21.725 ;
        RECT 80.095 21.725 80.745 21.925 ;
        RECT 81.060 21.925 81.260 22.990 ;
        RECT 82.545 21.925 82.745 22.990 ;
        RECT 81.060 21.725 81.705 21.925 ;
        RECT 80.095 21.635 80.385 21.725 ;
        RECT 81.415 21.635 81.705 21.725 ;
        RECT 82.095 21.725 82.745 21.925 ;
        RECT 83.060 21.925 83.260 22.990 ;
        RECT 84.545 21.925 84.745 22.990 ;
        RECT 83.060 21.725 83.705 21.925 ;
        RECT 82.095 21.635 82.385 21.725 ;
        RECT 83.415 21.635 83.705 21.725 ;
        RECT 84.095 21.725 84.745 21.925 ;
        RECT 85.060 21.925 85.260 22.990 ;
        RECT 86.545 21.925 86.745 22.990 ;
        RECT 85.060 21.725 85.705 21.925 ;
        RECT 84.095 21.635 84.385 21.725 ;
        RECT 85.415 21.635 85.705 21.725 ;
        RECT 86.095 21.725 86.745 21.925 ;
        RECT 87.060 21.925 87.260 22.990 ;
        RECT 88.545 21.925 88.745 22.990 ;
        RECT 87.060 21.725 87.705 21.925 ;
        RECT 86.095 21.635 86.385 21.725 ;
        RECT 87.415 21.635 87.705 21.725 ;
        RECT 88.095 21.725 88.745 21.925 ;
        RECT 89.060 21.925 89.260 22.990 ;
        RECT 90.545 21.925 90.745 22.990 ;
        RECT 89.060 21.725 89.705 21.925 ;
        RECT 88.095 21.635 88.385 21.725 ;
        RECT 89.415 21.635 89.705 21.725 ;
        RECT 90.095 21.725 90.745 21.925 ;
        RECT 91.060 21.925 91.260 22.990 ;
        RECT 92.545 21.925 92.745 22.990 ;
        RECT 91.060 21.725 91.705 21.925 ;
        RECT 90.095 21.635 90.385 21.725 ;
        RECT 91.415 21.635 91.705 21.725 ;
        RECT 92.095 21.725 92.745 21.925 ;
        RECT 93.060 21.925 93.260 22.990 ;
        RECT 94.545 21.925 94.745 22.990 ;
        RECT 93.060 21.725 93.705 21.925 ;
        RECT 92.095 21.635 92.385 21.725 ;
        RECT 93.415 21.635 93.705 21.725 ;
        RECT 94.095 21.725 94.745 21.925 ;
        RECT 95.060 21.925 95.260 22.990 ;
        RECT 96.545 21.925 96.745 22.990 ;
        RECT 95.060 21.725 95.705 21.925 ;
        RECT 94.095 21.635 94.385 21.725 ;
        RECT 95.415 21.635 95.705 21.725 ;
        RECT 96.095 21.725 96.745 21.925 ;
        RECT 97.060 21.925 97.260 22.990 ;
        RECT 98.545 21.925 98.745 22.990 ;
        RECT 97.060 21.725 97.705 21.925 ;
        RECT 96.095 21.635 96.385 21.725 ;
        RECT 97.415 21.635 97.705 21.725 ;
        RECT 98.095 21.725 98.745 21.925 ;
        RECT 99.060 21.925 99.260 22.990 ;
        RECT 100.545 21.925 100.745 22.990 ;
        RECT 99.060 21.725 99.705 21.925 ;
        RECT 98.095 21.635 98.385 21.725 ;
        RECT 99.415 21.635 99.705 21.725 ;
        RECT 100.095 21.725 100.745 21.925 ;
        RECT 101.060 21.925 101.260 22.990 ;
        RECT 102.545 21.925 102.745 22.990 ;
        RECT 101.060 21.725 101.705 21.925 ;
        RECT 100.095 21.635 100.385 21.725 ;
        RECT 101.415 21.635 101.705 21.725 ;
        RECT 102.095 21.725 102.745 21.925 ;
        RECT 103.060 21.925 103.260 22.990 ;
        RECT 104.545 21.925 104.745 22.990 ;
        RECT 103.060 21.725 103.705 21.925 ;
        RECT 102.095 21.635 102.385 21.725 ;
        RECT 103.415 21.635 103.705 21.725 ;
        RECT 104.095 21.725 104.745 21.925 ;
        RECT 105.060 21.925 105.260 22.990 ;
        RECT 106.545 21.925 106.745 22.990 ;
        RECT 105.060 21.725 105.705 21.925 ;
        RECT 104.095 21.635 104.385 21.725 ;
        RECT 105.415 21.635 105.705 21.725 ;
        RECT 106.095 21.725 106.745 21.925 ;
        RECT 107.060 21.925 107.260 22.990 ;
        RECT 108.545 21.925 108.745 22.990 ;
        RECT 107.060 21.725 107.705 21.925 ;
        RECT 106.095 21.635 106.385 21.725 ;
        RECT 107.415 21.635 107.705 21.725 ;
        RECT 108.095 21.725 108.745 21.925 ;
        RECT 109.060 21.925 109.260 22.990 ;
        RECT 110.545 21.925 110.745 22.990 ;
        RECT 109.060 21.725 109.705 21.925 ;
        RECT 108.095 21.635 108.385 21.725 ;
        RECT 109.415 21.635 109.705 21.725 ;
        RECT 110.095 21.725 110.745 21.925 ;
        RECT 111.060 21.925 111.260 22.990 ;
        RECT 112.545 21.925 112.745 22.990 ;
        RECT 111.060 21.725 111.705 21.925 ;
        RECT 110.095 21.635 110.385 21.725 ;
        RECT 111.415 21.635 111.705 21.725 ;
        RECT 112.095 21.725 112.745 21.925 ;
        RECT 113.060 21.925 113.260 22.990 ;
        RECT 114.545 21.925 114.745 22.990 ;
        RECT 113.060 21.725 113.705 21.925 ;
        RECT 112.095 21.635 112.385 21.725 ;
        RECT 113.415 21.635 113.705 21.725 ;
        RECT 114.095 21.725 114.745 21.925 ;
        RECT 115.060 21.925 115.260 22.990 ;
        RECT 116.545 21.925 116.745 22.990 ;
        RECT 115.060 21.725 115.705 21.925 ;
        RECT 114.095 21.635 114.385 21.725 ;
        RECT 115.415 21.635 115.705 21.725 ;
        RECT 116.095 21.725 116.745 21.925 ;
        RECT 117.060 21.925 117.260 22.990 ;
        RECT 118.545 21.925 118.745 22.990 ;
        RECT 117.060 21.725 117.705 21.925 ;
        RECT 116.095 21.635 116.385 21.725 ;
        RECT 117.415 21.635 117.705 21.725 ;
        RECT 118.095 21.725 118.745 21.925 ;
        RECT 119.060 21.925 119.260 22.990 ;
        RECT 120.545 21.925 120.745 22.990 ;
        RECT 119.060 21.725 119.705 21.925 ;
        RECT 118.095 21.635 118.385 21.725 ;
        RECT 119.415 21.635 119.705 21.725 ;
        RECT 120.095 21.725 120.745 21.925 ;
        RECT 121.060 21.925 121.260 22.990 ;
        RECT 122.545 21.925 122.745 22.990 ;
        RECT 121.060 21.725 121.705 21.925 ;
        RECT 120.095 21.635 120.385 21.725 ;
        RECT 121.415 21.635 121.705 21.725 ;
        RECT 122.095 21.725 122.745 21.925 ;
        RECT 123.060 21.925 123.260 22.990 ;
        RECT 124.545 21.925 124.745 22.990 ;
        RECT 123.060 21.725 123.705 21.925 ;
        RECT 122.095 21.635 122.385 21.725 ;
        RECT 123.415 21.635 123.705 21.725 ;
        RECT 124.095 21.725 124.745 21.925 ;
        RECT 125.060 21.925 125.260 22.990 ;
        RECT 126.545 21.925 126.745 22.990 ;
        RECT 125.060 21.725 125.705 21.925 ;
        RECT 124.095 21.635 124.385 21.725 ;
        RECT 125.415 21.635 125.705 21.725 ;
        RECT 126.095 21.725 126.745 21.925 ;
        RECT 127.060 21.925 127.260 22.990 ;
        RECT 128.545 21.925 128.745 22.990 ;
        RECT 127.060 21.725 127.705 21.925 ;
        RECT 126.095 21.635 126.385 21.725 ;
        RECT 127.415 21.635 127.705 21.725 ;
        RECT 128.095 21.725 128.745 21.925 ;
        RECT 129.060 21.925 129.260 22.990 ;
        RECT 130.545 21.925 130.745 22.990 ;
        RECT 129.060 21.725 129.705 21.925 ;
        RECT 128.095 21.635 128.385 21.725 ;
        RECT 129.415 21.635 129.705 21.725 ;
        RECT 130.095 21.725 130.745 21.925 ;
        RECT 131.060 21.925 131.260 22.990 ;
        RECT 132.545 21.925 132.745 22.990 ;
        RECT 131.060 21.725 131.705 21.925 ;
        RECT 130.095 21.635 130.385 21.725 ;
        RECT 131.415 21.635 131.705 21.725 ;
        RECT 132.095 21.725 132.745 21.925 ;
        RECT 132.095 21.635 132.385 21.725 ;
        RECT 1.755 21.135 2.045 21.425 ;
        RECT 3.755 21.135 4.045 21.425 ;
        RECT 5.755 21.135 6.045 21.425 ;
        RECT 7.755 21.135 8.045 21.425 ;
        RECT 9.755 21.135 10.045 21.425 ;
        RECT 11.755 21.135 12.045 21.425 ;
        RECT 13.755 21.135 14.045 21.425 ;
        RECT 15.755 21.135 16.045 21.425 ;
        RECT 17.755 21.135 18.045 21.425 ;
        RECT 19.755 21.135 20.045 21.425 ;
        RECT 21.755 21.135 22.045 21.425 ;
        RECT 23.755 21.135 24.045 21.425 ;
        RECT 25.755 21.135 26.045 21.425 ;
        RECT 27.755 21.135 28.045 21.425 ;
        RECT 29.755 21.135 30.045 21.425 ;
        RECT 31.755 21.135 32.045 21.425 ;
        RECT 33.755 21.135 34.045 21.425 ;
        RECT 35.755 21.135 36.045 21.425 ;
        RECT 37.755 21.135 38.045 21.425 ;
        RECT 39.755 21.135 40.045 21.425 ;
        RECT 41.755 21.135 42.045 21.425 ;
        RECT 43.755 21.135 44.045 21.425 ;
        RECT 45.755 21.135 46.045 21.425 ;
        RECT 47.755 21.135 48.045 21.425 ;
        RECT 49.755 21.135 50.045 21.425 ;
        RECT 51.755 21.135 52.045 21.425 ;
        RECT 53.755 21.135 54.045 21.425 ;
        RECT 55.755 21.135 56.045 21.425 ;
        RECT 57.755 21.135 58.045 21.425 ;
        RECT 59.755 21.135 60.045 21.425 ;
        RECT 61.755 21.135 62.045 21.425 ;
        RECT 63.755 21.135 64.045 21.425 ;
        RECT 65.755 21.135 66.045 21.425 ;
        RECT 67.755 21.135 68.045 21.425 ;
        RECT 69.755 21.135 70.045 21.425 ;
        RECT 71.755 21.135 72.045 21.425 ;
        RECT 73.755 21.135 74.045 21.425 ;
        RECT 75.755 21.135 76.045 21.425 ;
        RECT 77.755 21.135 78.045 21.425 ;
        RECT 79.755 21.135 80.045 21.425 ;
        RECT 81.755 21.135 82.045 21.425 ;
        RECT 83.755 21.135 84.045 21.425 ;
        RECT 85.755 21.135 86.045 21.425 ;
        RECT 87.755 21.135 88.045 21.425 ;
        RECT 89.755 21.135 90.045 21.425 ;
        RECT 91.755 21.135 92.045 21.425 ;
        RECT 93.755 21.135 94.045 21.425 ;
        RECT 95.755 21.135 96.045 21.425 ;
        RECT 97.755 21.135 98.045 21.425 ;
        RECT 99.755 21.135 100.045 21.425 ;
        RECT 101.755 21.135 102.045 21.425 ;
        RECT 103.755 21.135 104.045 21.425 ;
        RECT 105.755 21.135 106.045 21.425 ;
        RECT 107.755 21.135 108.045 21.425 ;
        RECT 109.755 21.135 110.045 21.425 ;
        RECT 111.755 21.135 112.045 21.425 ;
        RECT 113.755 21.135 114.045 21.425 ;
        RECT 115.755 21.135 116.045 21.425 ;
        RECT 117.755 21.135 118.045 21.425 ;
        RECT 119.755 21.135 120.045 21.425 ;
        RECT 121.755 21.135 122.045 21.425 ;
        RECT 123.755 21.135 124.045 21.425 ;
        RECT 125.755 21.135 126.045 21.425 ;
        RECT 127.755 21.135 128.045 21.425 ;
        RECT 129.755 21.135 130.045 21.425 ;
        RECT 131.755 21.135 132.045 21.425 ;
        RECT 1.800 20.495 2.000 21.135 ;
        RECT 3.800 20.495 4.000 21.135 ;
        RECT 5.800 20.495 6.000 21.135 ;
        RECT 7.800 20.495 8.000 21.135 ;
        RECT 9.800 20.495 10.000 21.135 ;
        RECT 11.800 20.495 12.000 21.135 ;
        RECT 13.800 20.495 14.000 21.135 ;
        RECT 15.800 20.495 16.000 21.135 ;
        RECT 17.800 20.495 18.000 21.135 ;
        RECT 19.800 20.495 20.000 21.135 ;
        RECT 21.800 20.495 22.000 21.135 ;
        RECT 23.800 20.495 24.000 21.135 ;
        RECT 25.800 20.495 26.000 21.135 ;
        RECT 27.800 20.495 28.000 21.135 ;
        RECT 29.800 20.495 30.000 21.135 ;
        RECT 31.800 20.495 32.000 21.135 ;
        RECT 33.800 20.495 34.000 21.135 ;
        RECT 35.800 20.495 36.000 21.135 ;
        RECT 37.800 20.495 38.000 21.135 ;
        RECT 39.800 20.495 40.000 21.135 ;
        RECT 41.800 20.495 42.000 21.135 ;
        RECT 43.800 20.495 44.000 21.135 ;
        RECT 45.800 20.495 46.000 21.135 ;
        RECT 47.800 20.495 48.000 21.135 ;
        RECT 49.800 20.495 50.000 21.135 ;
        RECT 51.800 20.495 52.000 21.135 ;
        RECT 53.800 20.495 54.000 21.135 ;
        RECT 55.800 20.495 56.000 21.135 ;
        RECT 57.800 20.495 58.000 21.135 ;
        RECT 59.800 20.495 60.000 21.135 ;
        RECT 61.800 20.495 62.000 21.135 ;
        RECT 63.800 20.495 64.000 21.135 ;
        RECT 65.800 20.495 66.000 21.135 ;
        RECT 67.800 20.495 68.000 21.135 ;
        RECT 69.800 20.495 70.000 21.135 ;
        RECT 71.800 20.495 72.000 21.135 ;
        RECT 73.800 20.495 74.000 21.135 ;
        RECT 75.800 20.495 76.000 21.135 ;
        RECT 77.800 20.495 78.000 21.135 ;
        RECT 79.800 20.495 80.000 21.135 ;
        RECT 81.800 20.495 82.000 21.135 ;
        RECT 83.800 20.495 84.000 21.135 ;
        RECT 85.800 20.495 86.000 21.135 ;
        RECT 87.800 20.495 88.000 21.135 ;
        RECT 89.800 20.495 90.000 21.135 ;
        RECT 91.800 20.495 92.000 21.135 ;
        RECT 93.800 20.495 94.000 21.135 ;
        RECT 95.800 20.495 96.000 21.135 ;
        RECT 97.800 20.495 98.000 21.135 ;
        RECT 99.800 20.495 100.000 21.135 ;
        RECT 101.800 20.495 102.000 21.135 ;
        RECT 103.800 20.495 104.000 21.135 ;
        RECT 105.800 20.495 106.000 21.135 ;
        RECT 107.800 20.495 108.000 21.135 ;
        RECT 109.800 20.495 110.000 21.135 ;
        RECT 111.800 20.495 112.000 21.135 ;
        RECT 113.800 20.495 114.000 21.135 ;
        RECT 115.800 20.495 116.000 21.135 ;
        RECT 117.800 20.495 118.000 21.135 ;
        RECT 119.800 20.495 120.000 21.135 ;
        RECT 121.800 20.495 122.000 21.135 ;
        RECT 123.800 20.495 124.000 21.135 ;
        RECT 125.800 20.495 126.000 21.135 ;
        RECT 127.800 20.495 128.000 21.135 ;
        RECT 129.800 20.495 130.000 21.135 ;
        RECT 131.800 20.495 132.000 21.135 ;
        RECT 1.800 20.295 2.670 20.495 ;
        RECT 3.800 20.295 4.670 20.495 ;
        RECT 5.800 20.295 6.670 20.495 ;
        RECT 7.800 20.295 8.670 20.495 ;
        RECT 9.800 20.295 10.670 20.495 ;
        RECT 11.800 20.295 12.670 20.495 ;
        RECT 13.800 20.295 14.670 20.495 ;
        RECT 15.800 20.295 16.670 20.495 ;
        RECT 17.800 20.295 18.670 20.495 ;
        RECT 19.800 20.295 20.670 20.495 ;
        RECT 21.800 20.295 22.670 20.495 ;
        RECT 23.800 20.295 24.670 20.495 ;
        RECT 25.800 20.295 26.670 20.495 ;
        RECT 27.800 20.295 28.670 20.495 ;
        RECT 29.800 20.295 30.670 20.495 ;
        RECT 31.800 20.295 32.670 20.495 ;
        RECT 33.800 20.295 34.670 20.495 ;
        RECT 35.800 20.295 36.670 20.495 ;
        RECT 37.800 20.295 38.670 20.495 ;
        RECT 39.800 20.295 40.670 20.495 ;
        RECT 41.800 20.295 42.670 20.495 ;
        RECT 43.800 20.295 44.670 20.495 ;
        RECT 45.800 20.295 46.670 20.495 ;
        RECT 47.800 20.295 48.670 20.495 ;
        RECT 49.800 20.295 50.670 20.495 ;
        RECT 51.800 20.295 52.670 20.495 ;
        RECT 53.800 20.295 54.670 20.495 ;
        RECT 55.800 20.295 56.670 20.495 ;
        RECT 57.800 20.295 58.670 20.495 ;
        RECT 59.800 20.295 60.670 20.495 ;
        RECT 61.800 20.295 62.670 20.495 ;
        RECT 63.800 20.295 64.670 20.495 ;
        RECT 65.800 20.295 66.670 20.495 ;
        RECT 67.800 20.295 68.670 20.495 ;
        RECT 69.800 20.295 70.670 20.495 ;
        RECT 71.800 20.295 72.670 20.495 ;
        RECT 73.800 20.295 74.670 20.495 ;
        RECT 75.800 20.295 76.670 20.495 ;
        RECT 77.800 20.295 78.670 20.495 ;
        RECT 79.800 20.295 80.670 20.495 ;
        RECT 81.800 20.295 82.670 20.495 ;
        RECT 83.800 20.295 84.670 20.495 ;
        RECT 85.800 20.295 86.670 20.495 ;
        RECT 87.800 20.295 88.670 20.495 ;
        RECT 89.800 20.295 90.670 20.495 ;
        RECT 91.800 20.295 92.670 20.495 ;
        RECT 93.800 20.295 94.670 20.495 ;
        RECT 95.800 20.295 96.670 20.495 ;
        RECT 97.800 20.295 98.670 20.495 ;
        RECT 99.800 20.295 100.670 20.495 ;
        RECT 101.800 20.295 102.670 20.495 ;
        RECT 103.800 20.295 104.670 20.495 ;
        RECT 105.800 20.295 106.670 20.495 ;
        RECT 107.800 20.295 108.670 20.495 ;
        RECT 109.800 20.295 110.670 20.495 ;
        RECT 111.800 20.295 112.670 20.495 ;
        RECT 113.800 20.295 114.670 20.495 ;
        RECT 115.800 20.295 116.670 20.495 ;
        RECT 117.800 20.295 118.670 20.495 ;
        RECT 119.800 20.295 120.670 20.495 ;
        RECT 121.800 20.295 122.670 20.495 ;
        RECT 123.800 20.295 124.670 20.495 ;
        RECT 125.800 20.295 126.670 20.495 ;
        RECT 127.800 20.295 128.670 20.495 ;
        RECT 129.800 20.295 130.670 20.495 ;
        RECT 131.800 20.295 132.670 20.495 ;
        RECT 2.470 14.645 2.670 20.295 ;
        RECT 4.470 14.645 4.670 20.295 ;
        RECT 6.470 14.645 6.670 20.295 ;
        RECT 8.470 14.645 8.670 20.295 ;
        RECT 10.470 14.645 10.670 20.295 ;
        RECT 12.470 14.645 12.670 20.295 ;
        RECT 14.470 14.645 14.670 20.295 ;
        RECT 16.470 14.645 16.670 20.295 ;
        RECT 18.470 14.645 18.670 20.295 ;
        RECT 20.470 14.645 20.670 20.295 ;
        RECT 22.470 14.645 22.670 20.295 ;
        RECT 24.470 14.645 24.670 20.295 ;
        RECT 26.470 14.645 26.670 20.295 ;
        RECT 28.470 14.645 28.670 20.295 ;
        RECT 30.470 14.645 30.670 20.295 ;
        RECT 32.470 14.645 32.670 20.295 ;
        RECT 34.470 14.645 34.670 20.295 ;
        RECT 36.470 14.645 36.670 20.295 ;
        RECT 38.470 14.645 38.670 20.295 ;
        RECT 40.470 14.645 40.670 20.295 ;
        RECT 42.470 14.645 42.670 20.295 ;
        RECT 44.470 14.645 44.670 20.295 ;
        RECT 46.470 14.645 46.670 20.295 ;
        RECT 48.470 14.645 48.670 20.295 ;
        RECT 50.470 14.645 50.670 20.295 ;
        RECT 52.470 14.645 52.670 20.295 ;
        RECT 54.470 14.645 54.670 20.295 ;
        RECT 56.470 14.645 56.670 20.295 ;
        RECT 58.470 14.645 58.670 20.295 ;
        RECT 60.470 14.645 60.670 20.295 ;
        RECT 62.470 14.645 62.670 20.295 ;
        RECT 64.470 14.645 64.670 20.295 ;
        RECT 66.470 14.645 66.670 20.295 ;
        RECT 68.470 14.645 68.670 20.295 ;
        RECT 70.470 14.645 70.670 20.295 ;
        RECT 72.470 14.645 72.670 20.295 ;
        RECT 74.470 14.645 74.670 20.295 ;
        RECT 76.470 14.645 76.670 20.295 ;
        RECT 78.470 14.645 78.670 20.295 ;
        RECT 80.470 14.645 80.670 20.295 ;
        RECT 82.470 14.645 82.670 20.295 ;
        RECT 84.470 14.645 84.670 20.295 ;
        RECT 86.470 14.645 86.670 20.295 ;
        RECT 88.470 14.645 88.670 20.295 ;
        RECT 90.470 14.645 90.670 20.295 ;
        RECT 92.470 14.645 92.670 20.295 ;
        RECT 94.470 14.645 94.670 20.295 ;
        RECT 96.470 14.645 96.670 20.295 ;
        RECT 98.470 14.645 98.670 20.295 ;
        RECT 100.470 14.645 100.670 20.295 ;
        RECT 102.470 14.645 102.670 20.295 ;
        RECT 104.470 14.645 104.670 20.295 ;
        RECT 106.470 14.645 106.670 20.295 ;
        RECT 108.470 14.645 108.670 20.295 ;
        RECT 110.470 14.645 110.670 20.295 ;
        RECT 112.470 14.645 112.670 20.295 ;
        RECT 114.470 14.645 114.670 20.295 ;
        RECT 116.470 14.645 116.670 20.295 ;
        RECT 118.470 14.645 118.670 20.295 ;
        RECT 120.470 14.645 120.670 20.295 ;
        RECT 122.470 14.645 122.670 20.295 ;
        RECT 124.470 14.645 124.670 20.295 ;
        RECT 126.470 14.645 126.670 20.295 ;
        RECT 128.470 14.645 128.670 20.295 ;
        RECT 130.470 14.645 130.670 20.295 ;
        RECT 132.470 14.645 132.670 20.295 ;
        RECT 2.460 14.055 2.680 14.645 ;
        RECT 4.460 14.055 4.680 14.645 ;
        RECT 6.460 14.055 6.680 14.645 ;
        RECT 8.460 14.055 8.680 14.645 ;
        RECT 10.460 14.055 10.680 14.645 ;
        RECT 12.460 14.055 12.680 14.645 ;
        RECT 14.460 14.055 14.680 14.645 ;
        RECT 16.460 14.055 16.680 14.645 ;
        RECT 18.460 14.055 18.680 14.645 ;
        RECT 20.460 14.055 20.680 14.645 ;
        RECT 22.460 14.055 22.680 14.645 ;
        RECT 24.460 14.055 24.680 14.645 ;
        RECT 26.460 14.055 26.680 14.645 ;
        RECT 28.460 14.055 28.680 14.645 ;
        RECT 30.460 14.055 30.680 14.645 ;
        RECT 32.460 14.055 32.680 14.645 ;
        RECT 34.460 14.055 34.680 14.645 ;
        RECT 36.460 14.055 36.680 14.645 ;
        RECT 38.460 14.055 38.680 14.645 ;
        RECT 40.460 14.055 40.680 14.645 ;
        RECT 42.460 14.055 42.680 14.645 ;
        RECT 44.460 14.055 44.680 14.645 ;
        RECT 46.460 14.055 46.680 14.645 ;
        RECT 48.460 14.055 48.680 14.645 ;
        RECT 50.460 14.055 50.680 14.645 ;
        RECT 52.460 14.055 52.680 14.645 ;
        RECT 54.460 14.055 54.680 14.645 ;
        RECT 56.460 14.055 56.680 14.645 ;
        RECT 58.460 14.055 58.680 14.645 ;
        RECT 60.460 14.055 60.680 14.645 ;
        RECT 62.460 14.055 62.680 14.645 ;
        RECT 64.460 14.055 64.680 14.645 ;
        RECT 66.460 14.055 66.680 14.645 ;
        RECT 68.460 14.055 68.680 14.645 ;
        RECT 70.460 14.055 70.680 14.645 ;
        RECT 72.460 14.055 72.680 14.645 ;
        RECT 74.460 14.055 74.680 14.645 ;
        RECT 76.460 14.055 76.680 14.645 ;
        RECT 78.460 14.055 78.680 14.645 ;
        RECT 80.460 14.055 80.680 14.645 ;
        RECT 82.460 14.055 82.680 14.645 ;
        RECT 84.460 14.055 84.680 14.645 ;
        RECT 86.460 14.055 86.680 14.645 ;
        RECT 88.460 14.055 88.680 14.645 ;
        RECT 90.460 14.055 90.680 14.645 ;
        RECT 92.460 14.055 92.680 14.645 ;
        RECT 94.460 14.055 94.680 14.645 ;
        RECT 96.460 14.055 96.680 14.645 ;
        RECT 98.460 14.055 98.680 14.645 ;
        RECT 100.460 14.055 100.680 14.645 ;
        RECT 102.460 14.055 102.680 14.645 ;
        RECT 104.460 14.055 104.680 14.645 ;
        RECT 106.460 14.055 106.680 14.645 ;
        RECT 108.460 14.055 108.680 14.645 ;
        RECT 110.460 14.055 110.680 14.645 ;
        RECT 112.460 14.055 112.680 14.645 ;
        RECT 114.460 14.055 114.680 14.645 ;
        RECT 116.460 14.055 116.680 14.645 ;
        RECT 118.460 14.055 118.680 14.645 ;
        RECT 120.460 14.055 120.680 14.645 ;
        RECT 122.460 14.055 122.680 14.645 ;
        RECT 124.460 14.055 124.680 14.645 ;
        RECT 126.460 14.055 126.680 14.645 ;
        RECT 128.460 14.055 128.680 14.645 ;
        RECT 130.460 14.055 130.680 14.645 ;
        RECT 132.460 14.055 132.680 14.645 ;
        RECT 1.120 11.545 1.340 12.135 ;
        RECT 3.120 11.545 3.340 12.135 ;
        RECT 5.120 11.545 5.340 12.135 ;
        RECT 7.120 11.545 7.340 12.135 ;
        RECT 9.120 11.545 9.340 12.135 ;
        RECT 11.120 11.545 11.340 12.135 ;
        RECT 13.120 11.545 13.340 12.135 ;
        RECT 15.120 11.545 15.340 12.135 ;
        RECT 17.120 11.545 17.340 12.135 ;
        RECT 19.120 11.545 19.340 12.135 ;
        RECT 21.120 11.545 21.340 12.135 ;
        RECT 23.120 11.545 23.340 12.135 ;
        RECT 25.120 11.545 25.340 12.135 ;
        RECT 27.120 11.545 27.340 12.135 ;
        RECT 29.120 11.545 29.340 12.135 ;
        RECT 31.120 11.545 31.340 12.135 ;
        RECT 33.120 11.545 33.340 12.135 ;
        RECT 35.120 11.545 35.340 12.135 ;
        RECT 37.120 11.545 37.340 12.135 ;
        RECT 39.120 11.545 39.340 12.135 ;
        RECT 41.120 11.545 41.340 12.135 ;
        RECT 43.120 11.545 43.340 12.135 ;
        RECT 45.120 11.545 45.340 12.135 ;
        RECT 47.120 11.545 47.340 12.135 ;
        RECT 49.120 11.545 49.340 12.135 ;
        RECT 51.120 11.545 51.340 12.135 ;
        RECT 53.120 11.545 53.340 12.135 ;
        RECT 55.120 11.545 55.340 12.135 ;
        RECT 57.120 11.545 57.340 12.135 ;
        RECT 59.120 11.545 59.340 12.135 ;
        RECT 61.120 11.545 61.340 12.135 ;
        RECT 63.120 11.545 63.340 12.135 ;
        RECT 65.120 11.545 65.340 12.135 ;
        RECT 67.120 11.545 67.340 12.135 ;
        RECT 69.120 11.545 69.340 12.135 ;
        RECT 71.120 11.545 71.340 12.135 ;
        RECT 73.120 11.545 73.340 12.135 ;
        RECT 75.120 11.545 75.340 12.135 ;
        RECT 77.120 11.545 77.340 12.135 ;
        RECT 79.120 11.545 79.340 12.135 ;
        RECT 81.120 11.545 81.340 12.135 ;
        RECT 83.120 11.545 83.340 12.135 ;
        RECT 85.120 11.545 85.340 12.135 ;
        RECT 87.120 11.545 87.340 12.135 ;
        RECT 89.120 11.545 89.340 12.135 ;
        RECT 91.120 11.545 91.340 12.135 ;
        RECT 93.120 11.545 93.340 12.135 ;
        RECT 95.120 11.545 95.340 12.135 ;
        RECT 97.120 11.545 97.340 12.135 ;
        RECT 99.120 11.545 99.340 12.135 ;
        RECT 101.120 11.545 101.340 12.135 ;
        RECT 103.120 11.545 103.340 12.135 ;
        RECT 105.120 11.545 105.340 12.135 ;
        RECT 107.120 11.545 107.340 12.135 ;
        RECT 109.120 11.545 109.340 12.135 ;
        RECT 111.120 11.545 111.340 12.135 ;
        RECT 113.120 11.545 113.340 12.135 ;
        RECT 115.120 11.545 115.340 12.135 ;
        RECT 117.120 11.545 117.340 12.135 ;
        RECT 119.120 11.545 119.340 12.135 ;
        RECT 121.120 11.545 121.340 12.135 ;
        RECT 123.120 11.545 123.340 12.135 ;
        RECT 125.120 11.545 125.340 12.135 ;
        RECT 127.120 11.545 127.340 12.135 ;
        RECT 129.120 11.545 129.340 12.135 ;
        RECT 131.120 11.545 131.340 12.135 ;
        RECT 1.130 5.895 1.330 11.545 ;
        RECT 3.130 5.895 3.330 11.545 ;
        RECT 5.130 5.895 5.330 11.545 ;
        RECT 7.130 5.895 7.330 11.545 ;
        RECT 9.130 5.895 9.330 11.545 ;
        RECT 11.130 5.895 11.330 11.545 ;
        RECT 13.130 5.895 13.330 11.545 ;
        RECT 15.130 5.895 15.330 11.545 ;
        RECT 17.130 5.895 17.330 11.545 ;
        RECT 19.130 5.895 19.330 11.545 ;
        RECT 21.130 5.895 21.330 11.545 ;
        RECT 23.130 5.895 23.330 11.545 ;
        RECT 25.130 5.895 25.330 11.545 ;
        RECT 27.130 5.895 27.330 11.545 ;
        RECT 29.130 5.895 29.330 11.545 ;
        RECT 31.130 5.895 31.330 11.545 ;
        RECT 33.130 5.895 33.330 11.545 ;
        RECT 35.130 5.895 35.330 11.545 ;
        RECT 37.130 5.895 37.330 11.545 ;
        RECT 39.130 5.895 39.330 11.545 ;
        RECT 41.130 5.895 41.330 11.545 ;
        RECT 43.130 5.895 43.330 11.545 ;
        RECT 45.130 5.895 45.330 11.545 ;
        RECT 47.130 5.895 47.330 11.545 ;
        RECT 49.130 5.895 49.330 11.545 ;
        RECT 51.130 5.895 51.330 11.545 ;
        RECT 53.130 5.895 53.330 11.545 ;
        RECT 55.130 5.895 55.330 11.545 ;
        RECT 57.130 5.895 57.330 11.545 ;
        RECT 59.130 5.895 59.330 11.545 ;
        RECT 61.130 5.895 61.330 11.545 ;
        RECT 63.130 5.895 63.330 11.545 ;
        RECT 65.130 5.895 65.330 11.545 ;
        RECT 67.130 5.895 67.330 11.545 ;
        RECT 69.130 5.895 69.330 11.545 ;
        RECT 71.130 5.895 71.330 11.545 ;
        RECT 73.130 5.895 73.330 11.545 ;
        RECT 75.130 5.895 75.330 11.545 ;
        RECT 77.130 5.895 77.330 11.545 ;
        RECT 79.130 5.895 79.330 11.545 ;
        RECT 81.130 5.895 81.330 11.545 ;
        RECT 83.130 5.895 83.330 11.545 ;
        RECT 85.130 5.895 85.330 11.545 ;
        RECT 87.130 5.895 87.330 11.545 ;
        RECT 89.130 5.895 89.330 11.545 ;
        RECT 91.130 5.895 91.330 11.545 ;
        RECT 93.130 5.895 93.330 11.545 ;
        RECT 95.130 5.895 95.330 11.545 ;
        RECT 97.130 5.895 97.330 11.545 ;
        RECT 99.130 5.895 99.330 11.545 ;
        RECT 101.130 5.895 101.330 11.545 ;
        RECT 103.130 5.895 103.330 11.545 ;
        RECT 105.130 5.895 105.330 11.545 ;
        RECT 107.130 5.895 107.330 11.545 ;
        RECT 109.130 5.895 109.330 11.545 ;
        RECT 111.130 5.895 111.330 11.545 ;
        RECT 113.130 5.895 113.330 11.545 ;
        RECT 115.130 5.895 115.330 11.545 ;
        RECT 117.130 5.895 117.330 11.545 ;
        RECT 119.130 5.895 119.330 11.545 ;
        RECT 121.130 5.895 121.330 11.545 ;
        RECT 123.130 5.895 123.330 11.545 ;
        RECT 125.130 5.895 125.330 11.545 ;
        RECT 127.130 5.895 127.330 11.545 ;
        RECT 129.130 5.895 129.330 11.545 ;
        RECT 131.130 5.895 131.330 11.545 ;
        RECT 1.130 5.695 2.000 5.895 ;
        RECT 3.130 5.695 4.000 5.895 ;
        RECT 5.130 5.695 6.000 5.895 ;
        RECT 7.130 5.695 8.000 5.895 ;
        RECT 9.130 5.695 10.000 5.895 ;
        RECT 11.130 5.695 12.000 5.895 ;
        RECT 13.130 5.695 14.000 5.895 ;
        RECT 15.130 5.695 16.000 5.895 ;
        RECT 17.130 5.695 18.000 5.895 ;
        RECT 19.130 5.695 20.000 5.895 ;
        RECT 21.130 5.695 22.000 5.895 ;
        RECT 23.130 5.695 24.000 5.895 ;
        RECT 25.130 5.695 26.000 5.895 ;
        RECT 27.130 5.695 28.000 5.895 ;
        RECT 29.130 5.695 30.000 5.895 ;
        RECT 31.130 5.695 32.000 5.895 ;
        RECT 33.130 5.695 34.000 5.895 ;
        RECT 35.130 5.695 36.000 5.895 ;
        RECT 37.130 5.695 38.000 5.895 ;
        RECT 39.130 5.695 40.000 5.895 ;
        RECT 41.130 5.695 42.000 5.895 ;
        RECT 43.130 5.695 44.000 5.895 ;
        RECT 45.130 5.695 46.000 5.895 ;
        RECT 47.130 5.695 48.000 5.895 ;
        RECT 49.130 5.695 50.000 5.895 ;
        RECT 51.130 5.695 52.000 5.895 ;
        RECT 53.130 5.695 54.000 5.895 ;
        RECT 55.130 5.695 56.000 5.895 ;
        RECT 57.130 5.695 58.000 5.895 ;
        RECT 59.130 5.695 60.000 5.895 ;
        RECT 61.130 5.695 62.000 5.895 ;
        RECT 63.130 5.695 64.000 5.895 ;
        RECT 65.130 5.695 66.000 5.895 ;
        RECT 67.130 5.695 68.000 5.895 ;
        RECT 69.130 5.695 70.000 5.895 ;
        RECT 71.130 5.695 72.000 5.895 ;
        RECT 73.130 5.695 74.000 5.895 ;
        RECT 75.130 5.695 76.000 5.895 ;
        RECT 77.130 5.695 78.000 5.895 ;
        RECT 79.130 5.695 80.000 5.895 ;
        RECT 81.130 5.695 82.000 5.895 ;
        RECT 83.130 5.695 84.000 5.895 ;
        RECT 85.130 5.695 86.000 5.895 ;
        RECT 87.130 5.695 88.000 5.895 ;
        RECT 89.130 5.695 90.000 5.895 ;
        RECT 91.130 5.695 92.000 5.895 ;
        RECT 93.130 5.695 94.000 5.895 ;
        RECT 95.130 5.695 96.000 5.895 ;
        RECT 97.130 5.695 98.000 5.895 ;
        RECT 99.130 5.695 100.000 5.895 ;
        RECT 101.130 5.695 102.000 5.895 ;
        RECT 103.130 5.695 104.000 5.895 ;
        RECT 105.130 5.695 106.000 5.895 ;
        RECT 107.130 5.695 108.000 5.895 ;
        RECT 109.130 5.695 110.000 5.895 ;
        RECT 111.130 5.695 112.000 5.895 ;
        RECT 113.130 5.695 114.000 5.895 ;
        RECT 115.130 5.695 116.000 5.895 ;
        RECT 117.130 5.695 118.000 5.895 ;
        RECT 119.130 5.695 120.000 5.895 ;
        RECT 121.130 5.695 122.000 5.895 ;
        RECT 123.130 5.695 124.000 5.895 ;
        RECT 125.130 5.695 126.000 5.895 ;
        RECT 127.130 5.695 128.000 5.895 ;
        RECT 129.130 5.695 130.000 5.895 ;
        RECT 131.130 5.695 132.000 5.895 ;
        RECT 1.800 5.055 2.000 5.695 ;
        RECT 3.800 5.055 4.000 5.695 ;
        RECT 5.800 5.055 6.000 5.695 ;
        RECT 7.800 5.055 8.000 5.695 ;
        RECT 9.800 5.055 10.000 5.695 ;
        RECT 11.800 5.055 12.000 5.695 ;
        RECT 13.800 5.055 14.000 5.695 ;
        RECT 15.800 5.055 16.000 5.695 ;
        RECT 17.800 5.055 18.000 5.695 ;
        RECT 19.800 5.055 20.000 5.695 ;
        RECT 21.800 5.055 22.000 5.695 ;
        RECT 23.800 5.055 24.000 5.695 ;
        RECT 25.800 5.055 26.000 5.695 ;
        RECT 27.800 5.055 28.000 5.695 ;
        RECT 29.800 5.055 30.000 5.695 ;
        RECT 31.800 5.055 32.000 5.695 ;
        RECT 33.800 5.055 34.000 5.695 ;
        RECT 35.800 5.055 36.000 5.695 ;
        RECT 37.800 5.055 38.000 5.695 ;
        RECT 39.800 5.055 40.000 5.695 ;
        RECT 41.800 5.055 42.000 5.695 ;
        RECT 43.800 5.055 44.000 5.695 ;
        RECT 45.800 5.055 46.000 5.695 ;
        RECT 47.800 5.055 48.000 5.695 ;
        RECT 49.800 5.055 50.000 5.695 ;
        RECT 51.800 5.055 52.000 5.695 ;
        RECT 53.800 5.055 54.000 5.695 ;
        RECT 55.800 5.055 56.000 5.695 ;
        RECT 57.800 5.055 58.000 5.695 ;
        RECT 59.800 5.055 60.000 5.695 ;
        RECT 61.800 5.055 62.000 5.695 ;
        RECT 63.800 5.055 64.000 5.695 ;
        RECT 65.800 5.055 66.000 5.695 ;
        RECT 67.800 5.055 68.000 5.695 ;
        RECT 69.800 5.055 70.000 5.695 ;
        RECT 71.800 5.055 72.000 5.695 ;
        RECT 73.800 5.055 74.000 5.695 ;
        RECT 75.800 5.055 76.000 5.695 ;
        RECT 77.800 5.055 78.000 5.695 ;
        RECT 79.800 5.055 80.000 5.695 ;
        RECT 81.800 5.055 82.000 5.695 ;
        RECT 83.800 5.055 84.000 5.695 ;
        RECT 85.800 5.055 86.000 5.695 ;
        RECT 87.800 5.055 88.000 5.695 ;
        RECT 89.800 5.055 90.000 5.695 ;
        RECT 91.800 5.055 92.000 5.695 ;
        RECT 93.800 5.055 94.000 5.695 ;
        RECT 95.800 5.055 96.000 5.695 ;
        RECT 97.800 5.055 98.000 5.695 ;
        RECT 99.800 5.055 100.000 5.695 ;
        RECT 101.800 5.055 102.000 5.695 ;
        RECT 103.800 5.055 104.000 5.695 ;
        RECT 105.800 5.055 106.000 5.695 ;
        RECT 107.800 5.055 108.000 5.695 ;
        RECT 109.800 5.055 110.000 5.695 ;
        RECT 111.800 5.055 112.000 5.695 ;
        RECT 113.800 5.055 114.000 5.695 ;
        RECT 115.800 5.055 116.000 5.695 ;
        RECT 117.800 5.055 118.000 5.695 ;
        RECT 119.800 5.055 120.000 5.695 ;
        RECT 121.800 5.055 122.000 5.695 ;
        RECT 123.800 5.055 124.000 5.695 ;
        RECT 125.800 5.055 126.000 5.695 ;
        RECT 127.800 5.055 128.000 5.695 ;
        RECT 129.800 5.055 130.000 5.695 ;
        RECT 131.800 5.055 132.000 5.695 ;
        RECT 1.755 4.765 2.045 5.055 ;
        RECT 3.755 4.765 4.045 5.055 ;
        RECT 5.755 4.765 6.045 5.055 ;
        RECT 7.755 4.765 8.045 5.055 ;
        RECT 9.755 4.765 10.045 5.055 ;
        RECT 11.755 4.765 12.045 5.055 ;
        RECT 13.755 4.765 14.045 5.055 ;
        RECT 15.755 4.765 16.045 5.055 ;
        RECT 17.755 4.765 18.045 5.055 ;
        RECT 19.755 4.765 20.045 5.055 ;
        RECT 21.755 4.765 22.045 5.055 ;
        RECT 23.755 4.765 24.045 5.055 ;
        RECT 25.755 4.765 26.045 5.055 ;
        RECT 27.755 4.765 28.045 5.055 ;
        RECT 29.755 4.765 30.045 5.055 ;
        RECT 31.755 4.765 32.045 5.055 ;
        RECT 33.755 4.765 34.045 5.055 ;
        RECT 35.755 4.765 36.045 5.055 ;
        RECT 37.755 4.765 38.045 5.055 ;
        RECT 39.755 4.765 40.045 5.055 ;
        RECT 41.755 4.765 42.045 5.055 ;
        RECT 43.755 4.765 44.045 5.055 ;
        RECT 45.755 4.765 46.045 5.055 ;
        RECT 47.755 4.765 48.045 5.055 ;
        RECT 49.755 4.765 50.045 5.055 ;
        RECT 51.755 4.765 52.045 5.055 ;
        RECT 53.755 4.765 54.045 5.055 ;
        RECT 55.755 4.765 56.045 5.055 ;
        RECT 57.755 4.765 58.045 5.055 ;
        RECT 59.755 4.765 60.045 5.055 ;
        RECT 61.755 4.765 62.045 5.055 ;
        RECT 63.755 4.765 64.045 5.055 ;
        RECT 65.755 4.765 66.045 5.055 ;
        RECT 67.755 4.765 68.045 5.055 ;
        RECT 69.755 4.765 70.045 5.055 ;
        RECT 71.755 4.765 72.045 5.055 ;
        RECT 73.755 4.765 74.045 5.055 ;
        RECT 75.755 4.765 76.045 5.055 ;
        RECT 77.755 4.765 78.045 5.055 ;
        RECT 79.755 4.765 80.045 5.055 ;
        RECT 81.755 4.765 82.045 5.055 ;
        RECT 83.755 4.765 84.045 5.055 ;
        RECT 85.755 4.765 86.045 5.055 ;
        RECT 87.755 4.765 88.045 5.055 ;
        RECT 89.755 4.765 90.045 5.055 ;
        RECT 91.755 4.765 92.045 5.055 ;
        RECT 93.755 4.765 94.045 5.055 ;
        RECT 95.755 4.765 96.045 5.055 ;
        RECT 97.755 4.765 98.045 5.055 ;
        RECT 99.755 4.765 100.045 5.055 ;
        RECT 101.755 4.765 102.045 5.055 ;
        RECT 103.755 4.765 104.045 5.055 ;
        RECT 105.755 4.765 106.045 5.055 ;
        RECT 107.755 4.765 108.045 5.055 ;
        RECT 109.755 4.765 110.045 5.055 ;
        RECT 111.755 4.765 112.045 5.055 ;
        RECT 113.755 4.765 114.045 5.055 ;
        RECT 115.755 4.765 116.045 5.055 ;
        RECT 117.755 4.765 118.045 5.055 ;
        RECT 119.755 4.765 120.045 5.055 ;
        RECT 121.755 4.765 122.045 5.055 ;
        RECT 123.755 4.765 124.045 5.055 ;
        RECT 125.755 4.765 126.045 5.055 ;
        RECT 127.755 4.765 128.045 5.055 ;
        RECT 129.755 4.765 130.045 5.055 ;
        RECT 131.755 4.765 132.045 5.055 ;
        RECT 1.415 4.465 1.705 4.555 ;
        RECT 1.055 4.265 1.705 4.465 ;
        RECT 2.095 4.465 2.385 4.555 ;
        RECT 3.415 4.465 3.705 4.555 ;
        RECT 2.095 4.265 2.740 4.465 ;
        RECT 1.055 3.200 1.255 4.265 ;
        RECT 2.540 3.200 2.740 4.265 ;
        RECT 3.055 4.265 3.705 4.465 ;
        RECT 4.095 4.465 4.385 4.555 ;
        RECT 5.415 4.465 5.705 4.555 ;
        RECT 4.095 4.265 4.740 4.465 ;
        RECT 3.055 3.200 3.255 4.265 ;
        RECT 4.540 3.200 4.740 4.265 ;
        RECT 5.055 4.265 5.705 4.465 ;
        RECT 6.095 4.465 6.385 4.555 ;
        RECT 7.415 4.465 7.705 4.555 ;
        RECT 6.095 4.265 6.740 4.465 ;
        RECT 5.055 3.200 5.255 4.265 ;
        RECT 6.540 3.200 6.740 4.265 ;
        RECT 7.055 4.265 7.705 4.465 ;
        RECT 8.095 4.465 8.385 4.555 ;
        RECT 9.415 4.465 9.705 4.555 ;
        RECT 8.095 4.265 8.740 4.465 ;
        RECT 7.055 3.200 7.255 4.265 ;
        RECT 8.540 3.200 8.740 4.265 ;
        RECT 9.055 4.265 9.705 4.465 ;
        RECT 10.095 4.465 10.385 4.555 ;
        RECT 11.415 4.465 11.705 4.555 ;
        RECT 10.095 4.265 10.740 4.465 ;
        RECT 9.055 3.200 9.255 4.265 ;
        RECT 10.540 3.200 10.740 4.265 ;
        RECT 11.055 4.265 11.705 4.465 ;
        RECT 12.095 4.465 12.385 4.555 ;
        RECT 13.415 4.465 13.705 4.555 ;
        RECT 12.095 4.265 12.740 4.465 ;
        RECT 11.055 3.200 11.255 4.265 ;
        RECT 12.540 3.200 12.740 4.265 ;
        RECT 13.055 4.265 13.705 4.465 ;
        RECT 14.095 4.465 14.385 4.555 ;
        RECT 15.415 4.465 15.705 4.555 ;
        RECT 14.095 4.265 14.740 4.465 ;
        RECT 13.055 3.200 13.255 4.265 ;
        RECT 14.540 3.200 14.740 4.265 ;
        RECT 15.055 4.265 15.705 4.465 ;
        RECT 16.095 4.465 16.385 4.555 ;
        RECT 17.415 4.465 17.705 4.555 ;
        RECT 16.095 4.265 16.740 4.465 ;
        RECT 15.055 3.200 15.255 4.265 ;
        RECT 16.540 3.200 16.740 4.265 ;
        RECT 17.055 4.265 17.705 4.465 ;
        RECT 18.095 4.465 18.385 4.555 ;
        RECT 19.415 4.465 19.705 4.555 ;
        RECT 18.095 4.265 18.740 4.465 ;
        RECT 17.055 3.200 17.255 4.265 ;
        RECT 18.540 3.200 18.740 4.265 ;
        RECT 19.055 4.265 19.705 4.465 ;
        RECT 20.095 4.465 20.385 4.555 ;
        RECT 21.415 4.465 21.705 4.555 ;
        RECT 20.095 4.265 20.740 4.465 ;
        RECT 19.055 3.200 19.255 4.265 ;
        RECT 20.540 3.200 20.740 4.265 ;
        RECT 21.055 4.265 21.705 4.465 ;
        RECT 22.095 4.465 22.385 4.555 ;
        RECT 23.415 4.465 23.705 4.555 ;
        RECT 22.095 4.265 22.740 4.465 ;
        RECT 21.055 3.200 21.255 4.265 ;
        RECT 22.540 3.200 22.740 4.265 ;
        RECT 23.055 4.265 23.705 4.465 ;
        RECT 24.095 4.465 24.385 4.555 ;
        RECT 25.415 4.465 25.705 4.555 ;
        RECT 24.095 4.265 24.740 4.465 ;
        RECT 23.055 3.200 23.255 4.265 ;
        RECT 24.540 3.200 24.740 4.265 ;
        RECT 25.055 4.265 25.705 4.465 ;
        RECT 26.095 4.465 26.385 4.555 ;
        RECT 27.415 4.465 27.705 4.555 ;
        RECT 26.095 4.265 26.740 4.465 ;
        RECT 25.055 3.200 25.255 4.265 ;
        RECT 26.540 3.200 26.740 4.265 ;
        RECT 27.055 4.265 27.705 4.465 ;
        RECT 28.095 4.465 28.385 4.555 ;
        RECT 29.415 4.465 29.705 4.555 ;
        RECT 28.095 4.265 28.740 4.465 ;
        RECT 27.055 3.200 27.255 4.265 ;
        RECT 28.540 3.200 28.740 4.265 ;
        RECT 29.055 4.265 29.705 4.465 ;
        RECT 30.095 4.465 30.385 4.555 ;
        RECT 31.415 4.465 31.705 4.555 ;
        RECT 30.095 4.265 30.740 4.465 ;
        RECT 29.055 3.200 29.255 4.265 ;
        RECT 30.540 3.200 30.740 4.265 ;
        RECT 31.055 4.265 31.705 4.465 ;
        RECT 32.095 4.465 32.385 4.555 ;
        RECT 33.415 4.465 33.705 4.555 ;
        RECT 32.095 4.265 32.740 4.465 ;
        RECT 31.055 3.200 31.255 4.265 ;
        RECT 32.540 3.200 32.740 4.265 ;
        RECT 33.055 4.265 33.705 4.465 ;
        RECT 34.095 4.465 34.385 4.555 ;
        RECT 35.415 4.465 35.705 4.555 ;
        RECT 34.095 4.265 34.740 4.465 ;
        RECT 33.055 3.200 33.255 4.265 ;
        RECT 34.540 3.200 34.740 4.265 ;
        RECT 35.055 4.265 35.705 4.465 ;
        RECT 36.095 4.465 36.385 4.555 ;
        RECT 37.415 4.465 37.705 4.555 ;
        RECT 36.095 4.265 36.740 4.465 ;
        RECT 35.055 3.200 35.255 4.265 ;
        RECT 36.540 3.200 36.740 4.265 ;
        RECT 37.055 4.265 37.705 4.465 ;
        RECT 38.095 4.465 38.385 4.555 ;
        RECT 39.415 4.465 39.705 4.555 ;
        RECT 38.095 4.265 38.740 4.465 ;
        RECT 37.055 3.200 37.255 4.265 ;
        RECT 38.540 3.200 38.740 4.265 ;
        RECT 39.055 4.265 39.705 4.465 ;
        RECT 40.095 4.465 40.385 4.555 ;
        RECT 41.415 4.465 41.705 4.555 ;
        RECT 40.095 4.265 40.740 4.465 ;
        RECT 39.055 3.200 39.255 4.265 ;
        RECT 40.540 3.200 40.740 4.265 ;
        RECT 41.055 4.265 41.705 4.465 ;
        RECT 42.095 4.465 42.385 4.555 ;
        RECT 43.415 4.465 43.705 4.555 ;
        RECT 42.095 4.265 42.740 4.465 ;
        RECT 41.055 3.200 41.255 4.265 ;
        RECT 42.540 3.200 42.740 4.265 ;
        RECT 43.055 4.265 43.705 4.465 ;
        RECT 44.095 4.465 44.385 4.555 ;
        RECT 45.415 4.465 45.705 4.555 ;
        RECT 44.095 4.265 44.740 4.465 ;
        RECT 43.055 3.200 43.255 4.265 ;
        RECT 44.540 3.200 44.740 4.265 ;
        RECT 45.055 4.265 45.705 4.465 ;
        RECT 46.095 4.465 46.385 4.555 ;
        RECT 47.415 4.465 47.705 4.555 ;
        RECT 46.095 4.265 46.740 4.465 ;
        RECT 45.055 3.200 45.255 4.265 ;
        RECT 46.540 3.200 46.740 4.265 ;
        RECT 47.055 4.265 47.705 4.465 ;
        RECT 48.095 4.465 48.385 4.555 ;
        RECT 49.415 4.465 49.705 4.555 ;
        RECT 48.095 4.265 48.740 4.465 ;
        RECT 47.055 3.200 47.255 4.265 ;
        RECT 48.540 3.200 48.740 4.265 ;
        RECT 49.055 4.265 49.705 4.465 ;
        RECT 50.095 4.465 50.385 4.555 ;
        RECT 51.415 4.465 51.705 4.555 ;
        RECT 50.095 4.265 50.740 4.465 ;
        RECT 49.055 3.200 49.255 4.265 ;
        RECT 50.540 3.200 50.740 4.265 ;
        RECT 51.055 4.265 51.705 4.465 ;
        RECT 52.095 4.465 52.385 4.555 ;
        RECT 53.415 4.465 53.705 4.555 ;
        RECT 52.095 4.265 52.740 4.465 ;
        RECT 51.055 3.200 51.255 4.265 ;
        RECT 52.540 3.200 52.740 4.265 ;
        RECT 53.055 4.265 53.705 4.465 ;
        RECT 54.095 4.465 54.385 4.555 ;
        RECT 55.415 4.465 55.705 4.555 ;
        RECT 54.095 4.265 54.740 4.465 ;
        RECT 53.055 3.200 53.255 4.265 ;
        RECT 54.540 3.200 54.740 4.265 ;
        RECT 55.055 4.265 55.705 4.465 ;
        RECT 56.095 4.465 56.385 4.555 ;
        RECT 57.415 4.465 57.705 4.555 ;
        RECT 56.095 4.265 56.740 4.465 ;
        RECT 55.055 3.200 55.255 4.265 ;
        RECT 56.540 3.200 56.740 4.265 ;
        RECT 57.055 4.265 57.705 4.465 ;
        RECT 58.095 4.465 58.385 4.555 ;
        RECT 59.415 4.465 59.705 4.555 ;
        RECT 58.095 4.265 58.740 4.465 ;
        RECT 57.055 3.200 57.255 4.265 ;
        RECT 58.540 3.200 58.740 4.265 ;
        RECT 59.055 4.265 59.705 4.465 ;
        RECT 60.095 4.465 60.385 4.555 ;
        RECT 61.415 4.465 61.705 4.555 ;
        RECT 60.095 4.265 60.740 4.465 ;
        RECT 59.055 3.200 59.255 4.265 ;
        RECT 60.540 3.200 60.740 4.265 ;
        RECT 61.055 4.265 61.705 4.465 ;
        RECT 62.095 4.465 62.385 4.555 ;
        RECT 63.415 4.465 63.705 4.555 ;
        RECT 62.095 4.265 62.740 4.465 ;
        RECT 61.055 3.200 61.255 4.265 ;
        RECT 62.540 3.200 62.740 4.265 ;
        RECT 63.055 4.265 63.705 4.465 ;
        RECT 64.095 4.465 64.385 4.555 ;
        RECT 65.415 4.465 65.705 4.555 ;
        RECT 64.095 4.265 64.740 4.465 ;
        RECT 63.055 3.200 63.255 4.265 ;
        RECT 64.540 3.200 64.740 4.265 ;
        RECT 65.055 4.265 65.705 4.465 ;
        RECT 66.095 4.465 66.385 4.555 ;
        RECT 67.415 4.465 67.705 4.555 ;
        RECT 66.095 4.265 66.740 4.465 ;
        RECT 65.055 3.200 65.255 4.265 ;
        RECT 66.540 3.200 66.740 4.265 ;
        RECT 67.055 4.265 67.705 4.465 ;
        RECT 68.095 4.465 68.385 4.555 ;
        RECT 69.415 4.465 69.705 4.555 ;
        RECT 68.095 4.265 68.740 4.465 ;
        RECT 67.055 3.200 67.255 4.265 ;
        RECT 68.540 3.200 68.740 4.265 ;
        RECT 69.055 4.265 69.705 4.465 ;
        RECT 70.095 4.465 70.385 4.555 ;
        RECT 71.415 4.465 71.705 4.555 ;
        RECT 70.095 4.265 70.740 4.465 ;
        RECT 69.055 3.200 69.255 4.265 ;
        RECT 70.540 3.200 70.740 4.265 ;
        RECT 71.055 4.265 71.705 4.465 ;
        RECT 72.095 4.465 72.385 4.555 ;
        RECT 73.415 4.465 73.705 4.555 ;
        RECT 72.095 4.265 72.740 4.465 ;
        RECT 71.055 3.200 71.255 4.265 ;
        RECT 72.540 3.200 72.740 4.265 ;
        RECT 73.055 4.265 73.705 4.465 ;
        RECT 74.095 4.465 74.385 4.555 ;
        RECT 75.415 4.465 75.705 4.555 ;
        RECT 74.095 4.265 74.740 4.465 ;
        RECT 73.055 3.200 73.255 4.265 ;
        RECT 74.540 3.200 74.740 4.265 ;
        RECT 75.055 4.265 75.705 4.465 ;
        RECT 76.095 4.465 76.385 4.555 ;
        RECT 77.415 4.465 77.705 4.555 ;
        RECT 76.095 4.265 76.740 4.465 ;
        RECT 75.055 3.200 75.255 4.265 ;
        RECT 76.540 3.200 76.740 4.265 ;
        RECT 77.055 4.265 77.705 4.465 ;
        RECT 78.095 4.465 78.385 4.555 ;
        RECT 79.415 4.465 79.705 4.555 ;
        RECT 78.095 4.265 78.740 4.465 ;
        RECT 77.055 3.200 77.255 4.265 ;
        RECT 78.540 3.200 78.740 4.265 ;
        RECT 79.055 4.265 79.705 4.465 ;
        RECT 80.095 4.465 80.385 4.555 ;
        RECT 81.415 4.465 81.705 4.555 ;
        RECT 80.095 4.265 80.740 4.465 ;
        RECT 79.055 3.200 79.255 4.265 ;
        RECT 80.540 3.200 80.740 4.265 ;
        RECT 81.055 4.265 81.705 4.465 ;
        RECT 82.095 4.465 82.385 4.555 ;
        RECT 83.415 4.465 83.705 4.555 ;
        RECT 82.095 4.265 82.740 4.465 ;
        RECT 81.055 3.200 81.255 4.265 ;
        RECT 82.540 3.200 82.740 4.265 ;
        RECT 83.055 4.265 83.705 4.465 ;
        RECT 84.095 4.465 84.385 4.555 ;
        RECT 85.415 4.465 85.705 4.555 ;
        RECT 84.095 4.265 84.740 4.465 ;
        RECT 83.055 3.200 83.255 4.265 ;
        RECT 84.540 3.200 84.740 4.265 ;
        RECT 85.055 4.265 85.705 4.465 ;
        RECT 86.095 4.465 86.385 4.555 ;
        RECT 87.415 4.465 87.705 4.555 ;
        RECT 86.095 4.265 86.740 4.465 ;
        RECT 85.055 3.200 85.255 4.265 ;
        RECT 86.540 3.200 86.740 4.265 ;
        RECT 87.055 4.265 87.705 4.465 ;
        RECT 88.095 4.465 88.385 4.555 ;
        RECT 89.415 4.465 89.705 4.555 ;
        RECT 88.095 4.265 88.740 4.465 ;
        RECT 87.055 3.200 87.255 4.265 ;
        RECT 88.540 3.200 88.740 4.265 ;
        RECT 89.055 4.265 89.705 4.465 ;
        RECT 90.095 4.465 90.385 4.555 ;
        RECT 91.415 4.465 91.705 4.555 ;
        RECT 90.095 4.265 90.740 4.465 ;
        RECT 89.055 3.200 89.255 4.265 ;
        RECT 90.540 3.200 90.740 4.265 ;
        RECT 91.055 4.265 91.705 4.465 ;
        RECT 92.095 4.465 92.385 4.555 ;
        RECT 93.415 4.465 93.705 4.555 ;
        RECT 92.095 4.265 92.740 4.465 ;
        RECT 91.055 3.200 91.255 4.265 ;
        RECT 92.540 3.200 92.740 4.265 ;
        RECT 93.055 4.265 93.705 4.465 ;
        RECT 94.095 4.465 94.385 4.555 ;
        RECT 95.415 4.465 95.705 4.555 ;
        RECT 94.095 4.265 94.740 4.465 ;
        RECT 93.055 3.200 93.255 4.265 ;
        RECT 94.540 3.200 94.740 4.265 ;
        RECT 95.055 4.265 95.705 4.465 ;
        RECT 96.095 4.465 96.385 4.555 ;
        RECT 97.415 4.465 97.705 4.555 ;
        RECT 96.095 4.265 96.740 4.465 ;
        RECT 95.055 3.200 95.255 4.265 ;
        RECT 96.540 3.200 96.740 4.265 ;
        RECT 97.055 4.265 97.705 4.465 ;
        RECT 98.095 4.465 98.385 4.555 ;
        RECT 99.415 4.465 99.705 4.555 ;
        RECT 98.095 4.265 98.740 4.465 ;
        RECT 97.055 3.200 97.255 4.265 ;
        RECT 98.540 3.200 98.740 4.265 ;
        RECT 99.055 4.265 99.705 4.465 ;
        RECT 100.095 4.465 100.385 4.555 ;
        RECT 101.415 4.465 101.705 4.555 ;
        RECT 100.095 4.265 100.740 4.465 ;
        RECT 99.055 3.200 99.255 4.265 ;
        RECT 100.540 3.200 100.740 4.265 ;
        RECT 101.055 4.265 101.705 4.465 ;
        RECT 102.095 4.465 102.385 4.555 ;
        RECT 103.415 4.465 103.705 4.555 ;
        RECT 102.095 4.265 102.740 4.465 ;
        RECT 101.055 3.200 101.255 4.265 ;
        RECT 102.540 3.200 102.740 4.265 ;
        RECT 103.055 4.265 103.705 4.465 ;
        RECT 104.095 4.465 104.385 4.555 ;
        RECT 105.415 4.465 105.705 4.555 ;
        RECT 104.095 4.265 104.740 4.465 ;
        RECT 103.055 3.200 103.255 4.265 ;
        RECT 104.540 3.200 104.740 4.265 ;
        RECT 105.055 4.265 105.705 4.465 ;
        RECT 106.095 4.465 106.385 4.555 ;
        RECT 107.415 4.465 107.705 4.555 ;
        RECT 106.095 4.265 106.740 4.465 ;
        RECT 105.055 3.200 105.255 4.265 ;
        RECT 106.540 3.200 106.740 4.265 ;
        RECT 107.055 4.265 107.705 4.465 ;
        RECT 108.095 4.465 108.385 4.555 ;
        RECT 109.415 4.465 109.705 4.555 ;
        RECT 108.095 4.265 108.740 4.465 ;
        RECT 107.055 3.200 107.255 4.265 ;
        RECT 108.540 3.200 108.740 4.265 ;
        RECT 109.055 4.265 109.705 4.465 ;
        RECT 110.095 4.465 110.385 4.555 ;
        RECT 111.415 4.465 111.705 4.555 ;
        RECT 110.095 4.265 110.740 4.465 ;
        RECT 109.055 3.200 109.255 4.265 ;
        RECT 110.540 3.200 110.740 4.265 ;
        RECT 111.055 4.265 111.705 4.465 ;
        RECT 112.095 4.465 112.385 4.555 ;
        RECT 113.415 4.465 113.705 4.555 ;
        RECT 112.095 4.265 112.740 4.465 ;
        RECT 111.055 3.200 111.255 4.265 ;
        RECT 112.540 3.200 112.740 4.265 ;
        RECT 113.055 4.265 113.705 4.465 ;
        RECT 114.095 4.465 114.385 4.555 ;
        RECT 115.415 4.465 115.705 4.555 ;
        RECT 114.095 4.265 114.740 4.465 ;
        RECT 113.055 3.200 113.255 4.265 ;
        RECT 114.540 3.200 114.740 4.265 ;
        RECT 115.055 4.265 115.705 4.465 ;
        RECT 116.095 4.465 116.385 4.555 ;
        RECT 117.415 4.465 117.705 4.555 ;
        RECT 116.095 4.265 116.740 4.465 ;
        RECT 115.055 3.200 115.255 4.265 ;
        RECT 116.540 3.200 116.740 4.265 ;
        RECT 117.055 4.265 117.705 4.465 ;
        RECT 118.095 4.465 118.385 4.555 ;
        RECT 119.415 4.465 119.705 4.555 ;
        RECT 118.095 4.265 118.740 4.465 ;
        RECT 117.055 3.200 117.255 4.265 ;
        RECT 118.540 3.200 118.740 4.265 ;
        RECT 119.055 4.265 119.705 4.465 ;
        RECT 120.095 4.465 120.385 4.555 ;
        RECT 121.415 4.465 121.705 4.555 ;
        RECT 120.095 4.265 120.740 4.465 ;
        RECT 119.055 3.200 119.255 4.265 ;
        RECT 120.540 3.200 120.740 4.265 ;
        RECT 121.055 4.265 121.705 4.465 ;
        RECT 122.095 4.465 122.385 4.555 ;
        RECT 123.415 4.465 123.705 4.555 ;
        RECT 122.095 4.265 122.740 4.465 ;
        RECT 121.055 3.200 121.255 4.265 ;
        RECT 122.540 3.200 122.740 4.265 ;
        RECT 123.055 4.265 123.705 4.465 ;
        RECT 124.095 4.465 124.385 4.555 ;
        RECT 125.415 4.465 125.705 4.555 ;
        RECT 124.095 4.265 124.740 4.465 ;
        RECT 123.055 3.200 123.255 4.265 ;
        RECT 124.540 3.200 124.740 4.265 ;
        RECT 125.055 4.265 125.705 4.465 ;
        RECT 126.095 4.465 126.385 4.555 ;
        RECT 127.415 4.465 127.705 4.555 ;
        RECT 126.095 4.265 126.740 4.465 ;
        RECT 125.055 3.200 125.255 4.265 ;
        RECT 126.540 3.200 126.740 4.265 ;
        RECT 127.055 4.265 127.705 4.465 ;
        RECT 128.095 4.465 128.385 4.555 ;
        RECT 129.415 4.465 129.705 4.555 ;
        RECT 128.095 4.265 128.740 4.465 ;
        RECT 127.055 3.200 127.255 4.265 ;
        RECT 128.540 3.200 128.740 4.265 ;
        RECT 129.055 4.265 129.705 4.465 ;
        RECT 130.095 4.465 130.385 4.555 ;
        RECT 131.415 4.465 131.705 4.555 ;
        RECT 130.095 4.265 130.740 4.465 ;
        RECT 129.055 3.200 129.255 4.265 ;
        RECT 130.540 3.200 130.740 4.265 ;
        RECT 131.055 4.265 131.705 4.465 ;
        RECT 132.095 4.465 132.385 4.555 ;
        RECT 132.095 4.265 132.740 4.465 ;
        RECT 131.055 3.200 131.255 4.265 ;
        RECT 132.540 3.200 132.740 4.265 ;
        RECT 1.010 2.910 1.300 3.200 ;
        RECT 2.500 2.910 2.790 3.200 ;
        RECT 3.010 2.910 3.300 3.200 ;
        RECT 4.500 2.910 4.790 3.200 ;
        RECT 5.010 2.910 5.300 3.200 ;
        RECT 6.500 2.910 6.790 3.200 ;
        RECT 7.010 2.910 7.300 3.200 ;
        RECT 8.500 2.910 8.790 3.200 ;
        RECT 9.010 2.910 9.300 3.200 ;
        RECT 10.500 2.910 10.790 3.200 ;
        RECT 11.010 2.910 11.300 3.200 ;
        RECT 12.500 2.910 12.790 3.200 ;
        RECT 13.010 2.910 13.300 3.200 ;
        RECT 14.500 2.910 14.790 3.200 ;
        RECT 15.010 2.910 15.300 3.200 ;
        RECT 16.500 2.910 16.790 3.200 ;
        RECT 17.010 2.910 17.300 3.200 ;
        RECT 18.500 2.910 18.790 3.200 ;
        RECT 19.010 2.910 19.300 3.200 ;
        RECT 20.500 2.910 20.790 3.200 ;
        RECT 21.010 2.910 21.300 3.200 ;
        RECT 22.500 2.910 22.790 3.200 ;
        RECT 23.010 2.910 23.300 3.200 ;
        RECT 24.500 2.910 24.790 3.200 ;
        RECT 25.010 2.910 25.300 3.200 ;
        RECT 26.500 2.910 26.790 3.200 ;
        RECT 27.010 2.910 27.300 3.200 ;
        RECT 28.500 2.910 28.790 3.200 ;
        RECT 29.010 2.910 29.300 3.200 ;
        RECT 30.500 2.910 30.790 3.200 ;
        RECT 31.010 2.910 31.300 3.200 ;
        RECT 32.500 2.910 32.790 3.200 ;
        RECT 33.010 2.910 33.300 3.200 ;
        RECT 34.500 2.910 34.790 3.200 ;
        RECT 35.010 2.910 35.300 3.200 ;
        RECT 36.500 2.910 36.790 3.200 ;
        RECT 37.010 2.910 37.300 3.200 ;
        RECT 38.500 2.910 38.790 3.200 ;
        RECT 39.010 2.910 39.300 3.200 ;
        RECT 40.500 2.910 40.790 3.200 ;
        RECT 41.010 2.910 41.300 3.200 ;
        RECT 42.500 2.910 42.790 3.200 ;
        RECT 43.010 2.910 43.300 3.200 ;
        RECT 44.500 2.910 44.790 3.200 ;
        RECT 45.010 2.910 45.300 3.200 ;
        RECT 46.500 2.910 46.790 3.200 ;
        RECT 47.010 2.910 47.300 3.200 ;
        RECT 48.500 2.910 48.790 3.200 ;
        RECT 49.010 2.910 49.300 3.200 ;
        RECT 50.500 2.910 50.790 3.200 ;
        RECT 51.010 2.910 51.300 3.200 ;
        RECT 52.500 2.910 52.790 3.200 ;
        RECT 53.010 2.910 53.300 3.200 ;
        RECT 54.500 2.910 54.790 3.200 ;
        RECT 55.010 2.910 55.300 3.200 ;
        RECT 56.500 2.910 56.790 3.200 ;
        RECT 57.010 2.910 57.300 3.200 ;
        RECT 58.500 2.910 58.790 3.200 ;
        RECT 59.010 2.910 59.300 3.200 ;
        RECT 60.500 2.910 60.790 3.200 ;
        RECT 61.010 2.910 61.300 3.200 ;
        RECT 62.500 2.910 62.790 3.200 ;
        RECT 63.010 2.910 63.300 3.200 ;
        RECT 64.500 2.910 64.790 3.200 ;
        RECT 65.010 2.910 65.300 3.200 ;
        RECT 66.500 2.910 66.790 3.200 ;
        RECT 67.010 2.910 67.300 3.200 ;
        RECT 68.500 2.910 68.790 3.200 ;
        RECT 69.010 2.910 69.300 3.200 ;
        RECT 70.500 2.910 70.790 3.200 ;
        RECT 71.010 2.910 71.300 3.200 ;
        RECT 72.500 2.910 72.790 3.200 ;
        RECT 73.010 2.910 73.300 3.200 ;
        RECT 74.500 2.910 74.790 3.200 ;
        RECT 75.010 2.910 75.300 3.200 ;
        RECT 76.500 2.910 76.790 3.200 ;
        RECT 77.010 2.910 77.300 3.200 ;
        RECT 78.500 2.910 78.790 3.200 ;
        RECT 79.010 2.910 79.300 3.200 ;
        RECT 80.500 2.910 80.790 3.200 ;
        RECT 81.010 2.910 81.300 3.200 ;
        RECT 82.500 2.910 82.790 3.200 ;
        RECT 83.010 2.910 83.300 3.200 ;
        RECT 84.500 2.910 84.790 3.200 ;
        RECT 85.010 2.910 85.300 3.200 ;
        RECT 86.500 2.910 86.790 3.200 ;
        RECT 87.010 2.910 87.300 3.200 ;
        RECT 88.500 2.910 88.790 3.200 ;
        RECT 89.010 2.910 89.300 3.200 ;
        RECT 90.500 2.910 90.790 3.200 ;
        RECT 91.010 2.910 91.300 3.200 ;
        RECT 92.500 2.910 92.790 3.200 ;
        RECT 93.010 2.910 93.300 3.200 ;
        RECT 94.500 2.910 94.790 3.200 ;
        RECT 95.010 2.910 95.300 3.200 ;
        RECT 96.500 2.910 96.790 3.200 ;
        RECT 97.010 2.910 97.300 3.200 ;
        RECT 98.500 2.910 98.790 3.200 ;
        RECT 99.010 2.910 99.300 3.200 ;
        RECT 100.500 2.910 100.790 3.200 ;
        RECT 101.010 2.910 101.300 3.200 ;
        RECT 102.500 2.910 102.790 3.200 ;
        RECT 103.010 2.910 103.300 3.200 ;
        RECT 104.500 2.910 104.790 3.200 ;
        RECT 105.010 2.910 105.300 3.200 ;
        RECT 106.500 2.910 106.790 3.200 ;
        RECT 107.010 2.910 107.300 3.200 ;
        RECT 108.500 2.910 108.790 3.200 ;
        RECT 109.010 2.910 109.300 3.200 ;
        RECT 110.500 2.910 110.790 3.200 ;
        RECT 111.010 2.910 111.300 3.200 ;
        RECT 112.500 2.910 112.790 3.200 ;
        RECT 113.010 2.910 113.300 3.200 ;
        RECT 114.500 2.910 114.790 3.200 ;
        RECT 115.010 2.910 115.300 3.200 ;
        RECT 116.500 2.910 116.790 3.200 ;
        RECT 117.010 2.910 117.300 3.200 ;
        RECT 118.500 2.910 118.790 3.200 ;
        RECT 119.010 2.910 119.300 3.200 ;
        RECT 120.500 2.910 120.790 3.200 ;
        RECT 121.010 2.910 121.300 3.200 ;
        RECT 122.500 2.910 122.790 3.200 ;
        RECT 123.010 2.910 123.300 3.200 ;
        RECT 124.500 2.910 124.790 3.200 ;
        RECT 125.010 2.910 125.300 3.200 ;
        RECT 126.500 2.910 126.790 3.200 ;
        RECT 127.010 2.910 127.300 3.200 ;
        RECT 128.500 2.910 128.790 3.200 ;
        RECT 129.010 2.910 129.300 3.200 ;
        RECT 130.500 2.910 130.790 3.200 ;
        RECT 131.010 2.910 131.300 3.200 ;
        RECT 132.500 2.910 132.790 3.200 ;
  END
END DAC2U128OUT4IN
END LIBRARY

