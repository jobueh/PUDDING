VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dac128module
  CLASS BLOCK ;
  FOREIGN dac128module ;
  ORIGIN 0.000 0.070 ;
  SIZE 133.800 BY 26.330 ;
  PIN VbiasP[1]
    ANTENNAGATEAREA 478.500000 ;
    ANTENNADIFFAREA 5.010000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 14.950 132.900 19.880 ;
    END
  END VbiasP[1]
  PIN Iout
    ANTENNADIFFAREA 66.047997 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 12.745 133.800 13.445 ;
    END
  END Iout
  PIN VbiasP[0]
    ANTENNAGATEAREA 478.500000 ;
    ANTENNADIFFAREA 5.010000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.900 6.310 132.900 11.240 ;
    END
  END VbiasP[0]
  PIN ON[64]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 130.030 23.715 130.320 26.190 ;
    END
  END ON[64]
  PIN ONB[64]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 129.480 23.715 129.770 26.190 ;
    END
  END ONB[64]
  PIN ON[65]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 128.030 23.715 128.320 26.190 ;
    END
  END ON[65]
  PIN ONB[65]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 127.480 23.715 127.770 26.190 ;
    END
  END ONB[65]
  PIN ON[66]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 126.030 23.715 126.320 26.190 ;
    END
  END ON[66]
  PIN ONB[66]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 125.480 23.715 125.770 26.190 ;
    END
  END ONB[66]
  PIN ON[67]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 124.030 23.715 124.320 26.190 ;
    END
  END ON[67]
  PIN ONB[67]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 123.480 23.715 123.770 26.190 ;
    END
  END ONB[67]
  PIN ON[68]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 122.030 23.715 122.320 26.190 ;
    END
  END ON[68]
  PIN ONB[68]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 121.480 23.715 121.770 26.190 ;
    END
  END ONB[68]
  PIN ON[69]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 120.030 23.715 120.320 26.190 ;
    END
  END ON[69]
  PIN ONB[69]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 119.480 23.715 119.770 26.190 ;
    END
  END ONB[69]
  PIN ON[70]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.030 23.715 118.320 26.190 ;
    END
  END ON[70]
  PIN ONB[70]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.480 23.715 117.770 26.190 ;
    END
  END ONB[70]
  PIN ON[71]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 116.030 23.715 116.320 26.190 ;
    END
  END ON[71]
  PIN ONB[71]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 115.480 23.715 115.770 26.190 ;
    END
  END ONB[71]
  PIN ON[72]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 114.030 23.715 114.320 26.190 ;
    END
  END ON[72]
  PIN ONB[72]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 113.480 23.715 113.770 26.190 ;
    END
  END ONB[72]
  PIN EN[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 132.030 23.715 132.320 26.190 ;
    END
  END EN[2]
  PIN ENB[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 131.480 23.715 131.770 26.190 ;
    END
  END ENB[2]
  PIN ON[73]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 112.030 23.715 112.320 26.190 ;
    END
  END ON[73]
  PIN ONB[73]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 111.480 23.715 111.770 26.190 ;
    END
  END ONB[73]
  PIN ON[74]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.030 23.715 110.320 26.190 ;
    END
  END ON[74]
  PIN ONB[74]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 109.480 23.715 109.770 26.190 ;
    END
  END ONB[74]
  PIN ON[75]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 108.030 23.715 108.320 26.190 ;
    END
  END ON[75]
  PIN ONB[75]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 107.480 23.715 107.770 26.190 ;
    END
  END ONB[75]
  PIN ON[76]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 106.030 23.715 106.320 26.190 ;
    END
  END ON[76]
  PIN ONB[76]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 105.480 23.715 105.770 26.190 ;
    END
  END ONB[76]
  PIN ON[77]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 104.030 23.715 104.320 26.190 ;
    END
  END ON[77]
  PIN ONB[77]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 103.480 23.715 103.770 26.190 ;
    END
  END ONB[77]
  PIN ON[78]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 102.030 23.715 102.320 26.190 ;
    END
  END ON[78]
  PIN ONB[78]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 101.480 23.715 101.770 26.190 ;
    END
  END ONB[78]
  PIN ON[79]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 100.030 23.715 100.320 26.190 ;
    END
  END ON[79]
  PIN ONB[79]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 99.480 23.715 99.770 26.190 ;
    END
  END ONB[79]
  PIN ON[80]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 98.030 23.715 98.320 26.190 ;
    END
  END ON[80]
  PIN ONB[80]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 97.480 23.715 97.770 26.190 ;
    END
  END ONB[80]
  PIN ON[81]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 96.030 23.715 96.320 26.190 ;
    END
  END ON[81]
  PIN ONB[81]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 95.480 23.715 95.770 26.190 ;
    END
  END ONB[81]
  PIN ON[82]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 94.030 23.715 94.320 26.190 ;
    END
  END ON[82]
  PIN ONB[82]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 93.480 23.715 93.770 26.190 ;
    END
  END ONB[82]
  PIN ON[83]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 92.030 23.715 92.320 26.190 ;
    END
  END ON[83]
  PIN ONB[83]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 91.480 23.715 91.770 26.190 ;
    END
  END ONB[83]
  PIN ON[84]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 90.030 23.715 90.320 26.190 ;
    END
  END ON[84]
  PIN ONB[84]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 89.480 23.715 89.770 26.190 ;
    END
  END ONB[84]
  PIN ON[85]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 88.030 23.715 88.320 26.190 ;
    END
  END ON[85]
  PIN ONB[85]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 87.480 23.715 87.770 26.190 ;
    END
  END ONB[85]
  PIN ON[86]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 86.030 23.715 86.320 26.190 ;
    END
  END ON[86]
  PIN ONB[86]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 85.480 23.715 85.770 26.190 ;
    END
  END ONB[86]
  PIN ON[87]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 84.030 23.715 84.320 26.190 ;
    END
  END ON[87]
  PIN ONB[87]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 83.480 23.715 83.770 26.190 ;
    END
  END ONB[87]
  PIN ON[88]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 82.030 23.715 82.320 26.190 ;
    END
  END ON[88]
  PIN ONB[88]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 81.480 23.715 81.770 26.190 ;
    END
  END ONB[88]
  PIN ON[89]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 80.030 23.715 80.320 26.190 ;
    END
  END ON[89]
  PIN ONB[89]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 79.480 23.715 79.770 26.190 ;
    END
  END ONB[89]
  PIN ON[90]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 78.030 23.715 78.320 26.190 ;
    END
  END ON[90]
  PIN ONB[90]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.480 23.715 77.770 26.190 ;
    END
  END ONB[90]
  PIN ON[91]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 76.030 23.715 76.320 26.190 ;
    END
  END ON[91]
  PIN ONB[91]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 75.480 23.715 75.770 26.190 ;
    END
  END ONB[91]
  PIN ON[92]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 74.030 23.715 74.320 26.190 ;
    END
  END ON[92]
  PIN ONB[92]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 73.480 23.715 73.770 26.190 ;
    END
  END ONB[92]
  PIN ON[93]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 72.030 23.715 72.320 26.190 ;
    END
  END ON[93]
  PIN ONB[93]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 71.480 23.715 71.770 26.190 ;
    END
  END ONB[93]
  PIN ON[94]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.030 23.715 70.320 26.190 ;
    END
  END ON[94]
  PIN ONB[94]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.480 23.715 69.770 26.190 ;
    END
  END ONB[94]
  PIN ON[95]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.030 23.715 68.320 26.190 ;
    END
  END ON[95]
  PIN ONB[95]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 67.480 23.715 67.770 26.190 ;
    END
  END ONB[95]
  PIN ON[96]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 66.030 23.715 66.320 26.190 ;
    END
  END ON[96]
  PIN ONB[96]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 65.480 23.715 65.770 26.190 ;
    END
  END ONB[96]
  PIN ON[97]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.030 23.715 64.320 26.190 ;
    END
  END ON[97]
  PIN ONB[97]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.480 23.715 63.770 26.190 ;
    END
  END ONB[97]
  PIN ON[98]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 62.030 23.715 62.320 26.190 ;
    END
  END ON[98]
  PIN ONB[98]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 61.480 23.715 61.770 26.190 ;
    END
  END ONB[98]
  PIN ON[99]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 60.030 23.715 60.320 26.190 ;
    END
  END ON[99]
  PIN ONB[99]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 59.480 23.715 59.770 26.190 ;
    END
  END ONB[99]
  PIN ON[100]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 58.030 23.715 58.320 26.190 ;
    END
  END ON[100]
  PIN ONB[100]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.480 23.715 57.770 26.190 ;
    END
  END ONB[100]
  PIN ON[101]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 56.030 23.715 56.320 26.190 ;
    END
  END ON[101]
  PIN ONB[101]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 55.480 23.715 55.770 26.190 ;
    END
  END ONB[101]
  PIN ON[102]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 54.030 23.715 54.320 26.190 ;
    END
  END ON[102]
  PIN ONB[102]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 53.480 23.715 53.770 26.190 ;
    END
  END ONB[102]
  PIN ON[103]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 52.030 23.715 52.320 26.190 ;
    END
  END ON[103]
  PIN ONB[103]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 51.480 23.715 51.770 26.190 ;
    END
  END ONB[103]
  PIN ON[104]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 50.030 23.715 50.320 26.190 ;
    END
  END ON[104]
  PIN ONB[104]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 49.480 23.715 49.770 26.190 ;
    END
  END ONB[104]
  PIN ON[105]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 48.030 23.715 48.320 26.190 ;
    END
  END ON[105]
  PIN ONB[105]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 47.480 23.715 47.770 26.190 ;
    END
  END ONB[105]
  PIN ON[106]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 46.030 23.715 46.320 26.190 ;
    END
  END ON[106]
  PIN ONB[106]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 45.480 23.715 45.770 26.190 ;
    END
  END ONB[106]
  PIN ON[107]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 44.030 23.715 44.320 26.190 ;
    END
  END ON[107]
  PIN ONB[107]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 43.480 23.715 43.770 26.190 ;
    END
  END ONB[107]
  PIN ON[108]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 42.030 23.715 42.320 26.190 ;
    END
  END ON[108]
  PIN ONB[108]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 41.480 23.715 41.770 26.190 ;
    END
  END ONB[108]
  PIN ON[109]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 40.030 23.715 40.320 26.190 ;
    END
  END ON[109]
  PIN ONB[109]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 39.480 23.715 39.770 26.190 ;
    END
  END ONB[109]
  PIN ON[110]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 38.030 23.715 38.320 26.190 ;
    END
  END ON[110]
  PIN ONB[110]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 37.480 23.715 37.770 26.190 ;
    END
  END ONB[110]
  PIN ON[111]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.030 23.715 36.320 26.190 ;
    END
  END ON[111]
  PIN ONB[111]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 35.480 23.715 35.770 26.190 ;
    END
  END ONB[111]
  PIN ON[112]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 34.030 23.715 34.320 26.190 ;
    END
  END ON[112]
  PIN ONB[112]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 33.480 23.715 33.770 26.190 ;
    END
  END ONB[112]
  PIN ON[113]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 32.030 23.715 32.320 26.190 ;
    END
  END ON[113]
  PIN ONB[113]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 31.480 23.715 31.770 26.190 ;
    END
  END ONB[113]
  PIN ON[114]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.030 23.715 30.320 26.190 ;
    END
  END ON[114]
  PIN ONB[114]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 29.480 23.715 29.770 26.190 ;
    END
  END ONB[114]
  PIN ON[115]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.030 23.715 28.320 26.190 ;
    END
  END ON[115]
  PIN ONB[115]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 27.480 23.715 27.770 26.190 ;
    END
  END ONB[115]
  PIN ON[116]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 26.030 23.715 26.320 26.190 ;
    END
  END ON[116]
  PIN ONB[116]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.480 23.715 25.770 26.190 ;
    END
  END ONB[116]
  PIN ON[117]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 24.030 23.715 24.320 26.190 ;
    END
  END ON[117]
  PIN ONB[117]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 23.480 23.715 23.770 26.190 ;
    END
  END ONB[117]
  PIN ON[118]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 22.030 23.715 22.320 26.190 ;
    END
  END ON[118]
  PIN ONB[118]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.480 23.715 21.770 26.190 ;
    END
  END ONB[118]
  PIN ON[119]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 20.030 23.715 20.320 26.190 ;
    END
  END ON[119]
  PIN ONB[119]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 19.480 23.715 19.770 26.190 ;
    END
  END ONB[119]
  PIN ON[120]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 18.030 23.715 18.320 26.190 ;
    END
  END ON[120]
  PIN ONB[120]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.480 23.715 17.770 26.190 ;
    END
  END ONB[120]
  PIN ON[121]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.030 23.715 16.320 26.190 ;
    END
  END ON[121]
  PIN ONB[121]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 15.480 23.715 15.770 26.190 ;
    END
  END ONB[121]
  PIN ON[122]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.030 23.715 14.320 26.190 ;
    END
  END ON[122]
  PIN ONB[122]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.480 23.715 13.770 26.190 ;
    END
  END ONB[122]
  PIN EN[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.030 23.715 2.320 26.190 ;
    END
  END EN[3]
  PIN ENB[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.480 23.715 1.770 26.190 ;
    END
  END ENB[3]
  PIN ON[123]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.030 23.715 12.320 26.190 ;
    END
  END ON[123]
  PIN ONB[123]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.480 23.715 11.770 26.190 ;
    END
  END ONB[123]
  PIN ON[124]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.030 23.715 10.320 26.190 ;
    END
  END ON[124]
  PIN ONB[124]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.480 23.715 9.770 26.190 ;
    END
  END ONB[124]
  PIN ON[125]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 8.030 23.715 8.320 26.190 ;
    END
  END ON[125]
  PIN ONB[125]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.480 23.715 7.770 26.190 ;
    END
  END ONB[125]
  PIN ON[126]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 6.030 23.715 6.320 26.190 ;
    END
  END ON[126]
  PIN ONB[126]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.480 23.715 5.770 26.190 ;
    END
  END ONB[126]
  PIN ON[127]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 4.030 23.715 4.320 26.190 ;
    END
  END ON[127]
  PIN ONB[127]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.480 23.715 3.770 26.190 ;
    END
  END ONB[127]
  PIN ON[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.480 0.000 3.770 2.475 ;
    END
  END ON[0]
  PIN ONB[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 4.030 0.000 4.320 2.475 ;
    END
  END ONB[0]
  PIN ON[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.480 0.000 5.770 2.475 ;
    END
  END ON[1]
  PIN ONB[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 6.030 0.000 6.320 2.475 ;
    END
  END ONB[1]
  PIN ON[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.480 0.000 7.770 2.475 ;
    END
  END ON[2]
  PIN ONB[2]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 8.030 0.000 8.320 2.475 ;
    END
  END ONB[2]
  PIN ON[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 9.480 0.000 9.770 2.475 ;
    END
  END ON[3]
  PIN ONB[3]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.030 0.000 10.320 2.475 ;
    END
  END ONB[3]
  PIN ON[4]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.480 0.000 11.770 2.475 ;
    END
  END ON[4]
  PIN ONB[4]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 12.030 0.000 12.320 2.475 ;
    END
  END ONB[4]
  PIN ON[5]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 13.480 0.000 13.770 2.475 ;
    END
  END ON[5]
  PIN ONB[5]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 14.030 0.000 14.320 2.475 ;
    END
  END ONB[5]
  PIN ON[6]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 15.480 0.000 15.770 2.475 ;
    END
  END ON[6]
  PIN EN[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.480 0.000 1.770 2.475 ;
    END
  END EN[0]
  PIN ENB[0]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 2.030 0.000 2.320 2.475 ;
    END
  END ENB[0]
  PIN ONB[6]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 16.030 0.000 16.320 2.475 ;
    END
  END ONB[6]
  PIN ON[7]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 17.480 0.000 17.770 2.475 ;
    END
  END ON[7]
  PIN ONB[7]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 18.030 0.000 18.320 2.475 ;
    END
  END ONB[7]
  PIN ON[8]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 19.480 0.000 19.770 2.475 ;
    END
  END ON[8]
  PIN ONB[8]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 20.030 0.000 20.320 2.475 ;
    END
  END ONB[8]
  PIN ON[9]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 21.480 0.000 21.770 2.475 ;
    END
  END ON[9]
  PIN ONB[9]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 22.030 0.000 22.320 2.475 ;
    END
  END ONB[9]
  PIN ON[10]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 23.480 0.000 23.770 2.475 ;
    END
  END ON[10]
  PIN ONB[10]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 24.030 0.000 24.320 2.475 ;
    END
  END ONB[10]
  PIN ON[11]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.480 0.000 25.770 2.475 ;
    END
  END ON[11]
  PIN ONB[11]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 26.030 0.000 26.320 2.475 ;
    END
  END ONB[11]
  PIN ON[12]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 27.480 0.000 27.770 2.475 ;
    END
  END ON[12]
  PIN ONB[12]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.030 0.000 28.320 2.475 ;
    END
  END ONB[12]
  PIN ON[13]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 29.480 0.000 29.770 2.475 ;
    END
  END ON[13]
  PIN ONB[13]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.030 0.000 30.320 2.475 ;
    END
  END ONB[13]
  PIN ON[14]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 31.480 0.000 31.770 2.475 ;
    END
  END ON[14]
  PIN ONB[14]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 32.030 0.000 32.320 2.475 ;
    END
  END ONB[14]
  PIN ON[15]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 33.480 0.000 33.770 2.475 ;
    END
  END ON[15]
  PIN ONB[15]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 34.030 0.000 34.320 2.475 ;
    END
  END ONB[15]
  PIN ON[16]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 35.480 0.000 35.770 2.475 ;
    END
  END ON[16]
  PIN ONB[16]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 36.030 0.000 36.320 2.475 ;
    END
  END ONB[16]
  PIN ON[17]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 37.480 0.000 37.770 2.475 ;
    END
  END ON[17]
  PIN ONB[17]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 38.030 0.000 38.320 2.475 ;
    END
  END ONB[17]
  PIN ON[18]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 39.480 0.000 39.770 2.475 ;
    END
  END ON[18]
  PIN ONB[18]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 40.030 0.000 40.320 2.475 ;
    END
  END ONB[18]
  PIN ON[19]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 41.480 0.000 41.770 2.475 ;
    END
  END ON[19]
  PIN ONB[19]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 42.030 0.000 42.320 2.475 ;
    END
  END ONB[19]
  PIN ON[20]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 43.480 0.000 43.770 2.475 ;
    END
  END ON[20]
  PIN ONB[20]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 44.030 0.000 44.320 2.475 ;
    END
  END ONB[20]
  PIN ON[21]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 45.480 0.000 45.770 2.475 ;
    END
  END ON[21]
  PIN ONB[21]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 46.030 0.000 46.320 2.475 ;
    END
  END ONB[21]
  PIN ON[22]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 47.480 0.000 47.770 2.475 ;
    END
  END ON[22]
  PIN ONB[22]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 48.030 0.000 48.320 2.475 ;
    END
  END ONB[22]
  PIN ON[23]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 49.480 0.000 49.770 2.475 ;
    END
  END ON[23]
  PIN ONB[23]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 50.030 0.000 50.320 2.475 ;
    END
  END ONB[23]
  PIN ON[24]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 51.480 0.000 51.770 2.475 ;
    END
  END ON[24]
  PIN ONB[24]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 52.030 0.000 52.320 2.475 ;
    END
  END ONB[24]
  PIN ON[25]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 53.480 0.000 53.770 2.475 ;
    END
  END ON[25]
  PIN ONB[25]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 54.030 0.000 54.320 2.475 ;
    END
  END ONB[25]
  PIN ON[26]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 55.480 0.000 55.770 2.475 ;
    END
  END ON[26]
  PIN ONB[26]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 56.030 0.000 56.320 2.475 ;
    END
  END ONB[26]
  PIN ON[27]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.480 0.000 57.770 2.475 ;
    END
  END ON[27]
  PIN ONB[27]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 58.030 0.000 58.320 2.475 ;
    END
  END ONB[27]
  PIN ON[28]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 59.480 0.000 59.770 2.475 ;
    END
  END ON[28]
  PIN ONB[28]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 60.030 0.000 60.320 2.475 ;
    END
  END ONB[28]
  PIN ON[29]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 61.480 0.000 61.770 2.475 ;
    END
  END ON[29]
  PIN ONB[29]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 62.030 0.000 62.320 2.475 ;
    END
  END ONB[29]
  PIN ON[30]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.480 0.000 63.770 2.475 ;
    END
  END ON[30]
  PIN ONB[30]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.030 0.000 64.320 2.475 ;
    END
  END ONB[30]
  PIN ON[31]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 65.480 0.000 65.770 2.475 ;
    END
  END ON[31]
  PIN ONB[31]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 66.030 0.000 66.320 2.475 ;
    END
  END ONB[31]
  PIN ON[33]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.480 0.000 69.770 2.475 ;
    END
  END ON[33]
  PIN ONB[33]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.030 0.000 70.320 2.475 ;
    END
  END ONB[33]
  PIN ON[32]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 67.480 0.000 67.770 2.475 ;
    END
  END ON[32]
  PIN ONB[32]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.030 0.000 68.320 2.475 ;
    END
  END ONB[32]
  PIN ON[34]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 71.480 0.000 71.770 2.475 ;
    END
  END ON[34]
  PIN ONB[34]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 72.030 0.000 72.320 2.475 ;
    END
  END ONB[34]
  PIN ON[35]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 73.480 0.000 73.770 2.475 ;
    END
  END ON[35]
  PIN ONB[35]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 74.030 0.000 74.320 2.475 ;
    END
  END ONB[35]
  PIN ON[36]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 75.480 0.000 75.770 2.475 ;
    END
  END ON[36]
  PIN ONB[36]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 76.030 0.000 76.320 2.475 ;
    END
  END ONB[36]
  PIN ON[37]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 77.480 0.000 77.770 2.475 ;
    END
  END ON[37]
  PIN ONB[37]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 78.030 0.000 78.320 2.475 ;
    END
  END ONB[37]
  PIN ON[38]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 79.480 0.000 79.770 2.475 ;
    END
  END ON[38]
  PIN ONB[38]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 80.030 0.000 80.320 2.475 ;
    END
  END ONB[38]
  PIN ON[39]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 81.480 0.000 81.770 2.475 ;
    END
  END ON[39]
  PIN ONB[39]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 82.030 0.000 82.320 2.475 ;
    END
  END ONB[39]
  PIN ON[40]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 83.480 0.000 83.770 2.475 ;
    END
  END ON[40]
  PIN ONB[40]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 84.030 0.000 84.320 2.475 ;
    END
  END ONB[40]
  PIN ON[41]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 85.480 0.000 85.770 2.475 ;
    END
  END ON[41]
  PIN ONB[41]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 86.030 0.000 86.320 2.475 ;
    END
  END ONB[41]
  PIN ON[42]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 87.480 0.000 87.770 2.475 ;
    END
  END ON[42]
  PIN ONB[42]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 88.030 0.000 88.320 2.475 ;
    END
  END ONB[42]
  PIN ON[43]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 89.480 0.000 89.770 2.475 ;
    END
  END ON[43]
  PIN ONB[43]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 90.030 0.000 90.320 2.475 ;
    END
  END ONB[43]
  PIN ON[44]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 91.480 0.000 91.770 2.475 ;
    END
  END ON[44]
  PIN ONB[44]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 92.030 0.000 92.320 2.475 ;
    END
  END ONB[44]
  PIN ON[45]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 93.480 0.000 93.770 2.475 ;
    END
  END ON[45]
  PIN ONB[45]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 94.030 0.000 94.320 2.475 ;
    END
  END ONB[45]
  PIN ON[46]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 95.480 0.000 95.770 2.475 ;
    END
  END ON[46]
  PIN ONB[46]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 96.030 0.000 96.320 2.475 ;
    END
  END ONB[46]
  PIN ON[47]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 97.480 0.000 97.770 2.475 ;
    END
  END ON[47]
  PIN ONB[47]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 98.030 0.000 98.320 2.475 ;
    END
  END ONB[47]
  PIN ON[48]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 99.480 0.000 99.770 2.475 ;
    END
  END ON[48]
  PIN ONB[48]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 100.030 0.000 100.320 2.475 ;
    END
  END ONB[48]
  PIN ON[49]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 101.480 0.000 101.770 2.475 ;
    END
  END ON[49]
  PIN ONB[49]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 102.030 0.000 102.320 2.475 ;
    END
  END ONB[49]
  PIN ON[50]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 103.480 0.000 103.770 2.475 ;
    END
  END ON[50]
  PIN ONB[50]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 104.030 0.000 104.320 2.475 ;
    END
  END ONB[50]
  PIN ON[51]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 105.480 0.000 105.770 2.475 ;
    END
  END ON[51]
  PIN ONB[51]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 106.030 0.000 106.320 2.475 ;
    END
  END ONB[51]
  PIN ON[52]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 107.480 0.000 107.770 2.475 ;
    END
  END ON[52]
  PIN ONB[52]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 108.030 0.000 108.320 2.475 ;
    END
  END ONB[52]
  PIN ON[53]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 109.480 0.000 109.770 2.475 ;
    END
  END ON[53]
  PIN ONB[53]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.030 0.000 110.320 2.475 ;
    END
  END ONB[53]
  PIN ON[54]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 111.480 0.000 111.770 2.475 ;
    END
  END ON[54]
  PIN ONB[54]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 112.030 0.000 112.320 2.475 ;
    END
  END ONB[54]
  PIN ON[55]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 113.480 0.000 113.770 2.475 ;
    END
  END ON[55]
  PIN ONB[55]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 114.030 0.000 114.320 2.475 ;
    END
  END ONB[55]
  PIN ON[56]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 115.480 0.000 115.770 2.475 ;
    END
  END ON[56]
  PIN ONB[56]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 116.030 0.000 116.320 2.475 ;
    END
  END ONB[56]
  PIN ON[57]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.480 0.000 117.770 2.475 ;
    END
  END ON[57]
  PIN ONB[57]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.030 0.000 118.320 2.475 ;
    END
  END ONB[57]
  PIN ON[58]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 119.480 0.000 119.770 2.475 ;
    END
  END ON[58]
  PIN ONB[58]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 120.030 0.000 120.320 2.475 ;
    END
  END ONB[58]
  PIN ON[59]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 121.480 0.000 121.770 2.475 ;
    END
  END ON[59]
  PIN ONB[59]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 122.030 0.000 122.320 2.475 ;
    END
  END ONB[59]
  PIN ON[60]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 123.480 0.000 123.770 2.475 ;
    END
  END ON[60]
  PIN ONB[60]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 124.030 0.000 124.320 2.475 ;
    END
  END ONB[60]
  PIN ON[61]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 125.480 0.000 125.770 2.475 ;
    END
  END ON[61]
  PIN ONB[61]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 126.030 0.000 126.320 2.475 ;
    END
  END ONB[61]
  PIN ON[62]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 127.480 0.000 127.770 2.475 ;
    END
  END ON[62]
  PIN ONB[62]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 128.030 0.000 128.320 2.475 ;
    END
  END ONB[62]
  PIN ON[63]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 129.480 0.000 129.770 2.475 ;
    END
  END ON[63]
  PIN ONB[63]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 130.030 0.000 130.320 2.475 ;
    END
  END ONB[63]
  PIN EN[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 131.480 0.000 131.770 2.475 ;
    END
  END EN[1]
  PIN ENB[1]
    ANTENNAGATEAREA 0.039000 ;
    PORT
      LAYER Metal2 ;
        RECT 132.030 0.000 132.320 2.475 ;
    END
  END ENB[1]
  PIN VcascP[1]
    ANTENNAGATEAREA 1.755000 ;
    ANTENNADIFFAREA 10.710000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.930 133.800 21.630 ;
    END
  END VcascP[1]
  PIN VcascP[0]
    ANTENNAGATEAREA 1.755000 ;
    ANTENNADIFFAREA 10.710000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 4.560 133.800 5.260 ;
    END
  END VcascP[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 0.000 14.380 133.800 26.190 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 0.000 0.000 133.800 11.810 ;
    END
  END VDD
  OBS
      LAYER GatPoly ;
        RECT 0.000 -0.070 133.800 26.260 ;
      LAYER Metal1 ;
        RECT 0.000 20.060 133.800 26.190 ;
        RECT 0.000 14.770 0.720 20.060 ;
        RECT 133.080 14.770 133.800 20.060 ;
        RECT 0.000 13.625 133.800 14.770 ;
        RECT 0.000 11.420 133.800 12.565 ;
        RECT 0.000 6.130 0.720 11.420 ;
        RECT 133.080 6.130 133.800 11.420 ;
        RECT 0.000 0.000 133.800 6.130 ;
      LAYER Metal2 ;
        RECT 0.005 23.505 1.270 26.190 ;
        RECT 2.530 23.505 3.270 26.190 ;
        RECT 4.530 23.505 5.270 26.190 ;
        RECT 6.530 23.505 7.270 26.190 ;
        RECT 8.530 23.505 9.270 26.190 ;
        RECT 10.530 23.505 11.270 26.190 ;
        RECT 12.530 23.505 13.270 26.190 ;
        RECT 14.530 23.505 15.270 26.190 ;
        RECT 16.530 23.505 17.270 26.190 ;
        RECT 18.530 23.505 19.270 26.190 ;
        RECT 20.530 23.505 21.270 26.190 ;
        RECT 22.530 23.505 23.270 26.190 ;
        RECT 24.530 23.505 25.270 26.190 ;
        RECT 26.530 23.505 27.270 26.190 ;
        RECT 28.530 23.505 29.270 26.190 ;
        RECT 30.530 23.505 31.270 26.190 ;
        RECT 32.530 23.505 33.270 26.190 ;
        RECT 34.530 23.505 35.270 26.190 ;
        RECT 36.530 23.505 37.270 26.190 ;
        RECT 38.530 23.505 39.270 26.190 ;
        RECT 40.530 23.505 41.270 26.190 ;
        RECT 42.530 23.505 43.270 26.190 ;
        RECT 44.530 23.505 45.270 26.190 ;
        RECT 46.530 23.505 47.270 26.190 ;
        RECT 48.530 23.505 49.270 26.190 ;
        RECT 50.530 23.505 51.270 26.190 ;
        RECT 52.530 23.505 53.270 26.190 ;
        RECT 54.530 23.505 55.270 26.190 ;
        RECT 56.530 23.505 57.270 26.190 ;
        RECT 58.530 23.505 59.270 26.190 ;
        RECT 60.530 23.505 61.270 26.190 ;
        RECT 62.530 23.505 63.270 26.190 ;
        RECT 64.530 23.505 65.270 26.190 ;
        RECT 66.530 23.505 67.270 26.190 ;
        RECT 68.530 23.505 69.270 26.190 ;
        RECT 70.530 23.505 71.270 26.190 ;
        RECT 72.530 23.505 73.270 26.190 ;
        RECT 74.530 23.505 75.270 26.190 ;
        RECT 76.530 23.505 77.270 26.190 ;
        RECT 78.530 23.505 79.270 26.190 ;
        RECT 80.530 23.505 81.270 26.190 ;
        RECT 82.530 23.505 83.270 26.190 ;
        RECT 84.530 23.505 85.270 26.190 ;
        RECT 86.530 23.505 87.270 26.190 ;
        RECT 88.530 23.505 89.270 26.190 ;
        RECT 90.530 23.505 91.270 26.190 ;
        RECT 92.530 23.505 93.270 26.190 ;
        RECT 94.530 23.505 95.270 26.190 ;
        RECT 96.530 23.505 97.270 26.190 ;
        RECT 98.530 23.505 99.270 26.190 ;
        RECT 100.530 23.505 101.270 26.190 ;
        RECT 102.530 23.505 103.270 26.190 ;
        RECT 104.530 23.505 105.270 26.190 ;
        RECT 106.530 23.505 107.270 26.190 ;
        RECT 108.530 23.505 109.270 26.190 ;
        RECT 110.530 23.505 111.270 26.190 ;
        RECT 112.530 23.505 113.270 26.190 ;
        RECT 114.530 23.505 115.270 26.190 ;
        RECT 116.530 23.505 117.270 26.190 ;
        RECT 118.530 23.505 119.270 26.190 ;
        RECT 120.530 23.505 121.270 26.190 ;
        RECT 122.530 23.505 123.270 26.190 ;
        RECT 124.530 23.505 125.270 26.190 ;
        RECT 126.530 23.505 127.270 26.190 ;
        RECT 128.530 23.505 129.270 26.190 ;
        RECT 130.530 23.505 131.270 26.190 ;
        RECT 132.530 23.505 133.795 26.190 ;
        RECT 0.005 2.685 133.795 23.505 ;
        RECT 0.005 0.000 1.270 2.685 ;
        RECT 2.530 0.000 3.270 2.685 ;
        RECT 4.530 0.000 5.270 2.685 ;
        RECT 6.530 0.000 7.270 2.685 ;
        RECT 8.530 0.000 9.270 2.685 ;
        RECT 10.530 0.000 11.270 2.685 ;
        RECT 12.530 0.000 13.270 2.685 ;
        RECT 14.530 0.000 15.270 2.685 ;
        RECT 16.530 0.000 17.270 2.685 ;
        RECT 18.530 0.000 19.270 2.685 ;
        RECT 20.530 0.000 21.270 2.685 ;
        RECT 22.530 0.000 23.270 2.685 ;
        RECT 24.530 0.000 25.270 2.685 ;
        RECT 26.530 0.000 27.270 2.685 ;
        RECT 28.530 0.000 29.270 2.685 ;
        RECT 30.530 0.000 31.270 2.685 ;
        RECT 32.530 0.000 33.270 2.685 ;
        RECT 34.530 0.000 35.270 2.685 ;
        RECT 36.530 0.000 37.270 2.685 ;
        RECT 38.530 0.000 39.270 2.685 ;
        RECT 40.530 0.000 41.270 2.685 ;
        RECT 42.530 0.000 43.270 2.685 ;
        RECT 44.530 0.000 45.270 2.685 ;
        RECT 46.530 0.000 47.270 2.685 ;
        RECT 48.530 0.000 49.270 2.685 ;
        RECT 50.530 0.000 51.270 2.685 ;
        RECT 52.530 0.000 53.270 2.685 ;
        RECT 54.530 0.000 55.270 2.685 ;
        RECT 56.530 0.000 57.270 2.685 ;
        RECT 58.530 0.000 59.270 2.685 ;
        RECT 60.530 0.000 61.270 2.685 ;
        RECT 62.530 0.000 63.270 2.685 ;
        RECT 64.530 0.000 65.270 2.685 ;
        RECT 66.530 0.000 67.270 2.685 ;
        RECT 68.530 0.000 69.270 2.685 ;
        RECT 70.530 0.000 71.270 2.685 ;
        RECT 72.530 0.000 73.270 2.685 ;
        RECT 74.530 0.000 75.270 2.685 ;
        RECT 76.530 0.000 77.270 2.685 ;
        RECT 78.530 0.000 79.270 2.685 ;
        RECT 80.530 0.000 81.270 2.685 ;
        RECT 82.530 0.000 83.270 2.685 ;
        RECT 84.530 0.000 85.270 2.685 ;
        RECT 86.530 0.000 87.270 2.685 ;
        RECT 88.530 0.000 89.270 2.685 ;
        RECT 90.530 0.000 91.270 2.685 ;
        RECT 92.530 0.000 93.270 2.685 ;
        RECT 94.530 0.000 95.270 2.685 ;
        RECT 96.530 0.000 97.270 2.685 ;
        RECT 98.530 0.000 99.270 2.685 ;
        RECT 100.530 0.000 101.270 2.685 ;
        RECT 102.530 0.000 103.270 2.685 ;
        RECT 104.530 0.000 105.270 2.685 ;
        RECT 106.530 0.000 107.270 2.685 ;
        RECT 108.530 0.000 109.270 2.685 ;
        RECT 110.530 0.000 111.270 2.685 ;
        RECT 112.530 0.000 113.270 2.685 ;
        RECT 114.530 0.000 115.270 2.685 ;
        RECT 116.530 0.000 117.270 2.685 ;
        RECT 118.530 0.000 119.270 2.685 ;
        RECT 120.530 0.000 121.270 2.685 ;
        RECT 122.530 0.000 123.270 2.685 ;
        RECT 124.530 0.000 125.270 2.685 ;
        RECT 126.530 0.000 127.270 2.685 ;
        RECT 128.530 0.000 129.270 2.685 ;
        RECT 130.530 0.000 131.270 2.685 ;
        RECT 132.530 0.000 133.795 2.685 ;
      LAYER Metal3 ;
        RECT 0.000 21.840 133.800 26.190 ;
        RECT 0.000 5.470 133.800 20.720 ;
        RECT 0.000 0.000 133.800 4.350 ;
      LAYER Metal4 ;
        RECT 0.000 0.000 133.800 26.190 ;
  END
END dac128module
END LIBRARY

