** sch_path: /foss/designs/PUDDING_dev_leardilap/analog/non_overlap/xschem/non_overlap_single_tran_sim.sch
**.subckt non_overlap_single_tran_sim
Vdd net1 GND 1.5
Vthermo thermo GND dc 0 ac 0 pulse(0, 1.5, 0, 100p, 100p, 10n, 20n, 5)
x1 thermo ON net1 GND ON_N non_overlap
**** begin user architecture code

.lib cornerMOSlv.lib mos_ff
.include sg13g2_stdcell.spice



.param temp=127
.control
save all
tran 50p 200n
meas tran tdelay TRIG v(thermo) VAl=0.9 FALl=1 TARG v(ON) VAl=0.9 RISE=1
write non_overlap_tran_logic.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  non_overlap.sym # of pins=5
** sym_path: /foss/designs/PUDDING_dev_leardilap/analog/non_overlap/xschem/non_overlap.sym
** sch_path: /foss/designs/PUDDING_dev_leardilap/analog/non_overlap/xschem/non_overlap.sch
.subckt non_overlap thermo ON VDD VSS ON_N
*.iopin VSS
*.ipin thermo
*.opin ON
*.opin ON_N
*.iopin VDD
x0 thermon thermo VDD VSS sg13g2_inv_1
x1 a1 thermo b2 VDD VSS sg13g2_nor2_1
x2 b1 a2 thermon VDD VSS sg13g2_nor2_1
x3 a2 a1 VDD VSS sg13g2_dlygate4sd3_1
x4 b2 b1 VDD VSS sg13g2_dlygate4sd3_1
x5 ON_N a2 VDD VSS sg13g2_buf_1
x6 ON b2 VDD VSS sg13g2_buf_1
.ends

.GLOBAL GND
.end
