* Extracted by KLayout with SG13G2 LVS runset on : 31/08/2025 07:57

.SUBCKT DAC2U128OUT4IN
M$1 \$536 \$537 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$2 \$1 \$536 \$537 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$3 \$2 \$3 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p PS=2.16u
+ PD=1.14u
M$4 \$1 \$2 \$3 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p PS=1.14u
+ PD=2.16u
M$5 \$538 \$539 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$6 \$1 \$538 \$539 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$7 \$4 \$5 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p PS=2.16u
+ PD=1.14u
M$8 \$1 \$4 \$5 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p PS=1.14u
+ PD=2.16u
M$9 \$540 \$541 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$10 \$1 \$540 \$541 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$11 \$6 \$7 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p PS=2.16u
+ PD=1.14u
M$12 \$1 \$6 \$7 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p PS=1.14u
+ PD=2.16u
M$13 \$542 \$543 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$14 \$1 \$542 \$543 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$15 \$8 \$9 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p PS=2.16u
+ PD=1.14u
M$16 \$1 \$8 \$9 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p PS=1.14u
+ PD=2.16u
M$17 \$10 \$11 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$18 \$1 \$10 \$11 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$19 \$544 \$545 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$20 \$1 \$544 \$545 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$21 \$12 \$13 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$22 \$1 \$12 \$13 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$23 \$546 \$547 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$24 \$1 \$546 \$547 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$25 \$14 \$15 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$26 \$1 \$14 \$15 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$27 \$548 \$549 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$28 \$1 \$548 \$549 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$29 \$16 \$17 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$30 \$1 \$16 \$17 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$31 \$550 \$551 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$32 \$1 \$550 \$551 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$33 \$18 \$19 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$34 \$1 \$18 \$19 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$35 \$552 \$553 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$36 \$1 \$552 \$553 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$37 \$20 \$21 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$38 \$1 \$20 \$21 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$39 \$554 \$555 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$40 \$1 \$554 \$555 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$41 \$556 \$557 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$42 \$1 \$556 \$557 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$43 \$22 \$23 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$44 \$1 \$22 \$23 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$45 \$558 \$559 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$46 \$1 \$558 \$559 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$47 \$24 \$25 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$48 \$1 \$24 \$25 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$49 \$26 \$27 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$50 \$1 \$26 \$27 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$51 \$560 \$561 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$52 \$1 \$560 \$561 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$53 \$562 \$563 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$54 \$1 \$562 \$563 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$55 \$28 \$29 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$56 \$1 \$28 \$29 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$57 \$564 \$565 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$58 \$1 \$564 \$565 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$59 \$30 \$31 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$60 \$1 \$30 \$31 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$61 \$32 \$33 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$62 \$1 \$32 \$33 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$63 \$566 \$567 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$64 \$1 \$566 \$567 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$65 \$34 \$35 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$66 \$1 \$34 \$35 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$67 \$568 \$569 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$68 \$1 \$568 \$569 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$69 \$570 \$571 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$70 \$1 \$570 \$571 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$71 \$36 \$37 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$72 \$1 \$36 \$37 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$73 \$572 \$573 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$74 \$1 \$572 \$573 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$75 \$38 \$39 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$76 \$1 \$38 \$39 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$77 \$574 \$575 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$78 \$1 \$574 \$575 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$79 \$40 \$41 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$80 \$1 \$40 \$41 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$81 \$576 \$577 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$82 \$1 \$576 \$577 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$83 \$42 \$43 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$84 \$1 \$42 \$43 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$85 \$44 \$45 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$86 \$1 \$44 \$45 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$87 \$578 \$579 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$88 \$1 \$578 \$579 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$89 \$46 \$47 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$90 \$1 \$46 \$47 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$91 \$580 \$581 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$92 \$1 \$580 \$581 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$93 \$48 \$49 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$94 \$1 \$48 \$49 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$95 \$582 \$583 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$96 \$1 \$582 \$583 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$97 \$584 \$585 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$98 \$1 \$584 \$585 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$99 \$50 \$51 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$100 \$1 \$50 \$51 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$101 \$586 \$587 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$102 \$1 \$586 \$587 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$103 \$52 \$53 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$104 \$1 \$52 \$53 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$105 \$54 \$55 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$106 \$1 \$54 \$55 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$107 \$588 \$589 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$108 \$1 \$588 \$589 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$109 \$590 \$591 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$110 \$1 \$590 \$591 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$111 \$56 \$57 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$112 \$1 \$56 \$57 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$113 \$58 \$59 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$114 \$1 \$58 \$59 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$115 \$592 \$593 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$116 \$1 \$592 \$593 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$117 \$594 \$595 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$118 \$1 \$594 \$595 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$119 \$60 \$61 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$120 \$1 \$60 \$61 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$121 \$62 \$63 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$122 \$1 \$62 \$63 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$123 \$596 \$597 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$124 \$1 \$596 \$597 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$125 \$598 \$599 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$126 \$1 \$598 \$599 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$127 \$64 \$65 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$128 \$1 \$64 \$65 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$129 \$600 \$601 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$130 \$1 \$600 \$601 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$131 \$66 \$67 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$132 \$1 \$66 \$67 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$133 \$68 \$69 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$134 \$1 \$68 \$69 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$135 \$602 \$603 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$136 \$1 \$602 \$603 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$137 \$604 \$605 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$138 \$1 \$604 \$605 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$139 \$70 \$71 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$140 \$1 \$70 \$71 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$141 \$72 \$73 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$142 \$1 \$72 \$73 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$143 \$606 \$607 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$144 \$1 \$606 \$607 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$145 \$608 \$609 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$146 \$1 \$608 \$609 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$147 \$74 \$75 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$148 \$1 \$74 \$75 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$149 \$610 \$611 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$150 \$1 \$610 \$611 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$151 \$76 \$77 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$152 \$1 \$76 \$77 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$153 \$78 \$79 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$154 \$1 \$78 \$79 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$155 \$612 \$613 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$156 \$1 \$612 \$613 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$157 \$80 \$81 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$158 \$1 \$80 \$81 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$159 \$614 \$615 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$160 \$1 \$614 \$615 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$161 \$616 \$617 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$162 \$1 \$616 \$617 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$163 \$82 \$83 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$164 \$1 \$82 \$83 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$165 \$618 \$619 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$166 \$1 \$618 \$619 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$167 \$84 \$85 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$168 \$1 \$84 \$85 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$169 \$86 \$87 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$170 \$1 \$86 \$87 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$171 \$620 \$621 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$172 \$1 \$620 \$621 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$173 \$622 \$623 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$174 \$1 \$622 \$623 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$175 \$88 \$89 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$176 \$1 \$88 \$89 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$177 \$90 \$91 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$178 \$1 \$90 \$91 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$179 \$624 \$625 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$180 \$1 \$624 \$625 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$181 \$92 \$93 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$182 \$1 \$92 \$93 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$183 \$626 \$627 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$184 \$1 \$626 \$627 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$185 \$628 \$629 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$186 \$1 \$628 \$629 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$187 \$94 \$95 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$188 \$1 \$94 \$95 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$189 \$630 \$631 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$190 \$1 \$630 \$631 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$191 \$96 \$97 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$192 \$1 \$96 \$97 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$193 \$98 \$99 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$194 \$1 \$98 \$99 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$195 \$632 \$633 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$196 \$1 \$632 \$633 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$197 \$634 \$635 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$198 \$1 \$634 \$635 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$199 \$100 \$101 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$200 \$1 \$100 \$101 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$201 \$636 \$637 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$202 \$1 \$636 \$637 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$203 \$102 \$103 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$204 \$1 \$102 \$103 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$205 \$104 \$105 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$206 \$1 \$104 \$105 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$207 \$638 \$639 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$208 \$1 \$638 \$639 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$209 \$106 \$107 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$210 \$1 \$106 \$107 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$211 \$640 \$641 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$212 \$1 \$640 \$641 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$213 \$108 \$109 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$214 \$1 \$108 \$109 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$215 \$642 \$643 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$216 \$1 \$642 \$643 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$217 \$644 \$645 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$218 \$1 \$644 \$645 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$219 \$110 \$111 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$220 \$1 \$110 \$111 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$221 \$112 \$113 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$222 \$1 \$112 \$113 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$223 \$646 \$647 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$224 \$1 \$646 \$647 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$225 \$648 \$649 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$226 \$1 \$648 \$649 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$227 \$114 \$115 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$228 \$1 \$114 \$115 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$229 \$116 \$117 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$230 \$1 \$116 \$117 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$231 \$650 \$651 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$232 \$1 \$650 \$651 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$233 \$652 \$653 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$234 \$1 \$652 \$653 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$235 \$118 \$119 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$236 \$1 \$118 \$119 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$237 \$120 \$121 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$238 \$1 \$120 \$121 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$239 \$654 \$655 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$240 \$1 \$654 \$655 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$241 \$656 \$657 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$242 \$1 \$656 \$657 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$243 \$122 \$123 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$244 \$1 \$122 \$123 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$245 \$658 \$659 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$246 \$1 \$658 \$659 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$247 \$124 \$125 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$248 \$1 \$124 \$125 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$249 \$126 \$127 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$250 \$1 \$126 \$127 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$251 \$660 \$661 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$252 \$1 \$660 \$661 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$253 \$128 \$129 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$254 \$1 \$128 \$129 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$255 \$662 \$663 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$256 \$1 \$662 \$663 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$257 \$130 \$131 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$258 \$1 \$130 \$131 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$259 \$664 \$665 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$260 \$1 \$664 \$665 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$261 \$132 \$133 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$262 \$1 \$132 \$133 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$263 \$666 \$667 \$1 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.162p AD=0.0855p
+ PS=2.16u PD=1.14u
M$264 \$1 \$666 \$667 \$1 sg13_lv_nmos L=0.52u W=0.15u AS=0.0855p AD=0.162p
+ PS=1.14u PD=2.16u
M$265 \$2 \$134 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$266 \$266 \$135 \$3 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$267 \$4 \$136 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$268 \$266 \$137 \$5 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$269 \$6 \$138 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$270 \$266 \$139 \$7 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$271 \$8 \$140 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$272 \$266 \$141 \$9 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$273 \$10 \$142 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$274 \$266 \$143 \$11 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$275 \$12 \$144 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$276 \$266 \$145 \$13 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$277 \$14 \$146 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$278 \$266 \$147 \$15 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$279 \$16 \$148 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$280 \$266 \$149 \$17 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$281 \$18 \$150 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$282 \$266 \$151 \$19 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$283 \$20 \$152 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$284 \$266 \$153 \$21 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$285 \$22 \$154 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$286 \$266 \$155 \$23 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$287 \$24 \$156 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$288 \$266 \$157 \$25 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$289 \$26 \$158 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$290 \$266 \$159 \$27 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$291 \$28 \$160 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$292 \$266 \$161 \$29 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$293 \$30 \$162 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$294 \$266 \$163 \$31 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$295 \$32 \$164 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$296 \$266 \$165 \$33 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$297 \$34 \$166 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$298 \$266 \$167 \$35 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$299 \$36 \$168 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$300 \$266 \$169 \$37 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$301 \$38 \$170 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$302 \$266 \$171 \$39 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$303 \$40 \$172 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$304 \$266 \$173 \$41 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$305 \$42 \$174 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$306 \$266 \$175 \$43 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$307 \$44 \$176 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$308 \$266 \$177 \$45 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$309 \$46 \$178 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$310 \$266 \$179 \$47 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$311 \$48 \$180 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$312 \$266 \$181 \$49 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$313 \$50 \$182 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$314 \$266 \$183 \$51 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$315 \$52 \$184 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$316 \$266 \$185 \$53 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$317 \$54 \$186 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$318 \$266 \$187 \$55 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$319 \$56 \$188 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$320 \$266 \$189 \$57 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$321 \$58 \$190 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$322 \$266 \$191 \$59 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$323 \$60 \$192 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$324 \$266 \$193 \$61 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$325 \$62 \$194 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$326 \$266 \$195 \$63 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$327 \$64 \$196 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$328 \$266 \$197 \$65 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$329 \$66 \$198 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$330 \$266 \$199 \$67 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$331 \$68 \$200 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$332 \$266 \$201 \$69 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$333 \$70 \$202 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$334 \$266 \$203 \$71 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$335 \$72 \$204 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$336 \$266 \$205 \$73 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$337 \$74 \$206 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$338 \$266 \$207 \$75 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$339 \$76 \$208 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$340 \$266 \$209 \$77 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$341 \$78 \$210 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$342 \$266 \$211 \$79 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$343 \$80 \$212 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$344 \$266 \$213 \$81 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$345 \$82 \$214 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$346 \$266 \$215 \$83 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$347 \$84 \$216 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$348 \$266 \$217 \$85 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$349 \$86 \$218 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$350 \$266 \$219 \$87 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$351 \$88 \$220 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$352 \$266 \$221 \$89 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$353 \$90 \$222 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$354 \$266 \$223 \$91 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$355 \$92 \$224 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$356 \$266 \$225 \$93 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$357 \$94 \$226 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$358 \$266 \$227 \$95 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$359 \$96 \$228 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$360 \$266 \$229 \$97 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$361 \$98 \$230 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$362 \$266 \$231 \$99 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$363 \$100 \$232 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$364 \$266 \$233 \$101 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$365 \$102 \$234 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$366 \$266 \$235 \$103 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$367 \$104 \$236 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$368 \$266 \$237 \$105 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$369 \$106 \$238 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$370 \$266 \$239 \$107 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$371 \$108 \$240 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$372 \$266 \$241 \$109 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$373 \$110 \$242 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$374 \$266 \$243 \$111 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$375 \$112 \$244 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$376 \$266 \$245 \$113 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$377 \$114 \$246 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$378 \$266 \$247 \$115 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$379 \$116 \$248 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$380 \$266 \$249 \$117 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$381 \$118 \$250 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$382 \$266 \$251 \$119 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$383 \$120 \$252 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$384 \$266 \$253 \$121 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$385 \$122 \$254 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$386 \$266 \$255 \$123 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$387 \$124 \$256 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$388 \$266 \$257 \$125 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$389 \$126 \$258 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$390 \$266 \$259 \$127 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$391 \$128 \$260 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$392 \$266 \$261 \$129 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$393 \$130 \$262 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$394 \$266 \$263 \$131 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$395 \$132 \$264 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$396 \$266 \$265 \$133 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$397 \$267 \$2 \$268 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$398 \$268 \$3 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$399 \$267 \$4 \$269 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$400 \$269 \$5 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$401 \$267 \$6 \$270 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$402 \$270 \$7 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$403 \$267 \$8 \$271 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$404 \$271 \$9 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$405 \$267 \$10 \$272 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$406 \$272 \$11 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$407 \$267 \$12 \$273 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$408 \$273 \$13 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$409 \$267 \$14 \$274 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$410 \$274 \$15 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$411 \$267 \$16 \$275 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$412 \$275 \$17 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$413 \$267 \$18 \$276 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$414 \$276 \$19 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$415 \$267 \$20 \$277 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$416 \$277 \$21 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$417 \$267 \$22 \$278 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$418 \$278 \$23 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$419 \$267 \$24 \$279 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$420 \$279 \$25 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$421 \$267 \$26 \$280 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$422 \$280 \$27 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$423 \$267 \$28 \$281 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$424 \$281 \$29 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$425 \$267 \$30 \$282 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$426 \$282 \$31 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$427 \$267 \$32 \$283 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$428 \$283 \$33 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$429 \$267 \$34 \$284 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$430 \$284 \$35 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$431 \$267 \$36 \$285 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$432 \$285 \$37 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$433 \$267 \$38 \$286 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$434 \$286 \$39 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$435 \$267 \$40 \$287 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$436 \$287 \$41 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$437 \$267 \$42 \$288 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$438 \$288 \$43 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$439 \$267 \$44 \$289 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$440 \$289 \$45 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$441 \$267 \$46 \$290 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$442 \$290 \$47 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$443 \$267 \$48 \$291 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$444 \$291 \$49 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$445 \$267 \$50 \$292 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$446 \$292 \$51 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$447 \$267 \$52 \$293 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$448 \$293 \$53 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$449 \$267 \$54 \$294 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$450 \$294 \$55 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$451 \$267 \$56 \$295 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$452 \$295 \$57 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$453 \$267 \$58 \$296 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$454 \$296 \$59 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$455 \$267 \$60 \$297 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$456 \$297 \$61 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$457 \$267 \$62 \$298 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$458 \$298 \$63 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$459 \$267 \$64 \$299 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$460 \$299 \$65 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$461 \$267 \$66 \$300 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$462 \$300 \$67 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$463 \$267 \$68 \$301 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$464 \$301 \$69 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$465 \$267 \$70 \$302 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$466 \$302 \$71 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$467 \$267 \$72 \$303 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$468 \$303 \$73 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$469 \$267 \$74 \$304 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$470 \$304 \$75 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$471 \$267 \$76 \$305 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$472 \$305 \$77 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$473 \$267 \$78 \$306 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$474 \$306 \$79 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$475 \$267 \$80 \$307 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$476 \$307 \$81 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$477 \$267 \$82 \$308 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$478 \$308 \$83 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$479 \$267 \$84 \$309 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$480 \$309 \$85 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$481 \$267 \$86 \$310 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$482 \$310 \$87 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$483 \$267 \$88 \$311 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$484 \$311 \$89 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$485 \$267 \$90 \$312 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$486 \$312 \$91 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$487 \$267 \$92 \$313 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$488 \$313 \$93 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$489 \$267 \$94 \$314 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$490 \$314 \$95 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$491 \$267 \$96 \$315 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$492 \$315 \$97 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$493 \$267 \$98 \$316 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$494 \$316 \$99 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$495 \$267 \$100 \$317 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$496 \$317 \$101 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$497 \$267 \$102 \$318 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$498 \$318 \$103 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$499 \$267 \$104 \$319 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$500 \$319 \$105 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$501 \$267 \$106 \$320 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$502 \$320 \$107 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$503 \$267 \$108 \$321 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$504 \$321 \$109 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$505 \$267 \$110 \$322 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$506 \$322 \$111 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$507 \$267 \$112 \$323 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$508 \$323 \$113 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$509 \$267 \$114 \$324 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$510 \$324 \$115 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$511 \$267 \$116 \$325 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$512 \$325 \$117 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$513 \$267 \$118 \$326 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$514 \$326 \$119 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$515 \$267 \$120 \$327 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$516 \$327 \$121 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$517 \$267 \$122 \$328 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$518 \$328 \$123 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$519 \$267 \$124 \$329 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$520 \$329 \$125 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$521 \$267 \$126 \$330 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$522 \$330 \$127 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$523 \$267 \$128 \$331 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$524 \$331 \$129 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$525 \$267 \$130 \$332 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$526 \$332 \$131 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$527 \$267 \$132 \$333 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$528 \$333 \$133 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$529 \$267 \$267 \$334 \$266 sg13_lv_pmos L=0.15u W=11.7u AS=3.978p AD=3.978p
+ PS=24.76u PD=24.76u
M$530 \$266 \$334 \$346 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$531 \$346 \$268 \$334 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$532 \$266 \$334 \$338 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$533 \$338 \$269 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$534 \$266 \$334 \$349 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$535 \$349 \$270 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$536 \$266 \$334 \$354 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$537 \$354 \$271 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$538 \$266 \$334 \$359 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$539 \$359 \$272 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$540 \$266 \$334 \$364 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$541 \$364 \$273 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$542 \$266 \$334 \$369 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$543 \$369 \$274 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$544 \$266 \$334 \$374 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$545 \$374 \$275 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$546 \$266 \$334 \$379 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$547 \$379 \$276 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$548 \$266 \$334 \$384 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$549 \$384 \$277 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$550 \$266 \$334 \$389 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$551 \$389 \$278 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$552 \$266 \$334 \$394 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$553 \$394 \$279 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$554 \$266 \$334 \$399 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$555 \$399 \$280 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$556 \$266 \$334 \$400 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$557 \$400 \$281 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$558 \$266 \$334 \$398 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$559 \$398 \$282 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$560 \$266 \$334 \$397 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$561 \$397 \$283 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$562 \$266 \$334 \$396 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$563 \$396 \$284 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$564 \$266 \$334 \$395 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$565 \$395 \$285 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$566 \$266 \$334 \$393 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$567 \$393 \$286 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$568 \$266 \$334 \$392 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$569 \$392 \$287 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$570 \$266 \$334 \$391 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$571 \$391 \$288 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$572 \$266 \$334 \$390 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$573 \$390 \$289 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$574 \$266 \$334 \$388 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$575 \$388 \$290 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$576 \$266 \$334 \$387 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$577 \$387 \$291 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$578 \$266 \$334 \$386 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$579 \$386 \$292 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$580 \$266 \$334 \$385 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$581 \$385 \$293 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$582 \$266 \$334 \$383 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$583 \$383 \$294 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$584 \$266 \$334 \$382 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$585 \$382 \$295 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$586 \$266 \$334 \$381 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$587 \$381 \$296 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$588 \$266 \$334 \$380 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$589 \$380 \$297 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$590 \$266 \$334 \$378 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$591 \$378 \$298 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$592 \$266 \$334 \$377 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$593 \$377 \$299 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$594 \$266 \$334 \$376 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$595 \$376 \$300 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$596 \$266 \$334 \$375 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$597 \$375 \$301 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$598 \$266 \$334 \$373 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$599 \$373 \$302 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$600 \$266 \$334 \$372 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$601 \$372 \$303 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$602 \$266 \$334 \$371 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$603 \$371 \$304 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$604 \$266 \$334 \$370 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$605 \$370 \$305 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$606 \$266 \$334 \$368 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$607 \$368 \$306 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$608 \$266 \$334 \$367 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$609 \$367 \$307 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$610 \$266 \$334 \$366 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$611 \$366 \$308 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$612 \$266 \$334 \$365 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$613 \$365 \$309 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$614 \$266 \$334 \$363 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$615 \$363 \$310 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$616 \$266 \$334 \$362 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$617 \$362 \$311 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$618 \$266 \$334 \$361 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$619 \$361 \$312 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$620 \$266 \$334 \$360 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$621 \$360 \$313 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$622 \$266 \$334 \$358 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$623 \$358 \$314 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$624 \$266 \$334 \$357 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$625 \$357 \$315 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$626 \$266 \$334 \$356 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$627 \$356 \$316 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$628 \$266 \$334 \$355 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$629 \$355 \$317 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$630 \$266 \$334 \$353 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$631 \$353 \$318 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$632 \$266 \$334 \$352 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$633 \$352 \$319 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$634 \$266 \$334 \$351 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$635 \$351 \$320 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$636 \$266 \$334 \$350 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$637 \$350 \$321 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$638 \$266 \$334 \$348 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$639 \$348 \$322 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$640 \$266 \$334 \$347 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$641 \$347 \$323 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$642 \$266 \$334 \$345 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$643 \$345 \$324 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$644 \$266 \$334 \$344 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$645 \$344 \$325 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$646 \$266 \$334 \$343 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$647 \$343 \$326 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$648 \$266 \$334 \$342 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$649 \$342 \$327 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$650 \$266 \$334 \$341 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$651 \$341 \$328 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$652 \$266 \$334 \$340 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$653 \$340 \$329 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$654 \$266 \$334 \$339 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$655 \$339 \$330 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$656 \$266 \$334 \$337 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$657 \$337 \$331 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$658 \$266 \$334 \$336 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$659 \$336 \$332 \$401 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$660 \$266 \$334 \$335 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.493p AD=0.20875p
+ PS=3.58u PD=1.75u
M$661 \$335 \$333 \$334 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.20875p AD=0.516p
+ PS=1.75u PD=3.26u
M$663 \$402 \$402 \$403 \$266 sg13_lv_pmos L=0.15u W=11.7u AS=3.978p AD=3.978p
+ PS=24.76u PD=24.76u
M$664 \$403 \$404 \$470 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$665 \$470 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$666 \$401 \$407 \$472 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$667 \$472 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$668 \$401 \$410 \$476 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$669 \$476 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$670 \$401 \$411 \$479 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$671 \$479 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$672 \$401 \$412 \$481 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$673 \$481 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$674 \$401 \$413 \$480 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$675 \$480 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$676 \$401 \$414 \$482 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$677 \$482 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$678 \$401 \$418 \$489 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$679 \$489 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$680 \$401 \$419 \$488 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$681 \$488 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$682 \$401 \$421 \$493 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$683 \$493 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$684 \$401 \$423 \$494 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$685 \$494 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$686 \$401 \$424 \$496 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$687 \$496 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$688 \$401 \$425 \$495 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$689 \$495 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$690 \$401 \$429 \$503 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$691 \$503 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$692 \$401 \$430 \$505 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$693 \$505 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$694 \$401 \$431 \$504 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$695 \$504 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$696 \$401 \$433 \$508 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$697 \$508 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$698 \$401 \$434 \$507 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$699 \$507 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$700 \$401 \$435 \$511 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$701 \$511 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$702 \$401 \$437 \$512 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$703 \$512 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$704 \$401 \$439 \$517 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$705 \$517 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$706 \$401 \$440 \$516 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$707 \$516 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$708 \$401 \$441 \$518 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$709 \$518 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$710 \$401 \$442 \$521 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$711 \$521 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$712 \$401 \$443 \$519 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$713 \$519 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$714 \$401 \$445 \$525 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$715 \$525 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$716 \$401 \$446 \$524 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$717 \$524 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$718 \$401 \$447 \$527 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$719 \$527 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$720 \$401 \$450 \$530 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$721 \$530 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$722 \$401 \$451 \$532 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$723 \$532 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$724 \$401 \$452 \$531 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$725 \$531 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$726 \$401 \$453 \$535 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$727 \$535 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$728 \$401 \$455 \$534 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$729 \$534 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$730 \$401 \$457 \$520 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$731 \$520 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$732 \$401 \$459 \$514 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$733 \$514 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$734 \$401 \$460 \$509 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$735 \$509 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$736 \$401 \$461 \$510 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$737 \$510 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$738 \$401 \$462 \$502 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$739 \$502 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$740 \$401 \$465 \$490 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$741 \$490 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$742 \$401 \$466 \$484 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$743 \$484 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$744 \$401 \$468 \$478 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$745 \$478 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$746 \$403 \$469 \$474 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$747 \$474 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$749 \$401 \$405 \$471 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$750 \$471 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$751 \$401 \$406 \$473 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$752 \$473 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$753 \$401 \$408 \$475 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$754 \$475 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$755 \$401 \$409 \$477 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$756 \$477 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$757 \$401 \$415 \$485 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$758 \$485 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$759 \$401 \$416 \$483 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$760 \$483 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$761 \$401 \$417 \$487 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$762 \$487 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$763 \$401 \$420 \$491 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$764 \$491 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$765 \$401 \$422 \$492 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$766 \$492 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$767 \$401 \$426 \$499 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$768 \$499 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$769 \$401 \$427 \$501 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$770 \$501 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$771 \$401 \$428 \$500 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$772 \$500 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$773 \$401 \$432 \$506 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$774 \$506 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$775 \$401 \$436 \$513 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$776 \$513 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$777 \$401 \$438 \$515 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$778 \$515 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$779 \$401 \$444 \$523 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$780 \$523 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$781 \$401 \$448 \$529 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$782 \$529 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$783 \$401 \$449 \$528 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$784 \$528 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$785 \$401 \$454 \$533 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$786 \$533 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$787 \$401 \$456 \$526 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$788 \$526 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$789 \$401 \$458 \$522 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$790 \$522 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$791 \$401 \$463 \$497 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$792 \$497 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$793 \$401 \$464 \$498 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$794 \$498 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$795 \$401 \$467 \$486 \$266 sg13_lv_pmos L=0.6u W=1.2u AS=0.516p AD=0.20875p
+ PS=3.26u PD=1.75u
M$796 \$486 \$403 \$266 \$266 sg13_lv_pmos L=5u W=1.45u AS=0.20875p AD=0.493p
+ PS=1.75u PD=3.58u
M$797 \$266 \$536 \$404 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$798 \$404 \$537 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$799 \$266 \$538 \$405 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$800 \$405 \$539 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$801 \$266 \$540 \$406 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$802 \$406 \$541 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$803 \$266 \$542 \$407 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$804 \$407 \$543 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$805 \$266 \$544 \$408 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$806 \$408 \$545 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$807 \$266 \$546 \$409 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$808 \$409 \$547 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$809 \$266 \$548 \$410 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$810 \$410 \$549 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$811 \$266 \$550 \$411 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$812 \$411 \$551 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$813 \$266 \$552 \$412 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$814 \$412 \$553 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$815 \$266 \$554 \$413 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$816 \$413 \$555 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$817 \$266 \$556 \$414 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$818 \$414 \$557 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$819 \$266 \$558 \$415 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$820 \$415 \$559 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$821 \$266 \$560 \$416 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$822 \$416 \$561 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$823 \$266 \$562 \$417 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$824 \$417 \$563 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$825 \$266 \$564 \$418 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$826 \$418 \$565 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$827 \$266 \$566 \$419 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$828 \$419 \$567 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$829 \$266 \$568 \$420 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$830 \$420 \$569 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$831 \$266 \$570 \$421 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$832 \$421 \$571 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$833 \$266 \$572 \$422 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$834 \$422 \$573 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$835 \$266 \$574 \$423 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$836 \$423 \$575 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$837 \$266 \$576 \$424 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$838 \$424 \$577 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$839 \$266 \$578 \$425 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$840 \$425 \$579 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$841 \$266 \$580 \$426 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$842 \$426 \$581 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$843 \$266 \$582 \$427 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$844 \$427 \$583 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$845 \$266 \$584 \$428 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$846 \$428 \$585 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$847 \$266 \$586 \$429 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$848 \$429 \$587 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$849 \$266 \$588 \$430 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$850 \$430 \$589 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$851 \$266 \$590 \$431 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$852 \$431 \$591 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$853 \$266 \$592 \$432 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$854 \$432 \$593 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$855 \$266 \$594 \$433 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$856 \$433 \$595 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$857 \$266 \$596 \$434 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$858 \$434 \$597 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$859 \$266 \$598 \$435 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$860 \$435 \$599 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$861 \$266 \$600 \$436 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$862 \$436 \$601 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$863 \$266 \$602 \$437 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$864 \$437 \$603 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$865 \$266 \$604 \$438 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$866 \$438 \$605 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$867 \$266 \$606 \$439 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$868 \$439 \$607 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$869 \$266 \$608 \$440 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$870 \$440 \$609 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$871 \$266 \$610 \$441 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$872 \$441 \$611 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$873 \$266 \$612 \$442 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$874 \$442 \$613 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$875 \$266 \$614 \$443 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$876 \$443 \$615 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$877 \$266 \$616 \$444 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$878 \$444 \$617 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$879 \$266 \$618 \$445 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$880 \$445 \$619 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$881 \$266 \$620 \$446 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$882 \$446 \$621 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$883 \$266 \$622 \$447 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$884 \$447 \$623 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$885 \$266 \$624 \$448 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$886 \$448 \$625 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$887 \$266 \$626 \$449 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$888 \$449 \$627 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$889 \$266 \$628 \$450 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$890 \$450 \$629 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$891 \$266 \$630 \$451 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$892 \$451 \$631 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$893 \$266 \$632 \$452 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$894 \$452 \$633 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$895 \$266 \$634 \$453 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$896 \$453 \$635 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$897 \$266 \$636 \$454 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$898 \$454 \$637 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$899 \$266 \$638 \$455 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$900 \$455 \$639 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$901 \$266 \$640 \$456 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$902 \$456 \$641 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$903 \$266 \$642 \$457 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$904 \$457 \$643 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$905 \$266 \$644 \$458 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$906 \$458 \$645 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$907 \$266 \$646 \$459 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$908 \$459 \$647 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$909 \$266 \$648 \$460 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$910 \$460 \$649 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$911 \$266 \$650 \$461 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$912 \$461 \$651 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$913 \$266 \$652 \$462 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$914 \$462 \$653 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$915 \$266 \$654 \$463 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$916 \$463 \$655 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$917 \$266 \$656 \$464 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$918 \$464 \$657 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$919 \$266 \$658 \$465 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$920 \$465 \$659 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$921 \$266 \$660 \$466 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$922 \$466 \$661 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$923 \$266 \$662 \$467 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$924 \$467 \$663 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$925 \$266 \$664 \$468 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$926 \$468 \$665 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$927 \$266 \$666 \$469 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$928 \$469 \$667 \$402 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
M$929 \$536 \$668 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$930 \$266 \$669 \$537 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$931 \$538 \$670 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$932 \$266 \$671 \$539 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$933 \$540 \$672 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$934 \$266 \$673 \$541 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$935 \$542 \$674 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$936 \$266 \$675 \$543 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$937 \$544 \$676 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$938 \$266 \$677 \$545 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$939 \$546 \$678 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$940 \$266 \$679 \$547 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$941 \$548 \$680 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$942 \$266 \$681 \$549 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$943 \$550 \$682 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$944 \$266 \$683 \$551 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$945 \$552 \$684 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$946 \$266 \$685 \$553 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$947 \$554 \$686 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$948 \$266 \$687 \$555 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$949 \$556 \$688 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$950 \$266 \$689 \$557 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$951 \$558 \$690 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$952 \$266 \$691 \$559 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$953 \$560 \$692 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$954 \$266 \$693 \$561 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$955 \$562 \$694 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$956 \$266 \$695 \$563 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$957 \$564 \$696 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$958 \$266 \$697 \$565 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$959 \$566 \$698 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$960 \$266 \$699 \$567 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$961 \$568 \$700 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$962 \$266 \$701 \$569 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$963 \$570 \$702 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$964 \$266 \$703 \$571 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$965 \$572 \$704 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$966 \$266 \$705 \$573 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$967 \$574 \$706 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$968 \$266 \$707 \$575 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$969 \$576 \$708 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$970 \$266 \$709 \$577 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$971 \$578 \$710 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$972 \$266 \$711 \$579 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$973 \$580 \$712 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$974 \$266 \$713 \$581 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$975 \$582 \$714 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$976 \$266 \$715 \$583 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$977 \$584 \$716 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$978 \$266 \$717 \$585 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$979 \$586 \$718 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$980 \$266 \$719 \$587 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$981 \$588 \$720 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$982 \$266 \$721 \$589 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$983 \$590 \$722 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$984 \$266 \$723 \$591 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$985 \$592 \$724 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$986 \$266 \$725 \$593 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$987 \$594 \$726 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$988 \$266 \$727 \$595 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$989 \$596 \$728 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$990 \$266 \$729 \$597 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$991 \$598 \$730 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$992 \$266 \$731 \$599 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$993 \$600 \$732 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$994 \$266 \$733 \$601 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$995 \$602 \$734 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$996 \$266 \$735 \$603 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$997 \$604 \$736 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$998 \$266 \$737 \$605 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$999 \$606 \$738 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1000 \$266 \$739 \$607 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1001 \$608 \$740 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1002 \$266 \$741 \$609 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1003 \$610 \$742 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1004 \$266 \$743 \$611 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1005 \$612 \$744 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1006 \$266 \$745 \$613 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1007 \$614 \$746 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1008 \$266 \$747 \$615 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1009 \$616 \$748 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1010 \$266 \$749 \$617 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1011 \$618 \$750 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1012 \$266 \$751 \$619 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1013 \$620 \$752 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1014 \$266 \$753 \$621 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1015 \$622 \$754 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1016 \$266 \$755 \$623 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1017 \$624 \$756 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1018 \$266 \$757 \$625 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1019 \$626 \$758 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1020 \$266 \$759 \$627 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1021 \$628 \$760 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1022 \$266 \$761 \$629 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1023 \$630 \$762 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1024 \$266 \$763 \$631 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1025 \$632 \$764 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1026 \$266 \$765 \$633 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1027 \$634 \$766 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1028 \$266 \$767 \$635 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1029 \$636 \$768 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1030 \$266 \$769 \$637 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1031 \$638 \$770 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1032 \$266 \$771 \$639 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1033 \$640 \$772 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1034 \$266 \$773 \$641 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1035 \$642 \$774 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1036 \$266 \$775 \$643 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1037 \$644 \$776 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1038 \$266 \$777 \$645 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1039 \$646 \$778 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1040 \$266 \$779 \$647 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1041 \$648 \$780 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1042 \$266 \$781 \$649 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1043 \$650 \$782 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1044 \$266 \$783 \$651 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1045 \$652 \$784 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1046 \$266 \$785 \$653 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1047 \$654 \$786 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1048 \$266 \$787 \$655 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1049 \$656 \$788 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1050 \$266 \$789 \$657 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1051 \$658 \$790 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1052 \$266 \$791 \$659 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1053 \$660 \$792 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1054 \$266 \$793 \$661 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1055 \$662 \$794 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1056 \$266 \$795 \$663 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1057 \$664 \$796 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1058 \$266 \$797 \$665 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
M$1059 \$666 \$798 \$266 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.1725p AD=0.057p
+ PS=1.75u PD=0.68u
M$1060 \$266 \$799 \$667 \$266 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.1725p
+ PS=0.68u PD=1.75u
.ENDS DAC2U128OUT4IN
